
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_rom_pc, property_invalid_dec_rom_pc, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [15:0] PC_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire \oc8051_golden_model_1.n1046 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire \oc8051_golden_model_1.n1063 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1214 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire \oc8051_golden_model_1.n1300 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1424 ;
  wire \oc8051_golden_model_1.n1425 ;
  wire [4:0] \oc8051_golden_model_1.n1430 ;
  wire \oc8051_golden_model_1.n1431 ;
  wire \oc8051_golden_model_1.n1439 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1456 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [8:0] \oc8051_golden_model_1.n1461 ;
  wire \oc8051_golden_model_1.n1462 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire \oc8051_golden_model_1.n1475 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [8:0] \oc8051_golden_model_1.n1496 ;
  wire \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [8:0] \oc8051_golden_model_1.n1593 ;
  wire \oc8051_golden_model_1.n1594 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [4:0] \oc8051_golden_model_1.n1597 ;
  wire \oc8051_golden_model_1.n1598 ;
  wire \oc8051_golden_model_1.n1605 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1622 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [8:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire [4:0] \oc8051_golden_model_1.n1630 ;
  wire \oc8051_golden_model_1.n1631 ;
  wire \oc8051_golden_model_1.n1638 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1655 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire [6:0] \oc8051_golden_model_1.n1748 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1879 ;
  wire [6:0] \oc8051_golden_model_1.n1880 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire \oc8051_golden_model_1.n1936 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire \oc8051_golden_model_1.n1953 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire \oc8051_golden_model_1.n2085 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire \oc8051_golden_model_1.n2102 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire \oc8051_golden_model_1.n2141 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire \oc8051_golden_model_1.n2200 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2444 ;
  wire \oc8051_golden_model_1.n2446 ;
  wire \oc8051_golden_model_1.n2452 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [7:0] \oc8051_golden_model_1.n2734 ;
  wire [6:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire \oc8051_golden_model_1.n2853 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire \oc8051_golden_model_1.n2875 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire [7:0] \oc8051_golden_model_1.n2914 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc_impl;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dec_rom_pc;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_rom_pc;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_43998_, rst);
  not (_14673_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_14684_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_14695_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _14684_);
  and (_14706_, _14695_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_14717_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _14684_);
  and (_14728_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _14684_);
  nor (_14739_, _14728_, _14717_);
  and (_14750_, _14739_, _14706_);
  nor (_14761_, _14750_, _14673_);
  and (_14772_, _14673_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_14783_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_14794_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _14783_);
  nor (_14805_, _14794_, _14772_);
  not (_14816_, _14805_);
  and (_14827_, _14816_, _14750_);
  or (_14838_, _14827_, _14761_);
  and (_24751_, _14838_, _43998_);
  nor (_14858_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_14869_, _14858_);
  and (_14880_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_14891_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_14902_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_14913_, _14902_);
  not (_14924_, _14794_);
  nor (_14945_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_14946_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_14957_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14946_);
  nor (_14968_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_14979_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_14990_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _14979_);
  nor (_15001_, _14990_, _14968_);
  nor (_15012_, _15001_, _14957_);
  not (_15023_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15034_, _14957_, _15023_);
  nor (_15045_, _15034_, _15012_);
  and (_15056_, _15045_, _14945_);
  not (_15067_, _15056_);
  and (_15078_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15089_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_15100_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15111_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _15100_);
  and (_15122_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_15133_, _15122_, _15089_);
  and (_15144_, _15133_, _15067_);
  nor (_15155_, _15144_, _14924_);
  not (_15166_, _14772_);
  nor (_15177_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_15188_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _14979_);
  nor (_15199_, _15188_, _15177_);
  nor (_15209_, _15199_, _14957_);
  not (_15220_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_15231_, _14957_, _15220_);
  nor (_15242_, _15231_, _15209_);
  and (_15253_, _15242_, _14945_);
  not (_15264_, _15253_);
  and (_15275_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_15286_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15297_, _15286_, _15275_);
  and (_15308_, _15297_, _15264_);
  nor (_15319_, _15308_, _15166_);
  nor (_15330_, _15319_, _15155_);
  nor (_15341_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_15352_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _14979_);
  nor (_15363_, _15352_, _15341_);
  nor (_15374_, _15363_, _14957_);
  not (_15385_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_15396_, _14957_, _15385_);
  nor (_15407_, _15396_, _15374_);
  and (_15418_, _15407_, _14945_);
  not (_15429_, _15418_);
  and (_15440_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_15451_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_15462_, _15451_, _15440_);
  and (_15473_, _15462_, _15429_);
  nor (_15484_, _15473_, _14816_);
  nor (_15495_, _15484_, _14858_);
  and (_15506_, _15495_, _15330_);
  nor (_15517_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_15528_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _14979_);
  nor (_15539_, _15528_, _15517_);
  nor (_15549_, _15539_, _14957_);
  not (_15560_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_15571_, _14957_, _15560_);
  nor (_15582_, _15571_, _15549_);
  and (_15593_, _15582_, _14945_);
  not (_15604_, _15593_);
  and (_15615_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_15626_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_15637_, _15626_, _15615_);
  and (_15648_, _15637_, _15604_);
  and (_15659_, _15648_, _14858_);
  nor (_15670_, _15659_, _15506_);
  not (_15681_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_15692_, _15681_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15703_, _15692_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15714_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_15725_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15736_, _15725_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15747_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_15758_, _15747_, _15714_);
  nor (_15769_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15780_, _15769_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_15791_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_15802_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15813_, _15692_, _15802_);
  and (_15824_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_15835_, _15824_, _15791_);
  and (_15846_, _15835_, _15758_);
  and (_15857_, _15769_, _15681_);
  and (_15868_, _15857_, _15582_);
  and (_15878_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15889_, _15878_, _15802_);
  and (_15900_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_15911_, _15878_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15922_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_15933_, _15922_, _15900_);
  not (_15944_, _15933_);
  nor (_15955_, _15944_, _15868_);
  and (_15966_, _15955_, _15846_);
  not (_15977_, _15966_);
  and (_15988_, _15977_, _15670_);
  not (_15999_, _15988_);
  nor (_16010_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16021_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _14979_);
  nor (_16032_, _16021_, _16010_);
  nor (_16043_, _16032_, _14957_);
  not (_16054_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_16065_, _14957_, _16054_);
  nor (_16076_, _16065_, _16043_);
  and (_16087_, _16076_, _14945_);
  not (_16098_, _16087_);
  and (_16109_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_16120_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_16131_, _16120_, _16109_);
  and (_16142_, _16131_, _16098_);
  nor (_16153_, _16142_, _14924_);
  nor (_16164_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_16175_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _14979_);
  nor (_16186_, _16175_, _16164_);
  nor (_16197_, _16186_, _14957_);
  not (_16208_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_16218_, _14957_, _16208_);
  nor (_16229_, _16218_, _16197_);
  and (_16240_, _16229_, _14945_);
  not (_16251_, _16240_);
  and (_16262_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_16273_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16284_, _16273_, _16262_);
  and (_16295_, _16284_, _16251_);
  nor (_16306_, _16295_, _15166_);
  nor (_16317_, _16306_, _16153_);
  nor (_16328_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_16339_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _14979_);
  nor (_16350_, _16339_, _16328_);
  nor (_16361_, _16350_, _14957_);
  not (_16372_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_16383_, _14957_, _16372_);
  nor (_16394_, _16383_, _16361_);
  and (_16405_, _16394_, _14945_);
  not (_16416_, _16405_);
  and (_16427_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_16438_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_16449_, _16438_, _16427_);
  and (_16460_, _16449_, _16416_);
  nor (_16471_, _16460_, _14816_);
  nor (_16482_, _16471_, _14858_);
  and (_16493_, _16482_, _16317_);
  nor (_16504_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_16515_, _14979_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_16526_, _16515_, _16504_);
  nor (_16537_, _16526_, _14957_);
  not (_16547_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_16558_, _14957_, _16547_);
  nor (_16569_, _16558_, _16537_);
  and (_16580_, _16569_, _14945_);
  not (_16591_, _16580_);
  and (_16602_, _15078_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_16613_, _15111_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_16624_, _16613_, _16602_);
  and (_16634_, _16624_, _16591_);
  and (_16645_, _16634_, _14858_);
  nor (_16656_, _16645_, _16493_);
  and (_16667_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_16689_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_16690_, _16689_, _16667_);
  and (_16701_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_16712_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_16723_, _16712_, _16701_);
  and (_16733_, _16723_, _16690_);
  and (_16744_, _16569_, _15857_);
  and (_16755_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_16766_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_16777_, _16766_, _16755_);
  not (_16788_, _16777_);
  nor (_16799_, _16788_, _16744_);
  and (_16810_, _16799_, _16733_);
  not (_16821_, _16810_);
  and (_16831_, _16821_, _16656_);
  and (_16842_, _16831_, _15999_);
  not (_16853_, _16842_);
  and (_16864_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_16875_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_16886_, _16875_, _16864_);
  and (_16897_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_16908_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_16918_, _16908_, _16897_);
  and (_16929_, _16918_, _16886_);
  and (_16940_, _16229_, _15857_);
  and (_16951_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_16962_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16973_, _16962_, _16951_);
  not (_16984_, _16973_);
  nor (_16995_, _16984_, _16940_);
  and (_17006_, _16995_, _16929_);
  not (_17016_, _17006_);
  and (_17027_, _17016_, _16656_);
  and (_17038_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17049_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17060_, _17049_, _17038_);
  and (_17071_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_17082_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_17093_, _17082_, _17071_);
  and (_17104_, _17093_, _17060_);
  and (_17114_, _15857_, _15242_);
  and (_17125_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_17136_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_17147_, _17136_, _17125_);
  not (_17158_, _17147_);
  nor (_17169_, _17158_, _17114_);
  and (_17180_, _17169_, _17104_);
  not (_17191_, _17180_);
  and (_17201_, _17191_, _15670_);
  and (_17212_, _17027_, _17201_);
  and (_17223_, _15977_, _17212_);
  nor (_17234_, _15988_, _17212_);
  nor (_17245_, _17234_, _17223_);
  and (_17256_, _17245_, _17027_);
  and (_17267_, _16831_, _15988_);
  and (_17278_, _15977_, _16656_);
  and (_17288_, _16821_, _15670_);
  nor (_17299_, _17288_, _17278_);
  nor (_17310_, _17299_, _17267_);
  and (_17321_, _17310_, _17256_);
  nor (_17332_, _17310_, _17256_);
  nor (_17343_, _17332_, _17321_);
  and (_17354_, _17343_, _17223_);
  nor (_17365_, _17354_, _17321_);
  nor (_17376_, _17365_, _16853_);
  and (_17386_, _16656_, _17191_);
  and (_17407_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_17408_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_17429_, _17408_, _17407_);
  and (_17430_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_17441_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_17452_, _17441_, _17430_);
  and (_17463_, _17452_, _17429_);
  and (_17474_, _16076_, _15857_);
  and (_17484_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_17495_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17506_, _17495_, _17484_);
  not (_17517_, _17506_);
  nor (_17528_, _17517_, _17474_);
  and (_17539_, _17528_, _17463_);
  not (_17550_, _17539_);
  and (_17561_, _17550_, _15670_);
  and (_17571_, _17561_, _17386_);
  and (_17582_, _17016_, _15670_);
  nor (_17593_, _17582_, _17386_);
  nor (_17604_, _17593_, _17212_);
  and (_17615_, _17604_, _17571_);
  nor (_17626_, _15988_, _17027_);
  nor (_17637_, _17626_, _17256_);
  and (_17648_, _17637_, _17615_);
  nor (_17659_, _17343_, _17223_);
  nor (_17669_, _17659_, _17354_);
  and (_17680_, _17669_, _17648_);
  nor (_17691_, _17669_, _17648_);
  nor (_17702_, _17691_, _17680_);
  not (_17713_, _17702_);
  and (_17724_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_17735_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_17746_, _17735_, _17724_);
  and (_17757_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_17767_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_17778_, _17767_, _17757_);
  and (_17789_, _17778_, _17746_);
  and (_17800_, _16394_, _15857_);
  and (_17811_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_17822_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17833_, _17822_, _17811_);
  not (_17844_, _17833_);
  nor (_17854_, _17844_, _17800_);
  and (_17865_, _17854_, _17789_);
  not (_17876_, _17865_);
  and (_17887_, _17876_, _16656_);
  and (_17898_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_17909_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_17920_, _17909_, _17898_);
  and (_17931_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_17942_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_17953_, _17942_, _17931_);
  and (_17963_, _17953_, _17920_);
  and (_17974_, _15857_, _15045_);
  and (_17985_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_17996_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_18007_, _17996_, _17985_);
  not (_18018_, _18007_);
  nor (_18029_, _18018_, _17974_);
  and (_18040_, _18029_, _17963_);
  not (_18051_, _18040_);
  and (_18062_, _18051_, _15670_);
  and (_18073_, _18062_, _17887_);
  and (_18083_, _17876_, _15670_);
  not (_18094_, _18083_);
  and (_18105_, _18051_, _16656_);
  and (_18116_, _18105_, _18094_);
  and (_18127_, _18116_, _17561_);
  nor (_18138_, _18127_, _18073_);
  and (_18149_, _17550_, _16656_);
  nor (_18160_, _18149_, _17201_);
  nor (_18171_, _18160_, _17571_);
  not (_18182_, _18171_);
  nor (_18193_, _18182_, _18138_);
  nor (_18203_, _17604_, _17571_);
  nor (_18214_, _18203_, _17615_);
  and (_18225_, _18214_, _18193_);
  nor (_18236_, _17637_, _17615_);
  nor (_18247_, _18236_, _17648_);
  and (_18258_, _18247_, _18225_);
  and (_18269_, _15703_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_18280_, _15736_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_18291_, _18280_, _18269_);
  and (_18302_, _15780_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_18312_, _15813_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_18323_, _18312_, _18302_);
  and (_18334_, _18323_, _18291_);
  and (_18345_, _15857_, _15407_);
  and (_18356_, _15889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18367_, _15911_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_18378_, _18367_, _18356_);
  not (_18389_, _18378_);
  nor (_18400_, _18389_, _18345_);
  and (_18411_, _18400_, _18334_);
  not (_18422_, _18411_);
  and (_18432_, _18422_, _16656_);
  and (_18443_, _18432_, _18083_);
  nor (_18454_, _18062_, _17887_);
  nor (_18465_, _18454_, _18073_);
  and (_18476_, _18465_, _18443_);
  nor (_18487_, _18116_, _17561_);
  nor (_18498_, _18487_, _18127_);
  and (_18509_, _18498_, _18476_);
  and (_18520_, _18182_, _18138_);
  nor (_18531_, _18520_, _18193_);
  and (_18541_, _18531_, _18509_);
  nor (_18552_, _18214_, _18193_);
  nor (_18563_, _18552_, _18225_);
  and (_18574_, _18563_, _18541_);
  nor (_18585_, _18247_, _18225_);
  nor (_18596_, _18585_, _18258_);
  and (_18607_, _18596_, _18574_);
  nor (_18618_, _18607_, _18258_);
  nor (_18629_, _18618_, _17713_);
  nor (_18640_, _18629_, _17680_);
  and (_18651_, _17365_, _16853_);
  nor (_18661_, _18651_, _17376_);
  not (_18672_, _18661_);
  nor (_18683_, _18672_, _18640_);
  or (_18694_, _18683_, _17267_);
  nor (_18705_, _18694_, _17376_);
  nor (_18716_, _18705_, _14913_);
  and (_18727_, _18705_, _14913_);
  nor (_18738_, _18727_, _18716_);
  not (_18749_, _18738_);
  and (_18760_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_18770_, _18672_, _18640_);
  nor (_18781_, _18770_, _18683_);
  and (_18792_, _18781_, _18760_);
  and (_18803_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_18814_, _18618_, _17713_);
  nor (_18825_, _18814_, _18629_);
  and (_18836_, _18825_, _18803_);
  nor (_18847_, _18825_, _18803_);
  nor (_18858_, _18847_, _18836_);
  not (_18869_, _18858_);
  and (_18879_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_18890_, _18596_, _18574_);
  nor (_18901_, _18890_, _18607_);
  and (_18912_, _18901_, _18879_);
  nor (_18923_, _18901_, _18879_);
  nor (_18934_, _18923_, _18912_);
  not (_18945_, _18934_);
  and (_18956_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_18967_, _18563_, _18541_);
  nor (_18978_, _18967_, _18574_);
  and (_18989_, _18978_, _18956_);
  nor (_18999_, _18978_, _18956_);
  nor (_19010_, _18999_, _18989_);
  not (_19021_, _19010_);
  and (_19032_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19043_, _18531_, _18509_);
  nor (_19054_, _19043_, _18541_);
  and (_19065_, _19054_, _19032_);
  and (_19076_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_19087_, _18498_, _18476_);
  nor (_19098_, _19087_, _18509_);
  and (_19109_, _19098_, _19076_);
  and (_19119_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_19130_, _18465_, _18443_);
  nor (_19141_, _19130_, _18476_);
  and (_19152_, _19141_, _19119_);
  nor (_19163_, _19098_, _19076_);
  nor (_19174_, _19163_, _19109_);
  and (_19185_, _19174_, _19152_);
  nor (_19196_, _19185_, _19109_);
  not (_19207_, _19196_);
  nor (_19218_, _19054_, _19032_);
  nor (_19228_, _19218_, _19065_);
  and (_19239_, _19228_, _19207_);
  nor (_19250_, _19239_, _19065_);
  nor (_19261_, _19250_, _19021_);
  nor (_19272_, _19261_, _18989_);
  nor (_19283_, _19272_, _18945_);
  nor (_19294_, _19283_, _18912_);
  nor (_19305_, _19294_, _18869_);
  nor (_19316_, _19305_, _18836_);
  nor (_19327_, _18781_, _18760_);
  nor (_19338_, _19327_, _18792_);
  not (_19348_, _19338_);
  nor (_19359_, _19348_, _19316_);
  nor (_19370_, _19359_, _18792_);
  nor (_19381_, _19370_, _18749_);
  nor (_19392_, _19381_, _18716_);
  not (_19403_, _19392_);
  and (_19414_, _19403_, _14891_);
  and (_19425_, _19414_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_19436_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_19447_, _19436_, _19425_);
  and (_19457_, _19447_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_19468_, _19457_, _14880_);
  and (_19479_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19490_, _19479_, _19468_);
  and (_19501_, _19468_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19512_, _19501_, _19490_);
  and (_26945_, _19512_, _43998_);
  nor (_19533_, _14750_, _14783_);
  and (_19544_, _14750_, _14783_);
  or (_19555_, _19544_, _19533_);
  and (_02688_, _19555_, _43998_);
  and (_19575_, _18422_, _15670_);
  and (_02889_, _19575_, _43998_);
  nor (_19596_, _18432_, _18083_);
  nor (_19607_, _19596_, _18443_);
  and (_03093_, _19607_, _43998_);
  nor (_19628_, _19141_, _19119_);
  nor (_19639_, _19628_, _19152_);
  and (_03304_, _19639_, _43998_);
  nor (_19660_, _19174_, _19152_);
  nor (_19671_, _19660_, _19185_);
  and (_03505_, _19671_, _43998_);
  nor (_19692_, _19228_, _19207_);
  nor (_19702_, _19692_, _19239_);
  and (_03706_, _19702_, _43998_);
  and (_19723_, _19250_, _19021_);
  nor (_19734_, _19723_, _19261_);
  and (_03907_, _19734_, _43998_);
  and (_19755_, _19272_, _18945_);
  nor (_19766_, _19755_, _19283_);
  and (_04108_, _19766_, _43998_);
  and (_19787_, _19294_, _18869_);
  nor (_19798_, _19787_, _19305_);
  and (_04309_, _19798_, _43998_);
  and (_19818_, _19348_, _19316_);
  nor (_19829_, _19818_, _19359_);
  and (_04423_, _19829_, _43998_);
  and (_19850_, _19370_, _18749_);
  nor (_19861_, _19850_, _19381_);
  and (_04536_, _19861_, _43998_);
  nor (_19882_, _19403_, _14891_);
  nor (_19893_, _19882_, _19414_);
  and (_04637_, _19893_, _43998_);
  and (_19914_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_19925_, _19914_, _19414_);
  nor (_19936_, _19925_, _19425_);
  and (_04738_, _19936_, _43998_);
  nor (_19956_, _19436_, _19425_);
  nor (_19967_, _19956_, _19447_);
  and (_04839_, _19967_, _43998_);
  and (_19988_, _14869_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_19999_, _19988_, _19447_);
  nor (_20010_, _19999_, _19457_);
  and (_04940_, _20010_, _43998_);
  nor (_20031_, _19457_, _14880_);
  nor (_20042_, _20031_, _19468_);
  and (_05041_, _20042_, _43998_);
  and (_20062_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _14684_);
  nor (_20073_, _20062_, _14695_);
  not (_20084_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_20095_, _14717_, _20084_);
  and (_20106_, _20095_, _20073_);
  and (_20117_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_20128_, _20117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20139_, _20117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20150_, _20139_, _20128_);
  and (_01042_, _20150_, _43998_);
  and (_01072_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _43998_);
  not (_20181_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_20192_, _16460_, _20181_);
  and (_20202_, _16142_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20213_, _20202_, _20192_);
  nor (_20224_, _20213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20235_, _16295_, _20181_);
  and (_20246_, _16634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_20257_, _20246_, _20235_);
  and (_20268_, _20257_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20279_, _20268_, _20224_);
  nor (_20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20301_, _20290_, _16810_);
  nor (_20312_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_20322_, _20312_, _20301_);
  not (_20333_, _20322_);
  and (_20344_, _15473_, _20181_);
  and (_20355_, _15144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20366_, _20355_, _20344_);
  nor (_20377_, _20366_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20388_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20399_, _15308_, _20181_);
  and (_20410_, _15648_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20421_, _20410_, _20399_);
  nor (_20431_, _20421_, _20388_);
  nor (_20442_, _20431_, _20377_);
  nor (_20453_, _20442_, _20333_);
  and (_20464_, _20442_, _20333_);
  nor (_20475_, _20464_, _20453_);
  and (_20486_, _20290_, _15966_);
  nor (_20497_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_20508_, _20497_, _20486_);
  not (_20519_, _20508_);
  nor (_20530_, _16460_, _20181_);
  nor (_20540_, _20530_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20551_, _16142_, _20181_);
  and (_20562_, _16295_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20573_, _20562_, _20551_);
  nor (_20584_, _20573_, _20388_);
  nor (_20595_, _20584_, _20540_);
  nor (_20606_, _20595_, _20519_);
  and (_20617_, _20595_, _20519_);
  nor (_20628_, _20617_, _20606_);
  not (_20639_, _20628_);
  nor (_20650_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_20660_, _20290_, _17006_);
  nor (_20671_, _20660_, _20650_);
  not (_20682_, _20671_);
  nor (_20693_, _15473_, _20181_);
  nor (_20704_, _20693_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20715_, _15144_, _20181_);
  and (_20726_, _15308_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20737_, _20726_, _20715_);
  nor (_20748_, _20737_, _20388_);
  nor (_20759_, _20748_, _20704_);
  nor (_20769_, _20759_, _20682_);
  and (_20780_, _20759_, _20682_);
  and (_20791_, _20213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20802_, _20791_);
  and (_20813_, _20290_, _17180_);
  nor (_20824_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  nor (_20835_, _20824_, _20813_);
  and (_20846_, _20835_, _20802_);
  and (_20857_, _20366_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20868_, _20857_);
  and (_20878_, _20290_, _17539_);
  nor (_20889_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_20900_, _20889_, _20878_);
  and (_20911_, _20900_, _20868_);
  nor (_20922_, _20900_, _20868_);
  nor (_20933_, _20922_, _20911_);
  not (_20944_, _20933_);
  and (_20955_, _20530_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20966_, _20955_);
  and (_20977_, _20290_, _18040_);
  nor (_20987_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_20998_, _20987_, _20977_);
  and (_21009_, _20998_, _20966_);
  and (_21020_, _20693_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21031_, _21020_);
  nor (_21042_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_21053_, _20290_, _17865_);
  nor (_21064_, _21053_, _21042_);
  nor (_21075_, _21064_, _21031_);
  not (_21086_, _21075_);
  nor (_21097_, _20998_, _20966_);
  nor (_21107_, _21097_, _21009_);
  and (_21118_, _21107_, _21086_);
  nor (_21129_, _21118_, _21009_);
  nor (_21140_, _21129_, _20944_);
  nor (_21151_, _21140_, _20911_);
  nor (_21162_, _20835_, _20802_);
  nor (_21173_, _21162_, _20846_);
  not (_21184_, _21173_);
  nor (_21195_, _21184_, _21151_);
  nor (_21205_, _21195_, _20846_);
  nor (_21216_, _21205_, _20780_);
  nor (_21227_, _21216_, _20769_);
  nor (_21238_, _21227_, _20639_);
  nor (_21249_, _21238_, _20606_);
  not (_21260_, _21249_);
  and (_21271_, _21260_, _20475_);
  or (_21282_, _21271_, _20453_);
  and (_21293_, _16634_, _15648_);
  or (_21304_, _21293_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_21315_, _20421_);
  and (_21325_, _20257_, _21315_);
  nor (_21336_, _20737_, _20573_);
  and (_21347_, _21336_, _21325_);
  or (_21358_, _21347_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21369_, _21358_, _21304_);
  and (_21380_, _21369_, _21282_);
  and (_21391_, _21380_, _20279_);
  nor (_21402_, _21260_, _20475_);
  or (_21413_, _21402_, _21271_);
  and (_21424_, _21413_, _21391_);
  nor (_21434_, _21391_, _20322_);
  nor (_21445_, _21434_, _21424_);
  not (_21456_, _21445_);
  and (_21467_, _21445_, _20279_);
  not (_21478_, _20442_);
  nor (_21489_, _21391_, _20519_);
  and (_21500_, _21227_, _20639_);
  nor (_21511_, _21500_, _21238_);
  and (_21522_, _21511_, _21391_);
  or (_21533_, _21522_, _21489_);
  and (_21543_, _21533_, _21478_);
  nor (_21554_, _21533_, _21478_);
  nor (_21565_, _21554_, _21543_);
  not (_21576_, _21565_);
  not (_21587_, _20595_);
  nor (_21598_, _21391_, _20682_);
  nor (_21620_, _20780_, _20769_);
  nor (_21632_, _21620_, _21205_);
  and (_21644_, _21620_, _21205_);
  or (_21656_, _21644_, _21632_);
  and (_21667_, _21656_, _21391_);
  or (_21679_, _21667_, _21598_);
  and (_21680_, _21679_, _21587_);
  nor (_21691_, _21679_, _21587_);
  not (_21702_, _20759_);
  and (_21713_, _21184_, _21151_);
  or (_21724_, _21713_, _21195_);
  and (_21735_, _21724_, _21391_);
  nor (_21746_, _21391_, _20835_);
  nor (_21757_, _21746_, _21735_);
  and (_21768_, _21757_, _21702_);
  and (_21778_, _21129_, _20944_);
  nor (_21789_, _21778_, _21140_);
  not (_21800_, _21789_);
  and (_21811_, _21800_, _21391_);
  nor (_21822_, _21391_, _20900_);
  nor (_21833_, _21822_, _21811_);
  and (_21844_, _21833_, _20802_);
  nor (_21855_, _21833_, _20802_);
  nor (_21866_, _21855_, _21844_);
  not (_21877_, _21866_);
  nor (_21887_, _21107_, _21086_);
  nor (_21898_, _21887_, _21118_);
  not (_21909_, _21898_);
  and (_21920_, _21909_, _21391_);
  nor (_21931_, _21391_, _20998_);
  nor (_21942_, _21931_, _21920_);
  and (_21953_, _21942_, _20868_);
  and (_21964_, _21391_, _21020_);
  nor (_21975_, _21964_, _21064_);
  and (_21986_, _21964_, _21064_);
  nor (_21996_, _21986_, _21975_);
  and (_22007_, _21996_, _20966_);
  nor (_22018_, _21996_, _20966_);
  nor (_22029_, _22018_, _22007_);
  nor (_22040_, _20290_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_22051_, _20290_, _18411_);
  nor (_22062_, _22051_, _22040_);
  nor (_22073_, _22062_, _21031_);
  not (_22084_, _22073_);
  and (_22095_, _22084_, _22029_);
  nor (_22105_, _22095_, _22007_);
  nor (_22116_, _21942_, _20868_);
  nor (_22127_, _22116_, _21953_);
  not (_22138_, _22127_);
  nor (_22149_, _22138_, _22105_);
  nor (_22160_, _22149_, _21953_);
  nor (_22171_, _22160_, _21877_);
  nor (_22192_, _22171_, _21844_);
  nor (_22193_, _21757_, _21702_);
  nor (_22204_, _22193_, _21768_);
  not (_22214_, _22204_);
  nor (_22225_, _22214_, _22192_);
  nor (_22236_, _22225_, _21768_);
  nor (_22247_, _22236_, _21691_);
  nor (_22258_, _22247_, _21680_);
  nor (_22269_, _22258_, _21576_);
  or (_22280_, _22269_, _21543_);
  or (_22291_, _22280_, _21467_);
  and (_22302_, _22291_, _21369_);
  nor (_22313_, _22302_, _21456_);
  and (_22324_, _21467_, _21369_);
  and (_22334_, _22324_, _22280_);
  or (_22345_, _22334_, _22313_);
  and (_01082_, _22345_, _43998_);
  or (_22366_, _21445_, _20279_);
  and (_22377_, _22366_, _22302_);
  and (_03050_, _22377_, _43998_);
  and (_03061_, _21391_, _43998_);
  and (_03082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _43998_);
  and (_03104_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _43998_);
  and (_03125_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _43998_);
  or (_22448_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_22449_, _20117_, rst);
  and (_03136_, _22449_, _22448_);
  not (_22470_, _22062_);
  and (_22481_, _22377_, _21020_);
  nor (_22492_, _22481_, _22470_);
  and (_22503_, _22481_, _22470_);
  or (_22514_, _22503_, _22492_);
  and (_03147_, _22514_, _43998_);
  nor (_22535_, _22084_, _22029_);
  or (_22545_, _22535_, _22095_);
  nand (_22556_, _22545_, _22377_);
  or (_22567_, _22377_, _21996_);
  and (_22578_, _22567_, _22556_);
  and (_03158_, _22578_, _43998_);
  and (_22599_, _22138_, _22105_);
  or (_22610_, _22599_, _22149_);
  nand (_22621_, _22610_, _22377_);
  or (_22632_, _22377_, _21942_);
  and (_22643_, _22632_, _22621_);
  and (_03169_, _22643_, _43998_);
  and (_22663_, _22160_, _21877_);
  or (_22674_, _22663_, _22171_);
  nand (_22685_, _22674_, _22377_);
  or (_22696_, _22377_, _21833_);
  and (_22707_, _22696_, _22685_);
  and (_03180_, _22707_, _43998_);
  and (_22728_, _22214_, _22192_);
  or (_22739_, _22728_, _22225_);
  nand (_22750_, _22739_, _22377_);
  or (_22761_, _22377_, _21757_);
  and (_22772_, _22761_, _22750_);
  and (_03191_, _22772_, _43998_);
  or (_22793_, _21691_, _21680_);
  and (_22804_, _22793_, _22236_);
  nor (_22815_, _22793_, _22236_);
  or (_22826_, _22815_, _22804_);
  nand (_22837_, _22826_, _22377_);
  or (_22848_, _22377_, _21679_);
  and (_22859_, _22848_, _22837_);
  and (_03202_, _22859_, _43998_);
  and (_22880_, _22258_, _21576_);
  or (_22891_, _22880_, _22269_);
  nand (_22902_, _22891_, _22377_);
  or (_22913_, _22377_, _21533_);
  and (_22923_, _22913_, _22902_);
  and (_03213_, _22923_, _43998_);
  not (_22944_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22955_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _14684_);
  and (_22966_, _22955_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_22977_, _22966_, _22944_);
  not (_22988_, _22977_);
  not (_22999_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_23010_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23021_, _23010_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_23032_, _23021_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_23043_, _23032_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_23054_, _23043_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_23065_, _23054_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23076_, _23065_, _22999_);
  and (_23087_, _23065_, _22999_);
  nor (_23098_, _23087_, _23076_);
  nor (_23119_, _23098_, _22988_);
  not (_23120_, _23119_);
  not (_23131_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23152_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _14684_);
  and (_23153_, _23152_, _22944_);
  and (_23164_, _23153_, _23131_);
  and (_23185_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_23186_, _23185_);
  and (_23197_, _22966_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_23218_, _23197_);
  not (_23219_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_23230_, _22955_, _23219_);
  and (_23251_, _23230_, _22944_);
  and (_23252_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_23263_, _23230_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23284_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_23285_, _23284_, _23252_);
  and (_23296_, _23285_, _23218_);
  and (_23316_, _23296_, _23186_);
  and (_23317_, _23316_, _23120_);
  not (_23328_, _23065_);
  nor (_23339_, _23054_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23350_, _23339_, _22988_);
  and (_23361_, _23350_, _23328_);
  not (_23372_, _23361_);
  and (_23383_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_23394_, _23383_, _23197_);
  and (_23405_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23416_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_23427_, _23416_, _23405_);
  and (_23438_, _23427_, _23394_);
  and (_23449_, _23438_, _23372_);
  nor (_23460_, _23449_, _23317_);
  not (_23471_, _23032_);
  nor (_23482_, _23021_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_23493_, _23482_, _22988_);
  and (_23504_, _23493_, _23471_);
  not (_23515_, _23504_);
  and (_23526_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or (_23537_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23548_, _23537_, _14684_);
  nor (_23559_, _23548_, _22955_);
  and (_23570_, _23559_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_23581_, _23570_, _23526_);
  and (_23592_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_23603_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_23614_, _23603_, _23592_);
  and (_23625_, _23614_, _23581_);
  and (_23636_, _23625_, _23515_);
  not (_23647_, _23636_);
  nor (_23658_, _23032_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_23669_, _23658_);
  nor (_23679_, _23043_, _22988_);
  and (_23690_, _23679_, _23669_);
  not (_23701_, _23690_);
  and (_23712_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_23723_, _23712_, _23197_);
  and (_23734_, _23559_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_23745_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_23756_, _23745_, _23734_);
  and (_23767_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  not (_23778_, _23767_);
  and (_23789_, _23778_, _23756_);
  and (_23800_, _23789_, _23723_);
  and (_23811_, _23800_, _23701_);
  nor (_23822_, _23811_, _23647_);
  nor (_23833_, _23043_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_23844_, _23833_);
  nor (_23855_, _23054_, _22988_);
  and (_23866_, _23855_, _23844_);
  not (_23877_, _23866_);
  and (_23888_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_23899_, _23888_, _23197_);
  and (_23910_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_23921_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_23932_, _23921_, _23910_);
  and (_23943_, _23932_, _23899_);
  and (_23954_, _23943_, _23877_);
  not (_23965_, _23954_);
  not (_23976_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23987_, _22977_, _23976_);
  and (_23998_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_24009_, _23998_, _23987_);
  and (_24020_, _23559_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  not (_24031_, _24020_);
  and (_24041_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24052_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_24063_, _24052_, _24041_);
  and (_24074_, _24063_, _24031_);
  and (_24085_, _24074_, _24009_);
  nor (_24096_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24107_, _24096_, _23010_);
  and (_24118_, _24107_, _22977_);
  and (_24129_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  nor (_24140_, _24129_, _24118_);
  and (_24151_, _23559_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  not (_24162_, _24151_);
  and (_24173_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24184_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24195_, _24184_, _24173_);
  and (_24206_, _24195_, _24162_);
  and (_24217_, _24206_, _24140_);
  nor (_24228_, _23010_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24239_, _24228_, _23021_);
  and (_24250_, _24239_, _22977_);
  and (_24261_, _23164_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24272_, _24261_, _24250_);
  and (_24283_, _23263_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24294_, _23251_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_24316_, _23559_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24328_, _24316_, _24294_);
  nor (_24340_, _24328_, _24283_);
  and (_24352_, _24340_, _24272_);
  and (_24364_, _24352_, _24217_);
  and (_24376_, _24364_, _24085_);
  and (_24388_, _24376_, _23965_);
  and (_24389_, _24388_, _23822_);
  nand (_24399_, _24389_, _23460_);
  and (_24410_, _22345_, _20106_);
  not (_24421_, _24410_);
  and (_24432_, _19512_, _14750_);
  not (_24443_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_24454_, _14695_, _24443_);
  and (_24465_, _24454_, _14739_);
  not (_24476_, _24465_);
  nor (_24487_, _16810_, _16634_);
  and (_24498_, _16810_, _16634_);
  nor (_24509_, _24498_, _24487_);
  not (_24520_, _15648_);
  nor (_24531_, _15966_, _24520_);
  nor (_24542_, _15966_, _15648_);
  and (_24553_, _15966_, _15648_);
  nor (_24564_, _24553_, _24542_);
  not (_24575_, _16295_);
  nor (_24586_, _17006_, _24575_);
  nor (_24597_, _17006_, _16295_);
  and (_24608_, _17006_, _16295_);
  nor (_24619_, _24608_, _24597_);
  not (_24630_, _15308_);
  and (_24641_, _17180_, _24630_);
  nor (_24652_, _24641_, _24619_);
  nor (_24663_, _24652_, _24586_);
  nor (_24674_, _24663_, _24564_);
  nor (_24685_, _24674_, _24531_);
  and (_24696_, _24663_, _24564_);
  nor (_24707_, _24696_, _24674_);
  not (_24718_, _24707_);
  and (_24729_, _24641_, _24619_);
  nor (_24740_, _24729_, _24652_);
  not (_24752_, _24740_);
  nor (_24763_, _17180_, _15308_);
  and (_24773_, _17180_, _15308_);
  nor (_24784_, _24773_, _24763_);
  not (_24795_, _24784_);
  and (_24806_, _17539_, _16142_);
  nor (_24817_, _17539_, _16142_);
  nor (_24828_, _24817_, _24806_);
  nor (_24839_, _18040_, _15144_);
  and (_24850_, _18040_, _15144_);
  nor (_24861_, _24850_, _24839_);
  nor (_24872_, _17865_, _16460_);
  and (_24883_, _17865_, _16460_);
  nor (_24894_, _24883_, _24872_);
  not (_24905_, _15473_);
  and (_24916_, _18411_, _24905_);
  nor (_24927_, _24916_, _24894_);
  not (_24938_, _16460_);
  nor (_24949_, _17865_, _24938_);
  nor (_24960_, _24949_, _24927_);
  nor (_24971_, _24960_, _24861_);
  not (_24982_, _15144_);
  nor (_24993_, _18040_, _24982_);
  nor (_25004_, _24993_, _24971_);
  nor (_25015_, _25004_, _24828_);
  and (_25026_, _25004_, _24828_);
  nor (_25037_, _25026_, _25015_);
  not (_25048_, _25037_);
  nor (_25059_, _18411_, _15473_);
  and (_25070_, _18411_, _15473_);
  nor (_25081_, _25070_, _25059_);
  not (_25092_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_25103_, _14957_, _25092_);
  not (_25114_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25124_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25135_, _25124_, _16526_);
  nor (_25146_, _25135_, _25114_);
  nor (_25157_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25168_, _25157_, _15199_);
  not (_25179_, _25168_);
  not (_25190_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25201_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25190_);
  and (_25212_, _25201_, _16186_);
  not (_25223_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25244_, _25223_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25245_, _25244_, _15539_);
  nor (_25256_, _25245_, _25212_);
  and (_25267_, _25256_, _25179_);
  and (_25288_, _25267_, _25146_);
  and (_25289_, _25124_, _16032_);
  nor (_25300_, _25289_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25321_, _25244_, _15001_);
  not (_25322_, _25321_);
  and (_25333_, _25201_, _16350_);
  and (_25344_, _25157_, _15363_);
  nor (_25355_, _25344_, _25333_);
  and (_25376_, _25355_, _25322_);
  and (_25377_, _25376_, _25300_);
  nor (_25388_, _25377_, _25288_);
  nor (_25399_, _25388_, _14957_);
  nor (_25410_, _25399_, _25103_);
  and (_25421_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25432_, _25421_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_25443_, _25432_);
  and (_25454_, _25443_, _25410_);
  and (_25465_, _25443_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_25476_, _25465_, _25454_);
  nor (_25486_, _25476_, _25081_);
  and (_25507_, _24960_, _24861_);
  nor (_25508_, _25507_, _24971_);
  and (_25519_, _24916_, _24894_);
  nor (_25530_, _25519_, _24927_);
  nor (_25541_, _25530_, _25508_);
  and (_25552_, _25541_, _25486_);
  and (_25563_, _25552_, _25048_);
  not (_25574_, _16142_);
  or (_25585_, _17539_, _25574_);
  and (_25596_, _17539_, _25574_);
  or (_25607_, _25004_, _25596_);
  and (_25618_, _25607_, _25585_);
  or (_25629_, _25618_, _25563_);
  and (_25640_, _25629_, _24795_);
  and (_25651_, _25640_, _24752_);
  and (_25662_, _25651_, _24718_);
  nor (_25683_, _25662_, _24685_);
  nor (_25684_, _25683_, _24509_);
  and (_25695_, _25683_, _24509_);
  nor (_25706_, _25695_, _25684_);
  nor (_25717_, _25706_, _24476_);
  not (_25728_, _25717_);
  not (_25739_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_25750_, _20062_, _25739_);
  and (_25761_, _25750_, _14739_);
  not (_25772_, _24509_);
  not (_25783_, _24564_);
  and (_25794_, _24763_, _24619_);
  nor (_25805_, _25794_, _24597_);
  nor (_25816_, _25805_, _25783_);
  not (_25826_, _24861_);
  and (_25837_, _25059_, _24894_);
  nor (_25848_, _25837_, _24872_);
  nor (_25859_, _25848_, _25826_);
  nor (_25880_, _25859_, _24839_);
  nor (_25881_, _25880_, _24828_);
  and (_25892_, _25880_, _24828_);
  nor (_25903_, _25892_, _25881_);
  not (_25914_, _25081_);
  nor (_25925_, _25476_, _25914_);
  and (_25936_, _25925_, _24894_);
  and (_25947_, _25848_, _25826_);
  nor (_25958_, _25947_, _25859_);
  and (_25969_, _25958_, _25936_);
  not (_25980_, _25969_);
  nor (_25991_, _25980_, _25903_);
  nor (_26002_, _25880_, _24806_);
  or (_26013_, _26002_, _24817_);
  or (_26024_, _26013_, _25991_);
  and (_26035_, _26024_, _24784_);
  and (_26046_, _26035_, _24619_);
  and (_26057_, _25805_, _25783_);
  nor (_26068_, _26057_, _25816_);
  and (_26079_, _26068_, _26046_);
  or (_26090_, _26079_, _25816_);
  nor (_26101_, _26090_, _24542_);
  nor (_26112_, _26101_, _25772_);
  and (_26123_, _26101_, _25772_);
  nor (_26134_, _26123_, _26112_);
  and (_26145_, _26134_, _25761_);
  nor (_26156_, _18411_, _17865_);
  and (_26166_, _26156_, _18051_);
  and (_26177_, _26166_, _17550_);
  and (_26188_, _26177_, _17191_);
  and (_26199_, _26188_, _17016_);
  and (_26210_, _26199_, _15977_);
  and (_26231_, _26210_, _25476_);
  not (_26232_, _25476_);
  and (_26243_, _15966_, _17006_);
  and (_26254_, _18411_, _17865_);
  and (_26265_, _26254_, _18040_);
  and (_26276_, _26265_, _17539_);
  and (_26287_, _26276_, _17180_);
  and (_26298_, _26287_, _26243_);
  and (_26309_, _26298_, _26232_);
  nor (_26320_, _26309_, _26231_);
  and (_26341_, _26320_, _16810_);
  not (_26342_, _26341_);
  and (_26353_, _14728_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26364_, _26353_, _24454_);
  not (_26375_, _26364_);
  nor (_26386_, _26320_, _16810_);
  nor (_26397_, _26386_, _26375_);
  and (_26408_, _26397_, _26342_);
  not (_26419_, _16634_);
  nor (_26430_, _25476_, _26419_);
  not (_26441_, _26430_);
  and (_26452_, _25476_, _16810_);
  and (_26463_, _26353_, _14706_);
  not (_26474_, _26463_);
  nor (_26484_, _26474_, _26452_);
  and (_26495_, _26484_, _26441_);
  not (_26506_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26517_, _14728_, _26506_);
  and (_26528_, _26517_, _25750_);
  not (_26539_, _26528_);
  nor (_26550_, _26539_, _24498_);
  and (_26561_, _26517_, _20073_);
  and (_26572_, _26561_, _24509_);
  nor (_26583_, _26572_, _26550_);
  not (_26594_, _26583_);
  nor (_26605_, _26594_, _26495_);
  not (_26616_, _26605_);
  nor (_26627_, _26616_, _26408_);
  and (_26638_, _25750_, _20095_);
  and (_26649_, _18040_, _17865_);
  nor (_26660_, _26649_, _17539_);
  and (_26671_, _26660_, _26638_);
  and (_26682_, _26671_, _17191_);
  nor (_26693_, _26682_, _17016_);
  and (_26704_, _26693_, _15966_);
  nor (_26715_, _26243_, _16810_);
  nor (_26726_, _26715_, _26671_);
  and (_26737_, _26726_, _25476_);
  nor (_26748_, _26737_, _26704_);
  and (_26759_, _26748_, _16821_);
  not (_26770_, _26638_);
  nor (_26791_, _26748_, _16821_);
  or (_26792_, _26791_, _26770_);
  nor (_26802_, _26792_, _26759_);
  and (_26813_, _26353_, _25750_);
  not (_26824_, _26813_);
  nor (_26835_, _26824_, _25476_);
  not (_26846_, _26835_);
  and (_26857_, _20095_, _14706_);
  and (_26868_, _26857_, _24487_);
  and (_26879_, _24454_, _20095_);
  and (_26890_, _26879_, _16810_);
  nor (_26901_, _26890_, _26868_);
  and (_26912_, _20073_, _14739_);
  not (_26923_, _26912_);
  nor (_26934_, _26923_, _16810_);
  not (_26946_, _26934_);
  and (_26957_, _26353_, _20073_);
  and (_26968_, _26957_, _18422_);
  and (_26979_, _26517_, _14695_);
  not (_26990_, _26979_);
  nor (_27001_, _26990_, _15966_);
  nor (_27012_, _27001_, _26968_);
  and (_27023_, _27012_, _26946_);
  and (_27034_, _27023_, _26901_);
  nand (_27045_, _27034_, _26846_);
  nor (_27056_, _27045_, _26802_);
  and (_27067_, _27056_, _26627_);
  not (_27088_, _27067_);
  nor (_27089_, _27088_, _26145_);
  and (_27100_, _27089_, _25728_);
  not (_27110_, _27100_);
  nor (_27121_, _27110_, _24432_);
  and (_27132_, _27121_, _24421_);
  not (_27143_, _27132_);
  or (_27154_, _27143_, _24399_);
  not (_27165_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_27176_, \oc8051_top_1.oc8051_decoder1.wr , _14684_);
  not (_27197_, _27176_);
  nor (_27198_, _27197_, _23153_);
  and (_27209_, _27198_, _27165_);
  not (_27220_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_27231_, _24399_, _27220_);
  and (_27242_, _27231_, _27209_);
  and (_27253_, _27242_, _27154_);
  nor (_27264_, _27198_, _27220_);
  not (_27275_, _25761_);
  nor (_27286_, _26112_, _24487_);
  nor (_27297_, _27286_, _27275_);
  not (_27308_, _27297_);
  and (_27319_, _16810_, _26419_);
  nor (_27330_, _27319_, _25684_);
  nor (_27341_, _27330_, _24476_);
  and (_27352_, _25476_, _15966_);
  and (_27363_, _27352_, _26693_);
  nor (_27374_, _27363_, _26452_);
  nor (_27385_, _25476_, _16810_);
  not (_27396_, _27385_);
  nor (_27416_, _27396_, _26704_);
  nor (_27417_, _27416_, _26770_);
  and (_27428_, _27417_, _27374_);
  not (_27439_, _27428_);
  and (_27450_, _26517_, _14706_);
  not (_27461_, _27450_);
  nor (_27472_, _27461_, _16810_);
  not (_27483_, _27472_);
  nor (_27494_, _26824_, _18411_);
  nor (_27505_, _27494_, _26671_);
  and (_27516_, _27505_, _27483_);
  nor (_27527_, _26923_, _25476_);
  not (_27538_, _27527_);
  and (_27549_, _27538_, _27516_);
  nor (_27560_, _25465_, _25410_);
  not (_27571_, _26561_);
  nor (_27582_, _27571_, _25454_);
  nor (_27593_, _27582_, _26528_);
  nor (_27604_, _27593_, _27560_);
  not (_27615_, _27604_);
  and (_27626_, _25432_, _25410_);
  and (_27637_, _26517_, _24454_);
  and (_27648_, _26857_, _25410_);
  nor (_27659_, _27648_, _27637_);
  nor (_27680_, _27659_, _27626_);
  and (_27681_, _26879_, _25476_);
  nand (_27692_, _26957_, _25465_);
  nor (_27703_, _27692_, _25410_);
  or (_27714_, _27703_, _27681_);
  nor (_27724_, _27714_, _27680_);
  and (_27735_, _27724_, _27615_);
  and (_27746_, _27735_, _27549_);
  and (_27757_, _27746_, _27439_);
  not (_27768_, _27757_);
  nor (_27779_, _27768_, _27341_);
  and (_27790_, _27779_, _27308_);
  nor (_27801_, _23954_, _23449_);
  not (_27812_, _23317_);
  and (_27823_, _23822_, _27812_);
  and (_27834_, _27823_, _27801_);
  not (_27845_, _24085_);
  nor (_27856_, _24352_, _24217_);
  and (_27867_, _27856_, _27845_);
  and (_27878_, _27867_, _27834_);
  nand (_27889_, _27878_, _27790_);
  and (_27900_, _27198_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_27911_, _27878_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_27922_, _27911_, _27900_);
  and (_27933_, _27922_, _27889_);
  or (_27944_, _27933_, _27264_);
  or (_27965_, _27944_, _27253_);
  and (_06731_, _27965_, _43998_);
  and (_27976_, _22514_, _20106_);
  not (_27987_, _27976_);
  and (_27998_, _19829_, _14750_);
  and (_28009_, _25476_, _25914_);
  nor (_28020_, _28009_, _25925_);
  not (_28031_, _28020_);
  nor (_28042_, _25761_, _24465_);
  nor (_28053_, _28042_, _28031_);
  nor (_28064_, _27461_, _25476_);
  not (_28075_, _28064_);
  nor (_28086_, _27571_, _25059_);
  nor (_28097_, _28086_, _26528_);
  or (_28108_, _28097_, _25070_);
  and (_28119_, _26353_, _25739_);
  not (_28130_, _28119_);
  nor (_28141_, _28130_, _17865_);
  and (_28152_, _27637_, _16821_);
  nor (_28163_, _28152_, _28141_);
  and (_28174_, _26857_, _25059_);
  and (_28185_, _26879_, _18411_);
  nor (_28196_, _28185_, _28174_);
  nor (_28207_, _26474_, _15473_);
  and (_28218_, _26364_, _18411_);
  nor (_28229_, _28218_, _28207_);
  nor (_28240_, _26912_, _26638_);
  nor (_28251_, _28240_, _18411_);
  not (_28262_, _28251_);
  and (_28273_, _28262_, _28229_);
  and (_28284_, _28273_, _28196_);
  and (_28295_, _28284_, _28163_);
  and (_28306_, _28295_, _28108_);
  and (_28317_, _28306_, _28075_);
  not (_28328_, _28317_);
  nor (_28339_, _28328_, _28053_);
  not (_28350_, _28339_);
  nor (_28361_, _28350_, _27998_);
  and (_28372_, _28361_, _27987_);
  not (_28383_, _28372_);
  or (_28404_, _28383_, _24399_);
  not (_28405_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_28416_, _24399_, _28405_);
  and (_28427_, _28416_, _27209_);
  and (_28438_, _28427_, _28404_);
  nor (_28449_, _27198_, _28405_);
  not (_28460_, _27790_);
  or (_28471_, _28460_, _24399_);
  and (_28482_, _28416_, _27900_);
  and (_28493_, _28482_, _28471_);
  or (_28504_, _28493_, _28449_);
  or (_28515_, _28504_, _28438_);
  and (_08963_, _28515_, _43998_);
  and (_28536_, _19861_, _14750_);
  not (_28547_, _28536_);
  and (_28558_, _22578_, _20106_);
  nor (_28569_, _26474_, _16460_);
  nor (_28590_, _26254_, _26156_);
  not (_28591_, _28590_);
  nor (_28602_, _28591_, _25476_);
  and (_28613_, _28591_, _25476_);
  nor (_28624_, _28613_, _28602_);
  and (_28635_, _28624_, _26364_);
  nor (_28646_, _28635_, _28569_);
  nor (_28657_, _26660_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_28668_, _28657_, _17876_);
  nor (_28679_, _28657_, _17876_);
  nor (_28690_, _28679_, _28668_);
  nor (_28701_, _28690_, _26770_);
  not (_28712_, _28701_);
  and (_28723_, _26561_, _24894_);
  nor (_28734_, _26539_, _24883_);
  not (_28745_, _28734_);
  and (_28756_, _26857_, _24872_);
  and (_28767_, _26879_, _17865_);
  nor (_28778_, _28767_, _28756_);
  nand (_28789_, _28778_, _28745_);
  nor (_28800_, _28789_, _28723_);
  nor (_28811_, _28130_, _18040_);
  not (_28832_, _28811_);
  nor (_28844_, _26923_, _17865_);
  nor (_28855_, _26990_, _18411_);
  nor (_28866_, _28855_, _28844_);
  and (_28877_, _28866_, _28832_);
  and (_28888_, _28877_, _28800_);
  and (_28899_, _28888_, _28712_);
  and (_28910_, _28899_, _28646_);
  nor (_28921_, _25059_, _24894_);
  or (_28932_, _28921_, _25837_);
  and (_28943_, _28932_, _25925_);
  nor (_28954_, _28932_, _25925_);
  or (_28965_, _28954_, _28943_);
  and (_28976_, _28965_, _25761_);
  not (_28987_, _25530_);
  and (_28998_, _28987_, _25486_);
  nor (_29009_, _28987_, _25486_);
  nor (_29020_, _29009_, _28998_);
  nor (_29031_, _29020_, _24476_);
  nor (_29042_, _29031_, _28976_);
  and (_29053_, _29042_, _28910_);
  not (_29064_, _29053_);
  nor (_29075_, _29064_, _28558_);
  and (_29086_, _29075_, _28547_);
  not (_29097_, _29086_);
  or (_29108_, _29097_, _24399_);
  not (_29119_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_29140_, _24399_, _29119_);
  and (_29141_, _29140_, _27209_);
  and (_29152_, _29141_, _29108_);
  nor (_29163_, _27198_, _29119_);
  and (_29174_, _24364_, _27845_);
  and (_29185_, _29174_, _27834_);
  or (_29196_, _29185_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29207_, _29196_, _27900_);
  nand (_29218_, _29185_, _27790_);
  and (_29228_, _29218_, _29207_);
  or (_29239_, _29228_, _29163_);
  or (_29250_, _29239_, _29152_);
  and (_08974_, _29250_, _43998_);
  and (_29271_, _19893_, _14750_);
  not (_29282_, _29271_);
  and (_29293_, _22643_, _20106_);
  nor (_29304_, _26474_, _15144_);
  and (_29315_, _26254_, _26232_);
  and (_29326_, _26156_, _25476_);
  nor (_29337_, _29326_, _29315_);
  nor (_29347_, _29337_, _18040_);
  and (_29358_, _29337_, _18040_);
  or (_29369_, _29358_, _26375_);
  nor (_29380_, _29369_, _29347_);
  nor (_29391_, _29380_, _29304_);
  not (_29402_, _28998_);
  and (_29413_, _29402_, _25508_);
  nor (_29424_, _29413_, _25552_);
  nor (_29435_, _29424_, _24476_);
  and (_29446_, _26561_, _24861_);
  nor (_29457_, _26539_, _24850_);
  not (_29468_, _29457_);
  and (_29479_, _26857_, _24839_);
  and (_29490_, _26879_, _18040_);
  nor (_29501_, _29490_, _29479_);
  nand (_29512_, _29501_, _29468_);
  nor (_29523_, _29512_, _29446_);
  nor (_29534_, _26990_, _17865_);
  not (_29545_, _29534_);
  nor (_29556_, _26923_, _18040_);
  nor (_29567_, _28130_, _17539_);
  nor (_29578_, _29567_, _29556_);
  and (_29589_, _29578_, _29545_);
  and (_29599_, _29589_, _29523_);
  not (_29610_, _29599_);
  nor (_29621_, _29610_, _29435_);
  nor (_29632_, _25958_, _25936_);
  nor (_29643_, _29632_, _27275_);
  and (_29654_, _29643_, _25980_);
  nor (_29665_, _28679_, _18040_);
  and (_29686_, _26649_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_29687_, _29686_, _29665_);
  nor (_29698_, _29687_, _26770_);
  nor (_29708_, _29698_, _29654_);
  and (_29719_, _29708_, _29621_);
  and (_29730_, _29719_, _29391_);
  not (_29741_, _29730_);
  nor (_29752_, _29741_, _29293_);
  and (_29763_, _29752_, _29282_);
  not (_29774_, _29763_);
  or (_29785_, _29774_, _24399_);
  not (_29796_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_29807_, _24399_, _29796_);
  and (_29818_, _29807_, _27209_);
  and (_29828_, _29818_, _29785_);
  nor (_29839_, _27198_, _29796_);
  nand (_29850_, _27834_, _24352_);
  nor (_29861_, _24217_, _24085_);
  or (_29872_, _29861_, _29850_);
  and (_29883_, _29872_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_29894_, _24217_);
  and (_29905_, _24352_, _29894_);
  and (_29916_, _29905_, _24085_);
  and (_29927_, _29916_, _28460_);
  and (_29947_, _24364_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_29948_, _29947_, _29927_);
  and (_29959_, _29948_, _27834_);
  or (_29970_, _29959_, _29883_);
  and (_29981_, _29970_, _27900_);
  or (_29992_, _29981_, _29839_);
  or (_30003_, _29992_, _29828_);
  and (_08985_, _30003_, _43998_);
  and (_30024_, _22707_, _20106_);
  not (_30035_, _30024_);
  and (_30046_, _19936_, _14750_);
  and (_30057_, _25980_, _25903_);
  nor (_30068_, _30057_, _25991_);
  and (_30079_, _30068_, _25761_);
  not (_30090_, _30079_);
  nor (_30101_, _25552_, _25048_);
  nor (_30112_, _30101_, _25563_);
  nor (_30122_, _30112_, _24476_);
  not (_30133_, _30122_);
  nor (_30144_, _26474_, _16142_);
  nor (_30155_, _26265_, _25476_);
  nor (_30166_, _26166_, _26232_);
  nor (_30177_, _30166_, _30155_);
  and (_30188_, _30177_, _17550_);
  not (_30199_, _30188_);
  nor (_30209_, _30177_, _17550_);
  nor (_30220_, _30209_, _26375_);
  and (_30231_, _30220_, _30199_);
  nor (_30252_, _30231_, _30144_);
  nor (_30253_, _26539_, _24806_);
  and (_30264_, _26561_, _24828_);
  nor (_30275_, _30264_, _30253_);
  not (_30286_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30296_, _26649_, _30286_);
  nor (_30307_, _30296_, _17550_);
  or (_30318_, _30307_, _26770_);
  or (_30329_, _30318_, _26660_);
  and (_30340_, _26857_, _24817_);
  and (_30351_, _26879_, _17539_);
  nor (_30362_, _30351_, _30340_);
  nor (_30373_, _28130_, _17180_);
  nor (_30383_, _26923_, _17539_);
  nor (_30394_, _26990_, _18040_);
  or (_30405_, _30394_, _30383_);
  nor (_30416_, _30405_, _30373_);
  and (_30427_, _30416_, _30362_);
  and (_30438_, _30427_, _30329_);
  and (_30449_, _30438_, _30275_);
  and (_30460_, _30449_, _30252_);
  and (_30470_, _30460_, _30133_);
  and (_30481_, _30470_, _30090_);
  not (_30492_, _30481_);
  nor (_30503_, _30492_, _30046_);
  and (_30514_, _30503_, _30035_);
  not (_30525_, _30514_);
  or (_30536_, _30525_, _24399_);
  not (_30547_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_30557_, _24399_, _30547_);
  and (_30578_, _30557_, _27209_);
  and (_30579_, _30578_, _30536_);
  nor (_30590_, _27198_, _30547_);
  and (_30601_, _29850_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_30612_, _29861_, _24352_);
  not (_30623_, _30612_);
  nor (_30634_, _30623_, _27790_);
  not (_30644_, _24352_);
  or (_30655_, _29861_, _30644_);
  nor (_30666_, _30655_, _30547_);
  or (_30677_, _30666_, _30634_);
  and (_30688_, _30677_, _27834_);
  or (_30699_, _30688_, _30601_);
  and (_30710_, _30699_, _27900_);
  or (_30721_, _30710_, _30590_);
  or (_30732_, _30721_, _30579_);
  and (_08996_, _30732_, _43998_);
  and (_30752_, _22772_, _20106_);
  not (_30763_, _30752_);
  and (_30774_, _19967_, _14750_);
  nor (_30785_, _25629_, _24784_);
  and (_30796_, _25629_, _24784_);
  nor (_30807_, _30796_, _30785_);
  and (_30817_, _30807_, _24465_);
  not (_30828_, _30817_);
  not (_30839_, _26035_);
  nor (_30850_, _26024_, _24784_);
  nor (_30861_, _30850_, _27275_);
  and (_30872_, _30861_, _30839_);
  not (_30883_, _30872_);
  and (_30894_, _26857_, _24763_);
  and (_30904_, _26879_, _17180_);
  nor (_30915_, _30904_, _30894_);
  nor (_30926_, _28130_, _17006_);
  not (_30937_, _30926_);
  and (_30948_, _30937_, _30915_);
  and (_30959_, _25476_, _17191_);
  nor (_30970_, _25476_, _15308_);
  or (_30981_, _30970_, _30959_);
  and (_30991_, _30981_, _26463_);
  and (_31002_, _26177_, _25476_);
  and (_31013_, _26276_, _26232_);
  nor (_31024_, _31013_, _31002_);
  nor (_31035_, _31024_, _17180_);
  and (_31056_, _31024_, _17180_);
  or (_31057_, _31056_, _26375_);
  nor (_31068_, _31057_, _31035_);
  nor (_31078_, _31068_, _30991_);
  nor (_31089_, _26671_, _17191_);
  not (_31100_, _31089_);
  nor (_31111_, _26682_, _26770_);
  and (_31122_, _31111_, _31100_);
  nor (_31133_, _26539_, _24773_);
  and (_31144_, _26561_, _24784_);
  nor (_31155_, _31144_, _31133_);
  nor (_31166_, _26923_, _17180_);
  nor (_31176_, _26990_, _17539_);
  nor (_31187_, _31176_, _31166_);
  nand (_31198_, _31187_, _31155_);
  nor (_31209_, _31198_, _31122_);
  and (_31220_, _31209_, _31078_);
  and (_31231_, _31220_, _30948_);
  and (_31242_, _31231_, _30883_);
  and (_31253_, _31242_, _30828_);
  not (_31263_, _31253_);
  nor (_31284_, _31263_, _30774_);
  and (_31285_, _31284_, _30763_);
  not (_31296_, _31285_);
  or (_31307_, _31296_, _24399_);
  not (_31318_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_31329_, _24399_, _31318_);
  and (_31340_, _31329_, _27209_);
  and (_31350_, _31340_, _31307_);
  nor (_31361_, _27198_, _31318_);
  not (_31372_, _27834_);
  and (_31383_, _24217_, _24085_);
  and (_31394_, _31383_, _30644_);
  nor (_31405_, _31383_, _30644_);
  nor (_31416_, _31405_, _31394_);
  or (_31427_, _31416_, _31372_);
  and (_31438_, _31427_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_31449_, _31394_);
  nor (_31459_, _31449_, _27790_);
  and (_31470_, _31405_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_31481_, _31470_, _31459_);
  and (_31492_, _31481_, _27834_);
  or (_31503_, _31492_, _31438_);
  and (_31514_, _31503_, _27900_);
  or (_31525_, _31514_, _31361_);
  or (_31536_, _31525_, _31350_);
  and (_09007_, _31536_, _43998_);
  and (_31557_, _20010_, _14750_);
  not (_31567_, _31557_);
  and (_31578_, _22859_, _20106_);
  nor (_31589_, _25476_, _16295_);
  and (_31600_, _25476_, _17016_);
  nor (_31611_, _31600_, _31589_);
  nor (_31622_, _31611_, _26474_);
  nor (_31633_, _26188_, _26232_);
  nor (_31644_, _26287_, _25476_);
  nor (_31655_, _31644_, _31633_);
  and (_31666_, _31655_, _17016_);
  nor (_31677_, _31655_, _17016_);
  or (_31687_, _31677_, _26375_);
  nor (_31698_, _31687_, _31666_);
  nor (_31709_, _31698_, _31622_);
  not (_31720_, _26737_);
  and (_31731_, _31720_, _26693_);
  nor (_31742_, _26737_, _26682_);
  nor (_31753_, _31742_, _17006_);
  nor (_31764_, _31753_, _31731_);
  nor (_31775_, _31764_, _26770_);
  nor (_31786_, _28130_, _15966_);
  and (_31797_, _26857_, _24597_);
  and (_31807_, _26879_, _17006_);
  nor (_31818_, _31807_, _31797_);
  nor (_31829_, _26539_, _24608_);
  and (_31840_, _26561_, _24619_);
  nor (_31861_, _31840_, _31829_);
  nor (_31862_, _26990_, _17180_);
  nor (_31873_, _26923_, _17006_);
  nor (_31884_, _31873_, _31862_);
  and (_31895_, _31884_, _31861_);
  nand (_31906_, _31895_, _31818_);
  nor (_31916_, _31906_, _31786_);
  not (_31927_, _31916_);
  nor (_31938_, _31927_, _31775_);
  nor (_31949_, _25640_, _24752_);
  nor (_31960_, _31949_, _25651_);
  nor (_31971_, _31960_, _24476_);
  nor (_31982_, _24763_, _24619_);
  or (_31993_, _31982_, _25794_);
  and (_32004_, _31993_, _30839_);
  not (_32015_, _32004_);
  nor (_32026_, _27275_, _26046_);
  and (_32036_, _32026_, _32015_);
  nor (_32047_, _32036_, _31971_);
  and (_32058_, _32047_, _31938_);
  and (_32069_, _32058_, _31709_);
  not (_32080_, _32069_);
  nor (_32091_, _32080_, _31578_);
  and (_32102_, _32091_, _31567_);
  not (_32113_, _32102_);
  or (_32124_, _32113_, _24399_);
  not (_32135_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_32145_, _24399_, _32135_);
  and (_32156_, _32145_, _27209_);
  and (_32167_, _32156_, _32124_);
  nor (_32178_, _27198_, _32135_);
  and (_32189_, _30644_, _24217_);
  nor (_32200_, _32189_, _29905_);
  or (_32211_, _32200_, _31372_);
  and (_32222_, _32211_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_32232_, _24217_, _27845_);
  and (_32243_, _32232_, _30644_);
  not (_32254_, _32243_);
  nor (_32265_, _32254_, _27790_);
  or (_32276_, _31394_, _29905_);
  and (_32287_, _32276_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_32298_, _32287_, _32265_);
  and (_32309_, _32298_, _27834_);
  or (_32320_, _32309_, _32222_);
  and (_32331_, _32320_, _27900_);
  or (_32342_, _32331_, _32178_);
  or (_32352_, _32342_, _32167_);
  and (_09018_, _32352_, _43998_);
  and (_32373_, _22923_, _20106_);
  not (_32384_, _32373_);
  and (_32395_, _20042_, _14750_);
  nor (_32406_, _25651_, _24718_);
  nor (_32417_, _32406_, _25662_);
  nor (_32428_, _32417_, _24476_);
  not (_32439_, _32428_);
  nor (_32450_, _26068_, _26046_);
  nor (_32461_, _32450_, _26079_);
  and (_32472_, _32461_, _25761_);
  nor (_32492_, _25476_, _24520_);
  or (_32493_, _32492_, _26474_);
  nor (_32504_, _32493_, _27352_);
  nor (_32515_, _25476_, _17016_);
  nand (_32526_, _32515_, _26287_);
  nand (_32537_, _26199_, _25476_);
  and (_32548_, _32537_, _32526_);
  nor (_32559_, _32548_, _15966_);
  not (_32570_, _32559_);
  and (_32581_, _32548_, _15966_);
  nor (_32592_, _32581_, _26375_);
  and (_32602_, _32592_, _32570_);
  nor (_32613_, _32602_, _32504_);
  nor (_32624_, _31731_, _15966_);
  and (_32635_, _31731_, _15966_);
  nor (_32646_, _32635_, _32624_);
  nor (_32657_, _32646_, _26770_);
  and (_32668_, _26561_, _24564_);
  nor (_32679_, _26539_, _24553_);
  not (_32690_, _32679_);
  and (_32701_, _26857_, _24542_);
  and (_32712_, _26879_, _15966_);
  nor (_32723_, _32712_, _32701_);
  nand (_32734_, _32723_, _32690_);
  nor (_32744_, _32734_, _32668_);
  nor (_32755_, _26990_, _17006_);
  not (_32766_, _32755_);
  nor (_32777_, _26923_, _15966_);
  nor (_32798_, _28130_, _16810_);
  nor (_32799_, _32798_, _32777_);
  and (_32810_, _32799_, _32766_);
  and (_32821_, _32810_, _32744_);
  not (_32832_, _32821_);
  nor (_32843_, _32832_, _32657_);
  and (_32854_, _32843_, _32613_);
  not (_32865_, _32854_);
  nor (_32875_, _32865_, _32472_);
  and (_32886_, _32875_, _32439_);
  not (_32897_, _32886_);
  nor (_32908_, _32897_, _32395_);
  and (_32919_, _32908_, _32384_);
  not (_32930_, _32919_);
  or (_32941_, _32930_, _24399_);
  not (_32952_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_32963_, _24399_, _32952_);
  and (_32974_, _32963_, _27209_);
  and (_32985_, _32974_, _32941_);
  nor (_32996_, _27198_, _32952_);
  not (_33006_, _27867_);
  nand (_33017_, _33006_, _27834_);
  and (_33028_, _33017_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_33039_, _27856_, _24085_);
  and (_33050_, _33039_, _28460_);
  nor (_33061_, _27856_, _32952_);
  or (_33072_, _33061_, _33050_);
  and (_33083_, _33072_, _27834_);
  or (_33094_, _33083_, _33028_);
  and (_33105_, _33094_, _27900_);
  or (_33115_, _33105_, _32996_);
  or (_33126_, _33115_, _32985_);
  and (_09029_, _33126_, _43998_);
  and (_33147_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_33158_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_33169_, _33158_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33180_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_33191_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_33202_, _33191_, _33180_);
  and (_33213_, _33158_, _14684_);
  and (_33224_, _33213_, _33202_);
  not (_33234_, _33224_);
  and (_33245_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33256_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33267_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_33278_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_33289_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_33300_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_33311_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33322_, _33311_, _33300_);
  and (_33333_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_33343_, _33311_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_33354_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_33365_, _33354_, _33333_);
  and (_33376_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33387_, _33376_, _33300_);
  and (_33398_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not (_33409_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33420_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _33409_);
  and (_33431_, _33420_, _33300_);
  and (_33442_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_33453_, _33442_, _33398_);
  nor (_33463_, _33311_, _33300_);
  and (_33474_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not (_33485_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_33496_, _33485_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33517_, _33496_, _33300_);
  and (_33518_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_33529_, _33518_, _33474_);
  and (_33540_, _33529_, _33453_);
  and (_33551_, _33540_, _33365_);
  nor (_33562_, _33551_, _33289_);
  and (_33573_, _33562_, _33278_);
  or (_33583_, _33573_, _33267_);
  and (_33594_, _33583_, _33256_);
  nor (_33605_, _33594_, _33245_);
  nor (_33616_, _33605_, _33234_);
  and (_33627_, _33202_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_33638_, _33627_, _33234_);
  nor (_33649_, _33638_, _33616_);
  and (_33660_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33671_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_33682_, _33289_);
  and (_33692_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_33703_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_33714_, _33703_, _33692_);
  and (_33725_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_33736_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_33747_, _33736_, _33725_);
  and (_33758_, _33747_, _33714_);
  and (_33769_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_33780_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_33791_, _33780_, _33769_);
  and (_33802_, _33791_, _33758_);
  and (_33812_, _33802_, _33682_);
  nor (_33823_, _33812_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_33834_, _33823_, _33671_);
  nor (_33845_, _33834_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_33856_, _33845_, _33660_);
  nor (_33867_, _33856_, _33234_);
  and (_33878_, _33202_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_33889_, _33878_, _33234_);
  nor (_33899_, _33889_, _33867_);
  and (_33910_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33921_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_33932_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_33943_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_33954_, _33943_, _33932_);
  and (_33965_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_33976_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_33986_, _33976_, _33965_);
  and (_33997_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_34008_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_34019_, _34008_, _33997_);
  and (_34040_, _34019_, _33986_);
  and (_34041_, _34040_, _33954_);
  nor (_34052_, _34041_, _33289_);
  and (_34063_, _34052_, _33278_);
  or (_34073_, _34063_, _33921_);
  and (_34084_, _34073_, _33256_);
  nor (_34095_, _34084_, _33910_);
  nor (_34106_, _34095_, _33234_);
  and (_34117_, _33202_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_34128_, _34117_, _33234_);
  nor (_34139_, _34128_, _34106_);
  nor (_34150_, _34139_, _33899_);
  and (_34160_, _34150_, _33649_);
  not (_34171_, _34160_);
  and (_34182_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34193_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34204_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_34215_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_34226_, _34215_, _34204_);
  and (_34237_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_34247_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34258_, _34247_, _34237_);
  and (_34269_, _34258_, _34226_);
  and (_34280_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34291_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_34312_, _34291_, _34280_);
  and (_34313_, _34312_, _34269_);
  nor (_34324_, _34313_, _33289_);
  and (_34334_, _34324_, _33278_);
  or (_34345_, _34334_, _34193_);
  and (_34356_, _34345_, _33256_);
  nor (_34367_, _34356_, _34182_);
  nor (_34378_, _34367_, _33234_);
  and (_34389_, _33202_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34400_, _34389_, _33234_);
  nor (_34411_, _34400_, _34378_);
  not (_34421_, _34411_);
  and (_34432_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34443_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34454_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_34465_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_34476_, _34465_, _34454_);
  and (_34487_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_34498_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34508_, _34498_, _34487_);
  and (_34519_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34530_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_34541_, _34530_, _34519_);
  and (_34552_, _34541_, _34508_);
  and (_34563_, _34552_, _34476_);
  nor (_34574_, _34563_, _33289_);
  and (_34585_, _34574_, _33278_);
  nor (_34595_, _34585_, _34443_);
  nor (_34606_, _34595_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34617_, _34606_, _34432_);
  nor (_34628_, _34617_, _33234_);
  and (_34639_, _33202_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34650_, _34639_, _33234_);
  nor (_34661_, _34650_, _34628_);
  and (_34672_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_34682_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_34693_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_34704_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34715_, _34704_, _34693_);
  and (_34726_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_34737_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_34748_, _34737_, _34726_);
  and (_34759_, _34748_, _34715_);
  and (_34769_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_34780_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_34791_, _34780_, _34769_);
  and (_34802_, _34791_, _34759_);
  nor (_34813_, _34802_, _33289_);
  and (_34824_, _34813_, _33278_);
  nor (_34835_, _34824_, _34682_);
  nor (_34846_, _34835_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34857_, _34846_, _34672_);
  nor (_34867_, _34857_, _33234_);
  and (_34878_, _33202_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34889_, _34878_, _33234_);
  nor (_34900_, _34889_, _34867_);
  and (_34911_, _34900_, _34661_);
  and (_34932_, _34911_, _34421_);
  nor (_34933_, _33289_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34944_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_34954_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_34965_, _34954_, _34944_);
  and (_34976_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_34987_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_34998_, _34987_, _34976_);
  and (_35009_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_35020_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_35031_, _35020_, _35009_);
  and (_35041_, _35031_, _34998_);
  and (_35052_, _35041_, _34965_);
  and (_35063_, _35052_, _34933_);
  nor (_35074_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _33278_);
  or (_35085_, _35074_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35096_, _35085_, _35063_);
  and (_35107_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_35118_, _35107_, _35096_);
  and (_35128_, _35118_, _33224_);
  and (_35139_, _33202_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_35150_, _35139_, _33234_);
  nor (_35161_, _35150_, _35128_);
  not (_35172_, _35161_);
  not (_35183_, _34661_);
  and (_35194_, _34900_, _35183_);
  and (_35205_, _35194_, _34411_);
  and (_35215_, _35205_, _35172_);
  nor (_35226_, _35215_, _34932_);
  nor (_35237_, _35226_, _34171_);
  not (_35248_, _35237_);
  nor (_35259_, _34661_, _34411_);
  and (_35270_, _35259_, _34900_);
  and (_35281_, _35270_, _35161_);
  and (_35292_, _35281_, _34160_);
  not (_35302_, _34900_);
  and (_35313_, _35302_, _34661_);
  and (_35324_, _35161_, _34411_);
  and (_35335_, _35324_, _35313_);
  and (_35346_, _35335_, _34160_);
  nor (_35357_, _35346_, _35292_);
  and (_35368_, _35357_, _35248_);
  nor (_35379_, _34900_, _34661_);
  and (_35389_, _35379_, _34411_);
  and (_35400_, _35389_, _34160_);
  and (_35411_, _35313_, _34411_);
  and (_35422_, _35411_, _35172_);
  and (_35433_, _35422_, _34160_);
  nor (_35444_, _35433_, _35400_);
  and (_35455_, _35172_, _33649_);
  and (_35466_, _35455_, _34150_);
  and (_35476_, _35313_, _34421_);
  and (_35487_, _35476_, _35466_);
  and (_35498_, _34911_, _34411_);
  and (_35509_, _35498_, _34160_);
  nor (_35520_, _35509_, _35487_);
  and (_35531_, _35520_, _35444_);
  and (_35542_, _35531_, _35368_);
  and (_35553_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35563_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35574_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_35585_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_35596_, _35585_, _35574_);
  and (_35607_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_35618_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_35640_, _35618_, _35607_);
  and (_35641_, _35640_, _35596_);
  and (_35662_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_35663_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_35685_, _35663_, _35662_);
  and (_35686_, _35685_, _35641_);
  nor (_35708_, _35686_, _33289_);
  and (_35709_, _35708_, _33278_);
  or (_35720_, _35709_, _35563_);
  and (_35731_, _35720_, _33256_);
  nor (_35741_, _35731_, _35553_);
  nor (_35752_, _35741_, _33234_);
  and (_35763_, _33202_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_35774_, _35763_, _33234_);
  nor (_35785_, _35774_, _35752_);
  not (_35796_, _35785_);
  not (_35807_, _33899_);
  and (_35818_, _33649_, _34139_);
  and (_35828_, _35818_, _35807_);
  and (_35839_, _35828_, _35796_);
  and (_35850_, _35476_, _35161_);
  and (_35861_, _35850_, _35839_);
  and (_35872_, _35270_, _35172_);
  or (_35883_, _35872_, _35422_);
  and (_35894_, _35883_, _35839_);
  nor (_35905_, _35894_, _35861_);
  and (_35915_, _35389_, _35172_);
  and (_35926_, _35785_, _33899_);
  and (_35937_, _35926_, _35818_);
  and (_35948_, _35937_, _35915_);
  and (_35959_, _35828_, _35785_);
  and (_35970_, _35959_, _34932_);
  nor (_35981_, _35970_, _35948_);
  and (_35992_, _35161_, _34160_);
  not (_36002_, _35992_);
  and (_36013_, _35259_, _35302_);
  nor (_36024_, _36013_, _35205_);
  nor (_36035_, _36024_, _36002_);
  not (_36046_, _36035_);
  and (_36057_, _36046_, _35981_);
  and (_36068_, _36057_, _35905_);
  and (_36079_, _36068_, _35542_);
  nor (_36090_, _36079_, _33169_);
  and (_36100_, _14684_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_36111_, _35970_, _36100_);
  and (_36122_, _36111_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_36133_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_36144_, _36100_, _36133_);
  and (_36155_, _36144_, _35270_);
  and (_36166_, _36155_, _35937_);
  or (_36177_, _36166_, _36122_);
  nor (_36187_, _36177_, _36090_);
  nor (_36198_, _36187_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36209_, _36198_, _33147_);
  and (_36220_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_36231_, _35959_, _35422_);
  not (_36242_, _34139_);
  and (_36253_, _33649_, _36242_);
  and (_36264_, _35796_, _33899_);
  and (_36274_, _36264_, _36253_);
  and (_36285_, _36274_, _35335_);
  nor (_36296_, _36285_, _36231_);
  not (_36307_, _33649_);
  and (_36318_, _35850_, _36307_);
  nor (_36329_, _36318_, _35970_);
  and (_36340_, _36329_, _36296_);
  and (_36350_, _35959_, _35335_);
  and (_36361_, _35828_, _35215_);
  nor (_36372_, _36361_, _36350_);
  and (_36383_, _36274_, _35281_);
  and (_36394_, _35389_, _35161_);
  and (_36405_, _36394_, _36274_);
  nor (_36416_, _36405_, _36383_);
  and (_36427_, _36416_, _36372_);
  and (_36437_, _36427_, _36340_);
  and (_36448_, _35937_, _34932_);
  and (_36459_, _36448_, _35161_);
  and (_36470_, _35172_, _34932_);
  and (_36481_, _35498_, _35172_);
  or (_36492_, _36481_, _36470_);
  and (_36503_, _36492_, _35937_);
  nor (_36514_, _36503_, _36459_);
  and (_36525_, _36013_, _35161_);
  and (_36535_, _36525_, _36274_);
  not (_36546_, _36535_);
  and (_36557_, _35324_, _34911_);
  and (_36568_, _36557_, _36274_);
  and (_36579_, _35476_, _35992_);
  nor (_36590_, _36579_, _36568_);
  and (_36601_, _36590_, _36546_);
  and (_36612_, _36601_, _36514_);
  and (_36622_, _36612_, _36437_);
  and (_36633_, _36274_, _35915_);
  and (_36644_, _36481_, _36274_);
  nor (_36655_, _36644_, _36633_);
  and (_36666_, _35324_, _35194_);
  and (_36677_, _36666_, _36274_);
  and (_36688_, _35937_, _35476_);
  nor (_36699_, _36688_, _36677_);
  and (_36709_, _36699_, _36655_);
  and (_36720_, _35476_, _35172_);
  and (_36731_, _35959_, _36720_);
  and (_36742_, _36394_, _35959_);
  nor (_36753_, _36742_, _36731_);
  and (_36764_, _35959_, _35872_);
  and (_36775_, _36666_, _35828_);
  nor (_36786_, _36775_, _36764_);
  and (_36796_, _36786_, _36753_);
  and (_36807_, _36796_, _36709_);
  and (_36818_, _35937_, _35389_);
  and (_36829_, _35828_, _35281_);
  nor (_36840_, _36829_, _36818_);
  not (_36851_, _36840_);
  or (_36862_, _36720_, _35422_);
  and (_36873_, _36862_, _36274_);
  nor (_36882_, _36873_, _36851_);
  not (_36889_, _36274_);
  nor (_36897_, _36889_, _35226_);
  and (_36905_, _35959_, _35915_);
  and (_36912_, _35959_, _35850_);
  nor (_36920_, _36912_, _36905_);
  not (_36928_, _36920_);
  nor (_36935_, _36928_, _36897_);
  and (_36942_, _36935_, _36882_);
  and (_36943_, _36942_, _36807_);
  and (_36944_, _36943_, _36622_);
  nor (_36948_, _36944_, _33169_);
  and (_36959_, _36100_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_36970_, _36959_, _35970_);
  not (_36981_, _36970_);
  and (_36992_, _35937_, _35194_);
  and (_37003_, _36992_, _36144_);
  not (_37014_, _36144_);
  nor (_37025_, _35172_, _34411_);
  and (_37036_, _37025_, _34911_);
  and (_37047_, _37036_, _35937_);
  and (_37058_, _36481_, _35937_);
  nor (_37069_, _37058_, _37047_);
  nor (_37080_, _37069_, _37014_);
  nor (_37091_, _37080_, _37003_);
  and (_37102_, _37091_, _36981_);
  not (_37113_, _37102_);
  nor (_37124_, _37113_, _36948_);
  nor (_37135_, _37124_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37146_, _37135_, _36220_);
  nor (_37157_, _37146_, _36209_);
  and (_37168_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37179_, _35926_, _36253_);
  and (_37189_, _37179_, _35335_);
  and (_37200_, _37179_, _35850_);
  nor (_37210_, _37200_, _37189_);
  and (_37216_, _37210_, _35905_);
  nor (_37227_, _37216_, _33169_);
  not (_37238_, _37227_);
  and (_37249_, _37200_, _14684_);
  and (_37260_, _37189_, _14684_);
  nor (_37271_, _37260_, _37249_);
  nor (_37282_, _37271_, _33158_);
  nor (_37293_, _37282_, _37003_);
  and (_37304_, _37293_, _37238_);
  nor (_37315_, _37304_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37326_, _37315_, _37168_);
  and (_37337_, _37326_, _43998_);
  and (_09579_, _37337_, _37157_);
  and (_37358_, _23954_, _23449_);
  not (_37369_, _23811_);
  nor (_37380_, _37369_, _23317_);
  and (_37391_, _37380_, _37358_);
  and (_37402_, _37391_, _29174_);
  and (_37413_, _27209_, _23636_);
  and (_37424_, _37413_, _37402_);
  nor (_37435_, _37424_, _22999_);
  not (_37446_, _37424_);
  and (_37457_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_37468_, _20106_, _14750_);
  and (_37479_, _25750_, _20084_);
  nor (_37490_, _26912_, _37479_);
  and (_37500_, _37490_, _37468_);
  nor (_37511_, _26979_, _28119_);
  and (_37522_, _37511_, _37500_);
  nor (_37532_, _37522_, _15966_);
  not (_37543_, _37532_);
  and (_37554_, _37543_, _32744_);
  and (_37564_, _37554_, _32613_);
  nor (_37575_, _37564_, _37446_);
  nor (_37586_, _37575_, _37457_);
  and (_37596_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_37607_, _37522_, _17006_);
  not (_37618_, _37607_);
  and (_37628_, _37618_, _31818_);
  and (_37639_, _37628_, _31861_);
  and (_37650_, _37639_, _31709_);
  nor (_37661_, _37650_, _37446_);
  nor (_37671_, _37661_, _37596_);
  and (_37682_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_37693_, _37522_, _17180_);
  not (_37703_, _37693_);
  and (_37714_, _37703_, _30915_);
  and (_37725_, _37714_, _31155_);
  and (_37736_, _37725_, _31078_);
  nor (_37747_, _37736_, _37446_);
  nor (_37758_, _37747_, _37682_);
  and (_37769_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_37780_, _37522_, _17539_);
  not (_37791_, _37780_);
  and (_37802_, _37791_, _30362_);
  and (_37813_, _37802_, _30275_);
  and (_37824_, _37813_, _30252_);
  nor (_37835_, _37824_, _37446_);
  nor (_37846_, _37835_, _37769_);
  and (_37857_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_37868_, _37522_, _18040_);
  not (_37879_, _37868_);
  and (_37890_, _37879_, _29523_);
  and (_37901_, _37890_, _29391_);
  nor (_37912_, _37901_, _37446_);
  nor (_37923_, _37912_, _37857_);
  and (_37934_, _37446_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_37945_, _37522_, _17865_);
  not (_37956_, _37945_);
  and (_37967_, _37956_, _28800_);
  and (_37978_, _37967_, _28646_);
  nor (_37989_, _37978_, _37446_);
  nor (_38000_, _37989_, _37934_);
  nor (_38011_, _37424_, _23976_);
  nor (_38022_, _37522_, _18411_);
  not (_38033_, _38022_);
  and (_38044_, _38033_, _28229_);
  and (_38055_, _38044_, _28196_);
  and (_38066_, _38055_, _28108_);
  not (_38077_, _38066_);
  and (_38088_, _38077_, _37424_);
  nor (_38099_, _38088_, _38011_);
  and (_38110_, _38099_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38121_, _38110_, _38000_);
  and (_38132_, _38121_, _37923_);
  and (_38143_, _38132_, _37846_);
  and (_38154_, _38143_, _37758_);
  and (_38165_, _38154_, _37671_);
  and (_38176_, _38165_, _37586_);
  and (_38187_, _38176_, _37435_);
  nor (_38198_, _38176_, _37435_);
  nor (_38209_, _38198_, _38187_);
  and (_38220_, _38209_, _22988_);
  nor (_38231_, _37424_, _23119_);
  not (_38242_, _38231_);
  nor (_38253_, _38242_, _38220_);
  or (_38263_, _37522_, _16810_);
  and (_38274_, _38263_, _26901_);
  and (_38285_, _38274_, _26627_);
  and (_38295_, _38285_, _37424_);
  or (_38306_, _38295_, _38253_);
  nor (_09600_, _38306_, rst);
  not (_38326_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38337_, _38099_, _38326_);
  nor (_38348_, _38099_, _38326_);
  nor (_38359_, _38348_, _38337_);
  and (_38369_, _38359_, _22988_);
  nor (_38380_, _38369_, _23987_);
  nor (_38391_, _38380_, _37424_);
  nor (_38401_, _38391_, _38088_);
  nand (_10726_, _38401_, _43998_);
  nor (_38422_, _38110_, _38000_);
  nor (_38433_, _38422_, _38121_);
  nor (_38444_, _38433_, _22977_);
  nor (_38455_, _38444_, _24118_);
  nor (_38463_, _38455_, _37424_);
  nor (_38464_, _38463_, _37989_);
  nand (_10737_, _38464_, _43998_);
  nor (_38465_, _38121_, _37923_);
  nor (_38466_, _38465_, _38132_);
  nor (_38467_, _38466_, _22977_);
  nor (_38468_, _38467_, _24250_);
  nor (_38469_, _38468_, _37424_);
  nor (_38470_, _38469_, _37912_);
  nand (_10748_, _38470_, _43998_);
  nor (_38471_, _38132_, _37846_);
  nor (_38472_, _38471_, _38143_);
  nor (_38473_, _38472_, _22977_);
  nor (_38474_, _38473_, _23504_);
  nor (_38475_, _38474_, _37424_);
  nor (_38476_, _38475_, _37835_);
  nor (_10759_, _38476_, rst);
  nor (_38477_, _38143_, _37758_);
  nor (_38478_, _38477_, _38154_);
  nor (_38479_, _38478_, _22977_);
  nor (_38480_, _38479_, _23690_);
  nor (_38481_, _38480_, _37424_);
  nor (_38482_, _38481_, _37747_);
  nor (_10770_, _38482_, rst);
  nor (_38483_, _38154_, _37671_);
  nor (_38484_, _38483_, _38165_);
  nor (_38485_, _38484_, _22977_);
  nor (_38486_, _38485_, _23866_);
  nor (_38487_, _38486_, _37424_);
  nor (_38488_, _38487_, _37661_);
  nor (_10781_, _38488_, rst);
  nor (_38489_, _38165_, _37586_);
  nor (_38490_, _38489_, _38176_);
  nor (_38491_, _38490_, _22977_);
  nor (_38492_, _38491_, _23361_);
  nor (_38493_, _38492_, _37424_);
  nor (_38494_, _38493_, _37575_);
  nor (_10792_, _38494_, rst);
  and (_38495_, _37413_, _30612_);
  nand (_38496_, _38495_, _37391_);
  nor (_38497_, _38496_, _27132_);
  and (_38498_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _14684_);
  and (_38499_, _38498_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38500_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38501_, _38500_, _38499_);
  or (_38502_, _38501_, _38497_);
  nor (_38503_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38504_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38505_, _38504_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38506_, _38505_, _38503_);
  nor (_38507_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38508_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38509_, _38508_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38510_, _38509_, _38507_);
  nor (_38511_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38512_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38513_, _38512_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38514_, _38513_, _38511_);
  not (_38515_, _38514_);
  nor (_38516_, _38515_, _27286_);
  nor (_38517_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38518_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38519_, _38518_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38520_, _38519_, _38517_);
  and (_38521_, _38520_, _38516_);
  nor (_38522_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38523_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38524_, _38523_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38525_, _38524_, _38522_);
  and (_38526_, _38525_, _38521_);
  and (_38527_, _38526_, _38510_);
  nor (_38528_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38529_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38530_, _38529_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38531_, _38530_, _38528_);
  and (_38532_, _38531_, _38527_);
  and (_38533_, _38532_, _38506_);
  nor (_38534_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38535_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38536_, _38535_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38537_, _38536_, _38534_);
  and (_38538_, _38537_, _38533_);
  nor (_38539_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38540_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38541_, _38540_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38542_, _38541_, _38539_);
  nor (_38543_, _38542_, _38538_);
  and (_38544_, _38542_, _38538_);
  or (_38545_, _38544_, _38543_);
  nor (_38546_, _38545_, _27275_);
  not (_38547_, _38546_);
  and (_38548_, _19798_, _14750_);
  and (_38549_, _25476_, _16295_);
  not (_38550_, _38549_);
  nor (_38551_, _16810_, _15473_);
  and (_38552_, _38551_, _26210_);
  and (_38553_, _38552_, _24938_);
  and (_38554_, _38553_, _24982_);
  and (_38555_, _38554_, _25574_);
  nor (_38556_, _38555_, _26232_);
  and (_38557_, _25476_, _15308_);
  nor (_38558_, _38557_, _38556_);
  and (_38559_, _38558_, _38550_);
  and (_38560_, _26298_, _16810_);
  and (_38561_, _16142_, _15144_);
  and (_38562_, _16460_, _15473_);
  and (_38563_, _38562_, _38561_);
  and (_38564_, _38563_, _38560_);
  and (_38565_, _16295_, _15308_);
  and (_38566_, _38565_, _38564_);
  nor (_38567_, _38566_, _25476_);
  not (_38568_, _38567_);
  and (_38569_, _38568_, _38559_);
  nor (_38570_, _25476_, _15648_);
  and (_38571_, _25476_, _15648_);
  nor (_38572_, _38571_, _38570_);
  and (_38573_, _38572_, _38569_);
  and (_38574_, _38573_, _26419_);
  nor (_38575_, _38573_, _26419_);
  nor (_38576_, _38575_, _38574_);
  and (_38577_, _38576_, _26364_);
  and (_38578_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38579_, _25476_, _26419_);
  nor (_38580_, _38579_, _27385_);
  nor (_38581_, _38580_, _26474_);
  nor (_38582_, _27461_, _17539_);
  nor (_38583_, _26923_, _16634_);
  or (_38584_, _38583_, _38582_);
  or (_38585_, _38584_, _38581_);
  nor (_38586_, _38585_, _38578_);
  not (_38587_, _38586_);
  nor (_38588_, _38587_, _38577_);
  not (_38589_, _38588_);
  nor (_38590_, _38589_, _38548_);
  and (_38591_, _38590_, _38547_);
  nand (_38592_, _38591_, _38499_);
  and (_38593_, _38592_, _43998_);
  and (_12736_, _38593_, _38502_);
  and (_38594_, _37413_, _29916_);
  and (_38595_, _38594_, _37391_);
  nor (_38596_, _38595_, _38499_);
  not (_38597_, _38596_);
  nand (_38598_, _38597_, _27132_);
  not (_38599_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_38600_, _38596_, _38599_);
  and (_38601_, _38600_, _43998_);
  and (_12757_, _38601_, _38598_);
  nor (_38602_, _38496_, _28372_);
  and (_38603_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38604_, _38603_, _38499_);
  or (_38605_, _38604_, _38602_);
  and (_38606_, _22377_, _20106_);
  not (_38607_, _38606_);
  and (_38608_, _38515_, _27286_);
  nor (_38609_, _38608_, _38516_);
  and (_38610_, _38609_, _25761_);
  nor (_38611_, _27385_, _26452_);
  not (_38612_, _38611_);
  nor (_38613_, _38612_, _26320_);
  nor (_38614_, _38613_, _24905_);
  and (_38615_, _38613_, _24905_);
  nor (_38616_, _38615_, _38614_);
  and (_38617_, _38616_, _26364_);
  nor (_38618_, _26923_, _15473_);
  and (_38619_, _19575_, _14750_);
  nor (_38620_, _27461_, _17180_);
  nor (_38621_, _26474_, _18411_);
  or (_38622_, _38621_, _38620_);
  or (_38623_, _38622_, _38619_);
  nor (_38624_, _38623_, _38618_);
  not (_38625_, _38624_);
  nor (_38626_, _38625_, _38617_);
  not (_38627_, _38626_);
  nor (_38628_, _38627_, _38610_);
  and (_38629_, _38628_, _38607_);
  nand (_38630_, _38629_, _38499_);
  and (_38631_, _38630_, _43998_);
  and (_13557_, _38631_, _38605_);
  nor (_38632_, _38496_, _29086_);
  and (_38633_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38634_, _38633_, _38499_);
  or (_38635_, _38634_, _38632_);
  nor (_38636_, _38520_, _38516_);
  nor (_38637_, _38636_, _38521_);
  and (_38638_, _38637_, _25761_);
  not (_38639_, _38638_);
  and (_38640_, _21391_, _20106_);
  nor (_38641_, _26923_, _16460_);
  and (_38642_, _38552_, _25476_);
  and (_38643_, _38560_, _15473_);
  and (_38644_, _38643_, _26232_);
  nor (_38645_, _38644_, _38642_);
  and (_38646_, _38645_, _16460_);
  nor (_38647_, _38645_, _16460_);
  or (_38648_, _38647_, _26375_);
  nor (_38649_, _38648_, _38646_);
  and (_38650_, _19607_, _14750_);
  nor (_38651_, _27461_, _17006_);
  nor (_38652_, _26474_, _17865_);
  or (_38653_, _38652_, _38651_);
  or (_38654_, _38653_, _38650_);
  or (_38655_, _38654_, _38649_);
  nor (_38656_, _38655_, _38641_);
  not (_38657_, _38656_);
  nor (_38658_, _38657_, _38640_);
  and (_38659_, _38658_, _38639_);
  nand (_38660_, _38659_, _38499_);
  and (_38661_, _38660_, _43998_);
  and (_13568_, _38661_, _38635_);
  nor (_38662_, _38496_, _29763_);
  and (_38663_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38664_, _38663_, _38499_);
  or (_38665_, _38664_, _38662_);
  nor (_38666_, _38525_, _38521_);
  nor (_38667_, _38666_, _38526_);
  and (_38668_, _38667_, _25761_);
  not (_38669_, _38668_);
  and (_38670_, _38643_, _16460_);
  and (_38671_, _38670_, _26232_);
  and (_38672_, _38553_, _25476_);
  nor (_38673_, _38672_, _38671_);
  and (_38674_, _38673_, _15144_);
  nor (_38675_, _38673_, _15144_);
  nor (_38676_, _38675_, _38674_);
  and (_38677_, _38676_, _26364_);
  not (_38678_, _38677_);
  nor (_38679_, _26474_, _18040_);
  and (_38680_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38681_, _38680_, _38679_);
  and (_38682_, _19639_, _14750_);
  nor (_38683_, _27461_, _15966_);
  nor (_38684_, _26923_, _15144_);
  or (_38685_, _38684_, _38683_);
  nor (_38686_, _38685_, _38682_);
  and (_38687_, _38686_, _38681_);
  and (_38688_, _38687_, _38678_);
  and (_38689_, _38688_, _38669_);
  nand (_38690_, _38689_, _38499_);
  and (_38691_, _38690_, _43998_);
  and (_13579_, _38691_, _38665_);
  nor (_38692_, _38496_, _30514_);
  and (_38693_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38694_, _38693_, _38499_);
  or (_38695_, _38694_, _38692_);
  nor (_38696_, _38526_, _38510_);
  not (_38697_, _38696_);
  nor (_38698_, _38527_, _27275_);
  and (_38699_, _38698_, _38697_);
  not (_38700_, _38699_);
  and (_38701_, _19671_, _14750_);
  nor (_38702_, _38554_, _25574_);
  not (_38703_, _38702_);
  and (_38704_, _38703_, _38556_);
  and (_38705_, _38670_, _15144_);
  nor (_38706_, _38705_, _16142_);
  nor (_38707_, _38706_, _38564_);
  nor (_38708_, _38707_, _25476_);
  nor (_38709_, _38708_, _38704_);
  nor (_38710_, _38709_, _26375_);
  nor (_38711_, _26923_, _16142_);
  nor (_38712_, _26474_, _17539_);
  and (_38713_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38714_, _38713_, _38712_);
  or (_38715_, _38714_, _27472_);
  nor (_38716_, _38715_, _38711_);
  not (_38717_, _38716_);
  nor (_38718_, _38717_, _38710_);
  not (_38719_, _38718_);
  nor (_38720_, _38719_, _38701_);
  and (_38721_, _38720_, _38700_);
  nand (_38722_, _38721_, _38499_);
  and (_38723_, _38722_, _43998_);
  and (_13590_, _38723_, _38695_);
  nor (_38724_, _38496_, _31285_);
  and (_38725_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38726_, _38725_, _38499_);
  or (_38727_, _38726_, _38724_);
  nor (_38728_, _38531_, _38527_);
  not (_38729_, _38728_);
  nor (_38730_, _38532_, _27275_);
  and (_38731_, _38730_, _38729_);
  not (_38732_, _38731_);
  and (_38733_, _19702_, _14750_);
  nor (_38735_, _38564_, _25476_);
  nor (_38738_, _38735_, _38556_);
  nor (_38739_, _38738_, _24630_);
  and (_38740_, _38738_, _24630_);
  nor (_38741_, _38740_, _38739_);
  and (_38742_, _38741_, _26364_);
  and (_38743_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38744_, _25476_, _17191_);
  or (_38745_, _38744_, _26474_);
  nor (_38746_, _38745_, _38557_);
  nor (_38747_, _27461_, _18411_);
  nor (_38748_, _26923_, _15308_);
  or (_38756_, _38748_, _38747_);
  or (_38762_, _38756_, _38746_);
  nor (_38768_, _38762_, _38743_);
  not (_38773_, _38768_);
  nor (_38774_, _38773_, _38742_);
  not (_38775_, _38774_);
  nor (_38776_, _38775_, _38733_);
  and (_38777_, _38776_, _38732_);
  nand (_38778_, _38777_, _38499_);
  and (_38779_, _38778_, _43998_);
  and (_13601_, _38779_, _38727_);
  nor (_38780_, _38496_, _32102_);
  and (_38781_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38782_, _38781_, _38499_);
  or (_38783_, _38782_, _38780_);
  nor (_38784_, _38532_, _38506_);
  nor (_38785_, _38784_, _38533_);
  and (_38786_, _38785_, _25761_);
  not (_38787_, _38786_);
  and (_38788_, _19734_, _14750_);
  and (_38789_, _38564_, _15308_);
  nor (_38790_, _38789_, _25476_);
  not (_38791_, _38790_);
  and (_38792_, _38791_, _38558_);
  and (_38793_, _38792_, _16295_);
  nor (_38794_, _38792_, _16295_);
  or (_38795_, _38794_, _38793_);
  and (_38796_, _38795_, _26364_);
  nor (_38797_, _32515_, _26474_);
  and (_38800_, _38797_, _38550_);
  nor (_38801_, _26923_, _16295_);
  nor (_38802_, _27461_, _17865_);
  and (_38803_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_38804_, _38803_, _38802_);
  nor (_38805_, _38804_, _38801_);
  not (_38806_, _38805_);
  nor (_38807_, _38806_, _38800_);
  not (_38808_, _38807_);
  nor (_38809_, _38808_, _38796_);
  not (_38810_, _38809_);
  nor (_38811_, _38810_, _38788_);
  and (_38812_, _38811_, _38787_);
  nand (_38813_, _38812_, _38499_);
  and (_38814_, _38813_, _43998_);
  and (_13612_, _38814_, _38783_);
  nor (_38815_, _38496_, _32919_);
  and (_38816_, _38496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38817_, _38816_, _38499_);
  or (_38818_, _38817_, _38815_);
  nor (_38819_, _38537_, _38533_);
  not (_38820_, _38819_);
  nor (_38821_, _38538_, _27275_);
  and (_38822_, _38821_, _38820_);
  not (_38823_, _38822_);
  and (_38824_, _19766_, _14750_);
  and (_38825_, _38569_, _15648_);
  nor (_38826_, _38569_, _15648_);
  nor (_38827_, _38826_, _38825_);
  nor (_38828_, _38827_, _26375_);
  and (_38829_, _20106_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38830_, _25476_, _15977_);
  or (_38831_, _38830_, _26474_);
  nor (_38832_, _38831_, _38571_);
  nor (_38833_, _27461_, _18040_);
  nor (_38834_, _26923_, _15648_);
  or (_38835_, _38834_, _38833_);
  or (_38836_, _38835_, _38832_);
  nor (_38838_, _38836_, _38829_);
  not (_38842_, _38838_);
  nor (_38848_, _38842_, _38828_);
  not (_38853_, _38848_);
  nor (_38860_, _38853_, _38824_);
  and (_38868_, _38860_, _38823_);
  nand (_38876_, _38868_, _38499_);
  and (_38877_, _38876_, _43998_);
  and (_13623_, _38877_, _38818_);
  nand (_38878_, _38597_, _28372_);
  not (_38879_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_38880_, _38596_, _38879_);
  and (_38881_, _38880_, _43998_);
  and (_13633_, _38881_, _38878_);
  nand (_38882_, _38597_, _29086_);
  not (_38883_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_38884_, _38596_, _38883_);
  and (_38885_, _38884_, _43998_);
  and (_13644_, _38885_, _38882_);
  nand (_38886_, _38597_, _29763_);
  not (_38887_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_38888_, _38596_, _38887_);
  and (_38889_, _38888_, _43998_);
  and (_13655_, _38889_, _38886_);
  nand (_38890_, _38597_, _30514_);
  or (_38891_, _38597_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38892_, _38891_, _43998_);
  and (_13666_, _38892_, _38890_);
  nand (_38893_, _38597_, _31285_);
  or (_38894_, _38597_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38895_, _38894_, _43998_);
  and (_13677_, _38895_, _38893_);
  nand (_38896_, _38597_, _32102_);
  or (_38897_, _38597_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38898_, _38897_, _43998_);
  and (_13688_, _38898_, _38896_);
  nand (_38899_, _38597_, _32919_);
  or (_38900_, _38597_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38901_, _38900_, _43998_);
  and (_13699_, _38901_, _38899_);
  and (_38902_, _23954_, _23822_);
  and (_38903_, _38902_, _23460_);
  and (_38904_, _38903_, _27900_);
  nor (_38905_, _33006_, _27790_);
  not (_38910_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38921_, _27867_, _38910_);
  or (_38923_, _38921_, _38905_);
  and (_38924_, _38923_, _38904_);
  nor (_38925_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38935_, _38925_);
  nand (_38942_, _38935_, _27790_);
  and (_38943_, _38925_, _38910_);
  not (_38944_, _23449_);
  and (_38945_, _38902_, _38944_);
  and (_38946_, _27900_, _27812_);
  and (_38947_, _38946_, _38945_);
  nor (_38948_, _38947_, _38943_);
  and (_38949_, _38948_, _38942_);
  and (_38950_, _27209_, _24376_);
  and (_38951_, _38950_, _38903_);
  or (_38952_, _38951_, _38949_);
  or (_38953_, _38952_, _38924_);
  nand (_38954_, _38951_, _38285_);
  and (_38955_, _38954_, _38953_);
  and (_16678_, _38955_, _43998_);
  not (_38956_, _38951_);
  not (_38957_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_38958_, _38904_, _29174_);
  nand (_38959_, _38958_, _38957_);
  and (_38960_, _38959_, _38956_);
  or (_38961_, _38958_, _28460_);
  and (_38962_, _38961_, _38960_);
  nor (_38963_, _38956_, _37978_);
  or (_38964_, _38963_, _38962_);
  and (_21609_, _38964_, _43998_);
  not (_38965_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38966_, _29916_, _38965_);
  or (_38967_, _38966_, _29927_);
  and (_38968_, _38967_, _38904_);
  or (_38969_, _19861_, _19829_);
  or (_38970_, _38969_, _19893_);
  or (_38971_, _38970_, _19936_);
  or (_38972_, _38971_, _20010_);
  or (_38973_, _38972_, _20042_);
  and (_38974_, _38973_, _14750_);
  or (_38975_, _27330_, _25683_);
  not (_38976_, _27319_);
  nand (_38977_, _38976_, _25683_);
  and (_38978_, _38977_, _24465_);
  and (_38979_, _38978_, _38975_);
  not (_38980_, _24487_);
  nand (_38981_, _26101_, _38980_);
  or (_38982_, _26101_, _24498_);
  and (_38983_, _25761_, _38982_);
  and (_38984_, _38983_, _38981_);
  and (_38985_, _38565_, _21293_);
  and (_38986_, _38563_, _20106_);
  nand (_38987_, _38986_, _38985_);
  nand (_38988_, _38987_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38989_, _38988_, _38984_);
  or (_38990_, _38989_, _38979_);
  or (_38991_, _38990_, _30774_);
  or (_38992_, _38991_, _24432_);
  or (_38993_, _38992_, _38974_);
  nor (_38994_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38995_, _38994_, _38904_);
  and (_38996_, _38995_, _38993_);
  or (_38997_, _38996_, _38968_);
  and (_38998_, _38997_, _38956_);
  nor (_38999_, _38956_, _37901_);
  or (_39000_, _38999_, _38998_);
  and (_21621_, _39000_, _43998_);
  not (_39001_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_39002_, _38904_, _30612_);
  nand (_39003_, _39002_, _39001_);
  and (_39004_, _39003_, _38956_);
  or (_39005_, _39002_, _28460_);
  and (_39006_, _39005_, _39004_);
  nor (_39007_, _38956_, _37824_);
  or (_39008_, _39007_, _39006_);
  and (_21633_, _39008_, _43998_);
  not (_39009_, _38947_);
  or (_39010_, _39009_, _31416_);
  and (_39011_, _39010_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_39012_, _31405_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39013_, _39012_, _31459_);
  and (_39014_, _39013_, _38904_);
  or (_39015_, _39014_, _39011_);
  and (_39016_, _39015_, _38956_);
  nor (_39017_, _38956_, _37736_);
  or (_39018_, _39017_, _39016_);
  and (_21645_, _39018_, _43998_);
  or (_39019_, _39009_, _32200_);
  and (_39020_, _39019_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_39021_, _39020_, _38951_);
  and (_39022_, _32276_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_39023_, _39022_, _32265_);
  and (_39024_, _39023_, _38904_);
  or (_39025_, _39024_, _39021_);
  nand (_39026_, _38951_, _37650_);
  and (_39027_, _39026_, _39025_);
  and (_21657_, _39027_, _43998_);
  nor (_39028_, _33039_, _30286_);
  or (_39029_, _39028_, _33050_);
  and (_39030_, _39029_, _38904_);
  and (_39031_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_39032_, _39031_, _26923_);
  and (_39033_, _39032_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_39034_, _25761_, _26024_);
  and (_39035_, _25629_, _24465_);
  or (_39036_, _39035_, _39034_);
  and (_39037_, _39036_, _39031_);
  nor (_39038_, _39037_, _39033_);
  nor (_39039_, _39038_, _38904_);
  or (_39040_, _39039_, _39030_);
  and (_39041_, _39040_, _38956_);
  nor (_39042_, _38956_, _37564_);
  or (_39043_, _39042_, _39041_);
  and (_21668_, _39043_, _43998_);
  not (_39044_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39045_, _38498_, _39044_);
  and (_39046_, _39045_, _38591_);
  nor (_39047_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39048_, _39047_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39049_, _24376_, _23636_);
  and (_39050_, _23965_, _23811_);
  and (_39051_, _39050_, _23460_);
  and (_39052_, _39051_, _39049_);
  and (_39053_, _39052_, _27209_);
  nor (_39054_, _39053_, _39048_);
  nor (_39055_, _39054_, _27132_);
  not (_39056_, _39045_);
  and (_39057_, _23811_, _23636_);
  and (_39058_, _39057_, _27801_);
  and (_39059_, _39058_, _38946_);
  and (_39060_, _39059_, _27867_);
  and (_39061_, _39060_, _27790_);
  not (_39062_, _39054_);
  nor (_39063_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_39064_, _39063_, _39062_);
  or (_39065_, _39064_, _39061_);
  and (_39066_, _39065_, _39056_);
  not (_39067_, _39066_);
  nor (_39068_, _39067_, _39055_);
  nor (_39069_, _39068_, _39046_);
  and (_22437_, _39069_, _43998_);
  and (_39070_, _39045_, _38629_);
  nor (_39071_, _39054_, _28372_);
  and (_39072_, _39059_, _24376_);
  and (_39073_, _39072_, _27790_);
  nor (_39074_, _39072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_39075_, _39074_, _39062_);
  or (_39076_, _39075_, _39073_);
  and (_39077_, _39076_, _39056_);
  not (_39078_, _39077_);
  nor (_39079_, _39078_, _39071_);
  nor (_39080_, _39079_, _39070_);
  and (_24305_, _39080_, _43998_);
  and (_39081_, _39045_, _38659_);
  nor (_39082_, _39054_, _29086_);
  and (_39083_, _39059_, _29174_);
  and (_39084_, _39083_, _27790_);
  nor (_39085_, _39083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_39086_, _39085_, _39062_);
  or (_39087_, _39086_, _39084_);
  and (_39088_, _39087_, _39056_);
  not (_39089_, _39088_);
  nor (_39090_, _39089_, _39082_);
  nor (_39091_, _39090_, _39081_);
  and (_24317_, _39091_, _43998_);
  nor (_39092_, _39056_, _38689_);
  and (_39093_, _39062_, _29763_);
  not (_39094_, _39059_);
  not (_39095_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_39096_, _29916_, _39095_);
  nor (_39097_, _39096_, _29927_);
  nor (_39098_, _39097_, _39094_);
  nor (_39099_, _39059_, _39095_);
  nor (_39100_, _39099_, _39062_);
  not (_39101_, _39100_);
  nor (_39102_, _39101_, _39098_);
  nor (_39103_, _39102_, _39045_);
  not (_39104_, _39103_);
  nor (_39105_, _39104_, _39093_);
  nor (_39106_, _39105_, _39092_);
  nor (_24329_, _39106_, rst);
  nor (_39107_, _39056_, _38721_);
  and (_39108_, _39062_, _30514_);
  not (_39109_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39110_, _30612_, _39109_);
  nor (_39111_, _39110_, _30634_);
  nor (_39112_, _39111_, _39094_);
  nor (_39113_, _39059_, _39109_);
  nor (_39114_, _39113_, _39062_);
  not (_39115_, _39114_);
  nor (_39116_, _39115_, _39112_);
  nor (_39117_, _39116_, _39045_);
  not (_39118_, _39117_);
  nor (_39126_, _39118_, _39108_);
  nor (_39137_, _39126_, _39107_);
  nor (_24341_, _39137_, rst);
  and (_39157_, _39045_, _38777_);
  nor (_39163_, _39054_, _31285_);
  and (_39173_, _39059_, _31394_);
  and (_39184_, _39173_, _27790_);
  nor (_39195_, _39173_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_39206_, _39195_, _39062_);
  or (_39217_, _39206_, _39184_);
  and (_39228_, _39217_, _39056_);
  not (_39239_, _39228_);
  nor (_39250_, _39239_, _39163_);
  nor (_39261_, _39250_, _39157_);
  and (_24353_, _39261_, _43998_);
  and (_39282_, _39045_, _38812_);
  nor (_39293_, _39054_, _32102_);
  and (_39304_, _39059_, _32243_);
  and (_39315_, _39304_, _27790_);
  nor (_39326_, _39304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_39331_, _39326_, _39062_);
  or (_39332_, _39331_, _39315_);
  and (_39333_, _39332_, _39056_);
  not (_39334_, _39333_);
  nor (_39335_, _39334_, _39293_);
  nor (_39336_, _39335_, _39282_);
  and (_24365_, _39336_, _43998_);
  and (_39337_, _39045_, _38868_);
  nor (_39338_, _39054_, _32919_);
  and (_39339_, _39059_, _33039_);
  and (_39340_, _39339_, _27790_);
  nor (_39341_, _39339_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_39342_, _39341_, _39062_);
  or (_39343_, _39342_, _39340_);
  and (_39344_, _39343_, _39056_);
  not (_39345_, _39344_);
  nor (_39346_, _39345_, _39338_);
  nor (_39347_, _39346_, _39337_);
  and (_24377_, _39347_, _43998_);
  and (_39348_, _39057_, _27812_);
  and (_39349_, _39348_, _37358_);
  and (_39350_, _39349_, _27867_);
  nand (_39351_, _39350_, _27790_);
  or (_39352_, _39350_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39353_, _39352_, _27900_);
  and (_39354_, _39353_, _39351_);
  and (_39355_, _37391_, _39049_);
  nand (_39356_, _39355_, _38285_);
  or (_39357_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39358_, _39357_, _27209_);
  and (_39359_, _39358_, _39356_);
  not (_39360_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39361_, _27198_, _39360_);
  or (_39362_, _39361_, rst);
  or (_39363_, _39362_, _39359_);
  or (_35629_, _39363_, _39354_);
  nor (_39364_, _38944_, _23317_);
  and (_39365_, _38902_, _39364_);
  and (_39366_, _39365_, _27867_);
  nand (_39367_, _39366_, _27790_);
  or (_39368_, _39366_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39369_, _39368_, _27900_);
  and (_39370_, _39369_, _39367_);
  and (_39371_, _39365_, _24376_);
  not (_39372_, _39371_);
  nor (_39373_, _39372_, _38285_);
  not (_39374_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39375_, _39371_, _39374_);
  or (_39376_, _39375_, _39373_);
  and (_39377_, _39376_, _27209_);
  nor (_39378_, _27198_, _39374_);
  or (_39379_, _39378_, rst);
  or (_39380_, _39379_, _39377_);
  or (_35651_, _39380_, _39370_);
  and (_39381_, _23965_, _23449_);
  and (_39382_, _39381_, _39348_);
  and (_39383_, _39382_, _27867_);
  nand (_39384_, _39383_, _27790_);
  or (_39385_, _39383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39386_, _39385_, _27900_);
  and (_39387_, _39386_, _39384_);
  and (_39388_, _39057_, _24388_);
  and (_39389_, _39388_, _39364_);
  not (_39390_, _39389_);
  nor (_39391_, _39390_, _38285_);
  not (_39392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39393_, _39389_, _39392_);
  or (_39394_, _39393_, _39391_);
  and (_39395_, _39394_, _27209_);
  nor (_39396_, _27198_, _39392_);
  or (_39397_, _39396_, rst);
  or (_39398_, _39397_, _39395_);
  or (_35674_, _39398_, _39387_);
  and (_39399_, _39381_, _27823_);
  not (_39400_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_39401_, _27867_, _39400_);
  or (_39402_, _39401_, _38905_);
  and (_39403_, _39402_, _39399_);
  nor (_39404_, _39399_, _39400_);
  or (_39405_, _39404_, _39403_);
  and (_39406_, _39405_, _27900_);
  and (_39407_, _39364_, _24389_);
  not (_39408_, _39407_);
  nor (_39409_, _39408_, _38285_);
  nor (_39410_, _39407_, _39400_);
  or (_39411_, _39410_, _39409_);
  and (_39412_, _39411_, _27209_);
  nor (_39413_, _27198_, _39400_);
  or (_39414_, _39413_, rst);
  or (_39415_, _39414_, _39412_);
  or (_35697_, _39415_, _39406_);
  or (_39416_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_39417_, _39355_, _27790_);
  and (_39418_, _39417_, _27900_);
  nand (_39419_, _39355_, _38066_);
  and (_39420_, _39419_, _27209_);
  or (_39421_, _39420_, _39418_);
  and (_39422_, _39421_, _39416_);
  not (_39423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39424_, _27198_, _39423_);
  or (_39425_, _39424_, rst);
  or (_41282_, _39425_, _39422_);
  and (_39426_, _39349_, _29174_);
  nand (_39427_, _39426_, _27790_);
  or (_39428_, _39426_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39429_, _39428_, _27900_);
  and (_39430_, _39429_, _39427_);
  nand (_39431_, _39355_, _37978_);
  or (_39432_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39433_, _39432_, _27209_);
  and (_39434_, _39433_, _39431_);
  not (_39435_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_39436_, _27198_, _39435_);
  or (_39437_, _39436_, rst);
  or (_39438_, _39437_, _39434_);
  or (_41284_, _39438_, _39430_);
  not (_39439_, _30655_);
  nand (_39440_, _39349_, _39439_);
  and (_39441_, _39440_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39442_, _24364_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39443_, _39442_, _29927_);
  and (_39444_, _39443_, _39349_);
  or (_39445_, _39444_, _39441_);
  and (_39446_, _39445_, _27900_);
  nand (_39447_, _39355_, _37901_);
  or (_39448_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39449_, _39448_, _27209_);
  and (_39450_, _39449_, _39447_);
  not (_39451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_39452_, _27198_, _39451_);
  or (_39453_, _39452_, rst);
  or (_39454_, _39453_, _39450_);
  or (_41286_, _39454_, _39446_);
  nand (_39455_, _39349_, _24352_);
  and (_39456_, _39455_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39457_, _39439_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39458_, _39457_, _30634_);
  and (_39459_, _39458_, _39349_);
  or (_39460_, _39459_, _39456_);
  and (_39461_, _39460_, _27900_);
  nand (_39462_, _39355_, _37824_);
  or (_39463_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39464_, _39463_, _27209_);
  and (_39465_, _39464_, _39462_);
  not (_39466_, _27198_);
  and (_39467_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39468_, _39467_, rst);
  or (_39469_, _39468_, _39465_);
  or (_41288_, _39469_, _39461_);
  and (_39470_, _39349_, _31394_);
  nand (_39471_, _39470_, _27790_);
  or (_39472_, _39470_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39473_, _39472_, _27900_);
  and (_39474_, _39473_, _39471_);
  nand (_39475_, _39355_, _37736_);
  or (_39476_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39477_, _39476_, _27209_);
  and (_39478_, _39477_, _39475_);
  and (_39479_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39480_, _39479_, rst);
  or (_39481_, _39480_, _39478_);
  or (_41290_, _39481_, _39474_);
  and (_39482_, _39349_, _32243_);
  nand (_39483_, _39482_, _27790_);
  or (_39484_, _39482_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39485_, _39484_, _27900_);
  and (_39486_, _39485_, _39483_);
  nand (_39487_, _39355_, _37650_);
  or (_39488_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39489_, _39488_, _27209_);
  and (_39490_, _39489_, _39487_);
  and (_39491_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39492_, _39491_, rst);
  or (_39493_, _39492_, _39490_);
  or (_41292_, _39493_, _39486_);
  nand (_39494_, _39349_, _33006_);
  and (_39495_, _39494_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_39496_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_39497_, _27856_, _39496_);
  or (_39498_, _39497_, _33050_);
  and (_39499_, _39498_, _39349_);
  or (_39500_, _39499_, _39495_);
  and (_39501_, _39500_, _27900_);
  nand (_39502_, _39355_, _37564_);
  or (_39503_, _39355_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39504_, _39503_, _27209_);
  and (_39505_, _39504_, _39502_);
  nor (_39506_, _27198_, _39496_);
  or (_39507_, _39506_, rst);
  or (_39508_, _39507_, _39505_);
  or (_41294_, _39508_, _39501_);
  nand (_39509_, _39371_, _27790_);
  or (_39510_, _39371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39511_, _39510_, _27900_);
  and (_39512_, _39511_, _39509_);
  and (_39513_, _39371_, _38077_);
  not (_39514_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39515_, _39371_, _39514_);
  or (_39516_, _39515_, _39513_);
  and (_39517_, _39516_, _27209_);
  nor (_39518_, _27198_, _39514_);
  or (_39519_, _39518_, rst);
  or (_39520_, _39519_, _39517_);
  or (_41295_, _39520_, _39512_);
  and (_39521_, _39365_, _29174_);
  nand (_39522_, _39521_, _27790_);
  or (_39523_, _39521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39524_, _39523_, _27900_);
  and (_39525_, _39524_, _39522_);
  nor (_39526_, _39372_, _37978_);
  not (_39527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_39528_, _39371_, _39527_);
  or (_39529_, _39528_, _39526_);
  and (_39530_, _39529_, _27209_);
  nor (_39531_, _27198_, _39527_);
  or (_39532_, _39531_, rst);
  or (_39533_, _39532_, _39530_);
  or (_41297_, _39533_, _39525_);
  and (_39534_, _39365_, _29916_);
  nand (_39535_, _39534_, _27790_);
  or (_39536_, _39534_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39537_, _39536_, _27900_);
  and (_39539_, _39537_, _39535_);
  nor (_39540_, _39372_, _37901_);
  not (_39541_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_39542_, _39371_, _39541_);
  or (_39543_, _39542_, _39540_);
  and (_39544_, _39543_, _27209_);
  nor (_39545_, _27198_, _39541_);
  or (_39546_, _39545_, rst);
  or (_39547_, _39546_, _39544_);
  or (_41299_, _39547_, _39539_);
  and (_39548_, _39365_, _30612_);
  nand (_39549_, _39548_, _27790_);
  or (_39550_, _39548_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39551_, _39550_, _27900_);
  and (_39552_, _39551_, _39549_);
  nor (_39553_, _39372_, _37824_);
  and (_39554_, _39372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39555_, _39554_, _39553_);
  and (_39556_, _39555_, _27209_);
  and (_39557_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39558_, _39557_, rst);
  or (_39559_, _39558_, _39556_);
  or (_41301_, _39559_, _39552_);
  and (_39560_, _39365_, _31394_);
  nand (_39561_, _39560_, _27790_);
  or (_39562_, _39560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39563_, _39562_, _27900_);
  and (_39564_, _39563_, _39561_);
  nor (_39565_, _39372_, _37736_);
  and (_39566_, _39372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39568_, _39566_, _39565_);
  and (_39572_, _39568_, _27209_);
  and (_39573_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39574_, _39573_, rst);
  or (_39575_, _39574_, _39572_);
  or (_41303_, _39575_, _39564_);
  and (_39576_, _39365_, _32243_);
  nand (_39577_, _39576_, _27790_);
  or (_39578_, _39576_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39579_, _39578_, _27900_);
  and (_39580_, _39579_, _39577_);
  nor (_39581_, _39372_, _37650_);
  and (_39582_, _39372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39583_, _39582_, _39581_);
  and (_39584_, _39583_, _27209_);
  and (_39585_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39586_, _39585_, rst);
  or (_39587_, _39586_, _39584_);
  or (_41305_, _39587_, _39580_);
  and (_39588_, _39365_, _33039_);
  nand (_39589_, _39588_, _27790_);
  or (_39590_, _39588_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39591_, _39590_, _27900_);
  and (_39592_, _39591_, _39589_);
  nor (_39593_, _39372_, _37564_);
  not (_39594_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_39595_, _39371_, _39594_);
  or (_39596_, _39595_, _39593_);
  and (_39597_, _39596_, _27209_);
  nor (_39598_, _27198_, _39594_);
  or (_39599_, _39598_, rst);
  or (_39600_, _39599_, _39597_);
  or (_41306_, _39600_, _39592_);
  and (_39601_, _39382_, _24376_);
  nand (_39602_, _39601_, _27790_);
  or (_39603_, _39601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39604_, _39603_, _27900_);
  and (_39605_, _39604_, _39602_);
  nor (_39606_, _39390_, _38066_);
  not (_39607_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39608_, _39389_, _39607_);
  or (_39609_, _39608_, _39606_);
  and (_39610_, _39609_, _27209_);
  nor (_39611_, _27198_, _39607_);
  or (_39612_, _39611_, rst);
  or (_39613_, _39612_, _39610_);
  or (_41308_, _39613_, _39605_);
  and (_39614_, _39382_, _29174_);
  nand (_39615_, _39614_, _27790_);
  or (_39616_, _39614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39617_, _39616_, _27900_);
  and (_39618_, _39617_, _39615_);
  nor (_39619_, _39390_, _37978_);
  not (_39620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_39621_, _39389_, _39620_);
  or (_39622_, _39621_, _39619_);
  and (_39623_, _39622_, _27209_);
  nor (_39624_, _27198_, _39620_);
  or (_39625_, _39624_, rst);
  or (_39626_, _39625_, _39623_);
  or (_41310_, _39626_, _39618_);
  and (_39627_, _39382_, _29916_);
  nand (_39628_, _39627_, _27790_);
  or (_39630_, _39627_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39637_, _39630_, _27900_);
  and (_39638_, _39637_, _39628_);
  nor (_39639_, _39390_, _37901_);
  not (_39640_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_39641_, _39389_, _39640_);
  or (_39642_, _39641_, _39639_);
  and (_39643_, _39642_, _27209_);
  nor (_39644_, _27198_, _39640_);
  or (_39645_, _39644_, rst);
  or (_39646_, _39645_, _39643_);
  or (_41312_, _39646_, _39638_);
  and (_39647_, _39382_, _30612_);
  nand (_39648_, _39647_, _27790_);
  or (_39649_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39650_, _39649_, _27900_);
  and (_39651_, _39650_, _39648_);
  nor (_39652_, _39390_, _37824_);
  and (_39653_, _39390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39654_, _39653_, _39652_);
  and (_39655_, _39654_, _27209_);
  and (_39656_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39657_, _39656_, rst);
  or (_39658_, _39657_, _39655_);
  or (_41314_, _39658_, _39651_);
  and (_39659_, _39382_, _31394_);
  nand (_39660_, _39659_, _27790_);
  or (_39661_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39662_, _39661_, _27900_);
  and (_39663_, _39662_, _39660_);
  nor (_39664_, _39390_, _37736_);
  and (_39665_, _39390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39666_, _39665_, _39664_);
  and (_39667_, _39666_, _27209_);
  and (_39668_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39669_, _39668_, rst);
  or (_39670_, _39669_, _39667_);
  or (_41316_, _39670_, _39663_);
  and (_39671_, _39382_, _32243_);
  nand (_39672_, _39671_, _27790_);
  or (_39673_, _39671_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39674_, _39673_, _27900_);
  and (_39675_, _39674_, _39672_);
  nor (_39676_, _39390_, _37650_);
  and (_39677_, _39390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39678_, _39677_, _39676_);
  and (_39679_, _39678_, _27209_);
  and (_39680_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39685_, _39680_, rst);
  or (_39686_, _39685_, _39679_);
  or (_41317_, _39686_, _39675_);
  and (_39687_, _39382_, _33039_);
  nand (_39688_, _39687_, _27790_);
  or (_39689_, _39687_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39690_, _39689_, _27900_);
  and (_39691_, _39690_, _39688_);
  nor (_39692_, _39390_, _37564_);
  not (_39693_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_39694_, _39389_, _39693_);
  or (_39695_, _39694_, _39692_);
  and (_39696_, _39695_, _27209_);
  nor (_39697_, _27198_, _39693_);
  or (_39698_, _39697_, rst);
  or (_39701_, _39698_, _39696_);
  or (_41319_, _39701_, _39691_);
  nand (_39709_, _27790_, _24376_);
  or (_39710_, _24376_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39711_, _39710_, _39399_);
  and (_39712_, _39711_, _39709_);
  not (_39713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39714_, _39399_, _39713_);
  or (_39715_, _39714_, _39712_);
  and (_39716_, _39715_, _27900_);
  nor (_39717_, _39408_, _38066_);
  nor (_39718_, _39407_, _39713_);
  or (_39719_, _39718_, _39717_);
  and (_39720_, _39719_, _27209_);
  nor (_39721_, _27198_, _39713_);
  or (_39722_, _39721_, rst);
  or (_39723_, _39722_, _39720_);
  or (_41321_, _39723_, _39716_);
  nand (_39724_, _29174_, _27790_);
  or (_39725_, _29174_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39726_, _39725_, _39399_);
  and (_39727_, _39726_, _39724_);
  not (_39728_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_39729_, _39399_, _39728_);
  or (_39730_, _39729_, _39727_);
  and (_39731_, _39730_, _27900_);
  nor (_39732_, _39408_, _37978_);
  nor (_39733_, _39407_, _39728_);
  or (_39734_, _39733_, _39732_);
  and (_39735_, _39734_, _27209_);
  nor (_39736_, _27198_, _39728_);
  or (_39737_, _39736_, rst);
  or (_39738_, _39737_, _39735_);
  or (_41323_, _39738_, _39731_);
  not (_39739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_39740_, _29916_, _39739_);
  or (_39741_, _39740_, _29927_);
  and (_39742_, _39741_, _39399_);
  nor (_39743_, _39399_, _39739_);
  or (_39744_, _39743_, _39742_);
  and (_39745_, _39744_, _27900_);
  nor (_39746_, _39408_, _37901_);
  nor (_39747_, _39407_, _39739_);
  or (_39748_, _39747_, _39746_);
  and (_39749_, _39748_, _27209_);
  nor (_39750_, _27198_, _39739_);
  or (_39751_, _39750_, rst);
  or (_39752_, _39751_, _39749_);
  or (_41325_, _39752_, _39745_);
  and (_39753_, _30623_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39754_, _39753_, _30634_);
  and (_39755_, _39754_, _39399_);
  not (_39756_, _39399_);
  and (_39757_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39758_, _39757_, _39755_);
  and (_39759_, _39758_, _27900_);
  nor (_39760_, _39408_, _37824_);
  and (_39761_, _39408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39762_, _39761_, _39760_);
  and (_39763_, _39762_, _27209_);
  and (_39764_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39765_, _39764_, rst);
  or (_39766_, _39765_, _39763_);
  or (_41327_, _39766_, _39759_);
  and (_39767_, _31449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39768_, _39767_, _31459_);
  and (_39769_, _39768_, _39399_);
  and (_39770_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39771_, _39770_, _39769_);
  and (_39772_, _39771_, _27900_);
  nor (_39773_, _39408_, _37736_);
  and (_39774_, _39408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39775_, _39774_, _39773_);
  and (_39776_, _39775_, _27209_);
  and (_39777_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39778_, _39777_, rst);
  or (_39779_, _39778_, _39776_);
  or (_41328_, _39779_, _39772_);
  and (_39780_, _32254_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39781_, _39780_, _32265_);
  and (_39782_, _39781_, _39399_);
  and (_39783_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39784_, _39783_, _39782_);
  and (_39785_, _39784_, _27900_);
  nor (_39786_, _39408_, _37650_);
  and (_39787_, _39408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39788_, _39787_, _39786_);
  and (_39789_, _39788_, _27209_);
  and (_39790_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39791_, _39790_, rst);
  or (_39792_, _39791_, _39789_);
  or (_41330_, _39792_, _39785_);
  not (_39793_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_39794_, _33039_, _39793_);
  or (_39795_, _39794_, _33050_);
  and (_39796_, _39795_, _39399_);
  nor (_39797_, _39399_, _39793_);
  or (_39798_, _39797_, _39796_);
  and (_39799_, _39798_, _27900_);
  nor (_39800_, _39408_, _37564_);
  nor (_39801_, _39407_, _39793_);
  or (_39802_, _39801_, _39800_);
  and (_39803_, _39802_, _27209_);
  nor (_39804_, _27198_, _39793_);
  or (_39805_, _39804_, rst);
  or (_39806_, _39805_, _39803_);
  or (_41332_, _39806_, _39799_);
  and (_39807_, _36503_, _36144_);
  and (_39808_, _36688_, _35161_);
  nor (_39809_, _39808_, _36764_);
  and (_39810_, _35937_, _36720_);
  nor (_39811_, _39810_, _36350_);
  and (_39812_, _39811_, _36920_);
  and (_39813_, _39812_, _39809_);
  not (_39814_, _36231_);
  and (_39815_, _36753_, _39814_);
  and (_39816_, _39815_, _36514_);
  and (_39817_, _39816_, _39813_);
  nor (_39818_, _39817_, _33169_);
  nor (_39819_, _39818_, _39807_);
  not (_39820_, _39819_);
  and (_39821_, _37326_, _37157_);
  not (_39822_, _38401_);
  and (_39823_, _39822_, _39821_);
  not (_39824_, _39823_);
  and (_39825_, _37326_, _36209_);
  and (_39826_, _39825_, _37146_);
  and (_39827_, _39826_, _35796_);
  not (_39828_, _36209_);
  and (_39829_, _37146_, _39828_);
  and (_39830_, _39829_, _37326_);
  nor (_39831_, _35785_, _24085_);
  and (_39832_, _35785_, _24085_);
  nor (_39833_, _39832_, _39831_);
  and (_39834_, _27176_, _23296_);
  not (_39835_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_39836_, _24364_, _39835_);
  and (_39837_, _39836_, _39834_);
  not (_39838_, _39837_);
  nor (_39839_, _39838_, _39833_);
  nor (_39840_, _38951_, _39001_);
  nor (_39841_, _39840_, _39007_);
  nor (_39842_, _39841_, _23647_);
  and (_39843_, _39841_, _23647_);
  nor (_39844_, _39843_, _39842_);
  and (_39845_, _39844_, _39839_);
  nor (_39846_, _39841_, _35785_);
  and (_39847_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_39848_, _39841_, _35796_);
  and (_39849_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_39850_, _39849_, _39847_);
  and (_39851_, _39841_, _35785_);
  and (_39852_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_39853_, _39841_, _35796_);
  and (_39854_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_39855_, _39854_, _39852_);
  and (_39856_, _39855_, _39850_);
  nor (_39857_, _39856_, _39845_);
  and (_39858_, _39845_, _38077_);
  nor (_39859_, _39858_, _39857_);
  not (_39860_, _39859_);
  and (_39861_, _39860_, _39830_);
  nor (_39862_, _37146_, _39828_);
  and (_39863_, _39862_, _37326_);
  not (_39864_, _33213_);
  and (_39865_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_39866_, _33682_, _33213_);
  not (_39867_, _39866_);
  and (_39868_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_39869_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_39870_, _39869_, _39868_);
  and (_39871_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_39872_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_39873_, _39872_, _39871_);
  and (_39874_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_39875_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_39876_, _39875_, _39874_);
  and (_39877_, _39876_, _39873_);
  and (_39878_, _39877_, _39870_);
  nor (_39879_, _39878_, _39867_);
  nor (_39880_, _39879_, _39865_);
  not (_39881_, _39880_);
  and (_39882_, _39881_, _39863_);
  or (_39883_, _39882_, _39861_);
  nor (_39884_, _39883_, _39827_);
  and (_39885_, _39884_, _39824_);
  nor (_39886_, _39885_, _39820_);
  and (_39887_, _36470_, _35937_);
  nor (_39888_, _37058_, _39887_);
  nor (_39889_, _39888_, _37014_);
  not (_39890_, _36905_);
  and (_39891_, _35313_, _37025_);
  and (_39892_, _39891_, _35937_);
  nor (_39893_, _39892_, _36764_);
  and (_39894_, _39893_, _39890_);
  and (_39895_, _39894_, _39814_);
  and (_39896_, _39891_, _35959_);
  not (_39897_, _39896_);
  and (_39898_, _39897_, _39888_);
  not (_39899_, _37047_);
  and (_39900_, _35379_, _35324_);
  and (_39901_, _39900_, _35959_);
  nor (_39902_, _39901_, _36731_);
  and (_39903_, _39902_, _39899_);
  and (_39904_, _39903_, _39898_);
  and (_39905_, _39904_, _39895_);
  and (_39906_, _39905_, _39811_);
  nor (_39907_, _39906_, _33169_);
  nor (_39908_, _39907_, _39889_);
  not (_39909_, _38306_);
  and (_39910_, _39909_, _39821_);
  not (_39911_, _39910_);
  and (_39912_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_39913_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_39914_, _39913_, _39912_);
  and (_39915_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_39916_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_39917_, _39916_, _39915_);
  and (_39918_, _39917_, _39914_);
  nor (_39919_, _39918_, _39845_);
  not (_39920_, _38285_);
  and (_39921_, _39845_, _39920_);
  nor (_39922_, _39921_, _39919_);
  not (_39923_, _39922_);
  and (_39924_, _39923_, _39829_);
  not (_39925_, _39924_);
  not (_39926_, _37326_);
  and (_39927_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_39928_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_39929_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_39930_, _39929_, _39928_);
  and (_39931_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_39932_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_39933_, _39932_, _39931_);
  and (_39934_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_39935_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_39936_, _39935_, _39934_);
  and (_39937_, _39936_, _39933_);
  and (_39938_, _39937_, _39930_);
  nor (_39939_, _39938_, _39867_);
  nor (_39940_, _39939_, _39927_);
  not (_39941_, _39940_);
  and (_39942_, _39941_, _39862_);
  nor (_39943_, _39942_, _39926_);
  and (_39944_, _39943_, _39925_);
  and (_39945_, _39944_, _39911_);
  not (_39946_, _39945_);
  nor (_39947_, _39946_, _39908_);
  not (_39948_, _37824_);
  and (_39949_, _39845_, _39948_);
  and (_39950_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_39951_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_39952_, _39951_, _39950_);
  and (_39953_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_39954_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_39955_, _39954_, _39953_);
  and (_39956_, _39955_, _39952_);
  nor (_39957_, _39956_, _39845_);
  nor (_39958_, _39957_, _39949_);
  not (_39959_, _39958_);
  and (_39960_, _39959_, _39830_);
  and (_39961_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_39962_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_39963_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_39964_, _39963_, _39962_);
  and (_39965_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_39966_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_39967_, _39966_, _39965_);
  and (_39968_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_39969_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_39970_, _39969_, _39968_);
  and (_39971_, _39970_, _39967_);
  and (_39972_, _39971_, _39964_);
  nor (_39973_, _39972_, _39867_);
  nor (_39974_, _39973_, _39961_);
  not (_39975_, _39974_);
  and (_39976_, _39975_, _39863_);
  nor (_39977_, _39976_, _39960_);
  not (_39978_, _38476_);
  and (_39979_, _39978_, _39821_);
  not (_39980_, _39841_);
  and (_39981_, _39826_, _39980_);
  nor (_39982_, _39981_, _39979_);
  and (_39983_, _39982_, _39977_);
  not (_39984_, _39983_);
  and (_39985_, _39984_, _39947_);
  nor (_39986_, _39985_, _39886_);
  and (_39987_, _23317_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_39988_, _39987_, _23647_);
  nor (_39989_, _24085_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_39990_, _39989_, _39988_);
  not (_39991_, _39990_);
  nor (_39992_, _39991_, _39986_);
  and (_39993_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_39994_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_39995_, _39994_, _39993_);
  and (_39996_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_39997_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_39998_, _39997_, _39996_);
  and (_39999_, _39998_, _39995_);
  nor (_40000_, _39999_, _39845_);
  not (_40001_, _37901_);
  and (_40002_, _39845_, _40001_);
  nor (_40003_, _40002_, _40000_);
  not (_40004_, _40003_);
  and (_40005_, _40004_, _39830_);
  not (_40006_, _40005_);
  and (_40007_, _39826_, _36242_);
  not (_40008_, _38470_);
  and (_40009_, _40008_, _39821_);
  and (_40010_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40011_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_40012_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40013_, _40012_, _40011_);
  and (_40014_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_40015_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_40016_, _40015_, _40014_);
  and (_40017_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40018_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_40019_, _40018_, _40017_);
  and (_40020_, _40019_, _40016_);
  and (_40021_, _40020_, _40013_);
  nor (_40022_, _40021_, _39867_);
  nor (_40023_, _40022_, _40010_);
  not (_40024_, _40023_);
  and (_40025_, _40024_, _39863_);
  or (_40026_, _40025_, _40009_);
  nor (_40027_, _40026_, _40007_);
  and (_40028_, _40027_, _40006_);
  nor (_40029_, _40028_, _39820_);
  and (_40030_, _39926_, _36209_);
  and (_40031_, _40030_, _37146_);
  not (_40032_, _40031_);
  not (_40033_, _37650_);
  and (_40034_, _39845_, _40033_);
  and (_40035_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_40036_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40037_, _40036_, _40035_);
  and (_40038_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_40039_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_40040_, _40039_, _40038_);
  and (_40041_, _40040_, _40037_);
  nor (_40042_, _40041_, _39845_);
  nor (_40043_, _40042_, _40034_);
  not (_40044_, _40043_);
  and (_40045_, _40044_, _39830_);
  and (_40046_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40047_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40048_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40049_, _40048_, _40047_);
  and (_40050_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40051_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40052_, _40051_, _40050_);
  and (_40053_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_40054_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_40055_, _40054_, _40053_);
  and (_40056_, _40055_, _40052_);
  and (_40057_, _40056_, _40049_);
  nor (_40058_, _40057_, _39867_);
  nor (_40059_, _40058_, _40046_);
  not (_40060_, _40059_);
  and (_40061_, _40060_, _39863_);
  nor (_40062_, _40061_, _40045_);
  and (_40063_, _40062_, _40032_);
  and (_40064_, _39926_, _37157_);
  not (_40065_, _38488_);
  and (_40066_, _40065_, _39821_);
  nor (_40067_, _40066_, _40064_);
  and (_40068_, _40067_, _40063_);
  not (_40069_, _40068_);
  and (_40070_, _39947_, _40069_);
  nor (_40071_, _40070_, _40029_);
  and (_40072_, _39987_, _23965_);
  nor (_40073_, _24352_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40074_, _40073_, _40072_);
  not (_40075_, _40074_);
  and (_40076_, _40075_, _40071_);
  nor (_40077_, _40076_, _39992_);
  not (_40078_, _39834_);
  and (_40079_, _39991_, _39986_);
  nor (_40080_, _40079_, _40078_);
  and (_40081_, _40080_, _40077_);
  and (_40082_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40083_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_40084_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_40085_, _40084_, _40083_);
  and (_40086_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40087_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40088_, _40087_, _40086_);
  and (_40089_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40090_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_40091_, _40090_, _40089_);
  and (_40092_, _40091_, _40088_);
  and (_40093_, _40092_, _40085_);
  nor (_40094_, _40093_, _39867_);
  nor (_40095_, _40094_, _40082_);
  not (_40096_, _40095_);
  and (_40097_, _40096_, _39863_);
  not (_40098_, _40097_);
  and (_40099_, _39829_, _39926_);
  and (_40100_, _39826_, _35807_);
  nor (_40101_, _40100_, _40099_);
  and (_40102_, _40101_, _40098_);
  not (_40103_, _38464_);
  and (_40104_, _40103_, _39821_);
  and (_40105_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_40106_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_40107_, _40106_, _40105_);
  and (_40108_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_40109_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40110_, _40109_, _40108_);
  and (_40111_, _40110_, _40107_);
  nor (_40112_, _40111_, _39845_);
  not (_40113_, _37978_);
  and (_40114_, _39845_, _40113_);
  nor (_40115_, _40114_, _40112_);
  not (_40116_, _40115_);
  and (_40117_, _40116_, _39830_);
  nor (_40118_, _40117_, _40104_);
  and (_40119_, _40118_, _40102_);
  nor (_40120_, _40119_, _39820_);
  and (_40121_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_40122_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_40123_, _40122_, _40121_);
  and (_40124_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_40125_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_40126_, _40125_, _40124_);
  nor (_40127_, _40126_, _40123_);
  nor (_40128_, _40127_, _39845_);
  not (_40129_, _37736_);
  and (_40130_, _39845_, _40129_);
  or (_40131_, _40130_, _40128_);
  and (_40132_, _40131_, _39830_);
  not (_40133_, _38482_);
  and (_40134_, _40133_, _39821_);
  or (_40135_, _40134_, _40030_);
  and (_40136_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40137_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_40138_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_40139_, _40138_, _40137_);
  and (_40140_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40141_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40142_, _40141_, _40140_);
  and (_40143_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40144_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_40145_, _40144_, _40143_);
  and (_40146_, _40145_, _40142_);
  and (_40147_, _40146_, _40139_);
  nor (_40148_, _40147_, _39867_);
  nor (_40149_, _40148_, _40136_);
  not (_40150_, _40149_);
  and (_40151_, _40150_, _39863_);
  not (_40152_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_40153_, _38951_, _40152_);
  or (_40154_, _40153_, _39017_);
  and (_40155_, _40154_, _39826_);
  or (_40156_, _40155_, _40151_);
  or (_40157_, _40156_, _40135_);
  or (_40158_, _40157_, _40132_);
  and (_40159_, _40158_, _39947_);
  nor (_40160_, _40159_, _40120_);
  and (_40161_, _39987_, _37369_);
  nor (_40162_, _24217_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40163_, _40162_, _40161_);
  nand (_40164_, _40163_, _40160_);
  or (_40165_, _40163_, _40160_);
  and (_40166_, _40165_, _40164_);
  not (_40167_, _40166_);
  nor (_40168_, _40075_, _40071_);
  not (_40169_, _40168_);
  and (_40170_, _39945_, _39820_);
  nor (_40171_, _39984_, _40170_);
  not (_40172_, _38494_);
  and (_40173_, _40172_, _39821_);
  not (_40174_, _40173_);
  and (_40175_, _39846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_40176_, _39848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_40177_, _40176_, _40175_);
  and (_40178_, _39851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_40179_, _39853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_40180_, _40179_, _40178_);
  and (_40181_, _40180_, _40177_);
  nor (_40182_, _40181_, _39845_);
  not (_40183_, _37564_);
  and (_40184_, _39845_, _40183_);
  nor (_40185_, _40184_, _40182_);
  not (_40186_, _40185_);
  and (_40187_, _40186_, _39830_);
  and (_40188_, _39864_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40189_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_40190_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_40191_, _40190_, _40189_);
  and (_40192_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_40193_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40194_, _40193_, _40192_);
  and (_40195_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40196_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_40197_, _40196_, _40195_);
  and (_40198_, _40197_, _40194_);
  and (_40199_, _40198_, _40191_);
  nor (_40200_, _40199_, _39867_);
  nor (_40201_, _40200_, _40188_);
  not (_40202_, _40201_);
  and (_40203_, _40202_, _39862_);
  or (_40204_, _40203_, _40030_);
  or (_40205_, _40204_, _40187_);
  nor (_40206_, _40205_, _40064_);
  and (_40207_, _40206_, _40174_);
  and (_40208_, _40207_, _40170_);
  nor (_40209_, _40208_, _40171_);
  nor (_40210_, _39987_, _23647_);
  and (_40211_, _39987_, _23449_);
  nor (_40212_, _40211_, _40210_);
  not (_40213_, _40212_);
  and (_40214_, _40213_, _40209_);
  nor (_40215_, _40213_, _40209_);
  nor (_40216_, _40215_, _40214_);
  and (_40217_, _40216_, _40169_);
  and (_40218_, _40217_, _40167_);
  and (_40219_, _40218_, _40081_);
  not (_40220_, _40071_);
  and (_40221_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40222_, _39986_);
  and (_40223_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_40224_, _40223_, _40221_);
  and (_40225_, _40224_, _40160_);
  not (_40226_, _40160_);
  not (_40227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40228_, _39986_, _40227_);
  and (_40229_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40230_, _40229_, _40228_);
  and (_40231_, _40230_, _40226_);
  or (_40232_, _40231_, _40225_);
  or (_40233_, _40232_, _40220_);
  not (_40234_, _40209_);
  and (_40235_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_40236_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_40237_, _40236_, _40235_);
  and (_40238_, _40237_, _40160_);
  not (_40239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40240_, _39986_, _40239_);
  and (_40241_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40242_, _40241_, _40240_);
  and (_40243_, _40242_, _40226_);
  or (_40244_, _40243_, _40238_);
  or (_40245_, _40244_, _40071_);
  and (_40246_, _40245_, _40234_);
  and (_40247_, _40246_, _40233_);
  or (_40248_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_40249_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40250_, _40249_, _40248_);
  and (_40251_, _40250_, _40160_);
  or (_40252_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_40254_, _39986_, _40253_);
  and (_40255_, _40254_, _40252_);
  and (_40256_, _40255_, _40226_);
  or (_40257_, _40256_, _40251_);
  or (_40258_, _40257_, _40220_);
  or (_40259_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_40260_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_40261_, _40260_, _40259_);
  and (_40262_, _40261_, _40160_);
  or (_40263_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_40264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_40265_, _39986_, _40264_);
  and (_40266_, _40265_, _40263_);
  and (_40267_, _40266_, _40226_);
  or (_40268_, _40267_, _40262_);
  or (_40269_, _40268_, _40071_);
  and (_40270_, _40269_, _40209_);
  and (_40271_, _40270_, _40258_);
  or (_40272_, _40271_, _40247_);
  or (_40273_, _40272_, _40219_);
  not (_40274_, _40219_);
  or (_40275_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_40276_, _40275_, _43998_);
  and (_41408_, _40276_, _40273_);
  nor (_40277_, _39990_, _40078_);
  nor (_40278_, _40163_, _40078_);
  and (_40279_, _40278_, _40277_);
  and (_40280_, _40212_, _39834_);
  nor (_40281_, _40074_, _40078_);
  and (_40282_, _40281_, _40280_);
  and (_40283_, _40282_, _40279_);
  and (_40284_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_40285_, _40284_, _25124_);
  nor (_40286_, _40285_, _27790_);
  nand (_40287_, _25124_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40288_, _16526_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40289_, _40288_, _40287_);
  nor (_40290_, _38285_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40291_, _40290_, _40289_);
  or (_40292_, _40291_, _40286_);
  and (_40293_, _40292_, _39834_);
  and (_40294_, _40293_, _40283_);
  not (_40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_40296_, _40283_, _40295_);
  or (_41418_, _40296_, _40294_);
  nor (_40297_, _40281_, _40280_);
  nor (_40298_, _40278_, _40277_);
  and (_40299_, _40298_, _39834_);
  and (_40300_, _40299_, _40297_);
  and (_40301_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25114_);
  and (_40302_, _40301_, _25157_);
  not (_40303_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40304_, _38066_, _40303_);
  or (_40305_, _15363_, _40303_);
  and (_40306_, _40305_, _40304_);
  or (_40307_, _40306_, _40302_);
  nand (_40308_, _40302_, _27790_);
  and (_40309_, _40308_, _40307_);
  and (_40310_, _40309_, _40300_);
  not (_40311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40312_, _40300_, _40311_);
  or (_41661_, _40312_, _40310_);
  nand (_40313_, _40301_, _25201_);
  nor (_40314_, _40313_, _27790_);
  nor (_40315_, _37978_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40316_, _40301_, _25223_);
  and (_40317_, _40301_, _25124_);
  or (_40318_, _40317_, _40284_);
  or (_40319_, _40318_, _40316_);
  and (_40320_, _40319_, _16350_);
  or (_40321_, _40320_, _40315_);
  or (_40322_, _40321_, _40314_);
  and (_40323_, _40322_, _40300_);
  not (_40324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40325_, _40300_, _40324_);
  or (_41666_, _40325_, _40323_);
  not (_40326_, _40300_);
  and (_40327_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_40328_, _40301_, _25244_);
  nor (_40329_, _40328_, _27790_);
  nor (_40330_, _37901_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40331_, _40301_, _25190_);
  or (_40332_, _40331_, _40318_);
  and (_40333_, _40332_, _15001_);
  or (_40334_, _40333_, _40330_);
  or (_40335_, _40334_, _40329_);
  and (_40336_, _40335_, _40300_);
  or (_41671_, _40336_, _40327_);
  and (_40337_, _40317_, _28460_);
  nor (_40338_, _37824_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40339_, _40316_, _40284_);
  or (_40340_, _40339_, _40331_);
  and (_40341_, _40340_, _16032_);
  or (_40342_, _40341_, _40338_);
  or (_40343_, _40342_, _40337_);
  and (_40344_, _40343_, _40300_);
  and (_40345_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_41676_, _40345_, _40344_);
  nand (_40346_, _40284_, _25157_);
  nor (_40347_, _40346_, _27790_);
  nor (_40348_, _37736_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40349_, _25157_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40350_, _15199_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40351_, _40350_, _40349_);
  or (_40352_, _40351_, _40348_);
  or (_40353_, _40352_, _40347_);
  and (_40354_, _40353_, _40300_);
  and (_40355_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_41681_, _40355_, _40354_);
  nand (_40356_, _40284_, _25201_);
  nor (_40357_, _40356_, _27790_);
  nor (_40358_, _37650_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40359_, _25201_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40360_, _16186_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40361_, _40360_, _40359_);
  or (_40362_, _40361_, _40358_);
  or (_40363_, _40362_, _40357_);
  and (_40364_, _40363_, _40300_);
  and (_40365_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_41686_, _40365_, _40364_);
  nand (_40366_, _40284_, _25244_);
  nor (_40367_, _40366_, _27790_);
  nor (_40368_, _37564_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40369_, _25244_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40370_, _15539_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40371_, _40370_, _40369_);
  or (_40372_, _40371_, _40368_);
  or (_40373_, _40372_, _40367_);
  and (_40374_, _40373_, _40300_);
  and (_40375_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_41692_, _40375_, _40374_);
  and (_40376_, _40300_, _40292_);
  and (_40377_, _40326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_41694_, _40377_, _40376_);
  and (_40378_, _40309_, _39834_);
  and (_40379_, _40277_, _40163_);
  and (_40380_, _40379_, _40297_);
  and (_40381_, _40380_, _40378_);
  not (_40382_, _40380_);
  and (_40383_, _40382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_41701_, _40383_, _40381_);
  and (_40384_, _40322_, _39834_);
  and (_40385_, _40380_, _40384_);
  and (_40386_, _40382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_41705_, _40386_, _40385_);
  and (_40387_, _40335_, _39834_);
  and (_40388_, _40380_, _40387_);
  and (_40389_, _40382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_41708_, _40389_, _40388_);
  and (_40390_, _40343_, _39834_);
  and (_40391_, _40380_, _40390_);
  not (_40392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_40393_, _40380_, _40392_);
  or (_41712_, _40393_, _40391_);
  and (_40394_, _40353_, _39834_);
  and (_40395_, _40380_, _40394_);
  not (_40396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_40397_, _40380_, _40396_);
  or (_41715_, _40397_, _40395_);
  and (_40398_, _40363_, _39834_);
  and (_40399_, _40380_, _40398_);
  not (_40400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40401_, _40380_, _40400_);
  or (_41719_, _40401_, _40399_);
  and (_40402_, _40373_, _39834_);
  and (_40403_, _40380_, _40402_);
  not (_40404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_40405_, _40380_, _40404_);
  or (_41722_, _40405_, _40403_);
  and (_40406_, _40380_, _40293_);
  and (_40407_, _40382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_41725_, _40407_, _40406_);
  and (_40408_, _40278_, _39990_);
  and (_40409_, _40408_, _40297_);
  and (_40410_, _40409_, _40378_);
  not (_40411_, _40409_);
  and (_40412_, _40411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41732_, _40412_, _40410_);
  and (_40413_, _40409_, _40384_);
  and (_40414_, _40411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41735_, _40414_, _40413_);
  and (_40415_, _40409_, _40387_);
  not (_40416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_40417_, _40409_, _40416_);
  or (_41739_, _40417_, _40415_);
  and (_40418_, _40409_, _40390_);
  and (_40419_, _40411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41742_, _40419_, _40418_);
  and (_40420_, _40409_, _40394_);
  not (_40421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_40422_, _40409_, _40421_);
  or (_41746_, _40422_, _40420_);
  and (_40423_, _40409_, _40398_);
  not (_40424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_40425_, _40409_, _40424_);
  or (_41749_, _40425_, _40423_);
  and (_40426_, _40409_, _40402_);
  not (_40427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_40428_, _40409_, _40427_);
  or (_41753_, _40428_, _40426_);
  and (_40429_, _40409_, _40293_);
  not (_40430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_40431_, _40409_, _40430_);
  or (_41756_, _40431_, _40429_);
  and (_40432_, _40297_, _40279_);
  and (_40433_, _40432_, _40378_);
  not (_40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_40435_, _40432_, _40434_);
  or (_41761_, _40435_, _40433_);
  and (_40436_, _40432_, _40384_);
  not (_40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_40438_, _40432_, _40437_);
  or (_41764_, _40438_, _40436_);
  and (_40439_, _40432_, _40387_);
  not (_40440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_40441_, _40432_, _40440_);
  or (_41768_, _40441_, _40439_);
  and (_40442_, _40432_, _40390_);
  not (_40443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_40444_, _40432_, _40443_);
  or (_41771_, _40444_, _40442_);
  and (_40445_, _40432_, _40394_);
  not (_40446_, _40432_);
  and (_40447_, _40446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_41775_, _40447_, _40445_);
  and (_40448_, _40432_, _40398_);
  and (_40449_, _40446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_41778_, _40449_, _40448_);
  and (_40450_, _40432_, _40402_);
  and (_40451_, _40446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_41782_, _40451_, _40450_);
  and (_40452_, _40432_, _40293_);
  nor (_40453_, _40432_, _40227_);
  or (_41784_, _40453_, _40452_);
  and (_40454_, _40281_, _40213_);
  and (_40455_, _40454_, _40298_);
  and (_40456_, _40455_, _40378_);
  not (_40457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_40458_, _40455_, _40457_);
  or (_41791_, _40458_, _40456_);
  and (_40459_, _40455_, _40384_);
  not (_40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_40461_, _40455_, _40460_);
  or (_41795_, _40461_, _40459_);
  and (_40462_, _40455_, _40387_);
  not (_40463_, _40455_);
  and (_40464_, _40463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_41798_, _40464_, _40462_);
  and (_40465_, _40455_, _40390_);
  not (_40466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_40467_, _40455_, _40466_);
  or (_41802_, _40467_, _40465_);
  and (_40468_, _40455_, _40394_);
  and (_40469_, _40463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_41805_, _40469_, _40468_);
  and (_40470_, _40455_, _40398_);
  and (_40471_, _40463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_41809_, _40471_, _40470_);
  and (_40472_, _40455_, _40402_);
  not (_40473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_40474_, _40455_, _40473_);
  or (_41812_, _40474_, _40472_);
  and (_40475_, _40455_, _40293_);
  and (_40476_, _40463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_41815_, _40476_, _40475_);
  and (_40477_, _40454_, _40379_);
  and (_40478_, _40477_, _40378_);
  not (_40479_, _40477_);
  and (_40480_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_41819_, _40480_, _40478_);
  and (_40481_, _40477_, _40384_);
  and (_40482_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_41823_, _40482_, _40481_);
  and (_40483_, _40477_, _40387_);
  and (_40485_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_41826_, _40485_, _40483_);
  and (_40496_, _40477_, _40390_);
  and (_40502_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_41830_, _40502_, _40496_);
  and (_40513_, _40477_, _40394_);
  not (_40515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_40516_, _40477_, _40515_);
  or (_41833_, _40516_, _40513_);
  and (_40517_, _40477_, _40398_);
  not (_40518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_40519_, _40477_, _40518_);
  or (_41837_, _40519_, _40517_);
  and (_40520_, _40477_, _40402_);
  and (_40521_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_41840_, _40521_, _40520_);
  and (_40522_, _40477_, _40293_);
  and (_40523_, _40479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_41843_, _40523_, _40522_);
  and (_40524_, _40454_, _40408_);
  and (_40525_, _40524_, _40378_);
  not (_40526_, _40524_);
  and (_40527_, _40526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41847_, _40527_, _40525_);
  and (_40528_, _40524_, _40384_);
  and (_40529_, _40526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41851_, _40529_, _40528_);
  and (_40530_, _40524_, _40387_);
  not (_40531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_40532_, _40524_, _40531_);
  or (_41854_, _40532_, _40530_);
  and (_40533_, _40524_, _40390_);
  and (_40534_, _40526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41858_, _40534_, _40533_);
  and (_40535_, _40524_, _40394_);
  not (_40536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_40537_, _40524_, _40536_);
  or (_41862_, _40537_, _40535_);
  and (_40538_, _40524_, _40398_);
  not (_40539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_40540_, _40524_, _40539_);
  or (_41865_, _40540_, _40538_);
  and (_40541_, _40524_, _40402_);
  and (_40544_, _40526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41869_, _40544_, _40541_);
  and (_40551_, _40524_, _40293_);
  not (_40552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_40553_, _40524_, _40552_);
  or (_41871_, _40553_, _40551_);
  and (_40558_, _40454_, _40279_);
  and (_40563_, _40558_, _40378_);
  not (_40564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_40565_, _40558_, _40564_);
  or (_41876_, _40565_, _40563_);
  and (_40572_, _40558_, _40384_);
  not (_40575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_40576_, _40558_, _40575_);
  or (_41879_, _40576_, _40572_);
  and (_40581_, _40558_, _40387_);
  not (_40586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_40587_, _40558_, _40586_);
  or (_41883_, _40587_, _40581_);
  and (_40589_, _40558_, _40390_);
  not (_40595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_40598_, _40558_, _40595_);
  or (_41886_, _40598_, _40589_);
  and (_40599_, _40558_, _40394_);
  not (_40605_, _40558_);
  and (_40609_, _40605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_41890_, _40609_, _40599_);
  and (_40610_, _40558_, _40398_);
  and (_40616_, _40605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_41893_, _40616_, _40610_);
  and (_40620_, _40558_, _40402_);
  not (_40621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_40626_, _40558_, _40621_);
  or (_41897_, _40626_, _40620_);
  and (_40631_, _40558_, _40293_);
  nor (_40632_, _40558_, _40239_);
  or (_41899_, _40632_, _40631_);
  and (_40639_, _40280_, _40074_);
  and (_40642_, _40639_, _40298_);
  and (_40643_, _40642_, _40378_);
  not (_40644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_40650_, _40642_, _40644_);
  or (_41906_, _40650_, _40643_);
  and (_40654_, _40642_, _40384_);
  not (_40655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_40661_, _40642_, _40655_);
  or (_41910_, _40661_, _40654_);
  and (_40665_, _40642_, _40387_);
  not (_40666_, _40642_);
  and (_40671_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_41913_, _40671_, _40665_);
  and (_40676_, _40642_, _40390_);
  and (_40677_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_41917_, _40677_, _40676_);
  and (_40686_, _40642_, _40394_);
  and (_40687_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_41920_, _40687_, _40686_);
  and (_40690_, _40642_, _40398_);
  and (_40696_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_41924_, _40696_, _40690_);
  and (_40698_, _40642_, _40402_);
  and (_40701_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_41927_, _40701_, _40698_);
  and (_40708_, _40642_, _40293_);
  and (_40709_, _40666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_41930_, _40709_, _40708_);
  and (_40717_, _40639_, _40379_);
  and (_40718_, _40717_, _40378_);
  not (_40719_, _40717_);
  and (_40720_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_41934_, _40720_, _40718_);
  and (_40721_, _40717_, _40384_);
  and (_40722_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_41938_, _40722_, _40721_);
  and (_40723_, _40717_, _40387_);
  and (_40724_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_41941_, _40724_, _40723_);
  and (_40725_, _40717_, _40390_);
  and (_40726_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_41945_, _40726_, _40725_);
  and (_40727_, _40717_, _40394_);
  not (_40728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_40729_, _40717_, _40728_);
  or (_41948_, _40729_, _40727_);
  and (_40730_, _40717_, _40398_);
  not (_40731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_40732_, _40717_, _40731_);
  or (_41952_, _40732_, _40730_);
  and (_40733_, _40717_, _40402_);
  and (_40734_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_41955_, _40734_, _40733_);
  and (_40735_, _40717_, _40293_);
  and (_40736_, _40719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_41958_, _40736_, _40735_);
  and (_40737_, _40639_, _40408_);
  and (_40738_, _40737_, _40378_);
  not (_40739_, _40737_);
  and (_40740_, _40739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_41962_, _40740_, _40738_);
  and (_40741_, _40737_, _40384_);
  and (_40742_, _40739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_41966_, _40742_, _40741_);
  and (_40743_, _40737_, _40387_);
  not (_40744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_40745_, _40737_, _40744_);
  or (_41968_, _40745_, _40743_);
  and (_40746_, _40737_, _40390_);
  not (_40747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_40748_, _40737_, _40747_);
  or (_41972_, _40748_, _40746_);
  and (_40749_, _40737_, _40394_);
  not (_40750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_40751_, _40737_, _40750_);
  or (_41975_, _40751_, _40749_);
  and (_40752_, _40737_, _40398_);
  not (_40753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_40754_, _40737_, _40753_);
  or (_41979_, _40754_, _40752_);
  and (_40755_, _40737_, _40402_);
  and (_40756_, _40739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_41983_, _40756_, _40755_);
  and (_40757_, _40737_, _40293_);
  nor (_40758_, _40737_, _40253_);
  or (_41986_, _40758_, _40757_);
  and (_40759_, _40639_, _40279_);
  and (_40760_, _40759_, _40378_);
  not (_40761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_40762_, _40759_, _40761_);
  or (_41991_, _40762_, _40760_);
  and (_40763_, _40759_, _40384_);
  not (_40764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_40765_, _40759_, _40764_);
  or (_41995_, _40765_, _40763_);
  and (_40766_, _40759_, _40387_);
  not (_40767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_40768_, _40759_, _40767_);
  or (_41999_, _40768_, _40766_);
  and (_40769_, _40759_, _40390_);
  not (_40770_, _40759_);
  and (_40771_, _40770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_42003_, _40771_, _40769_);
  and (_40772_, _40759_, _40394_);
  and (_40773_, _40770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_42007_, _40773_, _40772_);
  and (_40774_, _40759_, _40398_);
  and (_40775_, _40770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_42011_, _40775_, _40774_);
  and (_40776_, _40759_, _40402_);
  and (_40777_, _40770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_42015_, _40777_, _40776_);
  and (_40778_, _40759_, _40293_);
  not (_40779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_40780_, _40759_, _40779_);
  or (_42018_, _40780_, _40778_);
  and (_40781_, _40298_, _40282_);
  and (_40782_, _40781_, _40378_);
  not (_40783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_40784_, _40781_, _40783_);
  or (_42024_, _40784_, _40782_);
  and (_40785_, _40781_, _40384_);
  not (_40786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_40787_, _40781_, _40786_);
  or (_42028_, _40787_, _40785_);
  and (_40788_, _40781_, _40387_);
  not (_40789_, _40781_);
  and (_40790_, _40789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_42032_, _40790_, _40788_);
  and (_40791_, _40781_, _40390_);
  not (_40792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_40793_, _40781_, _40792_);
  or (_42036_, _40793_, _40791_);
  and (_40794_, _40781_, _40394_);
  and (_40795_, _40789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_42040_, _40795_, _40794_);
  and (_40796_, _40781_, _40398_);
  and (_40797_, _40789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_42044_, _40797_, _40796_);
  and (_40798_, _40781_, _40402_);
  not (_40799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_40800_, _40781_, _40799_);
  or (_42048_, _40800_, _40798_);
  and (_40801_, _40781_, _40293_);
  and (_40802_, _40789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_42051_, _40802_, _40801_);
  and (_40803_, _40379_, _40282_);
  and (_40804_, _40803_, _40378_);
  not (_40805_, _40803_);
  and (_40806_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_42056_, _40806_, _40804_);
  and (_40807_, _40803_, _40384_);
  and (_40808_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_42060_, _40808_, _40807_);
  and (_40809_, _40803_, _40387_);
  and (_40810_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_42064_, _40810_, _40809_);
  and (_40811_, _40803_, _40390_);
  and (_40812_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_42068_, _40812_, _40811_);
  and (_40813_, _40803_, _40394_);
  not (_40814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_40815_, _40803_, _40814_);
  or (_42072_, _40815_, _40813_);
  and (_40816_, _40803_, _40398_);
  not (_40817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_40818_, _40803_, _40817_);
  or (_42076_, _40818_, _40816_);
  and (_40819_, _40803_, _40402_);
  and (_40820_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_42080_, _40820_, _40819_);
  and (_40821_, _40803_, _40293_);
  and (_40822_, _40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_42083_, _40822_, _40821_);
  and (_40823_, _40408_, _40282_);
  and (_40824_, _40823_, _40378_);
  not (_40825_, _40823_);
  and (_40826_, _40825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_42088_, _40826_, _40824_);
  and (_40827_, _40823_, _40384_);
  and (_40828_, _40825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_42092_, _40828_, _40827_);
  and (_40829_, _40823_, _40387_);
  not (_40830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_40831_, _40823_, _40830_);
  or (_42096_, _40831_, _40829_);
  and (_40832_, _40823_, _40390_);
  and (_40833_, _40825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_42099_, _40833_, _40832_);
  and (_40834_, _40823_, _40394_);
  not (_40835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_40836_, _40823_, _40835_);
  or (_42103_, _40836_, _40834_);
  and (_40837_, _40823_, _40398_);
  not (_40838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_40839_, _40823_, _40838_);
  or (_42106_, _40839_, _40837_);
  and (_40840_, _40823_, _40402_);
  not (_40841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_40842_, _40823_, _40841_);
  or (_42110_, _40842_, _40840_);
  and (_40843_, _40823_, _40293_);
  nor (_40844_, _40823_, _40264_);
  or (_42113_, _40844_, _40843_);
  and (_40845_, _40378_, _40283_);
  not (_40846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_40847_, _40283_, _40846_);
  or (_42118_, _40847_, _40845_);
  and (_40848_, _40384_, _40283_);
  not (_40849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_40850_, _40283_, _40849_);
  or (_42122_, _40850_, _40848_);
  and (_40851_, _40387_, _40283_);
  not (_40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_40853_, _40283_, _40852_);
  or (_42126_, _40853_, _40851_);
  and (_40854_, _40390_, _40283_);
  not (_40855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_40856_, _40283_, _40855_);
  or (_42129_, _40856_, _40854_);
  and (_40857_, _40394_, _40283_);
  not (_40858_, _40283_);
  and (_40859_, _40858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_42133_, _40859_, _40857_);
  and (_40860_, _40398_, _40283_);
  and (_40861_, _40858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_42137_, _40861_, _40860_);
  and (_40862_, _40402_, _40283_);
  and (_40863_, _40858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_42141_, _40863_, _40862_);
  or (_40864_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_40865_, _39986_, _40311_);
  and (_40866_, _40865_, _40160_);
  and (_40867_, _40866_, _40864_);
  nor (_40868_, _39986_, _40434_);
  and (_40869_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_40870_, _40869_, _40868_);
  and (_40871_, _40870_, _40226_);
  or (_40872_, _40871_, _40867_);
  or (_40873_, _40872_, _40220_);
  or (_40874_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_40875_, _39986_, _40457_);
  and (_40876_, _40875_, _40160_);
  and (_40877_, _40876_, _40874_);
  nor (_40878_, _39986_, _40564_);
  and (_40879_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_40880_, _40879_, _40878_);
  and (_40881_, _40880_, _40226_);
  or (_40882_, _40881_, _40877_);
  or (_40883_, _40882_, _40071_);
  and (_40884_, _40883_, _40234_);
  and (_40885_, _40884_, _40873_);
  nand (_40886_, _39986_, _40644_);
  or (_40887_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_40888_, _40887_, _40886_);
  and (_40889_, _40888_, _40160_);
  and (_40890_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_40891_, _39986_, _40761_);
  or (_40892_, _40891_, _40890_);
  and (_40893_, _40892_, _40226_);
  or (_40894_, _40893_, _40889_);
  or (_40895_, _40894_, _40220_);
  nand (_40896_, _39986_, _40783_);
  or (_40897_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_40898_, _40897_, _40896_);
  and (_40899_, _40898_, _40160_);
  and (_40900_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_40901_, _39986_, _40846_);
  or (_40902_, _40901_, _40900_);
  and (_40903_, _40902_, _40226_);
  or (_40904_, _40903_, _40899_);
  or (_40905_, _40904_, _40071_);
  and (_40906_, _40905_, _40209_);
  and (_40907_, _40906_, _40895_);
  or (_40908_, _40907_, _40885_);
  or (_40909_, _40908_, _40219_);
  or (_40910_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_40911_, _40910_, _43998_);
  and (_43977_, _40911_, _40909_);
  or (_40912_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_40913_, _39986_, _40324_);
  and (_40914_, _40913_, _40160_);
  and (_40915_, _40914_, _40912_);
  nor (_40916_, _39986_, _40437_);
  and (_40917_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_40918_, _40917_, _40916_);
  and (_40919_, _40918_, _40226_);
  or (_40920_, _40919_, _40915_);
  or (_40921_, _40920_, _40220_);
  or (_40922_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_40923_, _39986_, _40460_);
  and (_40924_, _40923_, _40160_);
  and (_40925_, _40924_, _40922_);
  nor (_40926_, _39986_, _40575_);
  and (_40927_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_40928_, _40927_, _40926_);
  and (_40929_, _40928_, _40226_);
  or (_40930_, _40929_, _40925_);
  or (_40931_, _40930_, _40071_);
  and (_40932_, _40931_, _40234_);
  and (_40933_, _40932_, _40921_);
  nand (_40934_, _39986_, _40655_);
  or (_40935_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_40936_, _40935_, _40934_);
  and (_40937_, _40936_, _40160_);
  and (_40938_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_40939_, _39986_, _40764_);
  or (_40940_, _40939_, _40938_);
  and (_40941_, _40940_, _40226_);
  or (_40942_, _40941_, _40937_);
  or (_40943_, _40942_, _40220_);
  nand (_40944_, _39986_, _40786_);
  or (_40945_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_40946_, _40945_, _40944_);
  and (_40947_, _40946_, _40160_);
  and (_40948_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_40949_, _39986_, _40849_);
  or (_40950_, _40949_, _40948_);
  and (_40951_, _40950_, _40226_);
  or (_40952_, _40951_, _40947_);
  or (_40953_, _40952_, _40071_);
  and (_40954_, _40953_, _40209_);
  and (_40955_, _40954_, _40943_);
  or (_40956_, _40955_, _40933_);
  or (_40957_, _40956_, _40219_);
  or (_40958_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_40959_, _40958_, _43998_);
  and (_43979_, _40959_, _40957_);
  and (_40960_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_40961_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_40962_, _40961_, _40960_);
  and (_40963_, _40962_, _40160_);
  nor (_40964_, _39986_, _40440_);
  and (_40965_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_40966_, _40965_, _40964_);
  and (_40967_, _40966_, _40226_);
  or (_40968_, _40967_, _40963_);
  or (_40969_, _40968_, _40220_);
  and (_40970_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_40971_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_40972_, _40971_, _40970_);
  and (_40973_, _40972_, _40160_);
  nor (_40974_, _39986_, _40586_);
  and (_40975_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_40976_, _40975_, _40974_);
  and (_40977_, _40976_, _40226_);
  or (_40978_, _40977_, _40973_);
  or (_40979_, _40978_, _40071_);
  and (_40980_, _40979_, _40234_);
  and (_40981_, _40980_, _40969_);
  or (_40982_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_40983_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_40984_, _40983_, _40982_);
  and (_40985_, _40984_, _40160_);
  or (_40986_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_40987_, _39986_, _40744_);
  and (_40988_, _40987_, _40986_);
  and (_40989_, _40988_, _40226_);
  or (_40990_, _40989_, _40985_);
  or (_40991_, _40990_, _40220_);
  or (_40992_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_40993_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_40994_, _40993_, _40992_);
  and (_40995_, _40994_, _40160_);
  or (_40996_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_40997_, _39986_, _40830_);
  and (_40998_, _40997_, _40996_);
  and (_40999_, _40998_, _40226_);
  or (_41000_, _40999_, _40995_);
  or (_41001_, _41000_, _40071_);
  and (_41002_, _41001_, _40209_);
  and (_41003_, _41002_, _40991_);
  or (_41004_, _41003_, _40981_);
  or (_41005_, _41004_, _40219_);
  or (_41006_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41007_, _41006_, _43998_);
  and (_43980_, _41007_, _41005_);
  and (_41008_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41009_, _39986_, _40392_);
  or (_41010_, _41009_, _41008_);
  and (_41011_, _41010_, _40160_);
  nor (_41012_, _39986_, _40443_);
  and (_41013_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41014_, _41013_, _41012_);
  and (_41015_, _41014_, _40226_);
  or (_41016_, _41015_, _41011_);
  or (_41017_, _41016_, _40220_);
  or (_41018_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand (_41019_, _39986_, _40466_);
  and (_41020_, _41019_, _40160_);
  and (_41021_, _41020_, _41018_);
  nor (_41022_, _39986_, _40595_);
  and (_41023_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41024_, _41023_, _41022_);
  and (_41025_, _41024_, _40226_);
  or (_41026_, _41025_, _41021_);
  or (_41027_, _41026_, _40071_);
  and (_41028_, _41027_, _40234_);
  and (_41029_, _41028_, _41017_);
  or (_41030_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_41031_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_41032_, _41031_, _41030_);
  and (_41033_, _41032_, _40160_);
  or (_41034_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41035_, _39986_, _40747_);
  and (_41036_, _41035_, _41034_);
  and (_41037_, _41036_, _40226_);
  or (_41038_, _41037_, _41033_);
  or (_41039_, _41038_, _40220_);
  nand (_41040_, _39986_, _40792_);
  or (_41041_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41042_, _41041_, _41040_);
  and (_41043_, _41042_, _40160_);
  and (_41044_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_41045_, _39986_, _40855_);
  or (_41046_, _41045_, _41044_);
  and (_41047_, _41046_, _40226_);
  or (_41048_, _41047_, _41043_);
  or (_41049_, _41048_, _40071_);
  and (_41050_, _41049_, _40209_);
  and (_41051_, _41050_, _41039_);
  or (_41052_, _41051_, _41029_);
  or (_41053_, _41052_, _40219_);
  or (_41054_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41055_, _41054_, _43998_);
  and (_43982_, _41055_, _41053_);
  and (_41056_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41057_, _39986_, _40396_);
  or (_41058_, _41057_, _41056_);
  and (_41059_, _41058_, _40160_);
  or (_41060_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_41061_, _39986_, _40421_);
  and (_41062_, _41061_, _41060_);
  and (_41063_, _41062_, _40226_);
  or (_41064_, _41063_, _41059_);
  or (_41065_, _41064_, _40220_);
  and (_41066_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41067_, _39986_, _40515_);
  or (_41068_, _41067_, _41066_);
  and (_41069_, _41068_, _40160_);
  or (_41070_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_41071_, _39986_, _40536_);
  and (_41072_, _41071_, _41070_);
  and (_41073_, _41072_, _40226_);
  or (_41074_, _41073_, _41069_);
  or (_41075_, _41074_, _40071_);
  and (_41076_, _41075_, _40234_);
  and (_41077_, _41076_, _41065_);
  and (_41078_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41079_, _39986_, _40728_);
  or (_41080_, _41079_, _41078_);
  and (_41081_, _41080_, _40160_);
  or (_41082_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41083_, _39986_, _40750_);
  and (_41084_, _41083_, _41082_);
  and (_41085_, _41084_, _40226_);
  or (_41086_, _41085_, _41081_);
  or (_41087_, _41086_, _40220_);
  and (_41088_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41089_, _39986_, _40814_);
  or (_41090_, _41089_, _41088_);
  and (_41091_, _41090_, _40160_);
  or (_41092_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41093_, _39986_, _40835_);
  and (_41094_, _41093_, _41092_);
  and (_41095_, _41094_, _40226_);
  or (_41096_, _41095_, _41091_);
  or (_41097_, _41096_, _40071_);
  and (_41098_, _41097_, _40209_);
  and (_41099_, _41098_, _41087_);
  or (_41100_, _41099_, _41077_);
  or (_41101_, _41100_, _40219_);
  or (_41102_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41103_, _41102_, _43998_);
  and (_43984_, _41103_, _41101_);
  and (_41104_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41105_, _39986_, _40400_);
  or (_41106_, _41105_, _41104_);
  and (_41107_, _41106_, _40160_);
  or (_41108_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_41109_, _39986_, _40424_);
  and (_41110_, _41109_, _41108_);
  and (_41111_, _41110_, _40226_);
  or (_41112_, _41111_, _41107_);
  or (_41113_, _41112_, _40220_);
  and (_41114_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41115_, _39986_, _40518_);
  or (_41116_, _41115_, _41114_);
  and (_41117_, _41116_, _40160_);
  or (_41118_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_41119_, _39986_, _40539_);
  and (_41120_, _41119_, _41118_);
  and (_41121_, _41120_, _40226_);
  or (_41122_, _41121_, _41117_);
  or (_41123_, _41122_, _40071_);
  and (_41124_, _41123_, _40234_);
  and (_41125_, _41124_, _41113_);
  and (_41126_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41127_, _39986_, _40731_);
  or (_41128_, _41127_, _41126_);
  and (_41129_, _41128_, _40160_);
  or (_41130_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41131_, _39986_, _40753_);
  and (_41132_, _41131_, _41130_);
  and (_41133_, _41132_, _40226_);
  or (_41134_, _41133_, _41129_);
  or (_41135_, _41134_, _40220_);
  and (_41136_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41137_, _39986_, _40817_);
  or (_41138_, _41137_, _41136_);
  and (_41139_, _41138_, _40160_);
  or (_41140_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41141_, _39986_, _40838_);
  and (_41142_, _41141_, _41140_);
  and (_41143_, _41142_, _40226_);
  or (_41144_, _41143_, _41139_);
  or (_41145_, _41144_, _40071_);
  and (_41146_, _41145_, _40209_);
  and (_41147_, _41146_, _41135_);
  or (_41148_, _41147_, _41125_);
  or (_41149_, _41148_, _40219_);
  or (_41150_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41151_, _41150_, _43998_);
  and (_43986_, _41151_, _41149_);
  and (_41152_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41153_, _39986_, _40404_);
  or (_41154_, _41153_, _41152_);
  and (_41155_, _41154_, _40160_);
  or (_41156_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand (_41157_, _39986_, _40427_);
  and (_41158_, _41157_, _41156_);
  and (_41159_, _41158_, _40226_);
  or (_41160_, _41159_, _41155_);
  or (_41161_, _41160_, _40220_);
  or (_41162_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand (_41163_, _39986_, _40473_);
  and (_41164_, _41163_, _40160_);
  and (_41165_, _41164_, _41162_);
  nor (_41166_, _39986_, _40621_);
  and (_41167_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41168_, _41167_, _41166_);
  and (_41169_, _41168_, _40226_);
  or (_41170_, _41169_, _41165_);
  or (_41171_, _41170_, _40071_);
  and (_41172_, _41171_, _40234_);
  and (_41173_, _41172_, _41161_);
  or (_41174_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_41175_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_41176_, _41175_, _41174_);
  and (_41177_, _41176_, _40160_);
  or (_41178_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_41179_, _40222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_41180_, _41179_, _41178_);
  and (_41181_, _41180_, _40226_);
  or (_41182_, _41181_, _41177_);
  or (_41183_, _41182_, _40220_);
  nand (_41184_, _39986_, _40799_);
  or (_41185_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41186_, _41185_, _41184_);
  and (_41187_, _41186_, _40160_);
  or (_41188_, _39986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41189_, _39986_, _40841_);
  and (_41190_, _41189_, _41188_);
  and (_41191_, _41190_, _40226_);
  or (_41192_, _41191_, _41187_);
  or (_41193_, _41192_, _40071_);
  and (_41194_, _41193_, _40209_);
  and (_41195_, _41194_, _41183_);
  or (_41196_, _41195_, _41173_);
  or (_41197_, _41196_, _40219_);
  or (_41198_, _40274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41199_, _41198_, _43998_);
  and (_43988_, _41199_, _41197_);
  or (_41200_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41201_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41202_, _41201_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41203_, _41202_, _41200_);
  nand (_41204_, _41203_, _43998_);
  or (_41205_, \oc8051_gm_cxrom_1.cell0.data [7], _43998_);
  and (_43995_, _41205_, _41204_);
  or (_41206_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41207_, \oc8051_gm_cxrom_1.cell0.data [0], _41201_);
  nand (_41208_, _41207_, _41206_);
  nand (_41209_, _41208_, _43998_);
  or (_41210_, \oc8051_gm_cxrom_1.cell0.data [0], _43998_);
  and (_44001_, _41210_, _41209_);
  or (_41211_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41212_, \oc8051_gm_cxrom_1.cell0.data [1], _41201_);
  nand (_41213_, _41212_, _41211_);
  nand (_41214_, _41213_, _43998_);
  or (_41215_, \oc8051_gm_cxrom_1.cell0.data [1], _43998_);
  and (_44005_, _41215_, _41214_);
  or (_41216_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41217_, \oc8051_gm_cxrom_1.cell0.data [2], _41201_);
  nand (_41218_, _41217_, _41216_);
  nand (_41219_, _41218_, _43998_);
  or (_41220_, \oc8051_gm_cxrom_1.cell0.data [2], _43998_);
  and (_44009_, _41220_, _41219_);
  or (_41221_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41222_, \oc8051_gm_cxrom_1.cell0.data [3], _41201_);
  nand (_41223_, _41222_, _41221_);
  nand (_41224_, _41223_, _43998_);
  or (_41225_, \oc8051_gm_cxrom_1.cell0.data [3], _43998_);
  and (_44012_, _41225_, _41224_);
  or (_41226_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41227_, \oc8051_gm_cxrom_1.cell0.data [4], _41201_);
  nand (_41228_, _41227_, _41226_);
  nand (_41229_, _41228_, _43998_);
  or (_41230_, \oc8051_gm_cxrom_1.cell0.data [4], _43998_);
  and (_44016_, _41230_, _41229_);
  or (_41231_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41232_, \oc8051_gm_cxrom_1.cell0.data [5], _41201_);
  nand (_41233_, _41232_, _41231_);
  nand (_41234_, _41233_, _43998_);
  or (_41235_, \oc8051_gm_cxrom_1.cell0.data [5], _43998_);
  and (_44020_, _41235_, _41234_);
  or (_41236_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41237_, \oc8051_gm_cxrom_1.cell0.data [6], _41201_);
  nand (_41238_, _41237_, _41236_);
  nand (_41239_, _41238_, _43998_);
  or (_41240_, \oc8051_gm_cxrom_1.cell0.data [6], _43998_);
  and (_44023_, _41240_, _41239_);
  or (_41241_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41242_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41243_, _41242_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41244_, _41243_, _41241_);
  nand (_41245_, _41244_, _43998_);
  or (_41246_, \oc8051_gm_cxrom_1.cell1.data [7], _43998_);
  and (_44043_, _41246_, _41245_);
  or (_41247_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41248_, \oc8051_gm_cxrom_1.cell1.data [0], _41242_);
  nand (_41249_, _41248_, _41247_);
  nand (_41250_, _41249_, _43998_);
  or (_41251_, \oc8051_gm_cxrom_1.cell1.data [0], _43998_);
  and (_44049_, _41251_, _41250_);
  or (_41252_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41253_, \oc8051_gm_cxrom_1.cell1.data [1], _41242_);
  nand (_41254_, _41253_, _41252_);
  nand (_41255_, _41254_, _43998_);
  or (_41256_, \oc8051_gm_cxrom_1.cell1.data [1], _43998_);
  and (_44053_, _41256_, _41255_);
  or (_41257_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41258_, \oc8051_gm_cxrom_1.cell1.data [2], _41242_);
  nand (_41259_, _41258_, _41257_);
  nand (_41260_, _41259_, _43998_);
  or (_41261_, \oc8051_gm_cxrom_1.cell1.data [2], _43998_);
  and (_44056_, _41261_, _41260_);
  or (_41262_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41263_, \oc8051_gm_cxrom_1.cell1.data [3], _41242_);
  nand (_41264_, _41263_, _41262_);
  nand (_41265_, _41264_, _43998_);
  or (_41266_, \oc8051_gm_cxrom_1.cell1.data [3], _43998_);
  and (_44060_, _41266_, _41265_);
  or (_41267_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41268_, \oc8051_gm_cxrom_1.cell1.data [4], _41242_);
  nand (_41269_, _41268_, _41267_);
  nand (_41270_, _41269_, _43998_);
  or (_41271_, \oc8051_gm_cxrom_1.cell1.data [4], _43998_);
  and (_44063_, _41271_, _41270_);
  or (_41272_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41273_, \oc8051_gm_cxrom_1.cell1.data [5], _41242_);
  nand (_41274_, _41273_, _41272_);
  nand (_41275_, _41274_, _43998_);
  or (_41276_, \oc8051_gm_cxrom_1.cell1.data [5], _43998_);
  and (_44067_, _41276_, _41275_);
  or (_41277_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41278_, \oc8051_gm_cxrom_1.cell1.data [6], _41242_);
  nand (_41279_, _41278_, _41277_);
  nand (_41280_, _41279_, _43998_);
  or (_41281_, \oc8051_gm_cxrom_1.cell1.data [6], _43998_);
  and (_44071_, _41281_, _41280_);
  or (_41283_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41285_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41287_, _41285_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41289_, _41287_, _41283_);
  nand (_41291_, _41289_, _43998_);
  or (_41293_, \oc8051_gm_cxrom_1.cell2.data [7], _43998_);
  and (_44090_, _41293_, _41291_);
  or (_41296_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41298_, \oc8051_gm_cxrom_1.cell2.data [0], _41285_);
  nand (_41300_, _41298_, _41296_);
  nand (_41302_, _41300_, _43998_);
  or (_41304_, \oc8051_gm_cxrom_1.cell2.data [0], _43998_);
  and (_44097_, _41304_, _41302_);
  or (_41307_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41309_, \oc8051_gm_cxrom_1.cell2.data [1], _41285_);
  nand (_41311_, _41309_, _41307_);
  nand (_41313_, _41311_, _43998_);
  or (_41315_, \oc8051_gm_cxrom_1.cell2.data [1], _43998_);
  and (_44100_, _41315_, _41313_);
  or (_41318_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41320_, \oc8051_gm_cxrom_1.cell2.data [2], _41285_);
  nand (_41322_, _41320_, _41318_);
  nand (_41324_, _41322_, _43998_);
  or (_41326_, \oc8051_gm_cxrom_1.cell2.data [2], _43998_);
  and (_44104_, _41326_, _41324_);
  or (_41329_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41331_, \oc8051_gm_cxrom_1.cell2.data [3], _41285_);
  nand (_41333_, _41331_, _41329_);
  nand (_41334_, _41333_, _43998_);
  or (_41335_, \oc8051_gm_cxrom_1.cell2.data [3], _43998_);
  and (_00008_, _41335_, _41334_);
  or (_41336_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41337_, \oc8051_gm_cxrom_1.cell2.data [4], _41285_);
  nand (_41338_, _41337_, _41336_);
  nand (_41339_, _41338_, _43998_);
  or (_41340_, \oc8051_gm_cxrom_1.cell2.data [4], _43998_);
  and (_00009_, _41340_, _41339_);
  or (_41341_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41342_, \oc8051_gm_cxrom_1.cell2.data [5], _41285_);
  nand (_41343_, _41342_, _41341_);
  nand (_41344_, _41343_, _43998_);
  or (_41345_, \oc8051_gm_cxrom_1.cell2.data [5], _43998_);
  and (_00010_, _41345_, _41344_);
  or (_41346_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41347_, \oc8051_gm_cxrom_1.cell2.data [6], _41285_);
  nand (_41348_, _41347_, _41346_);
  nand (_41349_, _41348_, _43998_);
  or (_41350_, \oc8051_gm_cxrom_1.cell2.data [6], _43998_);
  and (_00013_, _41350_, _41349_);
  or (_41351_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_41352_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_41353_, _41352_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_41354_, _41353_, _41351_);
  nand (_41355_, _41354_, _43998_);
  or (_41356_, \oc8051_gm_cxrom_1.cell3.data [7], _43998_);
  and (_00030_, _41356_, _41355_);
  or (_41357_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41358_, \oc8051_gm_cxrom_1.cell3.data [0], _41352_);
  nand (_41359_, _41358_, _41357_);
  nand (_41360_, _41359_, _43998_);
  or (_41361_, \oc8051_gm_cxrom_1.cell3.data [0], _43998_);
  and (_00036_, _41361_, _41360_);
  or (_41362_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41363_, \oc8051_gm_cxrom_1.cell3.data [1], _41352_);
  nand (_41364_, _41363_, _41362_);
  nand (_41365_, _41364_, _43998_);
  or (_41366_, \oc8051_gm_cxrom_1.cell3.data [1], _43998_);
  and (_00039_, _41366_, _41365_);
  or (_41367_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41368_, \oc8051_gm_cxrom_1.cell3.data [2], _41352_);
  nand (_41369_, _41368_, _41367_);
  nand (_41370_, _41369_, _43998_);
  or (_41371_, \oc8051_gm_cxrom_1.cell3.data [2], _43998_);
  and (_00042_, _41371_, _41370_);
  or (_41372_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41373_, \oc8051_gm_cxrom_1.cell3.data [3], _41352_);
  nand (_41374_, _41373_, _41372_);
  nand (_41375_, _41374_, _43998_);
  or (_41376_, \oc8051_gm_cxrom_1.cell3.data [3], _43998_);
  and (_00045_, _41376_, _41375_);
  or (_41377_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41378_, \oc8051_gm_cxrom_1.cell3.data [4], _41352_);
  nand (_41379_, _41378_, _41377_);
  nand (_41380_, _41379_, _43998_);
  or (_41381_, \oc8051_gm_cxrom_1.cell3.data [4], _43998_);
  and (_00046_, _41381_, _41380_);
  or (_41382_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41383_, \oc8051_gm_cxrom_1.cell3.data [5], _41352_);
  nand (_41384_, _41383_, _41382_);
  nand (_41385_, _41384_, _43998_);
  or (_41386_, \oc8051_gm_cxrom_1.cell3.data [5], _43998_);
  and (_00050_, _41386_, _41385_);
  or (_41387_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41388_, \oc8051_gm_cxrom_1.cell3.data [6], _41352_);
  nand (_41389_, _41388_, _41387_);
  nand (_41390_, _41389_, _43998_);
  or (_41391_, \oc8051_gm_cxrom_1.cell3.data [6], _43998_);
  and (_00053_, _41391_, _41390_);
  or (_41392_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_41393_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_41394_, _41393_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_41395_, _41394_, _41392_);
  nand (_41396_, _41395_, _43998_);
  or (_41397_, \oc8051_gm_cxrom_1.cell4.data [7], _43998_);
  and (_00070_, _41397_, _41396_);
  or (_41398_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41399_, \oc8051_gm_cxrom_1.cell4.data [0], _41393_);
  nand (_41400_, _41399_, _41398_);
  nand (_41401_, _41400_, _43998_);
  or (_41402_, \oc8051_gm_cxrom_1.cell4.data [0], _43998_);
  and (_00075_, _41402_, _41401_);
  or (_41403_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41404_, \oc8051_gm_cxrom_1.cell4.data [1], _41393_);
  nand (_41405_, _41404_, _41403_);
  nand (_41406_, _41405_, _43998_);
  or (_41407_, \oc8051_gm_cxrom_1.cell4.data [1], _43998_);
  and (_00079_, _41407_, _41406_);
  or (_41409_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41410_, \oc8051_gm_cxrom_1.cell4.data [2], _41393_);
  nand (_41411_, _41410_, _41409_);
  nand (_41412_, _41411_, _43998_);
  or (_41413_, \oc8051_gm_cxrom_1.cell4.data [2], _43998_);
  and (_00082_, _41413_, _41412_);
  or (_41414_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41415_, \oc8051_gm_cxrom_1.cell4.data [3], _41393_);
  nand (_41416_, _41415_, _41414_);
  nand (_41417_, _41416_, _43998_);
  or (_41419_, \oc8051_gm_cxrom_1.cell4.data [3], _43998_);
  and (_00085_, _41419_, _41417_);
  or (_41420_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41421_, \oc8051_gm_cxrom_1.cell4.data [4], _41393_);
  nand (_41422_, _41421_, _41420_);
  nand (_41423_, _41422_, _43998_);
  or (_41424_, \oc8051_gm_cxrom_1.cell4.data [4], _43998_);
  and (_00088_, _41424_, _41423_);
  or (_41425_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41426_, \oc8051_gm_cxrom_1.cell4.data [5], _41393_);
  nand (_41427_, _41426_, _41425_);
  nand (_41428_, _41427_, _43998_);
  or (_41429_, \oc8051_gm_cxrom_1.cell4.data [5], _43998_);
  and (_00092_, _41429_, _41428_);
  or (_41430_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41431_, \oc8051_gm_cxrom_1.cell4.data [6], _41393_);
  nand (_41432_, _41431_, _41430_);
  nand (_41433_, _41432_, _43998_);
  or (_41434_, \oc8051_gm_cxrom_1.cell4.data [6], _43998_);
  and (_00095_, _41434_, _41433_);
  or (_41435_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_41436_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_41437_, _41436_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_41438_, _41437_, _41435_);
  nand (_41439_, _41438_, _43998_);
  or (_41440_, \oc8051_gm_cxrom_1.cell5.data [7], _43998_);
  and (_00112_, _41440_, _41439_);
  or (_41441_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41442_, \oc8051_gm_cxrom_1.cell5.data [0], _41436_);
  nand (_41443_, _41442_, _41441_);
  nand (_41444_, _41443_, _43998_);
  or (_41445_, \oc8051_gm_cxrom_1.cell5.data [0], _43998_);
  and (_00117_, _41445_, _41444_);
  or (_41446_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41447_, \oc8051_gm_cxrom_1.cell5.data [1], _41436_);
  nand (_41448_, _41447_, _41446_);
  nand (_41449_, _41448_, _43998_);
  or (_41450_, \oc8051_gm_cxrom_1.cell5.data [1], _43998_);
  and (_00121_, _41450_, _41449_);
  or (_41451_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41452_, \oc8051_gm_cxrom_1.cell5.data [2], _41436_);
  nand (_41453_, _41452_, _41451_);
  nand (_41454_, _41453_, _43998_);
  or (_41455_, \oc8051_gm_cxrom_1.cell5.data [2], _43998_);
  and (_00124_, _41455_, _41454_);
  or (_41456_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41457_, \oc8051_gm_cxrom_1.cell5.data [3], _41436_);
  nand (_41458_, _41457_, _41456_);
  nand (_41459_, _41458_, _43998_);
  or (_41460_, \oc8051_gm_cxrom_1.cell5.data [3], _43998_);
  and (_00127_, _41460_, _41459_);
  or (_41461_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41462_, \oc8051_gm_cxrom_1.cell5.data [4], _41436_);
  nand (_41463_, _41462_, _41461_);
  nand (_41464_, _41463_, _43998_);
  or (_41465_, \oc8051_gm_cxrom_1.cell5.data [4], _43998_);
  and (_00130_, _41465_, _41464_);
  or (_41466_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41467_, \oc8051_gm_cxrom_1.cell5.data [5], _41436_);
  nand (_41468_, _41467_, _41466_);
  nand (_41469_, _41468_, _43998_);
  or (_41470_, \oc8051_gm_cxrom_1.cell5.data [5], _43998_);
  and (_00134_, _41470_, _41469_);
  or (_41471_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41472_, \oc8051_gm_cxrom_1.cell5.data [6], _41436_);
  nand (_41473_, _41472_, _41471_);
  nand (_41474_, _41473_, _43998_);
  or (_41475_, \oc8051_gm_cxrom_1.cell5.data [6], _43998_);
  and (_00137_, _41475_, _41474_);
  or (_41476_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_41477_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_41478_, _41477_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_41479_, _41478_, _41476_);
  nand (_41480_, _41479_, _43998_);
  or (_41481_, \oc8051_gm_cxrom_1.cell6.data [7], _43998_);
  and (_00154_, _41481_, _41480_);
  or (_41482_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41483_, \oc8051_gm_cxrom_1.cell6.data [0], _41477_);
  nand (_41484_, _41483_, _41482_);
  nand (_41485_, _41484_, _43998_);
  or (_41486_, \oc8051_gm_cxrom_1.cell6.data [0], _43998_);
  and (_00159_, _41486_, _41485_);
  or (_41487_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41488_, \oc8051_gm_cxrom_1.cell6.data [1], _41477_);
  nand (_41489_, _41488_, _41487_);
  nand (_41490_, _41489_, _43998_);
  or (_41491_, \oc8051_gm_cxrom_1.cell6.data [1], _43998_);
  and (_00163_, _41491_, _41490_);
  or (_41492_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41493_, \oc8051_gm_cxrom_1.cell6.data [2], _41477_);
  nand (_41494_, _41493_, _41492_);
  nand (_41495_, _41494_, _43998_);
  or (_41496_, \oc8051_gm_cxrom_1.cell6.data [2], _43998_);
  and (_00166_, _41496_, _41495_);
  or (_41497_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41498_, \oc8051_gm_cxrom_1.cell6.data [3], _41477_);
  nand (_41499_, _41498_, _41497_);
  nand (_41500_, _41499_, _43998_);
  or (_41501_, \oc8051_gm_cxrom_1.cell6.data [3], _43998_);
  and (_00169_, _41501_, _41500_);
  or (_41502_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41503_, \oc8051_gm_cxrom_1.cell6.data [4], _41477_);
  nand (_41504_, _41503_, _41502_);
  nand (_41505_, _41504_, _43998_);
  or (_41506_, \oc8051_gm_cxrom_1.cell6.data [4], _43998_);
  and (_00172_, _41506_, _41505_);
  or (_41507_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41508_, \oc8051_gm_cxrom_1.cell6.data [5], _41477_);
  nand (_41509_, _41508_, _41507_);
  nand (_41510_, _41509_, _43998_);
  or (_41511_, \oc8051_gm_cxrom_1.cell6.data [5], _43998_);
  and (_00176_, _41511_, _41510_);
  or (_41512_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41513_, \oc8051_gm_cxrom_1.cell6.data [6], _41477_);
  nand (_41514_, _41513_, _41512_);
  nand (_41515_, _41514_, _43998_);
  or (_41516_, \oc8051_gm_cxrom_1.cell6.data [6], _43998_);
  and (_00179_, _41516_, _41515_);
  or (_41517_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_41518_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_41519_, _41518_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_41520_, _41519_, _41517_);
  nand (_41521_, _41520_, _43998_);
  or (_41522_, \oc8051_gm_cxrom_1.cell7.data [7], _43998_);
  and (_00196_, _41522_, _41521_);
  or (_41523_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41524_, \oc8051_gm_cxrom_1.cell7.data [0], _41518_);
  nand (_41525_, _41524_, _41523_);
  nand (_41526_, _41525_, _43998_);
  or (_41527_, \oc8051_gm_cxrom_1.cell7.data [0], _43998_);
  and (_00203_, _41527_, _41526_);
  or (_41528_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41529_, \oc8051_gm_cxrom_1.cell7.data [1], _41518_);
  nand (_41530_, _41529_, _41528_);
  nand (_41531_, _41530_, _43998_);
  or (_41532_, \oc8051_gm_cxrom_1.cell7.data [1], _43998_);
  and (_00206_, _41532_, _41531_);
  or (_41533_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41534_, \oc8051_gm_cxrom_1.cell7.data [2], _41518_);
  nand (_41535_, _41534_, _41533_);
  nand (_41536_, _41535_, _43998_);
  or (_41537_, \oc8051_gm_cxrom_1.cell7.data [2], _43998_);
  and (_00210_, _41537_, _41536_);
  or (_41538_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41539_, \oc8051_gm_cxrom_1.cell7.data [3], _41518_);
  nand (_41540_, _41539_, _41538_);
  nand (_41541_, _41540_, _43998_);
  or (_41542_, \oc8051_gm_cxrom_1.cell7.data [3], _43998_);
  and (_00213_, _41542_, _41541_);
  or (_41543_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41544_, \oc8051_gm_cxrom_1.cell7.data [4], _41518_);
  nand (_41545_, _41544_, _41543_);
  nand (_41546_, _41545_, _43998_);
  or (_41547_, \oc8051_gm_cxrom_1.cell7.data [4], _43998_);
  and (_00217_, _41547_, _41546_);
  or (_41548_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41549_, \oc8051_gm_cxrom_1.cell7.data [5], _41518_);
  nand (_41550_, _41549_, _41548_);
  nand (_41551_, _41550_, _43998_);
  or (_41552_, \oc8051_gm_cxrom_1.cell7.data [5], _43998_);
  and (_00221_, _41552_, _41551_);
  or (_41553_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41554_, \oc8051_gm_cxrom_1.cell7.data [6], _41518_);
  nand (_41555_, _41554_, _41553_);
  nand (_41556_, _41555_, _43998_);
  or (_41557_, \oc8051_gm_cxrom_1.cell7.data [6], _43998_);
  and (_00224_, _41557_, _41556_);
  or (_41558_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_41559_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_41560_, _41559_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_41561_, _41560_, _41558_);
  nand (_41562_, _41561_, _43998_);
  or (_41563_, \oc8051_gm_cxrom_1.cell8.data [7], _43998_);
  and (_00243_, _41563_, _41562_);
  or (_41564_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41565_, \oc8051_gm_cxrom_1.cell8.data [0], _41559_);
  nand (_41566_, _41565_, _41564_);
  nand (_41567_, _41566_, _43998_);
  or (_41568_, \oc8051_gm_cxrom_1.cell8.data [0], _43998_);
  and (_00249_, _41568_, _41567_);
  or (_41569_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41570_, \oc8051_gm_cxrom_1.cell8.data [1], _41559_);
  nand (_41571_, _41570_, _41569_);
  nand (_41572_, _41571_, _43998_);
  or (_41573_, \oc8051_gm_cxrom_1.cell8.data [1], _43998_);
  and (_00253_, _41573_, _41572_);
  or (_41574_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41575_, \oc8051_gm_cxrom_1.cell8.data [2], _41559_);
  nand (_41576_, _41575_, _41574_);
  nand (_41577_, _41576_, _43998_);
  or (_41578_, \oc8051_gm_cxrom_1.cell8.data [2], _43998_);
  and (_00256_, _41578_, _41577_);
  or (_41579_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41580_, \oc8051_gm_cxrom_1.cell8.data [3], _41559_);
  nand (_41581_, _41580_, _41579_);
  nand (_41582_, _41581_, _43998_);
  or (_41583_, \oc8051_gm_cxrom_1.cell8.data [3], _43998_);
  and (_00260_, _41583_, _41582_);
  or (_41584_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41585_, \oc8051_gm_cxrom_1.cell8.data [4], _41559_);
  nand (_41586_, _41585_, _41584_);
  nand (_41587_, _41586_, _43998_);
  or (_41588_, \oc8051_gm_cxrom_1.cell8.data [4], _43998_);
  and (_00263_, _41588_, _41587_);
  or (_41589_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41590_, \oc8051_gm_cxrom_1.cell8.data [5], _41559_);
  nand (_41591_, _41590_, _41589_);
  nand (_41592_, _41591_, _43998_);
  or (_41593_, \oc8051_gm_cxrom_1.cell8.data [5], _43998_);
  and (_00266_, _41593_, _41592_);
  or (_41594_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41595_, \oc8051_gm_cxrom_1.cell8.data [6], _41559_);
  nand (_41596_, _41595_, _41594_);
  nand (_41597_, _41596_, _43998_);
  or (_41598_, \oc8051_gm_cxrom_1.cell8.data [6], _43998_);
  and (_00270_, _41598_, _41597_);
  or (_41599_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_41600_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_41601_, _41600_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_41602_, _41601_, _41599_);
  nand (_41603_, _41602_, _43998_);
  or (_41604_, \oc8051_gm_cxrom_1.cell9.data [7], _43998_);
  and (_00287_, _41604_, _41603_);
  or (_41605_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41606_, \oc8051_gm_cxrom_1.cell9.data [0], _41600_);
  nand (_41607_, _41606_, _41605_);
  nand (_41608_, _41607_, _43998_);
  or (_41609_, \oc8051_gm_cxrom_1.cell9.data [0], _43998_);
  and (_00293_, _41609_, _41608_);
  or (_41610_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41611_, \oc8051_gm_cxrom_1.cell9.data [1], _41600_);
  nand (_41612_, _41611_, _41610_);
  nand (_41613_, _41612_, _43998_);
  or (_41614_, \oc8051_gm_cxrom_1.cell9.data [1], _43998_);
  and (_00296_, _41614_, _41613_);
  or (_41615_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41616_, \oc8051_gm_cxrom_1.cell9.data [2], _41600_);
  nand (_41617_, _41616_, _41615_);
  nand (_41618_, _41617_, _43998_);
  or (_41619_, \oc8051_gm_cxrom_1.cell9.data [2], _43998_);
  and (_00300_, _41619_, _41618_);
  or (_41620_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41621_, \oc8051_gm_cxrom_1.cell9.data [3], _41600_);
  nand (_41622_, _41621_, _41620_);
  nand (_41623_, _41622_, _43998_);
  or (_41624_, \oc8051_gm_cxrom_1.cell9.data [3], _43998_);
  and (_00303_, _41624_, _41623_);
  or (_41625_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41626_, \oc8051_gm_cxrom_1.cell9.data [4], _41600_);
  nand (_41627_, _41626_, _41625_);
  nand (_41628_, _41627_, _43998_);
  or (_41629_, \oc8051_gm_cxrom_1.cell9.data [4], _43998_);
  and (_00306_, _41629_, _41628_);
  or (_41630_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41631_, \oc8051_gm_cxrom_1.cell9.data [5], _41600_);
  nand (_41632_, _41631_, _41630_);
  nand (_41633_, _41632_, _43998_);
  or (_41634_, \oc8051_gm_cxrom_1.cell9.data [5], _43998_);
  and (_00309_, _41634_, _41633_);
  or (_41635_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41636_, \oc8051_gm_cxrom_1.cell9.data [6], _41600_);
  nand (_41637_, _41636_, _41635_);
  nand (_41638_, _41637_, _43998_);
  or (_41639_, \oc8051_gm_cxrom_1.cell9.data [6], _43998_);
  and (_00313_, _41639_, _41638_);
  or (_41640_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_41641_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_41642_, _41641_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_41643_, _41642_, _41640_);
  nand (_41644_, _41643_, _43998_);
  or (_41645_, \oc8051_gm_cxrom_1.cell10.data [7], _43998_);
  and (_00329_, _41645_, _41644_);
  or (_41646_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41647_, \oc8051_gm_cxrom_1.cell10.data [0], _41641_);
  nand (_41648_, _41647_, _41646_);
  nand (_41649_, _41648_, _43998_);
  or (_41650_, \oc8051_gm_cxrom_1.cell10.data [0], _43998_);
  and (_00335_, _41650_, _41649_);
  or (_41651_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41652_, \oc8051_gm_cxrom_1.cell10.data [1], _41641_);
  nand (_41653_, _41652_, _41651_);
  nand (_41654_, _41653_, _43998_);
  or (_41655_, \oc8051_gm_cxrom_1.cell10.data [1], _43998_);
  and (_00338_, _41655_, _41654_);
  or (_41656_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41657_, \oc8051_gm_cxrom_1.cell10.data [2], _41641_);
  nand (_41658_, _41657_, _41656_);
  nand (_41659_, _41658_, _43998_);
  or (_41660_, \oc8051_gm_cxrom_1.cell10.data [2], _43998_);
  and (_00342_, _41660_, _41659_);
  or (_41662_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41663_, \oc8051_gm_cxrom_1.cell10.data [3], _41641_);
  nand (_41664_, _41663_, _41662_);
  nand (_41665_, _41664_, _43998_);
  or (_41667_, \oc8051_gm_cxrom_1.cell10.data [3], _43998_);
  and (_00344_, _41667_, _41665_);
  or (_41668_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41669_, \oc8051_gm_cxrom_1.cell10.data [4], _41641_);
  nand (_41670_, _41669_, _41668_);
  nand (_41672_, _41670_, _43998_);
  or (_41673_, \oc8051_gm_cxrom_1.cell10.data [4], _43998_);
  and (_00348_, _41673_, _41672_);
  or (_41674_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41675_, \oc8051_gm_cxrom_1.cell10.data [5], _41641_);
  nand (_41677_, _41675_, _41674_);
  nand (_41678_, _41677_, _43998_);
  or (_41679_, \oc8051_gm_cxrom_1.cell10.data [5], _43998_);
  and (_00352_, _41679_, _41678_);
  or (_41680_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41682_, \oc8051_gm_cxrom_1.cell10.data [6], _41641_);
  nand (_41683_, _41682_, _41680_);
  nand (_41684_, _41683_, _43998_);
  or (_41685_, \oc8051_gm_cxrom_1.cell10.data [6], _43998_);
  and (_00356_, _41685_, _41684_);
  or (_41687_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_41688_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_41689_, _41688_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_41690_, _41689_, _41687_);
  nand (_41691_, _41690_, _43998_);
  or (_41693_, \oc8051_gm_cxrom_1.cell11.data [7], _43998_);
  and (_00378_, _41693_, _41691_);
  or (_41695_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41696_, \oc8051_gm_cxrom_1.cell11.data [0], _41688_);
  nand (_41697_, _41696_, _41695_);
  nand (_41698_, _41697_, _43998_);
  or (_41699_, \oc8051_gm_cxrom_1.cell11.data [0], _43998_);
  and (_00385_, _41699_, _41698_);
  or (_41700_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41702_, \oc8051_gm_cxrom_1.cell11.data [1], _41688_);
  nand (_41703_, _41702_, _41700_);
  nand (_41704_, _41703_, _43998_);
  or (_41706_, \oc8051_gm_cxrom_1.cell11.data [1], _43998_);
  and (_00389_, _41706_, _41704_);
  or (_41707_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41709_, \oc8051_gm_cxrom_1.cell11.data [2], _41688_);
  nand (_41710_, _41709_, _41707_);
  nand (_41711_, _41710_, _43998_);
  or (_41713_, \oc8051_gm_cxrom_1.cell11.data [2], _43998_);
  and (_00393_, _41713_, _41711_);
  or (_41714_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41716_, \oc8051_gm_cxrom_1.cell11.data [3], _41688_);
  nand (_41717_, _41716_, _41714_);
  nand (_41718_, _41717_, _43998_);
  or (_41720_, \oc8051_gm_cxrom_1.cell11.data [3], _43998_);
  and (_00397_, _41720_, _41718_);
  or (_41721_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41723_, \oc8051_gm_cxrom_1.cell11.data [4], _41688_);
  nand (_41724_, _41723_, _41721_);
  nand (_41726_, _41724_, _43998_);
  or (_41727_, \oc8051_gm_cxrom_1.cell11.data [4], _43998_);
  and (_00401_, _41727_, _41726_);
  or (_41728_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41729_, \oc8051_gm_cxrom_1.cell11.data [5], _41688_);
  nand (_41730_, _41729_, _41728_);
  nand (_41731_, _41730_, _43998_);
  or (_41733_, \oc8051_gm_cxrom_1.cell11.data [5], _43998_);
  and (_00405_, _41733_, _41731_);
  or (_41734_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_41736_, \oc8051_gm_cxrom_1.cell11.data [6], _41688_);
  nand (_41737_, _41736_, _41734_);
  nand (_41738_, _41737_, _43998_);
  or (_41740_, \oc8051_gm_cxrom_1.cell11.data [6], _43998_);
  and (_00409_, _41740_, _41738_);
  or (_41741_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_41743_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_41744_, _41743_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_41745_, _41744_, _41741_);
  nand (_41747_, _41745_, _43998_);
  or (_41748_, \oc8051_gm_cxrom_1.cell12.data [7], _43998_);
  and (_00431_, _41748_, _41747_);
  or (_41750_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41751_, \oc8051_gm_cxrom_1.cell12.data [0], _41743_);
  nand (_41752_, _41751_, _41750_);
  nand (_41754_, _41752_, _43998_);
  or (_41755_, \oc8051_gm_cxrom_1.cell12.data [0], _43998_);
  and (_00438_, _41755_, _41754_);
  or (_41757_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41758_, \oc8051_gm_cxrom_1.cell12.data [1], _41743_);
  nand (_41759_, _41758_, _41757_);
  nand (_41760_, _41759_, _43998_);
  or (_41762_, \oc8051_gm_cxrom_1.cell12.data [1], _43998_);
  and (_00442_, _41762_, _41760_);
  or (_41763_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41765_, \oc8051_gm_cxrom_1.cell12.data [2], _41743_);
  nand (_41766_, _41765_, _41763_);
  nand (_41767_, _41766_, _43998_);
  or (_41769_, \oc8051_gm_cxrom_1.cell12.data [2], _43998_);
  and (_00446_, _41769_, _41767_);
  or (_41770_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41772_, \oc8051_gm_cxrom_1.cell12.data [3], _41743_);
  nand (_41773_, _41772_, _41770_);
  nand (_41774_, _41773_, _43998_);
  or (_41776_, \oc8051_gm_cxrom_1.cell12.data [3], _43998_);
  and (_00450_, _41776_, _41774_);
  or (_41777_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41779_, \oc8051_gm_cxrom_1.cell12.data [4], _41743_);
  nand (_41780_, _41779_, _41777_);
  nand (_41781_, _41780_, _43998_);
  or (_41783_, \oc8051_gm_cxrom_1.cell12.data [4], _43998_);
  and (_00454_, _41783_, _41781_);
  or (_41785_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41786_, \oc8051_gm_cxrom_1.cell12.data [5], _41743_);
  nand (_41787_, _41786_, _41785_);
  nand (_41788_, _41787_, _43998_);
  or (_41789_, \oc8051_gm_cxrom_1.cell12.data [5], _43998_);
  and (_00458_, _41789_, _41788_);
  or (_41790_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_41792_, \oc8051_gm_cxrom_1.cell12.data [6], _41743_);
  nand (_41793_, _41792_, _41790_);
  nand (_41794_, _41793_, _43998_);
  or (_41796_, \oc8051_gm_cxrom_1.cell12.data [6], _43998_);
  and (_00462_, _41796_, _41794_);
  or (_41797_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_41799_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_41800_, _41799_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_41801_, _41800_, _41797_);
  nand (_41803_, _41801_, _43998_);
  or (_41804_, \oc8051_gm_cxrom_1.cell13.data [7], _43998_);
  and (_00484_, _41804_, _41803_);
  or (_41806_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41807_, \oc8051_gm_cxrom_1.cell13.data [0], _41799_);
  nand (_41808_, _41807_, _41806_);
  nand (_41810_, _41808_, _43998_);
  or (_41811_, \oc8051_gm_cxrom_1.cell13.data [0], _43998_);
  and (_00491_, _41811_, _41810_);
  or (_41813_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41814_, \oc8051_gm_cxrom_1.cell13.data [1], _41799_);
  nand (_41816_, _41814_, _41813_);
  nand (_41817_, _41816_, _43998_);
  or (_41818_, \oc8051_gm_cxrom_1.cell13.data [1], _43998_);
  and (_00495_, _41818_, _41817_);
  or (_41820_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41821_, \oc8051_gm_cxrom_1.cell13.data [2], _41799_);
  nand (_41822_, _41821_, _41820_);
  nand (_41824_, _41822_, _43998_);
  or (_41825_, \oc8051_gm_cxrom_1.cell13.data [2], _43998_);
  and (_00499_, _41825_, _41824_);
  or (_41827_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41828_, \oc8051_gm_cxrom_1.cell13.data [3], _41799_);
  nand (_41829_, _41828_, _41827_);
  nand (_41831_, _41829_, _43998_);
  or (_41832_, \oc8051_gm_cxrom_1.cell13.data [3], _43998_);
  and (_00503_, _41832_, _41831_);
  or (_41834_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41835_, \oc8051_gm_cxrom_1.cell13.data [4], _41799_);
  nand (_41836_, _41835_, _41834_);
  nand (_41838_, _41836_, _43998_);
  or (_41839_, \oc8051_gm_cxrom_1.cell13.data [4], _43998_);
  and (_00507_, _41839_, _41838_);
  or (_41841_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41842_, \oc8051_gm_cxrom_1.cell13.data [5], _41799_);
  nand (_41844_, _41842_, _41841_);
  nand (_41845_, _41844_, _43998_);
  or (_41846_, \oc8051_gm_cxrom_1.cell13.data [5], _43998_);
  and (_00511_, _41846_, _41845_);
  or (_41848_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_41849_, \oc8051_gm_cxrom_1.cell13.data [6], _41799_);
  nand (_41850_, _41849_, _41848_);
  nand (_41852_, _41850_, _43998_);
  or (_41853_, \oc8051_gm_cxrom_1.cell13.data [6], _43998_);
  and (_00515_, _41853_, _41852_);
  or (_41855_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_41856_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_41857_, _41856_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_41859_, _41857_, _41855_);
  nand (_41860_, _41859_, _43998_);
  or (_41861_, \oc8051_gm_cxrom_1.cell14.data [7], _43998_);
  and (_00537_, _41861_, _41860_);
  or (_41863_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41864_, \oc8051_gm_cxrom_1.cell14.data [0], _41856_);
  nand (_41866_, _41864_, _41863_);
  nand (_41867_, _41866_, _43998_);
  or (_41868_, \oc8051_gm_cxrom_1.cell14.data [0], _43998_);
  and (_00544_, _41868_, _41867_);
  or (_41870_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41872_, \oc8051_gm_cxrom_1.cell14.data [1], _41856_);
  nand (_41873_, _41872_, _41870_);
  nand (_41874_, _41873_, _43998_);
  or (_41875_, \oc8051_gm_cxrom_1.cell14.data [1], _43998_);
  and (_00548_, _41875_, _41874_);
  or (_41877_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41878_, \oc8051_gm_cxrom_1.cell14.data [2], _41856_);
  nand (_41880_, _41878_, _41877_);
  nand (_41881_, _41880_, _43998_);
  or (_41882_, \oc8051_gm_cxrom_1.cell14.data [2], _43998_);
  and (_00552_, _41882_, _41881_);
  or (_41884_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41885_, \oc8051_gm_cxrom_1.cell14.data [3], _41856_);
  nand (_41887_, _41885_, _41884_);
  nand (_41888_, _41887_, _43998_);
  or (_41889_, \oc8051_gm_cxrom_1.cell14.data [3], _43998_);
  and (_00556_, _41889_, _41888_);
  or (_41891_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41892_, \oc8051_gm_cxrom_1.cell14.data [4], _41856_);
  nand (_41894_, _41892_, _41891_);
  nand (_41895_, _41894_, _43998_);
  or (_41896_, \oc8051_gm_cxrom_1.cell14.data [4], _43998_);
  and (_00560_, _41896_, _41895_);
  or (_41898_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41900_, \oc8051_gm_cxrom_1.cell14.data [5], _41856_);
  nand (_41901_, _41900_, _41898_);
  nand (_41902_, _41901_, _43998_);
  or (_41903_, \oc8051_gm_cxrom_1.cell14.data [5], _43998_);
  and (_00564_, _41903_, _41902_);
  or (_41904_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_41905_, \oc8051_gm_cxrom_1.cell14.data [6], _41856_);
  nand (_41907_, _41905_, _41904_);
  nand (_41908_, _41907_, _43998_);
  or (_41909_, \oc8051_gm_cxrom_1.cell14.data [6], _43998_);
  and (_00568_, _41909_, _41908_);
  or (_41911_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_41912_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_41914_, _41912_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_41915_, _41914_, _41911_);
  or (_41916_, _41915_, rst);
  or (_41918_, \oc8051_gm_cxrom_1.cell15.data [7], _43998_);
  and (_00590_, _41918_, _41916_);
  or (_41919_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41921_, \oc8051_gm_cxrom_1.cell15.data [0], _41912_);
  and (_41922_, _41921_, _41919_);
  or (_41923_, _41922_, rst);
  or (_41925_, \oc8051_gm_cxrom_1.cell15.data [0], _43998_);
  and (_00597_, _41925_, _41923_);
  or (_41926_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41928_, \oc8051_gm_cxrom_1.cell15.data [1], _41912_);
  and (_41929_, _41928_, _41926_);
  or (_41931_, _41929_, rst);
  or (_41932_, \oc8051_gm_cxrom_1.cell15.data [1], _43998_);
  and (_00601_, _41932_, _41931_);
  or (_41933_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41935_, \oc8051_gm_cxrom_1.cell15.data [2], _41912_);
  and (_41936_, _41935_, _41933_);
  or (_41937_, _41936_, rst);
  or (_41939_, \oc8051_gm_cxrom_1.cell15.data [2], _43998_);
  and (_00605_, _41939_, _41937_);
  or (_41940_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41942_, \oc8051_gm_cxrom_1.cell15.data [3], _41912_);
  and (_41943_, _41942_, _41940_);
  or (_41944_, _41943_, rst);
  or (_41946_, \oc8051_gm_cxrom_1.cell15.data [3], _43998_);
  and (_00609_, _41946_, _41944_);
  or (_41947_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41949_, \oc8051_gm_cxrom_1.cell15.data [4], _41912_);
  and (_41950_, _41949_, _41947_);
  or (_41951_, _41950_, rst);
  or (_41953_, \oc8051_gm_cxrom_1.cell15.data [4], _43998_);
  and (_00613_, _41953_, _41951_);
  or (_41954_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41956_, \oc8051_gm_cxrom_1.cell15.data [5], _41912_);
  and (_41957_, _41956_, _41954_);
  or (_41959_, _41957_, rst);
  or (_41960_, \oc8051_gm_cxrom_1.cell15.data [5], _43998_);
  and (_00617_, _41960_, _41959_);
  or (_41961_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_41963_, \oc8051_gm_cxrom_1.cell15.data [6], _41912_);
  and (_41964_, _41963_, _41961_);
  or (_41965_, _41964_, rst);
  or (_41967_, \oc8051_gm_cxrom_1.cell15.data [6], _43998_);
  and (_00621_, _41967_, _41965_);
  nor (_04357_, _37304_, rst);
  and (_41969_, _33213_, _43998_);
  nand (_41970_, _41969_, _36013_);
  nor (_41971_, _35937_, _35828_);
  or (_04360_, _41971_, _41970_);
  not (_41973_, _34857_);
  and (_41974_, _41973_, _34617_);
  not (_41976_, _35118_);
  not (_41977_, _33605_);
  nor (_41978_, _41977_, _34095_);
  and (_41980_, _35741_, _33856_);
  and (_41981_, _41980_, _41978_);
  and (_41982_, _41981_, _41976_);
  and (_41984_, _41982_, _41974_);
  not (_41985_, _33856_);
  and (_41987_, _33605_, _34095_);
  and (_41988_, _41987_, _41985_);
  and (_41989_, _41988_, _35741_);
  and (_41990_, _34857_, _34617_);
  and (_41992_, _41990_, _34367_);
  and (_41993_, _41992_, _41989_);
  or (_41994_, _41993_, _41984_);
  not (_41996_, _34367_);
  and (_41997_, _41990_, _41996_);
  and (_41998_, _41997_, _41989_);
  nor (_42000_, _41976_, _34367_);
  nor (_42001_, _34857_, _34617_);
  and (_42002_, _42001_, _42000_);
  and (_42004_, _42002_, _41988_);
  nor (_42005_, _41976_, _33605_);
  and (_42006_, _42001_, _34367_);
  and (_42008_, _42006_, _42005_);
  or (_42009_, _42008_, _42004_);
  or (_42010_, _42009_, _41998_);
  not (_42012_, _34617_);
  and (_42013_, _34857_, _42012_);
  and (_42014_, _42013_, _42000_);
  not (_42016_, _35741_);
  and (_42017_, _41988_, _42016_);
  and (_42019_, _42017_, _42014_);
  and (_42020_, _35118_, _34367_);
  and (_42021_, _42020_, _42001_);
  and (_42022_, _41978_, _33856_);
  and (_42023_, _42022_, _42016_);
  and (_42025_, _42023_, _42021_);
  or (_42026_, _42025_, _42019_);
  or (_42027_, _42026_, _42010_);
  and (_42029_, _41974_, _41996_);
  and (_42030_, _41978_, _41985_);
  and (_42031_, _42030_, _35118_);
  or (_42033_, _42031_, _42005_);
  and (_42034_, _42033_, _42029_);
  nor (_42035_, _35118_, _34367_);
  and (_42037_, _42001_, _42035_);
  and (_42038_, _42037_, _41988_);
  and (_42039_, _42000_, _41974_);
  and (_42041_, _42039_, _42022_);
  or (_42042_, _42041_, _42038_);
  and (_42043_, _41987_, _41980_);
  and (_42045_, _42043_, _42014_);
  and (_42046_, _42013_, _42020_);
  and (_42047_, _42046_, _42043_);
  or (_42049_, _42047_, _42045_);
  and (_42050_, _42001_, _41996_);
  and (_42052_, _42043_, _42050_);
  or (_42053_, _42052_, _42049_);
  or (_42054_, _42053_, _42042_);
  or (_42055_, _42054_, _42034_);
  or (_42057_, _42055_, _42027_);
  and (_42058_, _42013_, _42035_);
  nor (_42059_, _42058_, _42016_);
  and (_42061_, _41987_, _33856_);
  not (_42062_, _42061_);
  nor (_42063_, _42062_, _42059_);
  not (_42065_, _42063_);
  and (_42066_, _42000_, _41990_);
  and (_42067_, _42043_, _42066_);
  and (_42069_, _41976_, _34367_);
  and (_42070_, _42013_, _42069_);
  and (_42071_, _42070_, _42043_);
  nor (_42073_, _42071_, _42067_);
  and (_42074_, _42073_, _42065_);
  and (_42075_, _42069_, _41974_);
  and (_42077_, _42043_, _42075_);
  or (_42078_, _42020_, _42035_);
  and (_42079_, _42043_, _41990_);
  and (_42081_, _42079_, _42078_);
  and (_42082_, _41974_, _34367_);
  and (_42084_, _42017_, _42082_);
  or (_42085_, _42084_, _42081_);
  nor (_42086_, _42085_, _42077_);
  nand (_42087_, _42086_, _42074_);
  or (_42089_, _42087_, _42057_);
  or (_42090_, _42089_, _41994_);
  and (_42091_, _42090_, _33224_);
  not (_42093_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42094_, _33202_, _14684_);
  and (_42095_, _42094_, _36133_);
  nor (_42097_, _42095_, _42093_);
  or (_42098_, _42097_, rst);
  or (_04363_, _42098_, _42091_);
  nand (_42100_, _34857_, _33158_);
  or (_42101_, _33158_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42102_, _42101_, _43998_);
  and (_04366_, _42102_, _42100_);
  and (_42104_, \oc8051_top_1.oc8051_sfr1.wait_data , _43998_);
  and (_42105_, _42104_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_42107_, _36992_, _36742_);
  and (_42108_, _36394_, _35839_);
  and (_42109_, _35937_, _35335_);
  and (_42111_, _35828_, _35915_);
  or (_42112_, _42111_, _42109_);
  or (_42114_, _42112_, _42108_);
  or (_42115_, _42114_, _42107_);
  not (_42116_, _36514_);
  and (_42117_, _37179_, _36525_);
  and (_42119_, _35839_, _35411_);
  and (_42120_, _42119_, _35161_);
  or (_42121_, _42120_, _42117_);
  or (_42123_, _42121_, _42116_);
  or (_42124_, _42123_, _42115_);
  and (_42125_, _42124_, _41969_);
  or (_04369_, _42125_, _42105_);
  and (_42127_, _35937_, _35422_);
  or (_42128_, _42127_, _35861_);
  and (_42130_, _35183_, _34411_);
  nor (_42131_, _35172_, _33649_);
  and (_42132_, _42131_, _42130_);
  and (_42134_, _42132_, _35302_);
  or (_42135_, _42134_, _35400_);
  and (_42136_, _36253_, _33899_);
  and (_42138_, _42136_, _36394_);
  or (_42139_, _42138_, _42135_);
  or (_42140_, _42139_, _42128_);
  and (_42142_, _42140_, _33213_);
  and (_42143_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42144_, \oc8051_top_1.oc8051_decoder1.state [0], _14684_);
  and (_42145_, _42144_, _42093_);
  not (_42146_, _37210_);
  and (_42147_, _42146_, _42145_);
  or (_42148_, _42147_, _42143_);
  or (_42149_, _42148_, _42142_);
  and (_04372_, _42149_, _43998_);
  and (_42150_, _42104_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nor (_42151_, _36557_, _35915_);
  nor (_42152_, _42151_, _33649_);
  nor (_42153_, _35161_, _33649_);
  and (_42154_, _42153_, _35498_);
  nor (_42155_, _42154_, _42152_);
  nand (_42156_, _42155_, _35520_);
  and (_42157_, _37179_, _36557_);
  nor (_42158_, _42151_, _36889_);
  or (_42159_, _42158_, _42157_);
  and (_42160_, _42136_, _36481_);
  or (_42161_, _42160_, _42159_);
  and (_42162_, _37179_, _36862_);
  and (_42163_, _36720_, _36307_);
  or (_42164_, _42163_, _42128_);
  or (_42165_, _42164_, _42162_);
  or (_42166_, _42165_, _42161_);
  or (_42167_, _42166_, _42156_);
  and (_42168_, _42167_, _41969_);
  or (_04375_, _42168_, _42150_);
  and (_42169_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42170_, _36285_, _33213_);
  or (_42171_, _42170_, _42169_);
  or (_42172_, _42171_, _42147_);
  and (_04378_, _42172_, _43998_);
  not (_42173_, _41971_);
  and (_42174_, _42173_, _36525_);
  nor (_42175_, _42174_, _42119_);
  not (_42176_, _42175_);
  and (_42177_, _42176_, _42145_);
  or (_42178_, _42177_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42179_, _36264_, _35818_);
  and (_42180_, _35959_, _35498_);
  nor (_42181_, _42180_, _42179_);
  nor (_42182_, _42181_, _35161_);
  not (_42183_, _33169_);
  and (_42184_, _42120_, _42183_);
  or (_42185_, _42184_, _42182_);
  and (_42186_, _42185_, _36133_);
  or (_42187_, _42186_, _42178_);
  or (_42188_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _14684_);
  and (_42189_, _42188_, _43998_);
  and (_04381_, _42189_, _42187_);
  and (_42190_, _42104_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_42191_, _42160_, _42111_);
  and (_42192_, _36481_, _34160_);
  and (_42193_, _36394_, _34160_);
  or (_42194_, _42193_, _42192_);
  or (_42195_, _42194_, _42191_);
  or (_42196_, _36633_, _35861_);
  or (_42197_, _36912_, _36731_);
  or (_42198_, _42197_, _42196_);
  and (_42199_, _42153_, _35389_);
  or (_42200_, _42154_, _42199_);
  or (_42201_, _42134_, _36405_);
  or (_42202_, _42201_, _42200_);
  or (_42203_, _42202_, _42198_);
  or (_42204_, _42203_, _42195_);
  and (_42205_, _42204_, _41969_);
  or (_04384_, _42205_, _42190_);
  and (_42206_, _42104_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nand (_42207_, _37179_, _36666_);
  nand (_42208_, _42207_, _36786_);
  not (_42209_, _42155_);
  and (_42210_, _35466_, _35389_);
  and (_42211_, _35992_, _42130_);
  or (_42212_, _42211_, _35292_);
  or (_42213_, _42212_, _42210_);
  or (_42214_, _42213_, _42209_);
  or (_42215_, _42214_, _42208_);
  nor (_42216_, _36829_, _35509_);
  nand (_42217_, _42216_, _36699_);
  and (_42218_, _42136_, _35281_);
  or (_42219_, _42218_, _42138_);
  and (_42220_, _42131_, _35270_);
  or (_42221_, _42220_, _42132_);
  and (_42222_, _35839_, _34911_);
  or (_42223_, _42222_, _42221_);
  or (_42224_, _42223_, _42219_);
  or (_42225_, _42224_, _42217_);
  or (_42226_, _42225_, _42161_);
  or (_42227_, _42226_, _42215_);
  and (_42228_, _42227_, _41969_);
  or (_04387_, _42228_, _42206_);
  and (_42229_, _42136_, _34932_);
  and (_42230_, _34932_, _34160_);
  and (_42231_, _42153_, _35411_);
  or (_42232_, _42231_, _42230_);
  or (_42233_, _42232_, _42229_);
  and (_42234_, _34932_, _36307_);
  or (_42235_, _42234_, _35433_);
  or (_42236_, _42235_, _42233_);
  and (_42237_, _42136_, _35422_);
  or (_42238_, _42237_, _42236_);
  and (_42239_, _42238_, _33213_);
  nand (_42240_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_42241_, _42240_, _37271_);
  or (_42242_, _42241_, _42239_);
  and (_04390_, _42242_, _43998_);
  or (_42243_, _36905_, _36405_);
  or (_42244_, _42158_, _36851_);
  or (_42245_, _42244_, _42243_);
  and (_42246_, _35259_, _35172_);
  and (_42247_, _42246_, _36274_);
  or (_42248_, _42247_, _36644_);
  and (_42249_, _36481_, _35959_);
  or (_42250_, _42249_, _36775_);
  or (_42251_, _42250_, _42248_);
  nand (_42252_, _36753_, _36296_);
  or (_42253_, _42252_, _42251_);
  or (_42254_, _42253_, _42245_);
  and (_42255_, _42153_, _35259_);
  or (_42256_, _42255_, _36318_);
  and (_42257_, _42179_, _35172_);
  and (_42258_, _42131_, _35411_);
  or (_42259_, _42258_, _42257_);
  or (_42260_, _42259_, _42135_);
  or (_42261_, _42260_, _42256_);
  and (_42262_, _42246_, _34160_);
  or (_42263_, _42262_, _35509_);
  or (_42264_, _42263_, _36579_);
  or (_42265_, _36361_, _35346_);
  or (_42266_, _42265_, _42264_);
  or (_42267_, _42266_, _42261_);
  or (_42268_, _42267_, _42209_);
  or (_42269_, _42268_, _42254_);
  and (_42270_, _42269_, _33213_);
  and (_42271_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42272_, _37058_, _36144_);
  or (_42273_, _42249_, _42257_);
  and (_42274_, _42273_, _36144_);
  or (_42275_, _42274_, _42147_);
  or (_42276_, _42275_, _42272_);
  or (_42277_, _42276_, _42271_);
  or (_42278_, _42277_, _42270_);
  and (_04393_, _42278_, _43998_);
  nor (_04453_, _36187_, rst);
  nor (_04455_, _37124_, rst);
  nand (_04458_, _42176_, _41969_);
  nand (_42279_, _41969_, _42119_);
  not (_42280_, _35937_);
  or (_42281_, _41970_, _42280_);
  and (_04461_, _42281_, _42279_);
  or (_42282_, _41998_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42283_, _42282_, _42084_);
  or (_42284_, _42283_, _41984_);
  and (_42285_, _42284_, _42095_);
  nor (_42286_, _42094_, _36133_);
  or (_42287_, _42286_, rst);
  or (_04464_, _42287_, _42285_);
  nand (_42288_, _35741_, _33158_);
  or (_42289_, _33158_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42290_, _42289_, _43998_);
  and (_04467_, _42290_, _42288_);
  nand (_42291_, _33856_, _33158_);
  or (_42292_, _33158_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42293_, _42292_, _43998_);
  and (_04470_, _42293_, _42291_);
  nand (_42294_, _34095_, _33158_);
  or (_42295_, _33158_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42296_, _42295_, _43998_);
  and (_04473_, _42296_, _42294_);
  nand (_42297_, _33605_, _33158_);
  or (_42298_, _33158_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42299_, _42298_, _43998_);
  and (_04476_, _42299_, _42297_);
  nand (_42300_, _41976_, _33158_);
  or (_42301_, _33158_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42302_, _42301_, _43998_);
  and (_04479_, _42302_, _42300_);
  nand (_42303_, _34367_, _33158_);
  or (_42304_, _33158_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42305_, _42304_, _43998_);
  and (_04482_, _42305_, _42303_);
  nand (_42306_, _34617_, _33158_);
  or (_42307_, _33158_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42308_, _42307_, _43998_);
  and (_04485_, _42308_, _42306_);
  or (_42309_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _14684_);
  and (_42310_, _42309_, _42178_);
  and (_42311_, _42136_, _36666_);
  or (_42312_, _42311_, _42127_);
  and (_42313_, _35466_, _35205_);
  nor (_42314_, _42220_, _42313_);
  not (_42315_, _42314_);
  or (_42316_, _42315_, _42312_);
  and (_42317_, _42153_, _35205_);
  or (_42318_, _42317_, _42234_);
  or (_42319_, _35498_, _35915_);
  and (_42320_, _42319_, _37179_);
  or (_42321_, _42320_, _42318_);
  or (_42322_, _42321_, _42316_);
  or (_42323_, _35433_, _35292_);
  or (_42324_, _36535_, _36035_);
  or (_42325_, _42324_, _42323_);
  and (_42326_, _42131_, _35205_);
  and (_42327_, _42131_, _36013_);
  or (_42328_, _42327_, _42326_);
  or (_42329_, _42328_, _35861_);
  or (_42330_, _42329_, _42233_);
  or (_42331_, _42330_, _42325_);
  and (_42332_, _42136_, _35215_);
  and (_42333_, _37179_, _35872_);
  and (_42334_, _36013_, _35172_);
  and (_42335_, _42334_, _37179_);
  or (_42336_, _42335_, _42333_);
  or (_42337_, _42336_, _42332_);
  or (_42338_, _42218_, _42117_);
  or (_42339_, _42237_, _42222_);
  or (_42340_, _42339_, _42338_);
  or (_42341_, _42340_, _42337_);
  or (_42342_, _42341_, _42331_);
  or (_42343_, _42342_, _42322_);
  and (_42344_, _42343_, _33213_);
  or (_42345_, _42344_, _42310_);
  and (_28812_, _42345_, _43998_);
  and (_42346_, _42104_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_42347_, _35194_, _35161_);
  and (_42348_, _35959_, _42347_);
  nor (_42349_, _42348_, _42221_);
  nand (_42350_, _42349_, _36416_);
  and (_42351_, _34661_, _34421_);
  and (_42352_, _42153_, _42351_);
  and (_42353_, _42352_, _35302_);
  nor (_42354_, _42353_, _35487_);
  not (_42355_, _42354_);
  or (_42356_, _42355_, _42312_);
  or (_42357_, _42356_, _42350_);
  or (_42358_, _42213_, _42121_);
  or (_42359_, _42358_, _42357_);
  not (_42360_, _35281_);
  nand (_42361_, _42360_, _35226_);
  or (_42362_, _42361_, _36862_);
  and (_42363_, _42362_, _37179_);
  or (_42364_, _42363_, _42359_);
  and (_42365_, _42364_, _41969_);
  or (_28814_, _42365_, _42346_);
  or (_42366_, _42265_, _42259_);
  or (_42367_, _42366_, _42254_);
  and (_42368_, _42367_, _33213_);
  and (_42369_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42370_, _42369_, _42276_);
  or (_42371_, _42370_, _42368_);
  and (_28816_, _42371_, _43998_);
  and (_42372_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42373_, _42372_, _42275_);
  and (_42374_, _36818_, _35161_);
  or (_42375_, _42374_, _35400_);
  or (_42376_, _42375_, _42264_);
  or (_42377_, _42376_, _42182_);
  and (_42378_, _42377_, _33213_);
  or (_42379_, _42378_, _42373_);
  and (_28818_, _42379_, _43998_);
  or (_42380_, _37200_, _42119_);
  and (_42381_, _42229_, _35172_);
  or (_42382_, _42381_, _42332_);
  or (_42383_, _42382_, _42380_);
  or (_42384_, _42231_, _35433_);
  or (_42385_, _42384_, _35237_);
  or (_42386_, _42385_, _42182_);
  or (_42387_, _42386_, _42383_);
  and (_42388_, _42136_, _36720_);
  or (_42389_, _42388_, _42117_);
  or (_42390_, _42335_, _37189_);
  or (_42391_, _42390_, _42320_);
  or (_42392_, _42391_, _42389_);
  and (_42393_, _37179_, _36394_);
  or (_42394_, _42339_, _42393_);
  or (_42395_, _42394_, _42318_);
  and (_42396_, _35872_, _35839_);
  and (_42397_, _35959_, _35215_);
  and (_42398_, _42334_, _36274_);
  or (_42399_, _42398_, _42397_);
  or (_42400_, _42399_, _42396_);
  and (_42401_, _37179_, _42347_);
  or (_42402_, _42262_, _42255_);
  or (_42403_, _42402_, _42401_);
  and (_42404_, _42229_, _35161_);
  or (_42405_, _42404_, _42333_);
  or (_42406_, _42405_, _42403_);
  or (_42407_, _42406_, _42400_);
  or (_42408_, _42407_, _42395_);
  or (_42409_, _42408_, _42392_);
  or (_42410_, _42409_, _42387_);
  and (_42411_, _42410_, _33213_);
  and (_42412_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42413_, _42177_, _37282_);
  or (_42414_, _42413_, _42412_);
  or (_42415_, _42414_, _42411_);
  and (_28820_, _42415_, _43998_);
  or (_42416_, _42247_, _36361_);
  or (_42417_, _42416_, _35894_);
  or (_42418_, _42417_, _36897_);
  or (_42419_, _42127_, _37200_);
  or (_42420_, _34150_, _36307_);
  and (_42421_, _42420_, _42334_);
  and (_42422_, _35839_, _42347_);
  or (_42423_, _42422_, _42421_);
  or (_42424_, _42423_, _42419_);
  or (_42425_, _42424_, _42385_);
  or (_42426_, _42425_, _42418_);
  or (_42427_, _42395_, _42392_);
  or (_42428_, _42427_, _42426_);
  and (_42429_, _42428_, _33213_);
  and (_42430_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42431_, _42430_, _42413_);
  or (_42432_, _42431_, _42429_);
  and (_28822_, _42432_, _43998_);
  and (_42433_, _42104_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_42434_, _35839_, _35915_);
  and (_42435_, _35839_, _35498_);
  and (_42436_, _42435_, _35172_);
  or (_42437_, _42436_, _42434_);
  not (_42438_, _39811_);
  or (_42439_, _42237_, _42438_);
  and (_42440_, _42420_, _36470_);
  or (_42441_, _42440_, _42381_);
  and (_42442_, _35839_, _36720_);
  and (_42443_, _36470_, _35839_);
  or (_42444_, _42443_, _42442_);
  or (_42445_, _42444_, _42441_);
  or (_42446_, _42445_, _42439_);
  or (_42447_, _42446_, _42437_);
  or (_42448_, _42243_, _42200_);
  or (_42449_, _42231_, _42134_);
  and (_42450_, _37179_, _35915_);
  or (_42451_, _42450_, _42160_);
  or (_42452_, _42451_, _42449_);
  or (_42453_, _42452_, _42448_);
  or (_42454_, _36231_, _35433_);
  or (_42455_, _42454_, _42194_);
  not (_42456_, _39809_);
  or (_42457_, _42196_, _42456_);
  or (_42458_, _42457_, _42455_);
  or (_42459_, _42458_, _42453_);
  or (_42460_, _42459_, _42447_);
  and (_42461_, _42460_, _41969_);
  or (_28824_, _42461_, _42433_);
  or (_42462_, _42211_, _42210_);
  or (_42463_, _42404_, _42396_);
  or (_42464_, _42463_, _42462_);
  or (_42465_, _42464_, _42208_);
  or (_42466_, _42465_, _42383_);
  or (_42467_, _42443_, _42450_);
  or (_42468_, _42436_, _42318_);
  or (_42469_, _42468_, _42467_);
  or (_42470_, _42132_, _35861_);
  or (_42471_, _42138_, _36677_);
  or (_42472_, _42471_, _42470_);
  nand (_42473_, _36372_, _35248_);
  or (_42474_, _42473_, _42472_);
  or (_42475_, _42474_, _42469_);
  or (_42476_, _42475_, _42466_);
  and (_42477_, _42476_, _41969_);
  and (_42478_, _42104_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_42479_, _33169_, _43998_);
  and (_42480_, _42479_, _37200_);
  or (_42481_, _42480_, _42478_);
  or (_28826_, _42481_, _42477_);
  not (_42482_, _36350_);
  nor (_42483_, _42332_, _36361_);
  and (_42484_, _42483_, _42482_);
  or (_42485_, _42237_, _42163_);
  and (_42486_, _35839_, _34932_);
  or (_42487_, _42317_, _42313_);
  or (_42488_, _42487_, _42486_);
  or (_42489_, _42488_, _42485_);
  nor (_42490_, _42138_, _39808_);
  nand (_42491_, _42490_, _35444_);
  nor (_42492_, _42491_, _42489_);
  nand (_42493_, _42492_, _42484_);
  and (_42494_, _35828_, _36720_);
  or (_42495_, _42494_, _42335_);
  or (_42496_, _42449_, _42389_);
  or (_42497_, _42496_, _42495_);
  or (_42498_, _42497_, _42161_);
  or (_42499_, _42498_, _42156_);
  or (_42500_, _42499_, _42493_);
  and (_42501_, _42500_, _33213_);
  and (_42502_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42503_, _42502_, _37249_);
  or (_42504_, _42503_, _42501_);
  and (_28828_, _42504_, _43998_);
  not (_42505_, _42483_);
  or (_42506_, _42505_, _42451_);
  or (_42507_, _42506_, _42495_);
  or (_42508_, _35509_, _35400_);
  or (_42509_, _42508_, _42435_);
  or (_42510_, _42509_, _42487_);
  or (_42511_, _42201_, _42438_);
  or (_42512_, _42511_, _42510_);
  or (_42513_, _42159_, _42209_);
  or (_42514_, _42513_, _42512_);
  or (_42515_, _42514_, _42507_);
  and (_42516_, _42515_, _33213_);
  and (_42517_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42518_, _42517_, _37260_);
  or (_42519_, _42518_, _42516_);
  and (_28830_, _42519_, _43998_);
  and (_42520_, _42104_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_42521_, _42108_, _36912_);
  nand (_42522_, _42521_, _39809_);
  not (_42523_, _35818_);
  or (_42524_, _35839_, _42523_);
  and (_42525_, _42524_, _36720_);
  or (_42526_, _42525_, _42467_);
  or (_42527_, _42526_, _42522_);
  or (_42528_, _42439_, _42236_);
  or (_42529_, _42528_, _42437_);
  or (_42530_, _42529_, _42527_);
  and (_42531_, _42530_, _41969_);
  or (_28833_, _42531_, _42520_);
  nor (_38734_, _34857_, rst);
  nor (_38736_, _39940_, rst);
  nor (_42532_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_42533_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_42534_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42535_, _42534_, _42533_);
  and (_42536_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_42537_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_42538_, _42537_, _42536_);
  and (_42539_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_42540_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_42541_, _42540_, _42539_);
  and (_42542_, _42541_, _42538_);
  and (_42543_, _42542_, _42535_);
  and (_42544_, _42543_, _33682_);
  nor (_42545_, _42544_, _42532_);
  nor (_42546_, _42545_, _39864_);
  nor (_42547_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nor (_42548_, _42547_, _42546_);
  and (_38737_, _42548_, _43998_);
  nor (_38749_, _35741_, rst);
  nor (_38750_, _33856_, rst);
  nor (_38751_, _34095_, rst);
  nor (_38752_, _33605_, rst);
  and (_38753_, _35118_, _43998_);
  nor (_38754_, _34367_, rst);
  nor (_38755_, _34617_, rst);
  nor (_38757_, _39880_, rst);
  nor (_38758_, _40095_, rst);
  nor (_38759_, _40023_, rst);
  nor (_38760_, _39974_, rst);
  nor (_38761_, _40149_, rst);
  nor (_38763_, _40059_, rst);
  nor (_38764_, _40201_, rst);
  nor (_42549_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_42550_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_42551_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42552_, _42551_, _42550_);
  and (_42553_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_42554_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_42555_, _42554_, _42553_);
  and (_42556_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_42557_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_42558_, _42557_, _42556_);
  and (_42559_, _42558_, _42555_);
  and (_42560_, _42559_, _42552_);
  and (_42561_, _42560_, _33682_);
  nor (_42562_, _42561_, _42549_);
  nor (_42563_, _42562_, _39864_);
  nor (_42564_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_42565_, _42564_, _42563_);
  and (_38765_, _42565_, _43998_);
  nor (_42566_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_42567_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_42568_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_42569_, _42568_, _42567_);
  and (_42570_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42571_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42572_, _42571_, _42570_);
  and (_42573_, _42572_, _42569_);
  and (_42574_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_42575_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42576_, _42575_, _42574_);
  and (_42577_, _42576_, _42573_);
  and (_42578_, _42577_, _33682_);
  nor (_42579_, _42578_, _42566_);
  nor (_42580_, _42579_, _39864_);
  nor (_42581_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nor (_42582_, _42581_, _42580_);
  and (_38766_, _42582_, _43998_);
  nor (_42583_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_42584_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_42585_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42586_, _42585_, _42584_);
  and (_42587_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_42588_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_42589_, _42588_, _42587_);
  and (_42590_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_42591_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_42592_, _42591_, _42590_);
  and (_42593_, _42592_, _42589_);
  and (_42594_, _42593_, _42586_);
  and (_42595_, _42594_, _33682_);
  nor (_42596_, _42595_, _42583_);
  nor (_42597_, _42596_, _39864_);
  nor (_42598_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nor (_42599_, _42598_, _42597_);
  and (_38767_, _42599_, _43998_);
  nor (_42600_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_42601_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_42602_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_42603_, _42602_, _42601_);
  and (_42604_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42605_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_42606_, _42605_, _42604_);
  and (_42607_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_42608_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42609_, _42608_, _42607_);
  and (_42610_, _42609_, _42606_);
  and (_42611_, _42610_, _42603_);
  and (_42612_, _42611_, _33682_);
  nor (_42613_, _42612_, _42600_);
  nor (_42614_, _42613_, _39864_);
  nor (_42615_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  nor (_42616_, _42615_, _42614_);
  and (_38769_, _42616_, _43998_);
  nor (_42617_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_42618_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_42619_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_42620_, _42619_, _42618_);
  and (_42621_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42622_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42623_, _42622_, _42621_);
  and (_42624_, _42623_, _42620_);
  and (_42625_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_42626_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42627_, _42626_, _42625_);
  and (_42628_, _42627_, _42624_);
  and (_42629_, _42628_, _33682_);
  nor (_42630_, _42629_, _42617_);
  nor (_42631_, _42630_, _39864_);
  nor (_42632_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  nor (_42633_, _42632_, _42631_);
  and (_38770_, _42633_, _43998_);
  nor (_42634_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_42635_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_42636_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42637_, _42636_, _42635_);
  and (_42638_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42639_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_42640_, _42639_, _42638_);
  and (_42641_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_42642_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_42643_, _42642_, _42641_);
  and (_42644_, _42643_, _42640_);
  and (_42645_, _42644_, _42637_);
  and (_42646_, _42645_, _33682_);
  nor (_42647_, _42646_, _42634_);
  nor (_42648_, _42647_, _39864_);
  nor (_42649_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  nor (_42650_, _42649_, _42648_);
  and (_38771_, _42650_, _43998_);
  nor (_42651_, _33682_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_42652_, _33343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42653_, _33517_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42654_, _42653_, _42652_);
  and (_42655_, _33387_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_42656_, _33431_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_42657_, _42656_, _42655_);
  and (_42658_, _33463_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_42659_, _33322_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42660_, _42659_, _42658_);
  and (_42661_, _42660_, _42657_);
  and (_42662_, _42661_, _42654_);
  and (_42663_, _42662_, _33682_);
  nor (_42664_, _42663_, _42651_);
  nor (_42665_, _42664_, _39864_);
  nor (_42666_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  nor (_42667_, _42666_, _42665_);
  and (_38772_, _42667_, _43998_);
  and (_42668_, _33224_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_42669_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_42670_, _42668_, _38540_);
  and (_42671_, _42670_, _43998_);
  and (_38798_, _42671_, _42669_);
  not (_42672_, _42668_);
  or (_42673_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _42668_, _43998_);
  and (_42674_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _43998_);
  or (_42675_, _42674_, _00000_);
  and (_38799_, _42675_, _42673_);
  nor (_38837_, _39945_, rst);
  and (_38839_, _40154_, _43998_);
  nor (_38840_, _39922_, rst);
  nor (_42676_, _39983_, _23647_);
  and (_42677_, _39983_, _23647_);
  nor (_42678_, _42677_, _42676_);
  nor (_42679_, _40207_, _38944_);
  and (_42680_, _40207_, _38944_);
  nor (_42681_, _42680_, _42679_);
  and (_42682_, _39945_, _27812_);
  nor (_42683_, _39945_, _27812_);
  or (_42684_, _42683_, _42682_);
  not (_42685_, _42684_);
  and (_42686_, _42685_, _42681_);
  nor (_42687_, _40068_, _23965_);
  and (_42688_, _40068_, _23965_);
  nor (_42689_, _42688_, _42687_);
  and (_42690_, _40158_, _23811_);
  nor (_42691_, _40158_, _23811_);
  nor (_42692_, _42691_, _42690_);
  and (_42693_, _42692_, _42689_);
  and (_42694_, _42693_, _42686_);
  and (_42695_, _42694_, _42678_);
  nor (_42696_, _40119_, _29894_);
  and (_42697_, _40119_, _29894_);
  or (_42698_, _42697_, _42696_);
  nor (_42699_, _42698_, _39466_);
  or (_42700_, _39885_, _24085_);
  nand (_42701_, _39885_, _24085_);
  and (_42702_, _42701_, _42700_);
  or (_42703_, _40028_, _24352_);
  nand (_42704_, _40028_, _24352_);
  and (_42705_, _42704_, _42703_);
  nor (_42706_, _42705_, _42702_);
  and (_42707_, _42706_, _42699_);
  and (_42708_, _42707_, _42695_);
  nor (_42709_, _23317_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_42710_, _42709_, _42708_);
  nor (_42711_, _36514_, _42144_);
  and (_42712_, _33006_, _27209_);
  and (_42713_, _42712_, _42711_);
  and (_42714_, _42713_, _42695_);
  nand (_42715_, _30112_, _25541_);
  nor (_42716_, _42715_, _30807_);
  and (_42717_, _42716_, _31960_);
  and (_42718_, _42717_, _32417_);
  and (_42719_, _39888_, _39899_);
  nor (_42720_, _42719_, _42144_);
  nor (_42721_, _42720_, _37003_);
  and (_42722_, _42721_, _28031_);
  and (_42723_, _42722_, _42718_);
  and (_42724_, _42723_, _25706_);
  and (_42725_, _42711_, _25410_);
  or (_42726_, _42711_, _34411_);
  and (_42727_, _42726_, _37003_);
  and (_42728_, _42727_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_42729_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_42730_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_42731_, _42730_, _42729_);
  nor (_42732_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_42733_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_42734_, _42733_, _42732_);
  and (_42735_, _42734_, _42731_);
  and (_42736_, _42735_, _36166_);
  or (_42737_, _42736_, _42728_);
  or (_42738_, _42737_, _42725_);
  nor (_42739_, _42738_, _42724_);
  not (_42740_, _42199_);
  nor (_42741_, _42388_, _36633_);
  and (_42742_, _42741_, _42740_);
  or (_42743_, _36470_, _35872_);
  or (_42744_, _42743_, _35215_);
  nand (_42745_, _42744_, _35937_);
  and (_42746_, _42745_, _42354_);
  nand (_42747_, _42746_, _42742_);
  nand (_42748_, _42747_, _42739_);
  nor (_42749_, _42109_, _42396_);
  nand (_42750_, _36992_, _35161_);
  and (_42751_, _42750_, _37069_);
  or (_42752_, _42751_, _42739_);
  and (_42753_, _42752_, _42749_);
  and (_42754_, _42753_, _42748_);
  or (_42755_, _42754_, _37014_);
  nor (_42756_, _42181_, _33169_);
  nor (_42757_, _42756_, _36111_);
  and (_42758_, _42757_, _42755_);
  or (_42759_, _38951_, _38935_);
  or (_42760_, _42759_, _38904_);
  and (_42761_, _42760_, _42727_);
  or (_42762_, _39048_, _39045_);
  nor (_42763_, _42762_, _39053_);
  nand (_42764_, _42763_, _39094_);
  and (_42765_, _42764_, _36166_);
  or (_42766_, _42765_, _42761_);
  or (_42767_, _42766_, _42758_);
  or (_42768_, _42767_, _42714_);
  nor (_42769_, _42768_, _42710_);
  nor (_42770_, _36122_, rst);
  and (_38844_, _42770_, _42769_);
  and (_38845_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _43998_);
  and (_38846_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _43998_);
  nor (_42771_, _33376_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_42772_, _42771_, _39864_);
  nor (_42773_, _42772_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_42774_, _42773_);
  and (_42775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_42776_, _42775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_42777_, _42776_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_42778_, _42777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_42779_, _42778_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_42780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_42781_, _42780_, _42779_);
  and (_42782_, _42781_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_42783_, _42782_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_42784_, _42783_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_42785_, _42784_, _42774_);
  and (_42786_, _42785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_42787_, _42786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_42788_, _42787_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_42789_, _42708_, _27812_);
  and (_42790_, _42789_, _27165_);
  and (_42791_, _42720_, _33006_);
  and (_42792_, _42791_, _27209_);
  and (_42793_, _42792_, _42695_);
  and (_42794_, _37003_, _34411_);
  and (_42795_, _42760_, _42794_);
  not (_42796_, _36111_);
  nand (_42797_, _42755_, _42796_);
  nor (_42798_, _42797_, _42756_);
  and (_42799_, _35937_, _35270_);
  and (_42800_, _42799_, _36144_);
  and (_42801_, _42764_, _42800_);
  or (_42802_, _42801_, _42798_);
  or (_42803_, _42802_, _42795_);
  or (_42804_, _42803_, _42793_);
  nor (_42805_, _42804_, _42790_);
  and (_42806_, _42787_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_42807_, _42806_, _42805_);
  and (_42808_, _42807_, _42788_);
  and (_42809_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_42810_, _42809_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_42811_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_42812_, _42811_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_42813_, _42812_, _42810_);
  and (_42814_, _42813_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_42815_, _42814_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_42816_, _42815_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_42817_, _42816_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_42818_, _42817_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_42819_, _42818_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_42820_, _42819_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_42821_, _42820_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_42822_, _42821_, _38540_);
  or (_42823_, _42821_, _38540_);
  and (_42824_, _42823_, _42822_);
  and (_42825_, _35937_, _42183_);
  and (_42826_, _42825_, _34932_);
  and (_42827_, _42354_, _42719_);
  not (_42828_, _36992_);
  and (_42829_, _42749_, _42828_);
  and (_42830_, _42829_, _42742_);
  and (_42831_, _42830_, _42827_);
  nor (_42832_, _42831_, _37014_);
  nor (_42833_, _42832_, _42826_);
  and (_42834_, _42827_, _42741_);
  nor (_42835_, _42834_, _37014_);
  not (_42836_, _42835_);
  and (_42837_, _42180_, _42183_);
  nor (_42838_, _42826_, _42837_);
  and (_42839_, _42838_, _36981_);
  and (_42840_, _42839_, _42836_);
  and (_42841_, _36144_, _42396_);
  nor (_42842_, _42841_, _42756_);
  not (_42843_, _42842_);
  and (_42844_, _42843_, _42840_);
  and (_42845_, _42844_, _42833_);
  and (_42846_, _42845_, _42824_);
  nor (_42847_, _36981_, _27132_);
  not (_42848_, _42841_);
  nor (_42849_, _42848_, _38591_);
  not (_42850_, _42179_);
  and (_42851_, _36557_, _35959_);
  nor (_42852_, _42851_, _42249_);
  and (_42853_, _42852_, _42850_);
  or (_42854_, _42853_, _33169_);
  nor (_42855_, _35785_, _33899_);
  and (_42856_, _42855_, _35818_);
  nand (_42857_, _42856_, _35872_);
  or (_42858_, _37014_, _42857_);
  and (_42859_, _42858_, _42854_);
  not (_42860_, _39887_);
  and (_42861_, _42852_, _42860_);
  and (_42862_, _42861_, _39899_);
  or (_42863_, _42862_, _33169_);
  nor (_42864_, _42835_, _36970_);
  and (_42865_, _42864_, _42863_);
  nor (_42866_, _39887_, _37047_);
  nor (_42867_, _42866_, _33169_);
  nor (_42868_, _42867_, _42832_);
  and (_42869_, _42868_, _42865_);
  and (_42870_, _42869_, _42859_);
  and (_42871_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_42872_, _42837_, _39941_);
  or (_42873_, _42872_, _42871_);
  or (_42874_, _42873_, _42849_);
  or (_42875_, _42874_, _42847_);
  or (_42876_, _42875_, _42846_);
  not (_42877_, _36122_);
  and (_42878_, _36448_, _42183_);
  nor (_42879_, _42837_, _42878_);
  and (_42880_, _42879_, _42877_);
  and (_42881_, _42880_, _42836_);
  and (_42882_, _42881_, _39941_);
  not (_42883_, _42881_);
  and (_42884_, _42883_, _42548_);
  nor (_42885_, _42884_, _42882_);
  not (_42886_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_42887_, _42885_, _42886_);
  not (_42888_, _42887_);
  and (_42889_, _42885_, _42886_);
  nor (_42890_, _42889_, _42887_);
  not (_42891_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_42892_, _42840_, _40201_);
  nor (_42893_, _42840_, _42667_);
  or (_42894_, _42893_, _42892_);
  nor (_42895_, _42894_, _42891_);
  and (_42896_, _42894_, _42891_);
  nor (_42897_, _42896_, _42895_);
  not (_42898_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_42899_, _42840_, _40059_);
  nor (_42900_, _42840_, _42650_);
  or (_42901_, _42900_, _42899_);
  nor (_42902_, _42901_, _42898_);
  and (_42903_, _42901_, _42898_);
  not (_42904_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_42905_, _42840_, _40149_);
  nor (_42906_, _42840_, _42633_);
  or (_42907_, _42906_, _42905_);
  or (_42908_, _42907_, _42904_);
  not (_42909_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_42910_, _42840_, _39974_);
  nor (_42911_, _42840_, _42616_);
  or (_42912_, _42911_, _42910_);
  nor (_42913_, _42912_, _42909_);
  and (_42914_, _42912_, _42909_);
  not (_42915_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_42916_, _42840_, _40023_);
  nor (_42917_, _42840_, _42599_);
  or (_42918_, _42917_, _42916_);
  nor (_42919_, _42918_, _42915_);
  not (_42920_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_42921_, _42840_, _40095_);
  nor (_42922_, _42840_, _42582_);
  or (_42923_, _42922_, _42921_);
  nor (_42924_, _42923_, _42920_);
  not (_42925_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_42926_, _42840_, _39880_);
  nor (_42927_, _42840_, _42565_);
  or (_42928_, _42927_, _42926_);
  nor (_42929_, _42928_, _42925_);
  and (_42930_, _42923_, _42920_);
  nor (_42931_, _42930_, _42924_);
  and (_42932_, _42931_, _42929_);
  nor (_42933_, _42932_, _42924_);
  not (_42934_, _42933_);
  and (_42935_, _42918_, _42915_);
  nor (_42936_, _42935_, _42919_);
  and (_42937_, _42936_, _42934_);
  nor (_42938_, _42937_, _42919_);
  nor (_42939_, _42938_, _42914_);
  or (_42940_, _42939_, _42913_);
  nand (_42941_, _42907_, _42904_);
  and (_42942_, _42941_, _42908_);
  nand (_42943_, _42942_, _42940_);
  and (_42944_, _42943_, _42908_);
  nor (_42945_, _42944_, _42903_);
  or (_42946_, _42945_, _42902_);
  and (_42947_, _42946_, _42897_);
  nor (_42948_, _42947_, _42895_);
  not (_42949_, _42948_);
  nand (_42950_, _42949_, _42890_);
  and (_42951_, _42950_, _42888_);
  and (_42952_, _42951_, _38512_);
  and (_42953_, _42952_, _38518_);
  and (_42954_, _42953_, _38523_);
  and (_42955_, _42954_, _38508_);
  and (_42956_, _42955_, _38529_);
  and (_42957_, _42956_, _38504_);
  and (_42958_, _42957_, _38535_);
  nor (_42959_, _42958_, _42885_);
  not (_42960_, _42885_);
  and (_42961_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_42962_, _42961_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_42963_, _42962_);
  nor (_42964_, _42963_, _42951_);
  and (_42965_, _42964_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_42966_, _42965_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_42967_, _42966_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_42968_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_42969_, _42968_, _42960_);
  nor (_42970_, _42969_, _42959_);
  or (_42971_, _42970_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_42972_, _42970_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_42973_, _42972_, _42971_);
  nor (_42974_, _42844_, _42833_);
  and (_42975_, _42974_, _42973_);
  or (_42976_, _42975_, _42876_);
  and (_42977_, _42976_, _42805_);
  or (_42978_, _42977_, _42808_);
  and (_38847_, _42978_, _43998_);
  and (_42979_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _43998_);
  and (_42980_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_42981_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_42982_, _33213_, _42981_);
  not (_42983_, _42982_);
  not (_42984_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_42985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_42986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_42987_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_42988_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_42989_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_42990_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_42991_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_42992_, _42991_, _42989_);
  and (_42993_, _42992_, _42990_);
  nor (_42994_, _42993_, _42989_);
  nor (_42995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_42996_, _42995_, _42988_);
  not (_42997_, _42996_);
  nor (_42998_, _42997_, _42994_);
  nor (_42999_, _42998_, _42988_);
  not (_43000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_43001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43004_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43005_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43007_, _43006_, _43005_);
  and (_43008_, _43007_, _43004_);
  and (_43009_, _43008_, _43003_);
  and (_43010_, _43009_, _43002_);
  and (_43011_, _43010_, _43001_);
  and (_43012_, _43011_, _43000_);
  and (_43013_, _43012_, _42999_);
  and (_43014_, _43013_, _42987_);
  and (_43015_, _43014_, _42986_);
  and (_43016_, _43015_, _42985_);
  and (_43017_, _43016_, _42984_);
  and (_43018_, _43017_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_43019_, _43017_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_43020_, _43019_, _43018_);
  nor (_43021_, _43016_, _42984_);
  or (_43022_, _43021_, _43017_);
  nor (_43023_, _43015_, _42985_);
  nor (_43024_, _43023_, _43016_);
  not (_43025_, _43024_);
  nor (_43026_, _43014_, _42986_);
  or (_43027_, _43026_, _43015_);
  nor (_43028_, _43013_, _42987_);
  nor (_43029_, _43028_, _43014_);
  not (_43030_, _43029_);
  and (_43031_, _43011_, _42999_);
  nor (_43032_, _43031_, _43000_);
  nor (_43033_, _43032_, _43013_);
  not (_43034_, _43033_);
  and (_43035_, _43010_, _42999_);
  nor (_43036_, _43035_, _43001_);
  nor (_43037_, _43036_, _43031_);
  not (_43038_, _43037_);
  and (_43039_, _42999_, _43009_);
  and (_43040_, _42999_, _43007_);
  and (_43041_, _43040_, _43004_);
  nor (_43042_, _43041_, _43003_);
  or (_43043_, _43042_, _43039_);
  nor (_43044_, _43040_, _43004_);
  or (_43045_, _43044_, _43041_);
  and (_43046_, _42999_, _43006_);
  nor (_43047_, _43046_, _43005_);
  nor (_43048_, _43047_, _43040_);
  not (_43049_, _43048_);
  not (_43050_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43051_, _42999_, _43050_);
  nor (_43052_, _42999_, _43050_);
  nor (_43053_, _43052_, _43051_);
  not (_43054_, _43053_);
  not (_43055_, _42049_);
  nor (_43056_, _42077_, _42008_);
  and (_43057_, _43056_, _43055_);
  and (_43058_, _43057_, _42074_);
  not (_43059_, _41989_);
  and (_43060_, _42001_, _42069_);
  nor (_43061_, _43060_, _42039_);
  nor (_43062_, _43061_, _43059_);
  and (_43063_, _42023_, _41997_);
  nor (_43064_, _43063_, _43062_);
  not (_43065_, _42023_);
  nor (_43066_, _42070_, _42002_);
  nor (_43067_, _43066_, _43065_);
  nor (_43068_, _43067_, _41993_);
  and (_43069_, _43068_, _43064_);
  and (_43070_, _43069_, _43058_);
  and (_43071_, _42039_, _41981_);
  or (_43072_, _43071_, _42081_);
  nor (_43073_, _43072_, _42025_);
  not (_43074_, _42043_);
  and (_43075_, _42035_, _41974_);
  nor (_43076_, _42006_, _43075_);
  nor (_43077_, _43076_, _43074_);
  not (_43078_, _42046_);
  nor (_43079_, _41989_, _42022_);
  nor (_43080_, _43079_, _43078_);
  nor (_43081_, _43080_, _43077_);
  and (_43082_, _43081_, _43073_);
  not (_43083_, _43075_);
  nor (_43084_, _42014_, _42075_);
  and (_43085_, _43084_, _43083_);
  nor (_43086_, _43085_, _33605_);
  not (_43087_, _43086_);
  and (_43088_, _41997_, _41982_);
  and (_43089_, _42066_, _41981_);
  nor (_43090_, _43089_, _43088_);
  and (_43091_, _42013_, _41996_);
  and (_43092_, _42031_, _43091_);
  and (_43093_, _41989_, _42075_);
  nor (_43094_, _43093_, _43092_);
  and (_43095_, _43094_, _43090_);
  and (_43096_, _43095_, _43087_);
  and (_43097_, _43096_, _43082_);
  and (_43098_, _43097_, _43070_);
  and (_43099_, _41974_, _41976_);
  and (_43100_, _43099_, _42030_);
  not (_43101_, _43100_);
  and (_43102_, _43060_, _42023_);
  not (_43103_, _43102_);
  and (_43104_, _42020_, _41974_);
  and (_43105_, _43104_, _42043_);
  and (_43106_, _42043_, _42039_);
  nor (_43107_, _43106_, _43105_);
  and (_43108_, _43107_, _43103_);
  and (_43109_, _42014_, _41981_);
  and (_43110_, _42037_, _42023_);
  nor (_43111_, _43110_, _43109_);
  and (_43112_, _42070_, _42017_);
  nor (_43113_, _43112_, _42034_);
  and (_43114_, _43113_, _43111_);
  and (_43115_, _43114_, _43108_);
  and (_43116_, _43115_, _43101_);
  and (_43117_, _42070_, _41981_);
  nor (_43118_, _43117_, _41989_);
  not (_43119_, _42070_);
  nor (_43120_, _42014_, _42021_);
  and (_43121_, _43120_, _43119_);
  nor (_43122_, _43121_, _43118_);
  not (_43123_, _43122_);
  not (_43124_, _42058_);
  nor (_43125_, _41988_, _42022_);
  nor (_43126_, _43125_, _43124_);
  and (_43127_, _43104_, _42022_);
  nor (_43128_, _43127_, _43126_);
  and (_43129_, _43128_, _43123_);
  and (_43130_, _42023_, _41992_);
  not (_43131_, _43130_);
  and (_43132_, _42039_, _42023_);
  and (_43133_, _42046_, _42017_);
  nor (_43134_, _43133_, _43132_);
  and (_43135_, _43134_, _43131_);
  and (_43136_, _42078_, _41974_);
  and (_43137_, _43136_, _41989_);
  nor (_43138_, _43084_, _43065_);
  nor (_43139_, _43138_, _43137_);
  and (_43140_, _43139_, _43135_);
  and (_43141_, _43140_, _43129_);
  and (_43142_, _43141_, _43116_);
  and (_43143_, _43142_, _43098_);
  not (_43144_, _43143_);
  nor (_43145_, _42992_, _42990_);
  nor (_43146_, _43145_, _42993_);
  nand (_43147_, _43146_, _43144_);
  nand (_43148_, _43134_, _43073_);
  or (_43149_, _42034_, _41993_);
  or (_43150_, _43149_, _43138_);
  or (_43151_, _43112_, _42067_);
  and (_43152_, _42058_, _42017_);
  or (_43153_, _43105_, _43152_);
  or (_43154_, _43153_, _43151_);
  or (_43155_, _43154_, _43150_);
  or (_43156_, _43155_, _43148_);
  nor (_43157_, _43156_, _43143_);
  not (_43158_, _43157_);
  nor (_43159_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43160_, _43159_, _42990_);
  and (_43161_, _43160_, _43158_);
  or (_43162_, _43146_, _43144_);
  and (_43163_, _43162_, _43147_);
  nand (_43164_, _43163_, _43161_);
  and (_43165_, _43164_, _43147_);
  not (_43166_, _43165_);
  and (_43167_, _42997_, _42994_);
  nor (_43168_, _43167_, _42998_);
  and (_43169_, _43168_, _43166_);
  and (_43170_, _43169_, _43054_);
  not (_43171_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43172_, _43051_, _43171_);
  or (_43173_, _43172_, _43046_);
  and (_43174_, _43173_, _43170_);
  and (_43175_, _43174_, _43049_);
  and (_43176_, _43175_, _43045_);
  and (_43177_, _43176_, _43043_);
  nor (_43178_, _43039_, _43002_);
  or (_43179_, _43178_, _43035_);
  and (_43180_, _43179_, _43177_);
  and (_43181_, _43180_, _43038_);
  and (_43182_, _43181_, _43034_);
  and (_43183_, _43182_, _43030_);
  and (_43184_, _43183_, _43027_);
  and (_43185_, _43184_, _43025_);
  and (_43186_, _43185_, _43022_);
  and (_43187_, _43186_, _43020_);
  nor (_43188_, _43186_, _43020_);
  or (_43189_, _43188_, _43187_);
  or (_43190_, _43189_, _42983_);
  or (_43191_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_43192_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_43193_, _43192_, _43191_);
  and (_43194_, _43193_, _43190_);
  or (_38849_, _43194_, _42980_);
  nor (_43195_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38850_, _43195_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38851_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _43998_);
  and (_43196_, \oc8051_top_1.oc8051_rom1.ea_int , _33180_);
  nand (_43197_, _43196_, _33213_);
  and (_38852_, _43197_, _38851_);
  and (_38854_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _43998_);
  nor (_43198_, _42773_, _39864_);
  or (_43199_, _43143_, _33485_);
  nor (_43200_, _43157_, _33409_);
  nand (_43201_, _43143_, _33485_);
  and (_43202_, _43201_, _43199_);
  nand (_43203_, _43202_, _43200_);
  and (_43204_, _43203_, _43199_);
  nor (_43205_, _43204_, _39864_);
  and (_43206_, _43205_, _33300_);
  nor (_43207_, _43205_, _33300_);
  nor (_43208_, _43207_, _43206_);
  nor (_43209_, _43208_, _43198_);
  and (_43210_, _33496_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43211_, _43210_, _43198_);
  and (_43212_, _43211_, _43156_);
  or (_43213_, _43212_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_43214_, _43213_, _43209_);
  and (_38855_, _43214_, _43998_);
  nor (_43215_, _34813_, _34574_);
  not (_43216_, _35708_);
  and (_43217_, _43216_, _34324_);
  and (_43218_, _43217_, _43215_);
  not (_43219_, _35052_);
  and (_43220_, _33224_, _43998_);
  and (_43221_, _43220_, _34041_);
  and (_43222_, _43221_, _43219_);
  nor (_43223_, _33562_, _33812_);
  and (_43224_, _43223_, _43222_);
  and (_38858_, _43224_, _43218_);
  nor (_43225_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_43226_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_43227_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38861_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _43998_);
  and (_43228_, _38861_, _43227_);
  or (_38859_, _43228_, _43226_);
  not (_43229_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_43230_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43231_, _43230_, _43229_);
  and (_43232_, _43230_, _43229_);
  nor (_43233_, _43232_, _43231_);
  not (_43234_, _43233_);
  and (_43235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43236_, _43235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43237_, _43235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43238_, _43237_, _43236_);
  or (_43239_, _43238_, _43230_);
  and (_43240_, _43239_, _43234_);
  nor (_43241_, _43231_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43242_, _43231_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_43243_, _43242_, _43241_);
  or (_43244_, _43236_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38863_, _43244_, _43998_);
  and (_43245_, _38863_, _43243_);
  and (_38862_, _43245_, _43240_);
  not (_43246_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_43247_, _42773_, _43246_);
  and (_43248_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_43249_, _43247_);
  and (_43250_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_43251_, _43250_, _43248_);
  and (_38864_, _43251_, _43998_);
  and (_43252_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43253_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_43254_, _43253_, _43252_);
  and (_38865_, _43254_, _43998_);
  and (_43255_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_43256_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43257_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _43256_);
  and (_43258_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_43259_, _43258_, _43255_);
  and (_38866_, _43259_, _43998_);
  and (_43260_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43261_, _43260_, _43257_);
  and (_38867_, _43261_, _43998_);
  or (_43262_, _43256_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38869_, _43262_, _43998_);
  not (_43263_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_43264_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_43265_, _43264_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43266_, _43256_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_43267_, _43266_, _43998_);
  and (_38870_, _43267_, _43265_);
  or (_43268_, _43256_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38871_, _43268_, _43998_);
  nor (_43269_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_43270_, _43269_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43271_, _43270_, _43998_);
  and (_43272_, _38861_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38872_, _43272_, _43271_);
  and (_43273_, _43246_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_43274_, _43273_, _43270_);
  and (_38873_, _43274_, _43998_);
  nand (_43275_, _43270_, _38591_);
  or (_43276_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_43277_, _43276_, _43998_);
  and (_38874_, _43277_, _43275_);
  and (_38875_, _37337_, _39828_);
  or (_43278_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_43279_, _42668_, _42925_);
  and (_43280_, _43279_, _43998_);
  and (_38906_, _43280_, _43278_);
  or (_43281_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_43282_, _42668_, _42920_);
  and (_43283_, _43282_, _43998_);
  and (_38907_, _43283_, _43281_);
  or (_43284_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_43285_, _42668_, _42915_);
  and (_43286_, _43285_, _43998_);
  and (_38908_, _43286_, _43284_);
  or (_43287_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_43288_, _42668_, _42909_);
  and (_43289_, _43288_, _43998_);
  and (_38909_, _43289_, _43287_);
  or (_43290_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_43291_, _42668_, _42904_);
  and (_43292_, _43291_, _43998_);
  and (_38911_, _43292_, _43290_);
  or (_43293_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_43294_, _42668_, _42898_);
  and (_43295_, _43294_, _43998_);
  and (_38912_, _43295_, _43293_);
  or (_43296_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_43297_, _42668_, _42891_);
  and (_43298_, _43297_, _43998_);
  and (_38913_, _43298_, _43296_);
  or (_43299_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_43300_, _42668_, _42886_);
  and (_43301_, _43300_, _43998_);
  and (_38914_, _43301_, _43299_);
  or (_43302_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_43303_, _42668_, _38512_);
  and (_43304_, _43303_, _43998_);
  and (_38915_, _43304_, _43302_);
  or (_43305_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_43306_, _42668_, _38518_);
  and (_43307_, _43306_, _43998_);
  and (_38916_, _43307_, _43305_);
  or (_43308_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_43309_, _42668_, _38523_);
  and (_43310_, _43309_, _43998_);
  and (_38917_, _43310_, _43308_);
  or (_43311_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_43312_, _42668_, _38508_);
  and (_43313_, _43312_, _43998_);
  and (_38918_, _43313_, _43311_);
  or (_43314_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_43315_, _42668_, _38529_);
  and (_43316_, _43315_, _43998_);
  and (_38919_, _43316_, _43314_);
  or (_43317_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_43318_, _42668_, _38504_);
  and (_43319_, _43318_, _43998_);
  and (_38920_, _43319_, _43317_);
  or (_43320_, _42668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_43321_, _42668_, _38535_);
  and (_43322_, _43321_, _43998_);
  and (_38922_, _43322_, _43320_);
  or (_43323_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_43324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _43998_);
  or (_43325_, _43324_, _00000_);
  and (_38926_, _43325_, _43323_);
  or (_43326_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_43327_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _43998_);
  or (_43328_, _43327_, _00000_);
  and (_38927_, _43328_, _43326_);
  or (_43329_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_43330_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _43998_);
  or (_43331_, _43330_, _00000_);
  and (_38928_, _43331_, _43329_);
  or (_43332_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_43333_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _43998_);
  or (_43334_, _43333_, _00000_);
  and (_38929_, _43334_, _43332_);
  or (_43335_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_43336_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _43998_);
  or (_43337_, _43336_, _00000_);
  and (_38930_, _43337_, _43335_);
  or (_43338_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_43339_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _43998_);
  or (_43340_, _43339_, _00000_);
  and (_38931_, _43340_, _43338_);
  or (_43341_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_43342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _43998_);
  or (_43343_, _43342_, _00000_);
  and (_38932_, _43343_, _43341_);
  or (_43344_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_43345_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _43998_);
  or (_43346_, _43345_, _00000_);
  and (_38933_, _43346_, _43344_);
  or (_43347_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_43348_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _43998_);
  or (_43349_, _43348_, _00000_);
  and (_38934_, _43349_, _43347_);
  or (_43350_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_43351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _43998_);
  or (_43352_, _43351_, _00000_);
  and (_38936_, _43352_, _43350_);
  or (_43353_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_43354_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _43998_);
  or (_43355_, _43354_, _00000_);
  and (_38937_, _43355_, _43353_);
  or (_43356_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_43357_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _43998_);
  or (_43358_, _43357_, _00000_);
  and (_38938_, _43358_, _43356_);
  or (_43359_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_43360_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _43998_);
  or (_43361_, _43360_, _00000_);
  and (_38939_, _43361_, _43359_);
  or (_43362_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_43363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _43998_);
  or (_43364_, _43363_, _00000_);
  and (_38940_, _43364_, _43362_);
  or (_43365_, _42672_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_43366_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _43998_);
  or (_43367_, _43366_, _00000_);
  and (_38941_, _43367_, _43365_);
  and (_43368_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_43369_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_43370_, _43369_, _43247_);
  or (_43371_, _43370_, _43368_);
  and (_39119_, _43371_, _43998_);
  and (_43372_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_43373_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_43374_, _43373_, _43372_);
  and (_39120_, _43374_, _43998_);
  and (_43375_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_43376_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_43377_, _43376_, _43375_);
  and (_39121_, _43377_, _43998_);
  and (_43378_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_43379_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_43380_, _43379_, _43378_);
  and (_39122_, _43380_, _43998_);
  and (_43381_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_43382_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_43383_, _43382_, _43247_);
  or (_43384_, _43383_, _43381_);
  and (_39123_, _43384_, _43998_);
  and (_43385_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_43386_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_43387_, _43386_, _43385_);
  and (_39124_, _43387_, _43998_);
  and (_43388_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_43389_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_43390_, _43389_, _43388_);
  and (_39125_, _43390_, _43998_);
  and (_43391_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_43392_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_43393_, _43392_, _43391_);
  and (_39127_, _43393_, _43998_);
  and (_43394_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_43395_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_43396_, _43395_, _43394_);
  and (_39128_, _43396_, _43998_);
  and (_43397_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_43398_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_43399_, _43398_, _43397_);
  and (_39129_, _43399_, _43998_);
  and (_43400_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_43401_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_43402_, _43401_, _43400_);
  and (_39130_, _43402_, _43998_);
  and (_43403_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_43404_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_43405_, _43404_, _43403_);
  and (_39131_, _43405_, _43998_);
  and (_43406_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_43407_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_43408_, _43407_, _43406_);
  and (_39132_, _43408_, _43998_);
  and (_43409_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_43410_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_43411_, _43410_, _43409_);
  and (_39133_, _43411_, _43998_);
  and (_43412_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_43413_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_43420_, _43413_, _43412_);
  and (_39134_, _43420_, _43998_);
  and (_43429_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_43437_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_43442_, _43437_, _43429_);
  and (_39135_, _43442_, _43998_);
  and (_43453_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_43460_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_43464_, _43460_, _43453_);
  and (_39136_, _43464_, _43998_);
  and (_43477_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_43482_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_43486_, _43482_, _43477_);
  and (_39138_, _43486_, _43998_);
  and (_43494_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_43503_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_43511_, _43503_, _43494_);
  and (_39139_, _43511_, _43998_);
  and (_43521_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_43527_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_43535_, _43527_, _43521_);
  and (_39140_, _43535_, _43998_);
  and (_43543_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_43551_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_43558_, _43551_, _43543_);
  and (_39141_, _43558_, _43998_);
  and (_43567_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_43575_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_43580_, _43575_, _43567_);
  and (_39142_, _43580_, _43998_);
  and (_43591_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_43598_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_43602_, _43598_, _43591_);
  and (_39143_, _43602_, _43998_);
  and (_43615_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_43620_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_43624_, _43620_, _43615_);
  and (_39144_, _43624_, _43998_);
  and (_43632_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_43633_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_43634_, _43633_, _43632_);
  and (_39145_, _43634_, _43998_);
  and (_43635_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_43636_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_43637_, _43636_, _43635_);
  and (_39146_, _43637_, _43998_);
  and (_43638_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_43639_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_43640_, _43639_, _43638_);
  and (_39147_, _43640_, _43998_);
  and (_43641_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_43642_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_43643_, _43642_, _43641_);
  and (_39148_, _43643_, _43998_);
  and (_43644_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_43645_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_43646_, _43645_, _43644_);
  and (_39149_, _43646_, _43998_);
  and (_43647_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_43648_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_43649_, _43648_, _43647_);
  and (_39150_, _43649_, _43998_);
  and (_43650_, _43247_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_43651_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_43652_, _43651_, _43650_);
  and (_39151_, _43652_, _43998_);
  nor (_39152_, _35785_, rst);
  nor (_39153_, _33899_, rst);
  nor (_39154_, _34139_, rst);
  nor (_39155_, _39841_, rst);
  nor (_39156_, _39859_, rst);
  nor (_39158_, _40115_, rst);
  nor (_39159_, _40003_, rst);
  nor (_39160_, _39958_, rst);
  and (_39161_, _40131_, _43998_);
  nor (_39162_, _40043_, rst);
  nor (_39164_, _40185_, rst);
  and (_39180_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _43998_);
  and (_39181_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _43998_);
  and (_39182_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _43998_);
  and (_39183_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _43998_);
  and (_39185_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _43998_);
  and (_39186_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _43998_);
  and (_39187_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _43998_);
  or (_43653_, _42769_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_43654_, _43653_, _43998_);
  and (_43655_, _42833_, _42842_);
  and (_43656_, _43655_, _42840_);
  or (_43657_, _43656_, _42841_);
  and (_43658_, _43657_, _28383_);
  and (_43659_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_43660_, _42837_, _42565_);
  and (_43661_, _42845_, _39881_);
  or (_43662_, _43661_, _43660_);
  or (_43663_, _43662_, _43659_);
  and (_43664_, _42928_, _42925_);
  nor (_43665_, _43664_, _42929_);
  and (_43666_, _43665_, _42974_);
  nor (_43667_, _43666_, _43663_);
  nand (_43668_, _43667_, _42805_);
  or (_43669_, _43668_, _43658_);
  and (_39188_, _43669_, _43654_);
  or (_43670_, _42769_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_43671_, _43670_, _43998_);
  and (_43672_, _43657_, _29097_);
  and (_43673_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_43674_, _42837_, _42582_);
  and (_43675_, _42845_, _40096_);
  or (_43676_, _43675_, _43674_);
  or (_43677_, _43676_, _43673_);
  or (_43678_, _43677_, _43672_);
  or (_43679_, _42931_, _42929_);
  nand (_43680_, _43679_, _42974_);
  or (_43681_, _43680_, _42932_);
  nand (_43682_, _43681_, _42805_);
  or (_43683_, _43682_, _43678_);
  and (_39189_, _43683_, _43671_);
  not (_43684_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_43685_, _42773_, _43684_);
  and (_43686_, _42773_, _43684_);
  nor (_43687_, _43686_, _43685_);
  or (_43688_, _43687_, _42769_);
  and (_43689_, _43688_, _43998_);
  and (_43690_, _43657_, _29774_);
  and (_43691_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43692_, _42837_, _42599_);
  and (_43693_, _42845_, _40024_);
  or (_43694_, _43693_, _43692_);
  or (_43695_, _43694_, _43691_);
  or (_43696_, _43695_, _43690_);
  nor (_43697_, _42936_, _42934_);
  nor (_43698_, _43697_, _42937_);
  nand (_43699_, _43698_, _42974_);
  nand (_43700_, _43699_, _42805_);
  or (_43701_, _43700_, _43696_);
  and (_39190_, _43701_, _43689_);
  and (_43702_, _43685_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_43703_, _43685_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_43704_, _43703_, _43702_);
  or (_43705_, _43704_, _42769_);
  and (_43706_, _43705_, _43998_);
  and (_43707_, _43657_, _30525_);
  and (_43708_, _42837_, _42616_);
  and (_43709_, _42845_, _39975_);
  or (_43710_, _43709_, _43708_);
  or (_43711_, _42914_, _42913_);
  or (_43712_, _43711_, _42938_);
  nand (_43713_, _43711_, _42938_);
  and (_43714_, _43713_, _42974_);
  and (_43715_, _43714_, _43712_);
  or (_43716_, _43715_, _43710_);
  or (_43717_, _43716_, _43707_);
  nand (_43718_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_43719_, _43718_, _42805_);
  or (_43720_, _43719_, _43717_);
  and (_39191_, _43720_, _43706_);
  and (_43721_, _42776_, _42774_);
  nor (_43722_, _43702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43723_, _43722_, _43721_);
  or (_43724_, _43723_, _42769_);
  and (_43725_, _43724_, _43998_);
  and (_43726_, _43657_, _31296_);
  and (_43727_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43728_, _42837_, _42633_);
  and (_43729_, _42845_, _40150_);
  or (_43730_, _43729_, _43728_);
  or (_43731_, _43730_, _43727_);
  or (_43732_, _43731_, _43726_);
  or (_43733_, _42942_, _42940_);
  and (_43734_, _43733_, _42943_);
  nand (_43735_, _43734_, _42974_);
  nand (_43736_, _43735_, _42805_);
  or (_43737_, _43736_, _43732_);
  and (_39192_, _43737_, _43725_);
  not (_43738_, _42777_);
  nor (_43739_, _43738_, _42773_);
  nor (_43740_, _43721_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43741_, _43740_, _43739_);
  or (_43742_, _43741_, _42769_);
  and (_43743_, _43742_, _43998_);
  and (_43744_, _43657_, _32113_);
  and (_43745_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43746_, _42837_, _42650_);
  and (_43747_, _42845_, _40060_);
  or (_43748_, _43747_, _43746_);
  or (_43749_, _43748_, _43745_);
  or (_43750_, _42902_, _42903_);
  or (_43751_, _43750_, _42944_);
  nand (_43752_, _43750_, _42944_);
  and (_43753_, _43752_, _42974_);
  and (_43754_, _43753_, _43751_);
  nor (_43755_, _43754_, _43749_);
  nand (_43756_, _43755_, _42805_);
  or (_43757_, _43756_, _43744_);
  and (_39193_, _43757_, _43743_);
  nor (_43758_, _43739_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43759_, _43739_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_43760_, _43759_, _43758_);
  or (_43761_, _43760_, _42769_);
  and (_43762_, _43761_, _43998_);
  not (_43763_, _42805_);
  nor (_43764_, _42946_, _42897_);
  nor (_43765_, _43764_, _42947_);
  and (_43766_, _43765_, _42974_);
  and (_43767_, _43657_, _32930_);
  and (_43768_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43769_, _42837_, _42667_);
  and (_43770_, _42845_, _40202_);
  or (_43771_, _43770_, _43769_);
  or (_43772_, _43771_, _43768_);
  or (_43773_, _43772_, _43767_);
  or (_43774_, _43773_, _43766_);
  or (_43775_, _43774_, _43763_);
  and (_39194_, _43775_, _43762_);
  nor (_43776_, _43759_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43777_, _43759_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_43778_, _43777_, _43776_);
  or (_43779_, _43778_, _42769_);
  and (_43780_, _43779_, _43998_);
  and (_43781_, _43657_, _27143_);
  and (_43782_, _36970_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43783_, _42837_, _42548_);
  and (_43784_, _42845_, _39941_);
  or (_43785_, _43784_, _43783_);
  or (_43786_, _43785_, _43782_);
  or (_43787_, _42949_, _42890_);
  and (_43788_, _42974_, _42950_);
  and (_43789_, _43788_, _43787_);
  or (_43790_, _43789_, _43786_);
  or (_43791_, _43790_, _43781_);
  or (_43792_, _43791_, _43763_);
  and (_39196_, _43792_, _43780_);
  or (_43793_, _43777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43795_, _43794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_43796_, _43795_, _43739_);
  and (_43797_, _43796_, _43793_);
  or (_43798_, _43797_, _42769_);
  and (_43799_, _43798_, _43998_);
  nor (_43800_, _36981_, _28372_);
  nor (_43801_, _42848_, _38629_);
  and (_43802_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43803_, _42837_, _39881_);
  or (_43804_, _43803_, _43802_);
  or (_43805_, _43804_, _43801_);
  and (_43806_, _42845_, _41996_);
  nor (_43807_, _42951_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43808_, _42951_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_43809_, _43808_, _43807_);
  and (_43810_, _43809_, _42960_);
  nor (_43811_, _43809_, _42960_);
  or (_43812_, _43811_, _43810_);
  and (_43813_, _43812_, _42974_);
  or (_43814_, _43813_, _43806_);
  or (_43815_, _43814_, _43805_);
  or (_43816_, _43815_, _43800_);
  or (_43817_, _43816_, _43763_);
  and (_39197_, _43817_, _43799_);
  nand (_43818_, _43796_, _43001_);
  or (_43819_, _43796_, _43001_);
  and (_43820_, _43819_, _43818_);
  or (_43821_, _43820_, _42769_);
  and (_43822_, _43821_, _43998_);
  and (_43823_, _42845_, _42012_);
  nor (_43824_, _42848_, _38659_);
  and (_43825_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_43826_, _42837_, _40096_);
  or (_43827_, _43826_, _43825_);
  or (_43828_, _43827_, _43824_);
  or (_43829_, _43828_, _43823_);
  nor (_43830_, _36981_, _29086_);
  or (_43831_, _43830_, _43829_);
  and (_43832_, _42952_, _42960_);
  nor (_43833_, _42951_, _38512_);
  and (_43834_, _43833_, _42885_);
  nor (_43835_, _43834_, _43832_);
  nand (_43836_, _43835_, _38518_);
  or (_43837_, _43835_, _38518_);
  and (_43838_, _43837_, _43836_);
  and (_43839_, _43838_, _42974_);
  or (_43840_, _43839_, _43763_);
  or (_43841_, _43840_, _43831_);
  and (_39198_, _43841_, _43822_);
  and (_43842_, _43795_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_43843_, _43842_, _43739_);
  and (_43844_, _43843_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_43845_, _43843_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_43846_, _43845_, _43844_);
  or (_43847_, _43846_, _42769_);
  and (_43848_, _43847_, _43998_);
  nor (_43849_, _36981_, _29763_);
  nor (_43850_, _42848_, _38689_);
  and (_43851_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43852_, _42837_, _40024_);
  or (_43853_, _43852_, _43851_);
  or (_43854_, _43853_, _43850_);
  and (_43855_, _42845_, _41973_);
  and (_43856_, _42953_, _42960_);
  and (_43857_, _43834_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_43858_, _43857_, _43856_);
  or (_43859_, _43858_, _38523_);
  nand (_43860_, _43858_, _38523_);
  and (_43861_, _43860_, _42974_);
  and (_43862_, _43861_, _43859_);
  or (_43863_, _43862_, _43855_);
  or (_43864_, _43863_, _43854_);
  or (_43865_, _43864_, _43849_);
  or (_43866_, _43865_, _43763_);
  and (_39199_, _43866_, _43848_);
  nor (_43867_, _43844_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43868_, _42781_, _42774_);
  and (_43869_, _43868_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43870_, _43869_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_43871_, _43870_, _43867_);
  or (_43872_, _43871_, _42769_);
  and (_43873_, _43872_, _43998_);
  nor (_43874_, _36981_, _30514_);
  nor (_43875_, _42848_, _38721_);
  and (_43876_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43877_, _42837_, _39975_);
  or (_43878_, _43877_, _43876_);
  or (_43879_, _43878_, _43875_);
  nor (_43880_, _42817_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_43881_, _43880_, _42818_);
  and (_43882_, _43881_, _42845_);
  and (_43883_, _42964_, _42885_);
  and (_43884_, _42954_, _42960_);
  nor (_43885_, _43884_, _43883_);
  and (_43886_, _43885_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_43887_, _43885_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_43888_, _43887_, _43886_);
  and (_43889_, _43888_, _42974_);
  or (_43890_, _43889_, _43882_);
  or (_43891_, _43890_, _43879_);
  or (_43892_, _43891_, _43874_);
  or (_43893_, _43892_, _43763_);
  and (_39200_, _43893_, _43873_);
  and (_43894_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43895_, _43894_, _43844_);
  nor (_43896_, _43870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_43897_, _43896_, _43895_);
  or (_43898_, _43897_, _42769_);
  and (_43899_, _43898_, _43998_);
  nor (_43900_, _42848_, _38777_);
  and (_43901_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_43902_, _42837_, _40150_);
  or (_43903_, _43902_, _43901_);
  or (_43904_, _43903_, _43900_);
  and (_43905_, _42814_, _42962_);
  and (_43906_, _43905_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_43907_, _43906_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_43908_, _43907_, _42819_);
  and (_43909_, _43908_, _42845_);
  and (_43910_, _42965_, _42885_);
  and (_43911_, _42955_, _42960_);
  nor (_43912_, _43911_, _43910_);
  and (_43913_, _43912_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_43914_, _43912_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_43915_, _43914_, _43913_);
  and (_43916_, _43915_, _42974_);
  or (_43917_, _43916_, _43909_);
  or (_43918_, _43917_, _43904_);
  nor (_43919_, _36981_, _31285_);
  or (_43920_, _43919_, _43763_);
  or (_43921_, _43920_, _43918_);
  and (_39201_, _43921_, _43899_);
  and (_43922_, _43895_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43923_, _43895_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43924_, _43923_, _43922_);
  or (_43925_, _43924_, _42769_);
  and (_43926_, _43925_, _43998_);
  and (_43927_, _42966_, _42885_);
  and (_43928_, _42956_, _42960_);
  nor (_43929_, _43928_, _43927_);
  and (_43930_, _43929_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43931_, _43929_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_43932_, _43931_, _43930_);
  and (_43933_, _43932_, _42974_);
  nor (_43934_, _42819_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43935_, _43934_, _42820_);
  and (_43936_, _43935_, _42845_);
  nor (_43937_, _36981_, _32102_);
  nor (_43938_, _42848_, _38812_);
  and (_43939_, _42837_, _40060_);
  and (_43940_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_43941_, _43940_, _43939_);
  or (_43942_, _43941_, _43938_);
  or (_43943_, _43942_, _43937_);
  or (_43944_, _43943_, _43936_);
  or (_43945_, _43944_, _43933_);
  or (_43946_, _43945_, _43763_);
  and (_39202_, _43946_, _43926_);
  nor (_43947_, _43922_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_43948_, _43947_, _42787_);
  or (_43949_, _43948_, _42769_);
  and (_43950_, _43949_, _43998_);
  nor (_43951_, _42967_, _42960_);
  nor (_43952_, _42957_, _42885_);
  nor (_43953_, _43952_, _43951_);
  nand (_43954_, _43953_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_43955_, _43953_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43956_, _43955_, _42974_);
  and (_43957_, _43956_, _43954_);
  or (_43958_, _42820_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43959_, _43958_, _42821_);
  and (_43960_, _43959_, _42845_);
  nor (_43961_, _36981_, _32919_);
  nor (_43962_, _42848_, _38868_);
  and (_43963_, _42870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_43964_, _42837_, _40202_);
  or (_43965_, _43964_, _43963_);
  or (_43966_, _43965_, _43962_);
  or (_43967_, _43966_, _43961_);
  or (_43968_, _43967_, _43960_);
  or (_43969_, _43968_, _43957_);
  or (_43970_, _43969_, _43763_);
  and (_39203_, _43970_, _43950_);
  and (_43971_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_43972_, _43160_, _43158_);
  nor (_43973_, _43972_, _43161_);
  or (_43974_, _43973_, _42983_);
  or (_43975_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_43976_, _43975_, _43192_);
  and (_43978_, _43976_, _43974_);
  or (_39204_, _43978_, _43971_);
  or (_43981_, _43163_, _43161_);
  and (_43983_, _43981_, _43164_);
  or (_43985_, _43983_, _42983_);
  or (_43987_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_43989_, _43987_, _43192_);
  and (_43990_, _43989_, _43985_);
  and (_43991_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39205_, _43991_, _43990_);
  nor (_43992_, _43168_, _43166_);
  nor (_43993_, _43992_, _43169_);
  or (_43994_, _43993_, _42983_);
  or (_43996_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43997_, _43996_, _43192_);
  and (_43999_, _43997_, _43994_);
  and (_44000_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_39207_, _44000_, _43999_);
  and (_44002_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_44003_, _43169_, _43054_);
  nor (_44004_, _44003_, _43170_);
  or (_44006_, _44004_, _42983_);
  or (_44007_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_44008_, _44007_, _43192_);
  and (_44010_, _44008_, _44006_);
  or (_39208_, _44010_, _44002_);
  and (_44011_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_44013_, _43173_, _43170_);
  nor (_44014_, _44013_, _43174_);
  or (_44015_, _44014_, _42983_);
  or (_44017_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_44018_, _44017_, _43192_);
  and (_44019_, _44018_, _44015_);
  or (_39209_, _44019_, _44011_);
  and (_44021_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_44022_, _43174_, _43049_);
  nor (_44024_, _44022_, _43175_);
  or (_44025_, _44024_, _42983_);
  or (_44026_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_44027_, _44026_, _43192_);
  and (_44028_, _44027_, _44025_);
  or (_39210_, _44028_, _44021_);
  nor (_44029_, _43175_, _43045_);
  nor (_44030_, _44029_, _43176_);
  or (_44031_, _44030_, _42983_);
  or (_44032_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_44033_, _44032_, _43192_);
  and (_44034_, _44033_, _44031_);
  and (_44035_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39211_, _44035_, _44034_);
  nor (_44036_, _43176_, _43043_);
  nor (_44037_, _44036_, _43177_);
  or (_44038_, _44037_, _42983_);
  or (_44039_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_44040_, _44039_, _43192_);
  and (_44041_, _44040_, _44038_);
  and (_44042_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_39212_, _44042_, _44041_);
  and (_44044_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_44046_, _43179_, _43177_);
  nor (_44047_, _44046_, _43180_);
  or (_44048_, _44047_, _42983_);
  or (_44050_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_44051_, _44050_, _43192_);
  and (_44052_, _44051_, _44048_);
  or (_39213_, _44052_, _44044_);
  nor (_44054_, _43180_, _43038_);
  nor (_44055_, _44054_, _43181_);
  or (_44057_, _44055_, _42983_);
  or (_44058_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_44059_, _44058_, _43192_);
  and (_44061_, _44059_, _44057_);
  and (_44062_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39214_, _44062_, _44061_);
  or (_44064_, _43181_, _43034_);
  nor (_44065_, _43182_, _42983_);
  and (_44066_, _44065_, _44064_);
  nor (_44068_, _42982_, _38523_);
  or (_44069_, _44068_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_44070_, _44069_, _44066_);
  or (_44072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _33180_);
  and (_44073_, _44072_, _43998_);
  and (_39215_, _44073_, _44070_);
  nor (_44074_, _43182_, _43030_);
  nor (_44075_, _44074_, _43183_);
  or (_44076_, _44075_, _42983_);
  or (_44077_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_44078_, _44077_, _43192_);
  and (_44079_, _44078_, _44076_);
  and (_44080_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39216_, _44080_, _44079_);
  nor (_44081_, _43183_, _43027_);
  nor (_44082_, _44081_, _43184_);
  or (_44083_, _44082_, _42983_);
  or (_44084_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_44085_, _44084_, _43192_);
  and (_44086_, _44085_, _44083_);
  and (_44087_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39218_, _44087_, _44086_);
  nor (_44088_, _43184_, _43025_);
  nor (_44089_, _44088_, _43185_);
  or (_44091_, _44089_, _42983_);
  or (_44092_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_44094_, _44092_, _43192_);
  and (_44095_, _44094_, _44091_);
  and (_44096_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39219_, _44096_, _44095_);
  nor (_44098_, _43185_, _43022_);
  nor (_44099_, _44098_, _43186_);
  or (_44101_, _44099_, _42983_);
  or (_44102_, _42982_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_44103_, _44102_, _43192_);
  and (_44105_, _44103_, _44101_);
  and (_44106_, _42979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39220_, _44106_, _44105_);
  and (_39221_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _43998_);
  and (_39222_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _43998_);
  and (_39223_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _43998_);
  and (_39224_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _43998_);
  and (_39225_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _43998_);
  and (_39226_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _43998_);
  and (_39227_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _43998_);
  nor (_00011_, _43157_, _39864_);
  nand (_00012_, _00011_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00014_, _00011_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00015_, _00014_, _43192_);
  and (_39229_, _00015_, _00012_);
  or (_00016_, _43202_, _43200_);
  and (_00017_, _00016_, _43203_);
  or (_00018_, _00017_, _39864_);
  or (_00019_, _33213_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00020_, _00019_, _43192_);
  and (_39230_, _00020_, _00018_);
  and (_00021_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00022_, _43369_, _38861_);
  or (_39246_, _00022_, _00021_);
  and (_00023_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00024_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00025_, _00024_, _38861_);
  or (_39247_, _00025_, _00023_);
  and (_00026_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00027_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00028_, _00027_, _38861_);
  or (_39248_, _00028_, _00026_);
  and (_00029_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00031_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00032_, _00031_, _38861_);
  or (_39249_, _00032_, _00029_);
  and (_00034_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00035_, _43382_, _38861_);
  or (_39251_, _00035_, _00034_);
  and (_00037_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00038_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00040_, _00038_, _38861_);
  or (_39252_, _00040_, _00037_);
  and (_00041_, _43225_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00043_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00044_, _00043_, _38861_);
  or (_39253_, _00044_, _00041_);
  and (_39254_, _43233_, _43998_);
  nor (_39255_, _43243_, rst);
  and (_39256_, _43239_, _43998_);
  and (_00047_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00048_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00049_, _00048_, _00047_);
  and (_39257_, _00049_, _43998_);
  and (_00051_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00052_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00054_, _00052_, _00051_);
  and (_39258_, _00054_, _43998_);
  and (_00055_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00056_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00057_, _00056_, _00055_);
  and (_39259_, _00057_, _43998_);
  and (_00058_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00059_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00060_, _00059_, _00058_);
  and (_39260_, _00060_, _43998_);
  and (_00061_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00062_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00063_, _00062_, _00061_);
  and (_39262_, _00063_, _43998_);
  and (_00064_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00065_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00066_, _00065_, _00064_);
  and (_39263_, _00066_, _43998_);
  and (_00067_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00068_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00069_, _00068_, _00067_);
  and (_39264_, _00069_, _43998_);
  and (_00071_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00073_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00074_, _00073_, _00071_);
  and (_39265_, _00074_, _43998_);
  and (_00076_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00077_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00078_, _00077_, _00076_);
  and (_39266_, _00078_, _43998_);
  and (_00080_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00081_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00083_, _00081_, _00080_);
  and (_39267_, _00083_, _43998_);
  and (_00084_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00086_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00087_, _00086_, _00084_);
  and (_39268_, _00087_, _43998_);
  and (_00089_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00090_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00091_, _00090_, _00089_);
  and (_39269_, _00091_, _43998_);
  and (_00093_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00094_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00096_, _00094_, _00093_);
  and (_39270_, _00096_, _43998_);
  and (_00097_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00098_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00099_, _00098_, _00097_);
  and (_39271_, _00099_, _43998_);
  and (_00100_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00101_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00102_, _00101_, _00100_);
  and (_39272_, _00102_, _43998_);
  and (_00103_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00104_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00105_, _00104_, _00103_);
  and (_39273_, _00105_, _43998_);
  and (_00106_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00107_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00108_, _00107_, _00106_);
  and (_39274_, _00108_, _43998_);
  and (_00109_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00110_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00111_, _00110_, _00109_);
  and (_39275_, _00111_, _43998_);
  and (_00113_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00115_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00116_, _00115_, _00113_);
  and (_39276_, _00116_, _43998_);
  and (_00118_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00119_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00120_, _00119_, _00118_);
  and (_39277_, _00120_, _43998_);
  and (_00122_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00123_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00125_, _00123_, _00122_);
  and (_39278_, _00125_, _43998_);
  and (_00126_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00128_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00129_, _00128_, _00126_);
  and (_39279_, _00129_, _43998_);
  and (_00131_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00132_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00133_, _00132_, _00131_);
  and (_39280_, _00133_, _43998_);
  and (_00135_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00136_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00138_, _00136_, _00135_);
  and (_39281_, _00138_, _43998_);
  and (_00139_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00140_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00141_, _00140_, _00139_);
  and (_39283_, _00141_, _43998_);
  and (_00142_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00143_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00144_, _00143_, _00142_);
  and (_39284_, _00144_, _43998_);
  and (_00145_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00146_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00147_, _00146_, _00145_);
  and (_39285_, _00147_, _43998_);
  and (_00148_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00149_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00150_, _00149_, _00148_);
  and (_39286_, _00150_, _43998_);
  and (_00151_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00152_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00153_, _00152_, _00151_);
  and (_39287_, _00153_, _43998_);
  and (_00155_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00157_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00158_, _00157_, _00155_);
  and (_39288_, _00158_, _43998_);
  and (_00160_, _43247_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00161_, _43249_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00162_, _00161_, _00160_);
  and (_39289_, _00162_, _43998_);
  and (_00164_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00165_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00167_, _00165_, _00164_);
  and (_39290_, _00167_, _43998_);
  and (_00168_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00170_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00171_, _00170_, _00168_);
  and (_39291_, _00171_, _43998_);
  and (_00173_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00174_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00175_, _00174_, _00173_);
  and (_39292_, _00175_, _43998_);
  and (_00177_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00178_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00180_, _00178_, _00177_);
  and (_39294_, _00180_, _43998_);
  and (_00181_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00182_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00183_, _00182_, _00181_);
  and (_39295_, _00183_, _43998_);
  and (_00184_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00185_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00186_, _00185_, _00184_);
  and (_39296_, _00186_, _43998_);
  and (_00187_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00188_, _43257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00189_, _00188_, _00187_);
  and (_39297_, _00189_, _43998_);
  and (_00190_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00191_, _39859_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00192_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00193_, _00192_, _43256_);
  and (_00194_, _00193_, _00191_);
  or (_00195_, _00194_, _00190_);
  and (_39298_, _00195_, _43998_);
  and (_00197_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00198_, _40115_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00200_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00201_, _00200_, _43256_);
  and (_00202_, _00201_, _00198_);
  or (_00204_, _00202_, _00197_);
  and (_39299_, _00204_, _43998_);
  and (_00205_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00207_, _40003_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00208_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00209_, _00208_, _43256_);
  and (_00211_, _00209_, _00207_);
  or (_00212_, _00211_, _00205_);
  and (_39300_, _00212_, _43998_);
  and (_00214_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00215_, _39958_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00216_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00218_, _00216_, _43256_);
  and (_00219_, _00218_, _00215_);
  or (_00220_, _00219_, _00214_);
  and (_39301_, _00220_, _43998_);
  and (_00222_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00223_, _40131_, _43263_);
  or (_00225_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00226_, _00225_, _43256_);
  and (_00227_, _00226_, _00223_);
  or (_00228_, _00227_, _00222_);
  and (_39302_, _00228_, _43998_);
  and (_00229_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00230_, _40043_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00231_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00232_, _00231_, _43256_);
  and (_00233_, _00232_, _00230_);
  or (_00234_, _00233_, _00229_);
  and (_39303_, _00234_, _43998_);
  and (_00235_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00236_, _40185_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00237_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00238_, _00237_, _43256_);
  and (_00239_, _00238_, _00236_);
  or (_00240_, _00239_, _00235_);
  and (_39305_, _00240_, _43998_);
  and (_00241_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00242_, _39922_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00244_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00245_, _00244_, _43256_);
  and (_00247_, _00245_, _00242_);
  or (_00248_, _00247_, _00241_);
  and (_39306_, _00248_, _43998_);
  and (_00250_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00251_, _00250_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00252_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _43256_);
  and (_00254_, _00252_, _43998_);
  and (_39307_, _00254_, _00251_);
  and (_00255_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00257_, _00255_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00258_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _43256_);
  and (_00259_, _00258_, _43998_);
  and (_39308_, _00259_, _00257_);
  and (_00261_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00262_, _00261_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00264_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _43256_);
  and (_00265_, _00264_, _43998_);
  and (_39309_, _00265_, _00262_);
  and (_00267_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00268_, _00267_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00269_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _43256_);
  and (_00271_, _00269_, _43998_);
  and (_39310_, _00271_, _00268_);
  and (_00272_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00273_, _00272_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00274_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _43256_);
  and (_00275_, _00274_, _43998_);
  and (_39311_, _00275_, _00273_);
  and (_00276_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00277_, _00276_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00278_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _43256_);
  and (_00279_, _00278_, _43998_);
  and (_39312_, _00279_, _00277_);
  and (_00280_, _43263_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00281_, _00280_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00282_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _43256_);
  and (_00283_, _00282_, _43998_);
  and (_39313_, _00283_, _00281_);
  nand (_00284_, _43270_, _28372_);
  or (_00285_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00286_, _00285_, _43998_);
  and (_39314_, _00286_, _00284_);
  nand (_00288_, _43270_, _29086_);
  or (_00289_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00291_, _00289_, _43998_);
  and (_39316_, _00291_, _00288_);
  nand (_00292_, _43270_, _29763_);
  or (_00294_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00295_, _00294_, _43998_);
  and (_39317_, _00295_, _00292_);
  nand (_00297_, _43270_, _30514_);
  or (_00298_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00299_, _00298_, _43998_);
  and (_39318_, _00299_, _00297_);
  nand (_00301_, _43270_, _31285_);
  or (_00302_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00304_, _00302_, _43998_);
  and (_39319_, _00304_, _00301_);
  nand (_00305_, _43270_, _32102_);
  or (_00307_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00308_, _00307_, _43998_);
  and (_39320_, _00308_, _00305_);
  nand (_00310_, _43270_, _32919_);
  or (_00311_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00312_, _00311_, _43998_);
  and (_39321_, _00312_, _00310_);
  nand (_00314_, _43270_, _27132_);
  or (_00315_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00316_, _00315_, _43998_);
  and (_39322_, _00316_, _00314_);
  nand (_00317_, _43270_, _38629_);
  or (_00318_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00319_, _00318_, _43998_);
  and (_39323_, _00319_, _00317_);
  nand (_00320_, _43270_, _38659_);
  or (_00321_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00322_, _00321_, _43998_);
  and (_39324_, _00322_, _00320_);
  nand (_00323_, _43270_, _38689_);
  or (_00324_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00325_, _00324_, _43998_);
  and (_39325_, _00325_, _00323_);
  nand (_00326_, _43270_, _38721_);
  or (_00327_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00328_, _00327_, _43998_);
  and (_39327_, _00328_, _00326_);
  nand (_00330_, _43270_, _38777_);
  or (_00331_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00333_, _00331_, _43998_);
  and (_39328_, _00333_, _00330_);
  nand (_00334_, _43270_, _38812_);
  or (_00336_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00337_, _00336_, _43998_);
  and (_39329_, _00337_, _00334_);
  nand (_00339_, _43270_, _38868_);
  or (_00340_, _43270_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00341_, _00340_, _43998_);
  and (_39330_, _00341_, _00339_);
  nor (_39538_, _39819_, rst);
  nor (_00343_, _40207_, _40068_);
  nor (_00345_, _39984_, _39945_);
  not (_00346_, _00345_);
  nor (_00347_, _00346_, _40158_);
  and (_00349_, _00347_, _00343_);
  and (_00350_, _00349_, _39048_);
  and (_00351_, _40158_, _40068_);
  and (_00353_, _00351_, _39983_);
  nor (_00354_, _40207_, _39945_);
  and (_00355_, _00354_, _00353_);
  not (_00357_, _40028_);
  nor (_00358_, _39091_, _39080_);
  and (_00359_, _39091_, _39080_);
  nor (_00360_, _00359_, _00358_);
  nor (_00361_, _39137_, _39106_);
  and (_00362_, _39137_, _39106_);
  nor (_00363_, _00362_, _00361_);
  nor (_00364_, _00363_, _00360_);
  and (_00365_, _00363_, _00360_);
  nor (_00366_, _00365_, _00364_);
  nor (_00367_, _39336_, _39261_);
  and (_00368_, _39336_, _39261_);
  nor (_00369_, _00368_, _00367_);
  not (_00370_, _39069_);
  nor (_00371_, _39347_, _00370_);
  and (_00372_, _39347_, _00370_);
  nor (_00373_, _00372_, _00371_);
  nor (_00374_, _00373_, _00369_);
  and (_00375_, _00373_, _00369_);
  or (_00376_, _00375_, _00374_);
  or (_00377_, _00376_, _00366_);
  nand (_00379_, _00376_, _00366_);
  and (_00380_, _00379_, _00377_);
  or (_00382_, _00380_, _00357_);
  and (_00383_, _39885_, _40119_);
  or (_00384_, _40028_, _39018_);
  and (_00386_, _00384_, _00383_);
  and (_00387_, _00386_, _00382_);
  not (_00388_, _40119_);
  nor (_00390_, _39885_, _00388_);
  and (_00391_, _00357_, _39027_);
  and (_00392_, _40028_, _38964_);
  or (_00394_, _00392_, _00391_);
  and (_00395_, _00394_, _00390_);
  nor (_00396_, _39885_, _40119_);
  and (_00398_, _00396_, _00357_);
  and (_00399_, _00398_, _38955_);
  and (_00400_, _00396_, _40028_);
  and (_00402_, _00400_, _39008_);
  or (_00403_, _00402_, _00399_);
  or (_00404_, _00403_, _00395_);
  or (_00406_, _00357_, _39000_);
  and (_00407_, _39885_, _00388_);
  or (_00408_, _40028_, _39043_);
  and (_00410_, _00408_, _00407_);
  and (_00411_, _00410_, _00406_);
  or (_00412_, _00411_, _00404_);
  or (_00413_, _00412_, _00387_);
  and (_00414_, _00413_, _00355_);
  and (_00415_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_00416_, _00415_, _40028_);
  and (_00417_, _00383_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00418_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_00419_, _00396_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00420_, _00419_, _00418_);
  or (_00421_, _00420_, _00417_);
  or (_00422_, _00421_, _00416_);
  and (_00423_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00424_, _00423_, _00357_);
  and (_00425_, _00396_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00426_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00427_, _00383_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_00428_, _00427_, _00426_);
  or (_00429_, _00428_, _00425_);
  or (_00430_, _00429_, _00424_);
  and (_00432_, _00430_, _00422_);
  or (_00433_, _00432_, _40207_);
  not (_00435_, _40207_);
  and (_00436_, _35992_, _35194_);
  not (_00437_, _00436_);
  nor (_00439_, _36905_, _36568_);
  and (_00440_, _00439_, _00437_);
  and (_00441_, _00440_, _42155_);
  and (_00443_, _00441_, _42484_);
  and (_00444_, _35205_, _36307_);
  nor (_00445_, _00444_, _36383_);
  and (_00447_, _00445_, _42216_);
  and (_00448_, _00447_, _42314_);
  and (_00449_, _00448_, _36807_);
  and (_00451_, _00449_, _00443_);
  nor (_00452_, _00451_, _33169_);
  and (_00453_, _42672_, p3in_reg[5]);
  and (_00455_, _42668_, p3_in[5]);
  or (_00456_, _00455_, _00453_);
  or (_00457_, _00456_, _00452_);
  not (_00459_, _00452_);
  or (_00460_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00461_, _00460_, _00457_);
  and (_00463_, _00461_, _00390_);
  or (_00464_, _00463_, _40028_);
  and (_00465_, _42672_, p3in_reg[4]);
  and (_00466_, _42668_, p3_in[4]);
  or (_00467_, _00466_, _00465_);
  or (_00468_, _00467_, _00452_);
  or (_00469_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00470_, _00469_, _00468_);
  and (_00471_, _00470_, _00383_);
  and (_00472_, _42672_, p3in_reg[6]);
  and (_00473_, _42668_, p3_in[6]);
  or (_00474_, _00473_, _00472_);
  or (_00475_, _00474_, _00452_);
  nand (_00476_, _00452_, _39793_);
  and (_00477_, _00476_, _00475_);
  and (_00478_, _00477_, _00407_);
  and (_00479_, _42672_, p3in_reg[7]);
  and (_00480_, _42668_, p3_in[7]);
  or (_00481_, _00480_, _00479_);
  or (_00482_, _00481_, _00452_);
  nand (_00483_, _00452_, _39400_);
  and (_00485_, _00483_, _00482_);
  and (_00486_, _00485_, _00396_);
  or (_00488_, _00486_, _00478_);
  or (_00489_, _00488_, _00471_);
  or (_00490_, _00489_, _00464_);
  and (_00492_, _42672_, p3in_reg[1]);
  and (_00493_, _42668_, p3_in[1]);
  or (_00494_, _00493_, _00492_);
  or (_00496_, _00494_, _00452_);
  nand (_00497_, _00452_, _39728_);
  and (_00498_, _00497_, _00496_);
  and (_00500_, _00498_, _00390_);
  or (_00501_, _00500_, _00357_);
  and (_00502_, _42672_, p3in_reg[3]);
  and (_00504_, _42668_, p3_in[3]);
  or (_00505_, _00504_, _00502_);
  or (_00506_, _00505_, _00452_);
  or (_00508_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00509_, _00508_, _00506_);
  and (_00510_, _00509_, _00396_);
  and (_00512_, _42672_, p3in_reg[2]);
  and (_00513_, _42668_, p3_in[2]);
  or (_00514_, _00513_, _00512_);
  or (_00516_, _00514_, _00452_);
  nand (_00517_, _00452_, _39739_);
  and (_00518_, _00517_, _00516_);
  and (_00519_, _00518_, _00407_);
  and (_00520_, _42672_, p3in_reg[0]);
  and (_00521_, _42668_, p3_in[0]);
  or (_00522_, _00521_, _00520_);
  or (_00523_, _00522_, _00452_);
  nand (_00524_, _00452_, _39713_);
  and (_00525_, _00524_, _00523_);
  and (_00526_, _00525_, _00383_);
  or (_00527_, _00526_, _00519_);
  or (_00528_, _00527_, _00510_);
  or (_00529_, _00528_, _00501_);
  and (_00530_, _00529_, _00490_);
  or (_00531_, _00530_, _00435_);
  and (_00532_, _40158_, _40069_);
  and (_00533_, _00532_, _00345_);
  and (_00534_, _00533_, _00531_);
  and (_00535_, _00534_, _00433_);
  nor (_00536_, _40207_, _40069_);
  nor (_00538_, _00346_, _00536_);
  nor (_00539_, _00538_, _00355_);
  nor (_00541_, _00539_, _27165_);
  and (_00542_, _00541_, _42708_);
  and (_00543_, _42672_, p1in_reg[5]);
  and (_00545_, _42668_, p1_in[5]);
  or (_00546_, _00545_, _00543_);
  or (_00547_, _00546_, _00452_);
  or (_00549_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00550_, _00549_, _00547_);
  and (_00551_, _00550_, _00390_);
  or (_00553_, _00551_, _40028_);
  and (_00554_, _42672_, p1in_reg[4]);
  and (_00555_, _42668_, p1_in[4]);
  or (_00557_, _00555_, _00554_);
  or (_00558_, _00557_, _00452_);
  or (_00559_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00561_, _00559_, _00558_);
  and (_00562_, _00561_, _00383_);
  and (_00563_, _42672_, p1in_reg[6]);
  and (_00565_, _42668_, p1_in[6]);
  or (_00566_, _00565_, _00563_);
  or (_00567_, _00566_, _00452_);
  nand (_00569_, _00452_, _39594_);
  and (_00570_, _00569_, _00567_);
  and (_00571_, _00570_, _00407_);
  and (_00572_, _42672_, p1in_reg[7]);
  and (_00573_, _42668_, p1_in[7]);
  or (_00574_, _00573_, _00572_);
  or (_00575_, _00574_, _00452_);
  nand (_00576_, _00452_, _39374_);
  and (_00577_, _00576_, _00575_);
  and (_00578_, _00577_, _00396_);
  or (_00579_, _00578_, _00571_);
  or (_00580_, _00579_, _00562_);
  or (_00581_, _00580_, _00553_);
  and (_00582_, _40207_, _39946_);
  and (_00583_, _00582_, _00353_);
  and (_00584_, _42672_, p1in_reg[1]);
  and (_00585_, _42668_, p1_in[1]);
  or (_00586_, _00585_, _00584_);
  or (_00587_, _00586_, _00452_);
  nand (_00588_, _00452_, _39527_);
  and (_00589_, _00588_, _00587_);
  and (_00591_, _00589_, _00390_);
  or (_00592_, _00591_, _00357_);
  and (_00594_, _42672_, p1in_reg[0]);
  and (_00595_, _42668_, p1_in[0]);
  or (_00596_, _00595_, _00594_);
  or (_00598_, _00596_, _00452_);
  nand (_00599_, _00452_, _39514_);
  and (_00600_, _00599_, _00598_);
  and (_00602_, _00600_, _00383_);
  and (_00603_, _42672_, p1in_reg[2]);
  and (_00604_, _42668_, p1_in[2]);
  or (_00606_, _00604_, _00603_);
  or (_00607_, _00606_, _00452_);
  nand (_00608_, _00452_, _39541_);
  and (_00610_, _00608_, _00607_);
  and (_00611_, _00610_, _00407_);
  and (_00612_, _42672_, p1in_reg[3]);
  and (_00614_, _42668_, p1_in[3]);
  or (_00615_, _00614_, _00612_);
  or (_00616_, _00615_, _00452_);
  or (_00618_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00619_, _00618_, _00616_);
  and (_00620_, _00619_, _00396_);
  or (_00622_, _00620_, _00611_);
  or (_00623_, _00622_, _00602_);
  or (_00624_, _00623_, _00592_);
  and (_00625_, _00624_, _00583_);
  and (_00626_, _00625_, _00581_);
  and (_00627_, _42672_, p0in_reg[0]);
  and (_00628_, _42668_, p0_in[0]);
  or (_00629_, _00628_, _00627_);
  or (_00630_, _00629_, _00452_);
  nand (_00631_, _00452_, _39423_);
  and (_00632_, _00631_, _00630_);
  and (_00633_, _00632_, _00383_);
  or (_00634_, _00633_, _00357_);
  and (_00635_, _42672_, p0in_reg[2]);
  and (_00636_, _42668_, p0_in[2]);
  or (_00637_, _00636_, _00635_);
  or (_00638_, _00637_, _00452_);
  nand (_00639_, _00452_, _39451_);
  and (_00640_, _00639_, _00638_);
  and (_00641_, _00640_, _00407_);
  and (_00642_, _42672_, p0in_reg[1]);
  and (_00643_, _42668_, p0_in[1]);
  or (_00644_, _00643_, _00642_);
  or (_00645_, _00644_, _00452_);
  nand (_00646_, _00452_, _39435_);
  and (_00647_, _00646_, _00645_);
  and (_00648_, _00647_, _00390_);
  and (_00649_, _42672_, p0in_reg[3]);
  and (_00650_, _42668_, p0_in[3]);
  or (_00651_, _00650_, _00649_);
  or (_00652_, _00651_, _00452_);
  or (_00653_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00654_, _00653_, _00652_);
  and (_00655_, _00654_, _00396_);
  or (_00656_, _00655_, _00648_);
  or (_00657_, _00656_, _00641_);
  or (_00658_, _00657_, _00634_);
  nor (_00659_, _40158_, _40069_);
  and (_00660_, _00659_, _40207_);
  and (_00661_, _00660_, _00345_);
  and (_00662_, _42672_, p0in_reg[4]);
  and (_00663_, _42668_, p0_in[4]);
  or (_00664_, _00663_, _00662_);
  or (_00665_, _00664_, _00452_);
  or (_00666_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00667_, _00666_, _00665_);
  and (_00668_, _00667_, _00383_);
  or (_00669_, _00668_, _40028_);
  and (_00670_, _42672_, p0in_reg[6]);
  and (_00671_, _42668_, p0_in[6]);
  or (_00672_, _00671_, _00670_);
  or (_00673_, _00672_, _00452_);
  nand (_00674_, _00452_, _39496_);
  and (_00675_, _00674_, _00673_);
  and (_00676_, _00675_, _00407_);
  and (_00677_, _42672_, p0in_reg[5]);
  and (_00678_, _42668_, p0_in[5]);
  or (_00679_, _00678_, _00677_);
  or (_00680_, _00679_, _00452_);
  or (_00681_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_00682_, _00681_, _00680_);
  and (_00683_, _00682_, _00390_);
  and (_00684_, _42672_, p0in_reg[7]);
  and (_00685_, _42668_, p0_in[7]);
  or (_00686_, _00685_, _00684_);
  or (_00687_, _00686_, _00452_);
  nand (_00688_, _00452_, _39360_);
  and (_00689_, _00688_, _00687_);
  and (_00690_, _00689_, _00396_);
  or (_00691_, _00690_, _00683_);
  or (_00692_, _00691_, _00676_);
  or (_00693_, _00692_, _00669_);
  and (_00694_, _00693_, _00661_);
  and (_00695_, _00694_, _00658_);
  or (_00696_, _00695_, _00626_);
  and (_00697_, _42672_, p2in_reg[2]);
  and (_00698_, _42668_, p2_in[2]);
  or (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, _00452_);
  nand (_00701_, _00452_, _39640_);
  and (_00702_, _00701_, _00700_);
  and (_00703_, _00702_, _00407_);
  or (_00704_, _00703_, _00357_);
  and (_00705_, _42672_, p2in_reg[3]);
  and (_00706_, _42668_, p2_in[3]);
  or (_00707_, _00706_, _00705_);
  or (_00708_, _00707_, _00452_);
  or (_00709_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00710_, _00709_, _00708_);
  and (_00711_, _00710_, _00396_);
  and (_00712_, _42672_, p2in_reg[1]);
  and (_00713_, _42668_, p2_in[1]);
  or (_00714_, _00713_, _00712_);
  or (_00715_, _00714_, _00452_);
  nand (_00716_, _00452_, _39620_);
  and (_00717_, _00716_, _00715_);
  and (_00718_, _00717_, _00390_);
  and (_00719_, _42672_, p2in_reg[0]);
  and (_00720_, _42668_, p2_in[0]);
  or (_00721_, _00720_, _00719_);
  or (_00722_, _00721_, _00452_);
  nand (_00723_, _00452_, _39607_);
  and (_00724_, _00723_, _00722_);
  and (_00725_, _00724_, _00383_);
  or (_00726_, _00725_, _00718_);
  or (_00727_, _00726_, _00711_);
  or (_00728_, _00727_, _00704_);
  and (_00729_, _00345_, _40207_);
  nor (_00730_, _40158_, _40068_);
  and (_00731_, _00730_, _00729_);
  and (_00732_, _42672_, p2in_reg[6]);
  and (_00733_, _42668_, p2_in[6]);
  or (_00734_, _00733_, _00732_);
  or (_00735_, _00734_, _00452_);
  nand (_00736_, _00452_, _39693_);
  and (_00737_, _00736_, _00735_);
  and (_00738_, _00737_, _00407_);
  or (_00739_, _00738_, _40028_);
  and (_00740_, _42672_, p2in_reg[4]);
  and (_00741_, _42668_, p2_in[4]);
  or (_00742_, _00741_, _00740_);
  or (_00743_, _00742_, _00452_);
  or (_00744_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00745_, _00744_, _00743_);
  and (_00746_, _00745_, _00383_);
  and (_00747_, _42672_, p2in_reg[5]);
  and (_00748_, _42668_, p2_in[5]);
  or (_00749_, _00748_, _00747_);
  or (_00750_, _00749_, _00452_);
  or (_00751_, _00459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00752_, _00751_, _00750_);
  and (_00753_, _00752_, _00390_);
  and (_00754_, _42672_, p2in_reg[7]);
  and (_00755_, _42668_, p2_in[7]);
  or (_00756_, _00755_, _00754_);
  or (_00757_, _00756_, _00452_);
  nand (_00758_, _00452_, _39392_);
  and (_00759_, _00758_, _00757_);
  and (_00760_, _00759_, _00396_);
  or (_00761_, _00760_, _00753_);
  or (_00762_, _00761_, _00746_);
  or (_00763_, _00762_, _00739_);
  and (_00764_, _00763_, _00731_);
  and (_00765_, _00764_, _00728_);
  and (_00766_, _00383_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00767_, _00766_, _00357_);
  and (_00768_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00769_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00770_, _00396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00771_, _00770_, _00769_);
  or (_00772_, _00771_, _00768_);
  or (_00773_, _00772_, _00767_);
  and (_00774_, _00383_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00775_, _00774_, _40028_);
  and (_00776_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00777_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00778_, _00396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_00779_, _00778_, _00777_);
  or (_00780_, _00779_, _00776_);
  or (_00781_, _00780_, _00775_);
  and (_00782_, _00781_, _00349_);
  and (_00783_, _00782_, _00773_);
  or (_00784_, _00783_, _00765_);
  or (_00785_, _00784_, _00696_);
  or (_00786_, _00785_, _00542_);
  or (_00787_, _00786_, _00535_);
  or (_00788_, _00787_, _00414_);
  nand (_00789_, _00542_, _27790_);
  nand (_00790_, _00789_, _00788_);
  nor (_00791_, _00790_, _00350_);
  or (_00792_, _00357_, _39080_);
  or (_00793_, _40028_, _39261_);
  and (_00794_, _00793_, _00383_);
  and (_00795_, _00794_, _00792_);
  or (_00796_, _40028_, _39336_);
  or (_00797_, _00357_, _39091_);
  and (_00798_, _00797_, _00390_);
  and (_00799_, _00798_, _00796_);
  and (_00800_, _00398_, _39069_);
  not (_00801_, _00400_);
  nor (_00802_, _00801_, _39137_);
  or (_00803_, _00802_, _00800_);
  or (_00804_, _00803_, _00799_);
  or (_00805_, _40028_, _39347_);
  nand (_00806_, _40028_, _39106_);
  and (_00807_, _00806_, _00407_);
  and (_00808_, _00807_, _00805_);
  or (_00809_, _00808_, _00804_);
  or (_00810_, _00809_, _00795_);
  and (_00811_, _00810_, _00350_);
  and (_00812_, _00729_, _00459_);
  not (_00813_, _38950_);
  or (_00814_, _00539_, _00813_);
  nor (_00815_, _00814_, _00812_);
  and (_00816_, _00815_, _42695_);
  or (_00817_, _00816_, _00811_);
  or (_00818_, _00817_, _00791_);
  and (_00819_, _00390_, _40113_);
  or (_00820_, _00819_, _00357_);
  and (_00821_, _00407_, _40001_);
  and (_00822_, _00396_, _39948_);
  and (_00823_, _00383_, _38077_);
  or (_00824_, _00823_, _00822_);
  or (_00825_, _00824_, _00821_);
  or (_00826_, _00825_, _00820_);
  and (_00827_, _00390_, _40033_);
  or (_00828_, _00827_, _40028_);
  and (_00829_, _00407_, _40183_);
  and (_00830_, _00396_, _39920_);
  and (_00831_, _00383_, _40129_);
  or (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00829_);
  or (_00834_, _00833_, _00828_);
  nand (_00835_, _00834_, _00826_);
  nand (_00836_, _00835_, _00816_);
  and (_00837_, _00836_, _43998_);
  and (_39567_, _00837_, _00818_);
  and (_00838_, _39983_, _40028_);
  and (_00839_, _00838_, _00383_);
  and (_00840_, _00839_, _00351_);
  and (_00841_, _00840_, _00354_);
  and (_00842_, _00841_, _38935_);
  and (_00843_, _00661_, _00400_);
  and (_00844_, _00843_, _38499_);
  nor (_00845_, _00844_, _00842_);
  nor (_00846_, _00845_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00847_, _00839_, _00730_);
  and (_00848_, _00847_, _00354_);
  and (_00849_, _00848_, _42762_);
  not (_00850_, _00398_);
  and (_00851_, _00850_, _38946_);
  and (_00852_, _00851_, _42695_);
  or (_00853_, _00852_, _00849_);
  or (_00854_, _00853_, _42710_);
  or (_00855_, _00854_, _00846_);
  and (_00856_, _00582_, _00659_);
  and (_00857_, _00838_, _00407_);
  and (_00858_, _00857_, _00856_);
  and (_00859_, _00858_, _38499_);
  nor (_00860_, _00859_, rst);
  and (_39569_, _00860_, _00855_);
  not (_00861_, _00859_);
  and (_00862_, _00856_, _00839_);
  and (_00863_, _00862_, _00689_);
  and (_00864_, _00840_, _00582_);
  and (_00865_, _00864_, _00577_);
  and (_00866_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_00867_, _00866_, _00865_);
  or (_00868_, _00867_, _00863_);
  and (_00869_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00870_, _00838_, _00390_);
  and (_00871_, _00870_, _00856_);
  and (_00872_, _00871_, _39909_);
  or (_00873_, _00872_, _00869_);
  or (_00874_, _00873_, _00868_);
  and (_00875_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_00876_, _00839_, _00532_);
  and (_00877_, _00876_, _00354_);
  and (_00878_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_00879_, _00847_, _00582_);
  and (_00880_, _00879_, _00759_);
  or (_00881_, _00880_, _00878_);
  and (_00882_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00883_, _00876_, _00582_);
  and (_00884_, _00883_, _00485_);
  or (_00885_, _00884_, _00882_);
  or (_00886_, _00885_, _00881_);
  or (_00887_, _00886_, _00875_);
  nor (_00888_, _00887_, _00874_);
  nor (_00889_, _00888_, _00855_);
  and (_00890_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_00891_, _00890_, _00889_);
  and (_00892_, _00891_, _00861_);
  nor (_00893_, _00861_, _27132_);
  or (_00894_, _00893_, _00892_);
  and (_39570_, _00894_, _43998_);
  and (_00895_, _00841_, _00380_);
  and (_00896_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00897_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00898_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00899_, _00898_, _00897_);
  or (_00900_, _00899_, _00896_);
  and (_00901_, _00871_, _39822_);
  and (_00902_, _00862_, _00632_);
  or (_00903_, _00902_, _00901_);
  or (_00904_, _00903_, _00900_);
  and (_00905_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00906_, _00864_, _00600_);
  and (_00907_, _00879_, _00724_);
  or (_00908_, _00907_, _00906_);
  and (_00909_, _00883_, _00525_);
  or (_00910_, _00909_, _00908_);
  or (_00911_, _00910_, _00905_);
  or (_00912_, _00911_, _00904_);
  or (_00913_, _00912_, _00855_);
  or (_00914_, _00913_, _00895_);
  and (_00915_, _00850_, _42695_);
  and (_00916_, _00915_, _38946_);
  nor (_00917_, _00916_, _42790_);
  and (_00918_, _00848_, _39048_);
  and (_00919_, _00848_, _39045_);
  not (_00920_, _00919_);
  and (_00921_, _00920_, _00845_);
  nor (_00922_, _00921_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_00923_, _00922_, _00918_);
  and (_00924_, _00923_, _00917_);
  or (_00925_, _00924_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_00926_, _00925_, _00914_);
  or (_00927_, _00926_, _00859_);
  nand (_00928_, _00859_, _28372_);
  and (_00929_, _00928_, _43998_);
  and (_39629_, _00929_, _00927_);
  and (_00930_, _00862_, _00647_);
  and (_00931_, _00864_, _00589_);
  and (_00932_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_00933_, _00932_, _00931_);
  or (_00934_, _00933_, _00930_);
  and (_00935_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00936_, _00871_, _40103_);
  or (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _00934_);
  and (_00939_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_00940_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00941_, _00879_, _00717_);
  or (_00942_, _00941_, _00940_);
  and (_00943_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00944_, _00883_, _00498_);
  or (_00945_, _00944_, _00943_);
  or (_00946_, _00945_, _00942_);
  or (_00947_, _00946_, _00939_);
  nor (_00948_, _00947_, _00938_);
  nor (_00949_, _00948_, _00855_);
  and (_00950_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_00951_, _00950_, _00949_);
  and (_00952_, _00951_, _00861_);
  nor (_00953_, _00861_, _29086_);
  or (_00954_, _00953_, _00952_);
  and (_39631_, _00954_, _43998_);
  and (_00955_, _00862_, _00640_);
  and (_00956_, _00864_, _00610_);
  and (_00957_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_00958_, _00957_, _00956_);
  or (_00959_, _00958_, _00955_);
  and (_00960_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00961_, _00871_, _40008_);
  or (_00962_, _00961_, _00960_);
  or (_00963_, _00962_, _00959_);
  and (_00964_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_00965_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00966_, _00879_, _00702_);
  or (_00967_, _00966_, _00965_);
  and (_00968_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00969_, _00883_, _00518_);
  or (_00970_, _00969_, _00968_);
  or (_00971_, _00970_, _00967_);
  or (_00972_, _00971_, _00964_);
  nor (_00973_, _00972_, _00963_);
  nor (_00974_, _00973_, _00855_);
  and (_00975_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_00976_, _00975_, _00974_);
  and (_00977_, _00976_, _00861_);
  nor (_00978_, _00861_, _29763_);
  or (_00979_, _00978_, _00977_);
  and (_39632_, _00979_, _43998_);
  and (_00980_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00981_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00982_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_00983_, _00982_, _00981_);
  or (_00984_, _00983_, _00980_);
  and (_00985_, _00871_, _39978_);
  and (_00986_, _00862_, _00654_);
  or (_00987_, _00986_, _00985_);
  or (_00988_, _00987_, _00984_);
  and (_00989_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_00990_, _00864_, _00619_);
  and (_00991_, _00879_, _00710_);
  or (_00992_, _00991_, _00990_);
  and (_00993_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00994_, _00883_, _00509_);
  or (_00995_, _00994_, _00993_);
  or (_00996_, _00995_, _00992_);
  or (_00997_, _00996_, _00989_);
  nor (_00998_, _00997_, _00988_);
  nor (_00999_, _00998_, _00855_);
  and (_01000_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_01001_, _01000_, _00999_);
  and (_01002_, _01001_, _00861_);
  nor (_01003_, _00861_, _30514_);
  or (_01004_, _01003_, _01002_);
  and (_39633_, _01004_, _43998_);
  and (_01005_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01006_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01007_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_01008_, _01007_, _01006_);
  or (_01009_, _01008_, _01005_);
  and (_01010_, _00871_, _40133_);
  and (_01011_, _00862_, _00667_);
  or (_01012_, _01011_, _01010_);
  or (_01013_, _01012_, _01009_);
  and (_01014_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_01015_, _00864_, _00561_);
  and (_01016_, _00879_, _00745_);
  or (_01017_, _01016_, _01015_);
  and (_01018_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01019_, _00883_, _00470_);
  or (_01020_, _01019_, _01018_);
  or (_01021_, _01020_, _01017_);
  or (_01022_, _01021_, _01014_);
  nor (_01023_, _01022_, _01013_);
  nor (_01024_, _01023_, _00855_);
  and (_01025_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_01026_, _01025_, _01024_);
  and (_01027_, _01026_, _00861_);
  nor (_01028_, _00861_, _31285_);
  or (_01029_, _01028_, _01027_);
  and (_39634_, _01029_, _43998_);
  and (_01030_, _00862_, _00682_);
  and (_01031_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01032_, _00879_, _00752_);
  or (_01033_, _01032_, _01031_);
  or (_01034_, _01033_, _01030_);
  and (_01035_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01036_, _00871_, _40065_);
  or (_01037_, _01036_, _01035_);
  or (_01038_, _01037_, _01034_);
  and (_01039_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01040_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01041_, _00883_, _00461_);
  or (_01043_, _01041_, _01040_);
  and (_01044_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01045_, _00864_, _00550_);
  or (_01046_, _01045_, _01044_);
  or (_01047_, _01046_, _01043_);
  or (_01048_, _01047_, _01039_);
  nor (_01049_, _01048_, _01038_);
  nor (_01050_, _01049_, _00855_);
  and (_01051_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_01052_, _01051_, _01050_);
  and (_01053_, _01052_, _00861_);
  nor (_01054_, _00861_, _32102_);
  or (_01055_, _01054_, _01053_);
  and (_39635_, _01055_, _43998_);
  and (_01056_, _00862_, _00675_);
  and (_01057_, _00864_, _00570_);
  and (_01058_, _00841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_01059_, _01058_, _01057_);
  or (_01060_, _01059_, _01056_);
  and (_01061_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01062_, _00871_, _40172_);
  or (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _01060_);
  and (_01065_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_01066_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01067_, _00879_, _00737_);
  or (_01068_, _01067_, _01066_);
  and (_01069_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01070_, _00883_, _00477_);
  or (_01071_, _01070_, _01069_);
  or (_01073_, _01071_, _01068_);
  or (_01074_, _01073_, _01065_);
  nor (_01075_, _01074_, _01064_);
  nor (_01076_, _01075_, _00855_);
  and (_01077_, _00855_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_01078_, _01077_, _01076_);
  and (_01079_, _01078_, _00861_);
  nor (_01080_, _00861_, _32919_);
  or (_01081_, _01080_, _01079_);
  and (_39636_, _01081_, _43998_);
  and (_39681_, _40219_, _43998_);
  and (_39682_, _40292_, _43998_);
  nor (_39684_, _40028_, rst);
  and (_39699_, _40309_, _43998_);
  and (_39700_, _40322_, _43998_);
  and (_39702_, _40335_, _43998_);
  and (_39703_, _40343_, _43998_);
  and (_39704_, _40353_, _43998_);
  and (_39705_, _40363_, _43998_);
  and (_39706_, _40373_, _43998_);
  nor (_39707_, _39885_, rst);
  nor (_39708_, _40119_, rst);
  not (_01083_, _41561_);
  nor (_01084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01085_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01086_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01085_);
  nor (_01087_, _01086_, _01084_);
  nor (_01088_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01089_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01085_);
  nor (_01090_, _01089_, _01088_);
  nor (_01091_, _01090_, _01087_);
  not (_01092_, _01091_);
  nor (_01093_, _43687_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01094_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01085_);
  nor (_01095_, _01094_, _01093_);
  and (_01096_, _01095_, _01092_);
  nor (_01097_, _01095_, _01092_);
  nor (_01098_, _01097_, _01096_);
  nor (_01099_, _43704_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01100_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01085_);
  nor (_01101_, _01100_, _01099_);
  not (_01102_, _01101_);
  nor (_01103_, _01102_, _01096_);
  and (_01104_, _01102_, _01096_);
  nor (_01105_, _01104_, _01103_);
  nor (_01106_, _01105_, _01098_);
  not (_01107_, _01090_);
  and (_01108_, _01107_, _01087_);
  and (_01109_, _01108_, _01106_);
  and (_01110_, _01109_, _01083_);
  not (_01111_, _41643_);
  and (_01112_, _01090_, _01087_);
  and (_01113_, _01106_, _01112_);
  and (_01114_, _01113_, _01111_);
  not (_01115_, _41602_);
  nor (_01116_, _01107_, _01087_);
  and (_01117_, _01116_, _01106_);
  and (_01118_, _01117_, _01115_);
  or (_01119_, _01118_, _01114_);
  or (_01120_, _01119_, _01110_);
  not (_01121_, _41438_);
  and (_01122_, _01102_, _01098_);
  and (_01123_, _01122_, _01116_);
  and (_01124_, _01123_, _01121_);
  not (_01125_, _41479_);
  and (_01126_, _01122_, _01112_);
  and (_01127_, _01126_, _01125_);
  or (_01128_, _01127_, _01124_);
  not (_01129_, _41395_);
  and (_01130_, _01122_, _01108_);
  and (_01131_, _01130_, _01129_);
  not (_01132_, _41520_);
  and (_01133_, _01095_, _01091_);
  and (_01134_, _01102_, _01133_);
  and (_01135_, _01134_, _01132_);
  not (_01136_, _41354_);
  and (_01137_, _01102_, _01097_);
  and (_01138_, _01137_, _01136_);
  or (_01139_, _01138_, _01135_);
  and (_01140_, _01101_, _01133_);
  and (_01141_, _01140_, _41915_);
  not (_01142_, _41690_);
  and (_01143_, _01101_, _01097_);
  and (_01144_, _01143_, _01142_);
  or (_01145_, _01144_, _01141_);
  or (_01146_, _01145_, _01139_);
  or (_01147_, _01146_, _01131_);
  or (_01148_, _01147_, _01128_);
  not (_01149_, _41289_);
  not (_01150_, _01098_);
  and (_01151_, _01105_, _01150_);
  and (_01152_, _01151_, _01112_);
  and (_01153_, _01152_, _01149_);
  not (_01154_, _41859_);
  and (_01155_, _01103_, _01112_);
  and (_01156_, _01155_, _01154_);
  not (_01157_, _41801_);
  and (_01158_, _01116_, _01103_);
  and (_01159_, _01158_, _01157_);
  or (_01160_, _01159_, _01156_);
  not (_01161_, _41745_);
  and (_01162_, _01108_, _01103_);
  and (_01163_, _01162_, _01161_);
  or (_01164_, _01163_, _01160_);
  or (_01165_, _01164_, _01153_);
  not (_01166_, _41203_);
  and (_01167_, _01151_, _01108_);
  and (_01168_, _01167_, _01166_);
  not (_01169_, _41244_);
  and (_01170_, _01151_, _01116_);
  and (_01171_, _01170_, _01169_);
  or (_01172_, _01171_, _01168_);
  or (_01173_, _01172_, _01165_);
  or (_01174_, _01173_, _01148_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01174_, _01120_);
  and (_01175_, _01167_, _01154_);
  and (_01176_, _01155_, _01161_);
  and (_01177_, _01158_, _01142_);
  or (_01178_, _01177_, _01176_);
  or (_01179_, _01178_, _01175_);
  and (_01180_, _01170_, _41915_);
  and (_01181_, _01117_, _01132_);
  or (_01182_, _01181_, _01180_);
  or (_01183_, _01182_, _01179_);
  and (_01184_, _01126_, _01129_);
  and (_01185_, _01123_, _01136_);
  or (_01186_, _01185_, _01184_);
  and (_01187_, _01134_, _01121_);
  or (_01188_, _01187_, _01186_);
  and (_01189_, _01137_, _01169_);
  and (_01190_, _01109_, _01125_);
  or (_01191_, _01190_, _01189_);
  or (_01192_, _01191_, _01188_);
  or (_01193_, _01192_, _01183_);
  and (_01194_, _01140_, _01157_);
  and (_01195_, _01152_, _01166_);
  and (_01196_, _01130_, _01149_);
  or (_01197_, _01196_, _01195_);
  and (_01198_, _01113_, _01083_);
  and (_01199_, _01143_, _01115_);
  and (_01200_, _01162_, _01111_);
  or (_01201_, _01200_, _01199_);
  or (_01202_, _01201_, _01198_);
  or (_01203_, _01202_, _01197_);
  or (_01204_, _01203_, _01194_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01204_, _01193_);
  and (_01205_, _01167_, _41915_);
  and (_01206_, _01113_, _01115_);
  and (_01207_, _01109_, _01132_);
  or (_01208_, _01207_, _01206_);
  or (_01209_, _01208_, _01205_);
  and (_01210_, _01130_, _01136_);
  and (_01211_, _01143_, _01111_);
  and (_01212_, _01134_, _01125_);
  or (_01213_, _01212_, _01211_);
  and (_01214_, _01140_, _01154_);
  and (_01215_, _01137_, _01149_);
  or (_01216_, _01215_, _01214_);
  or (_01217_, _01216_, _01213_);
  or (_01218_, _01217_, _01210_);
  and (_01219_, _01126_, _01121_);
  and (_01220_, _01123_, _01129_);
  or (_01221_, _01220_, _01219_);
  or (_01222_, _01221_, _01218_);
  and (_01223_, _01170_, _01166_);
  and (_01224_, _01155_, _01157_);
  and (_01225_, _01162_, _01142_);
  and (_01226_, _01158_, _01161_);
  or (_01227_, _01226_, _01225_);
  or (_01228_, _01227_, _01224_);
  or (_01229_, _01228_, _01223_);
  and (_01230_, _01117_, _01083_);
  and (_01231_, _01152_, _01169_);
  or (_01232_, _01231_, _01230_);
  or (_01233_, _01232_, _01229_);
  or (_01234_, _01233_, _01222_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01234_, _01209_);
  and (_01235_, _01167_, _01157_);
  and (_01236_, _01152_, _41915_);
  and (_01237_, _01109_, _01121_);
  or (_01238_, _01237_, _01236_);
  or (_01239_, _01238_, _01235_);
  and (_01240_, _01130_, _01169_);
  and (_01241_, _01134_, _01129_);
  and (_01242_, _01140_, _01161_);
  or (_01243_, _01242_, _01241_);
  and (_01244_, _01137_, _01166_);
  and (_01245_, _01143_, _01083_);
  or (_01246_, _01245_, _01244_);
  or (_01247_, _01246_, _01243_);
  or (_01248_, _01247_, _01240_);
  and (_01249_, _01123_, _01149_);
  and (_01250_, _01126_, _01136_);
  or (_01251_, _01250_, _01249_);
  or (_01252_, _01251_, _01248_);
  and (_01253_, _01113_, _01132_);
  and (_01254_, _01162_, _01115_);
  and (_01255_, _01158_, _01111_);
  and (_01256_, _01155_, _01142_);
  or (_01257_, _01256_, _01255_);
  or (_01258_, _01257_, _01254_);
  or (_01259_, _01258_, _01253_);
  and (_01260_, _01117_, _01125_);
  and (_01261_, _01170_, _01154_);
  or (_01262_, _01261_, _01260_);
  or (_01263_, _01262_, _01259_);
  or (_01264_, _01263_, _01252_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01264_, _01239_);
  not (_01265_, _41607_);
  and (_01266_, _01117_, _01265_);
  not (_01267_, _41648_);
  and (_01268_, _01113_, _01267_);
  not (_01269_, _41566_);
  and (_01270_, _01109_, _01269_);
  or (_01271_, _01270_, _01268_);
  or (_01272_, _01271_, _01266_);
  not (_01273_, _41443_);
  and (_01274_, _01123_, _01273_);
  not (_01275_, _41484_);
  and (_01276_, _01126_, _01275_);
  or (_01277_, _01276_, _01274_);
  not (_01278_, _41400_);
  and (_01279_, _01130_, _01278_);
  not (_01280_, _41525_);
  and (_01281_, _01134_, _01280_);
  not (_01282_, _41359_);
  and (_01283_, _01137_, _01282_);
  or (_01284_, _01283_, _01281_);
  and (_01285_, _01140_, _41922_);
  not (_01286_, _41697_);
  and (_01287_, _01143_, _01286_);
  or (_01288_, _01287_, _01285_);
  or (_01289_, _01288_, _01284_);
  or (_01290_, _01289_, _01279_);
  or (_01291_, _01290_, _01277_);
  not (_01292_, _41752_);
  and (_01293_, _01162_, _01292_);
  not (_01294_, _41808_);
  and (_01295_, _01158_, _01294_);
  not (_01296_, _41866_);
  and (_01297_, _01155_, _01296_);
  or (_01298_, _01297_, _01295_);
  or (_01299_, _01298_, _01293_);
  not (_01300_, _41300_);
  and (_01301_, _01152_, _01300_);
  or (_01302_, _01301_, _01299_);
  not (_01303_, _41208_);
  and (_01304_, _01167_, _01303_);
  not (_01305_, _41249_);
  and (_01306_, _01170_, _01305_);
  or (_01307_, _01306_, _01304_);
  or (_01308_, _01307_, _01302_);
  or (_01309_, _01308_, _01291_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01309_, _01272_);
  not (_01310_, _41612_);
  and (_01311_, _01117_, _01310_);
  not (_01312_, _41653_);
  and (_01313_, _01113_, _01312_);
  not (_01314_, _41571_);
  and (_01315_, _01109_, _01314_);
  or (_01316_, _01315_, _01313_);
  or (_01317_, _01316_, _01311_);
  not (_01318_, _41489_);
  and (_01319_, _01126_, _01318_);
  not (_01320_, _41448_);
  and (_01321_, _01123_, _01320_);
  or (_01322_, _01321_, _01319_);
  not (_01323_, _41405_);
  and (_01324_, _01130_, _01323_);
  not (_01325_, _41530_);
  and (_01326_, _01134_, _01325_);
  not (_01327_, _41364_);
  and (_01328_, _01137_, _01327_);
  or (_01329_, _01328_, _01326_);
  and (_01330_, _01140_, _41929_);
  not (_01331_, _41703_);
  and (_01332_, _01143_, _01331_);
  or (_01333_, _01332_, _01330_);
  or (_01334_, _01333_, _01329_);
  or (_01335_, _01334_, _01324_);
  or (_01336_, _01335_, _01322_);
  not (_01337_, _41759_);
  and (_01338_, _01162_, _01337_);
  not (_01339_, _41816_);
  and (_01340_, _01158_, _01339_);
  not (_01341_, _41873_);
  and (_01342_, _01155_, _01341_);
  or (_01343_, _01342_, _01340_);
  or (_01344_, _01343_, _01338_);
  not (_01345_, _41311_);
  and (_01346_, _01152_, _01345_);
  or (_01347_, _01346_, _01344_);
  not (_01348_, _41213_);
  and (_01349_, _01167_, _01348_);
  not (_01350_, _41254_);
  and (_01351_, _01170_, _01350_);
  or (_01352_, _01351_, _01349_);
  or (_01353_, _01352_, _01347_);
  or (_01354_, _01353_, _01336_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01354_, _01317_);
  not (_01355_, _41617_);
  and (_01356_, _01117_, _01355_);
  not (_01357_, _41658_);
  and (_01358_, _01113_, _01357_);
  not (_01359_, _41576_);
  and (_01360_, _01109_, _01359_);
  or (_01361_, _01360_, _01358_);
  or (_01362_, _01361_, _01356_);
  not (_01363_, _41494_);
  and (_01364_, _01126_, _01363_);
  not (_01365_, _41453_);
  and (_01366_, _01123_, _01365_);
  or (_01367_, _01366_, _01364_);
  not (_01368_, _41411_);
  and (_01369_, _01130_, _01368_);
  not (_01370_, _41535_);
  and (_01371_, _01134_, _01370_);
  not (_01372_, _41369_);
  and (_01373_, _01137_, _01372_);
  or (_01374_, _01373_, _01371_);
  and (_01375_, _01140_, _41936_);
  not (_01376_, _41710_);
  and (_01377_, _01143_, _01376_);
  or (_01378_, _01377_, _01375_);
  or (_01379_, _01378_, _01374_);
  or (_01380_, _01379_, _01369_);
  or (_01381_, _01380_, _01367_);
  not (_01382_, _41766_);
  and (_01383_, _01162_, _01382_);
  not (_01384_, _41822_);
  and (_01385_, _01158_, _01384_);
  not (_01386_, _41880_);
  and (_01387_, _01155_, _01386_);
  or (_01388_, _01387_, _01385_);
  or (_01389_, _01388_, _01383_);
  not (_01390_, _41322_);
  and (_01391_, _01152_, _01390_);
  or (_01392_, _01391_, _01389_);
  not (_01393_, _41218_);
  and (_01394_, _01167_, _01393_);
  not (_01395_, _41259_);
  and (_01396_, _01170_, _01395_);
  or (_01397_, _01396_, _01394_);
  or (_01398_, _01397_, _01392_);
  or (_01399_, _01398_, _01381_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01399_, _01362_);
  not (_01400_, _41581_);
  and (_01401_, _01109_, _01400_);
  not (_01402_, _41664_);
  and (_01403_, _01113_, _01402_);
  not (_01404_, _41622_);
  and (_01405_, _01117_, _01404_);
  or (_01406_, _01405_, _01403_);
  or (_01407_, _01406_, _01401_);
  not (_01408_, _41499_);
  and (_01409_, _01126_, _01408_);
  not (_01410_, _41458_);
  and (_01411_, _01123_, _01410_);
  or (_01412_, _01411_, _01409_);
  not (_01413_, _41416_);
  and (_01414_, _01130_, _01413_);
  not (_01415_, _41540_);
  and (_01416_, _01134_, _01415_);
  not (_01417_, _41374_);
  and (_01418_, _01137_, _01417_);
  or (_01419_, _01418_, _01416_);
  and (_01420_, _01140_, _41943_);
  not (_01421_, _41717_);
  and (_01422_, _01143_, _01421_);
  or (_01423_, _01422_, _01420_);
  or (_01424_, _01423_, _01419_);
  or (_01425_, _01424_, _01414_);
  or (_01426_, _01425_, _01412_);
  not (_01427_, _41333_);
  and (_01428_, _01152_, _01427_);
  not (_01429_, _41773_);
  and (_01430_, _01162_, _01429_);
  not (_01431_, _41829_);
  and (_01432_, _01158_, _01431_);
  not (_01433_, _41887_);
  and (_01434_, _01155_, _01433_);
  or (_01435_, _01434_, _01432_);
  or (_01436_, _01435_, _01430_);
  or (_01437_, _01436_, _01428_);
  not (_01438_, _41223_);
  and (_01439_, _01167_, _01438_);
  not (_01440_, _41264_);
  and (_01441_, _01170_, _01440_);
  or (_01442_, _01441_, _01439_);
  or (_01443_, _01442_, _01437_);
  or (_01444_, _01443_, _01426_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01444_, _01407_);
  not (_01445_, _41586_);
  and (_01446_, _01109_, _01445_);
  not (_01447_, _41338_);
  and (_01448_, _01152_, _01447_);
  not (_01449_, _41627_);
  and (_01450_, _01117_, _01449_);
  or (_01451_, _01450_, _01448_);
  or (_01452_, _01451_, _01446_);
  not (_01453_, _41504_);
  and (_01454_, _01126_, _01453_);
  not (_01455_, _41379_);
  and (_01456_, _01137_, _01455_);
  not (_01457_, _41545_);
  and (_01458_, _01134_, _01457_);
  or (_01459_, _01458_, _01456_);
  and (_01460_, _01140_, _41950_);
  not (_01461_, _41724_);
  and (_01462_, _01143_, _01461_);
  or (_01463_, _01462_, _01460_);
  or (_01464_, _01463_, _01459_);
  or (_01465_, _01464_, _01454_);
  not (_01466_, _41463_);
  and (_01467_, _01123_, _01466_);
  not (_01468_, _41422_);
  and (_01469_, _01130_, _01468_);
  or (_01470_, _01469_, _01467_);
  or (_01471_, _01470_, _01465_);
  not (_01472_, _41670_);
  and (_01473_, _01113_, _01472_);
  not (_01474_, _41894_);
  and (_01475_, _01155_, _01474_);
  not (_01476_, _41836_);
  and (_01477_, _01158_, _01476_);
  not (_01478_, _41780_);
  and (_01479_, _01162_, _01478_);
  or (_01480_, _01479_, _01477_);
  or (_01481_, _01480_, _01475_);
  or (_01482_, _01481_, _01473_);
  not (_01483_, _41228_);
  and (_01484_, _01167_, _01483_);
  not (_01485_, _41269_);
  and (_01486_, _01170_, _01485_);
  or (_01487_, _01486_, _01484_);
  or (_01488_, _01487_, _01482_);
  or (_01489_, _01488_, _01471_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01489_, _01452_);
  not (_01490_, _41632_);
  and (_01491_, _01117_, _01490_);
  not (_01492_, _41677_);
  and (_01493_, _01113_, _01492_);
  not (_01494_, _41591_);
  and (_01495_, _01109_, _01494_);
  or (_01496_, _01495_, _01493_);
  or (_01497_, _01496_, _01491_);
  not (_01498_, _41509_);
  and (_01499_, _01126_, _01498_);
  not (_01500_, _41550_);
  and (_01501_, _01134_, _01500_);
  not (_01502_, _41384_);
  and (_01503_, _01137_, _01502_);
  or (_01504_, _01503_, _01501_);
  and (_01505_, _01140_, _41957_);
  not (_01506_, _41730_);
  and (_01507_, _01143_, _01506_);
  or (_01508_, _01507_, _01505_);
  or (_01509_, _01508_, _01504_);
  or (_01510_, _01509_, _01499_);
  not (_01511_, _41468_);
  and (_01512_, _01123_, _01511_);
  not (_01513_, _41427_);
  and (_01514_, _01130_, _01513_);
  or (_01515_, _01514_, _01512_);
  or (_01516_, _01515_, _01510_);
  not (_01517_, _41343_);
  and (_01518_, _01152_, _01517_);
  not (_01519_, _41844_);
  and (_01520_, _01158_, _01519_);
  not (_01521_, _41901_);
  and (_01522_, _01155_, _01521_);
  not (_01523_, _41787_);
  and (_01524_, _01162_, _01523_);
  or (_01525_, _01524_, _01522_);
  or (_01526_, _01525_, _01520_);
  or (_01527_, _01526_, _01518_);
  not (_01528_, _41233_);
  and (_01529_, _01167_, _01528_);
  not (_01530_, _41274_);
  and (_01531_, _01170_, _01530_);
  or (_01532_, _01531_, _01529_);
  or (_01533_, _01532_, _01527_);
  or (_01534_, _01533_, _01516_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01534_, _01497_);
  not (_01535_, _41637_);
  and (_01536_, _01117_, _01535_);
  not (_01537_, _41683_);
  and (_01538_, _01113_, _01537_);
  not (_01539_, _41596_);
  and (_01540_, _01109_, _01539_);
  or (_01541_, _01540_, _01538_);
  or (_01542_, _01541_, _01536_);
  not (_01543_, _41514_);
  and (_01544_, _01126_, _01543_);
  not (_01545_, _41473_);
  and (_01546_, _01123_, _01545_);
  or (_01547_, _01546_, _01544_);
  not (_01548_, _41432_);
  and (_01549_, _01130_, _01548_);
  not (_01550_, _41555_);
  and (_01551_, _01134_, _01550_);
  not (_01552_, _41389_);
  and (_01553_, _01137_, _01552_);
  or (_01554_, _01553_, _01551_);
  and (_01555_, _01140_, _41964_);
  not (_01556_, _41737_);
  and (_01557_, _01143_, _01556_);
  or (_01558_, _01557_, _01555_);
  or (_01559_, _01558_, _01554_);
  or (_01560_, _01559_, _01549_);
  or (_01561_, _01560_, _01547_);
  not (_01562_, _41348_);
  and (_01563_, _01152_, _01562_);
  not (_01564_, _41850_);
  and (_01565_, _01158_, _01564_);
  not (_01566_, _41907_);
  and (_01567_, _01155_, _01566_);
  not (_01568_, _41793_);
  and (_01569_, _01162_, _01568_);
  or (_01570_, _01569_, _01567_);
  or (_01571_, _01570_, _01565_);
  or (_01572_, _01571_, _01563_);
  not (_01573_, _41238_);
  and (_01574_, _01167_, _01573_);
  not (_01575_, _41279_);
  and (_01576_, _01170_, _01575_);
  or (_01577_, _01576_, _01574_);
  or (_01578_, _01577_, _01572_);
  or (_01579_, _01578_, _01561_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01579_, _01542_);
  and (_01580_, _01117_, _01280_);
  and (_01581_, _01170_, _41922_);
  and (_01582_, _01152_, _01303_);
  or (_01583_, _01582_, _01581_);
  or (_01584_, _01583_, _01580_);
  and (_01585_, _01126_, _01278_);
  and (_01586_, _01143_, _01265_);
  and (_01587_, _01140_, _01294_);
  or (_01588_, _01587_, _01586_);
  and (_01589_, _01134_, _01273_);
  and (_01590_, _01137_, _01305_);
  or (_01591_, _01590_, _01589_);
  or (_01592_, _01591_, _01588_);
  or (_01593_, _01592_, _01585_);
  and (_01594_, _01123_, _01282_);
  and (_01595_, _01130_, _01300_);
  or (_01596_, _01595_, _01594_);
  or (_01597_, _01596_, _01593_);
  and (_01598_, _01113_, _01269_);
  and (_01599_, _01162_, _01267_);
  and (_01600_, _01155_, _01292_);
  and (_01601_, _01158_, _01286_);
  or (_01602_, _01601_, _01600_);
  or (_01603_, _01602_, _01599_);
  or (_01604_, _01603_, _01598_);
  and (_01605_, _01167_, _01296_);
  and (_01606_, _01109_, _01275_);
  or (_01607_, _01606_, _01605_);
  or (_01608_, _01607_, _01604_);
  or (_01609_, _01608_, _01597_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01609_, _01584_);
  and (_01610_, _01170_, _41929_);
  and (_01611_, _01167_, _01341_);
  and (_01612_, _01109_, _01318_);
  or (_01613_, _01612_, _01611_);
  or (_01614_, _01613_, _01610_);
  and (_01615_, _01123_, _01327_);
  and (_01616_, _01143_, _01310_);
  and (_01617_, _01134_, _01320_);
  or (_01618_, _01617_, _01616_);
  and (_01619_, _01140_, _01339_);
  and (_01620_, _01137_, _01350_);
  or (_01621_, _01620_, _01619_);
  or (_01622_, _01621_, _01618_);
  or (_01623_, _01622_, _01615_);
  and (_01624_, _01130_, _01345_);
  and (_01625_, _01126_, _01323_);
  or (_01626_, _01625_, _01624_);
  or (_01627_, _01626_, _01623_);
  and (_01628_, _01117_, _01325_);
  and (_01629_, _01158_, _01331_);
  and (_01630_, _01155_, _01337_);
  and (_01631_, _01162_, _01312_);
  or (_01632_, _01631_, _01630_);
  or (_01633_, _01632_, _01629_);
  or (_01634_, _01633_, _01628_);
  and (_01635_, _01113_, _01314_);
  and (_01636_, _01152_, _01348_);
  or (_01637_, _01636_, _01635_);
  or (_01638_, _01637_, _01634_);
  or (_01639_, _01638_, _01627_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01639_, _01614_);
  and (_01640_, _01158_, _01376_);
  and (_01641_, _01155_, _01382_);
  or (_01642_, _01641_, _01640_);
  and (_01643_, _01167_, _01386_);
  or (_01644_, _01643_, _01642_);
  and (_01645_, _01117_, _01370_);
  and (_01646_, _01170_, _41936_);
  or (_01647_, _01646_, _01645_);
  or (_01648_, _01647_, _01644_);
  and (_01649_, _01134_, _01365_);
  and (_01650_, _01123_, _01372_);
  and (_01651_, _01126_, _01368_);
  or (_01652_, _01651_, _01650_);
  or (_01653_, _01652_, _01649_);
  and (_01654_, _01137_, _01395_);
  and (_01655_, _01109_, _01363_);
  or (_01656_, _01655_, _01654_);
  or (_01657_, _01656_, _01653_);
  or (_01658_, _01657_, _01648_);
  and (_01659_, _01140_, _01384_);
  and (_01660_, _01152_, _01393_);
  and (_01661_, _01130_, _01390_);
  or (_01662_, _01661_, _01660_);
  and (_01663_, _01113_, _01359_);
  and (_01664_, _01143_, _01355_);
  and (_01665_, _01162_, _01357_);
  or (_01666_, _01665_, _01664_);
  or (_01667_, _01666_, _01663_);
  or (_01668_, _01667_, _01662_);
  or (_01669_, _01668_, _01659_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01669_, _01658_);
  and (_01670_, _01158_, _01421_);
  and (_01671_, _01155_, _01429_);
  or (_01672_, _01671_, _01670_);
  and (_01673_, _01167_, _01433_);
  or (_01674_, _01673_, _01672_);
  and (_01675_, _01113_, _01400_);
  and (_01676_, _01170_, _41943_);
  or (_01677_, _01676_, _01675_);
  or (_01678_, _01677_, _01674_);
  and (_01679_, _01134_, _01410_);
  and (_01680_, _01123_, _01417_);
  and (_01681_, _01126_, _01413_);
  or (_01682_, _01681_, _01680_);
  or (_01683_, _01682_, _01679_);
  and (_01684_, _01137_, _01440_);
  and (_01685_, _01109_, _01408_);
  or (_01686_, _01685_, _01684_);
  or (_01687_, _01686_, _01683_);
  or (_01688_, _01687_, _01678_);
  and (_01689_, _01140_, _01431_);
  and (_01690_, _01152_, _01438_);
  and (_01691_, _01130_, _01427_);
  or (_01692_, _01691_, _01690_);
  and (_01693_, _01117_, _01415_);
  and (_01694_, _01143_, _01404_);
  and (_01695_, _01162_, _01402_);
  or (_01696_, _01695_, _01694_);
  or (_01697_, _01696_, _01693_);
  or (_01698_, _01697_, _01692_);
  or (_01699_, _01698_, _01689_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01699_, _01688_);
  and (_01700_, _01158_, _01461_);
  and (_01701_, _01155_, _01478_);
  or (_01702_, _01701_, _01700_);
  and (_01703_, _01167_, _01474_);
  or (_01704_, _01703_, _01702_);
  and (_01705_, _01113_, _01445_);
  and (_01706_, _01170_, _41950_);
  or (_01707_, _01706_, _01705_);
  or (_01708_, _01707_, _01704_);
  and (_01709_, _01134_, _01466_);
  and (_01710_, _01123_, _01455_);
  and (_01711_, _01126_, _01468_);
  or (_01712_, _01711_, _01710_);
  or (_01713_, _01712_, _01709_);
  and (_01714_, _01137_, _01485_);
  and (_01715_, _01109_, _01453_);
  or (_01716_, _01715_, _01714_);
  or (_01717_, _01716_, _01713_);
  or (_01718_, _01717_, _01708_);
  and (_01719_, _01140_, _01476_);
  and (_01720_, _01152_, _01483_);
  and (_01721_, _01130_, _01447_);
  or (_01722_, _01721_, _01720_);
  and (_01723_, _01117_, _01457_);
  and (_01724_, _01143_, _01449_);
  and (_01725_, _01162_, _01472_);
  or (_01726_, _01725_, _01724_);
  or (_01727_, _01726_, _01723_);
  or (_01728_, _01727_, _01722_);
  or (_01729_, _01728_, _01719_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01729_, _01718_);
  and (_01730_, _01158_, _01506_);
  and (_01731_, _01155_, _01523_);
  or (_01732_, _01731_, _01730_);
  and (_01733_, _01167_, _01521_);
  or (_01734_, _01733_, _01732_);
  and (_01735_, _01113_, _01494_);
  and (_01736_, _01170_, _41957_);
  or (_01737_, _01736_, _01735_);
  or (_01738_, _01737_, _01734_);
  and (_01739_, _01134_, _01511_);
  and (_01740_, _01123_, _01502_);
  and (_01741_, _01126_, _01513_);
  or (_01742_, _01741_, _01740_);
  or (_01743_, _01742_, _01739_);
  and (_01744_, _01137_, _01530_);
  and (_01745_, _01109_, _01498_);
  or (_01746_, _01745_, _01744_);
  or (_01747_, _01746_, _01743_);
  or (_01748_, _01747_, _01738_);
  and (_01749_, _01140_, _01519_);
  and (_01750_, _01152_, _01528_);
  and (_01751_, _01130_, _01517_);
  or (_01752_, _01751_, _01750_);
  and (_01753_, _01117_, _01500_);
  and (_01754_, _01143_, _01490_);
  and (_01755_, _01162_, _01492_);
  or (_01756_, _01755_, _01754_);
  or (_01757_, _01756_, _01753_);
  or (_01758_, _01757_, _01752_);
  or (_01759_, _01758_, _01749_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01759_, _01748_);
  and (_01760_, _01167_, _01566_);
  and (_01761_, _01170_, _41964_);
  and (_01762_, _01152_, _01573_);
  or (_01763_, _01762_, _01761_);
  or (_01764_, _01763_, _01760_);
  and (_01765_, _01123_, _01552_);
  and (_01766_, _01126_, _01548_);
  or (_01767_, _01766_, _01765_);
  and (_01768_, _01130_, _01562_);
  and (_01769_, _01134_, _01545_);
  and (_01770_, _01137_, _01575_);
  or (_01771_, _01770_, _01769_);
  and (_01772_, _01143_, _01535_);
  and (_01773_, _01140_, _01564_);
  or (_01774_, _01773_, _01772_);
  or (_01775_, _01774_, _01771_);
  or (_01776_, _01775_, _01768_);
  or (_01777_, _01776_, _01767_);
  and (_01778_, _01117_, _01550_);
  and (_01779_, _01113_, _01539_);
  or (_01780_, _01779_, _01778_);
  and (_01781_, _01109_, _01543_);
  and (_01782_, _01155_, _01568_);
  and (_01783_, _01162_, _01537_);
  and (_01784_, _01158_, _01556_);
  or (_01785_, _01784_, _01783_);
  or (_01786_, _01785_, _01782_);
  or (_01787_, _01786_, _01781_);
  or (_01788_, _01787_, _01780_);
  or (_01789_, _01788_, _01777_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01789_, _01764_);
  and (_01790_, _01113_, _01265_);
  and (_01791_, _01170_, _01303_);
  and (_01792_, _01117_, _01269_);
  or (_01793_, _01792_, _01791_);
  or (_01794_, _01793_, _01790_);
  and (_01795_, _01123_, _01278_);
  and (_01796_, _01134_, _01275_);
  and (_01797_, _01137_, _01300_);
  or (_01798_, _01797_, _01796_);
  and (_01799_, _01143_, _01267_);
  and (_01800_, _01140_, _01296_);
  or (_01801_, _01800_, _01799_);
  or (_01802_, _01801_, _01798_);
  or (_01803_, _01802_, _01795_);
  and (_01804_, _01126_, _01273_);
  and (_01805_, _01130_, _01282_);
  or (_01806_, _01805_, _01804_);
  or (_01807_, _01806_, _01803_);
  and (_01808_, _01109_, _01280_);
  and (_01809_, _01155_, _01294_);
  and (_01810_, _01158_, _01292_);
  and (_01811_, _01162_, _01286_);
  or (_01812_, _01811_, _01810_);
  or (_01813_, _01812_, _01809_);
  or (_01814_, _01813_, _01808_);
  and (_01815_, _01167_, _41922_);
  and (_01816_, _01152_, _01305_);
  or (_01817_, _01816_, _01815_);
  or (_01818_, _01817_, _01814_);
  or (_01819_, _01818_, _01807_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01819_, _01794_);
  and (_01820_, _01152_, _01350_);
  and (_01821_, _01170_, _01348_);
  and (_01822_, _01113_, _01310_);
  or (_01823_, _01822_, _01821_);
  or (_01824_, _01823_, _01820_);
  and (_01825_, _01123_, _01323_);
  and (_01826_, _01134_, _01318_);
  and (_01827_, _01140_, _01341_);
  or (_01828_, _01827_, _01826_);
  and (_01829_, _01137_, _01345_);
  and (_01830_, _01143_, _01312_);
  or (_01831_, _01830_, _01829_);
  or (_01832_, _01831_, _01828_);
  or (_01833_, _01832_, _01825_);
  and (_01834_, _01126_, _01320_);
  and (_01835_, _01130_, _01327_);
  or (_01836_, _01835_, _01834_);
  or (_01837_, _01836_, _01833_);
  and (_01838_, _01117_, _01314_);
  and (_01839_, _01155_, _01339_);
  and (_01840_, _01158_, _01337_);
  and (_01841_, _01162_, _01331_);
  or (_01842_, _01841_, _01840_);
  or (_01843_, _01842_, _01839_);
  or (_01844_, _01843_, _01838_);
  and (_01845_, _01167_, _41929_);
  and (_01846_, _01109_, _01325_);
  or (_01847_, _01846_, _01845_);
  or (_01848_, _01847_, _01844_);
  or (_01849_, _01848_, _01837_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01849_, _01824_);
  and (_01850_, _01167_, _41936_);
  and (_01851_, _01113_, _01355_);
  and (_01852_, _01109_, _01370_);
  or (_01853_, _01852_, _01851_);
  or (_01854_, _01853_, _01850_);
  and (_01855_, _01130_, _01372_);
  and (_01856_, _01143_, _01357_);
  and (_01857_, _01134_, _01363_);
  or (_01858_, _01857_, _01856_);
  and (_01859_, _01140_, _01386_);
  and (_01860_, _01137_, _01390_);
  or (_01861_, _01860_, _01859_);
  or (_01862_, _01861_, _01858_);
  or (_01863_, _01862_, _01855_);
  and (_01864_, _01126_, _01365_);
  and (_01865_, _01123_, _01368_);
  or (_01866_, _01865_, _01864_);
  or (_01867_, _01866_, _01863_);
  and (_01868_, _01170_, _01393_);
  and (_01869_, _01155_, _01384_);
  and (_01870_, _01162_, _01376_);
  and (_01871_, _01158_, _01382_);
  or (_01872_, _01871_, _01870_);
  or (_01873_, _01872_, _01869_);
  or (_01874_, _01873_, _01868_);
  and (_01875_, _01117_, _01359_);
  and (_01876_, _01152_, _01395_);
  or (_01877_, _01876_, _01875_);
  or (_01878_, _01877_, _01874_);
  or (_01879_, _01878_, _01867_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01879_, _01854_);
  and (_01880_, _01167_, _41943_);
  and (_01881_, _01170_, _01438_);
  and (_01882_, _01109_, _01415_);
  or (_01883_, _01882_, _01881_);
  or (_01884_, _01883_, _01880_);
  and (_01885_, _01123_, _01413_);
  and (_01886_, _01130_, _01417_);
  or (_01887_, _01886_, _01885_);
  and (_01888_, _01126_, _01410_);
  and (_01889_, _01134_, _01408_);
  and (_01890_, _01140_, _01433_);
  or (_01891_, _01890_, _01889_);
  and (_01892_, _01137_, _01427_);
  and (_01893_, _01143_, _01402_);
  or (_01894_, _01893_, _01892_);
  or (_01895_, _01894_, _01891_);
  or (_01896_, _01895_, _01888_);
  or (_01897_, _01896_, _01887_);
  and (_01898_, _01113_, _01404_);
  and (_01899_, _01155_, _01431_);
  and (_01900_, _01158_, _01429_);
  and (_01901_, _01162_, _01421_);
  or (_01902_, _01901_, _01900_);
  or (_01903_, _01902_, _01899_);
  or (_01904_, _01903_, _01898_);
  and (_01905_, _01152_, _01440_);
  and (_01906_, _01117_, _01400_);
  or (_01907_, _01906_, _01905_);
  or (_01908_, _01907_, _01904_);
  or (_01909_, _01908_, _01897_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01909_, _01884_);
  and (_01910_, _01113_, _01449_);
  and (_01911_, _01167_, _41950_);
  and (_01912_, _01170_, _01483_);
  or (_01913_, _01912_, _01911_);
  or (_01914_, _01913_, _01910_);
  and (_01915_, _01123_, _01468_);
  and (_01916_, _01134_, _01453_);
  and (_01917_, _01137_, _01447_);
  or (_01918_, _01917_, _01916_);
  and (_01919_, _01140_, _01474_);
  and (_01920_, _01143_, _01472_);
  or (_01921_, _01920_, _01919_);
  or (_01922_, _01921_, _01918_);
  or (_01923_, _01922_, _01915_);
  and (_01924_, _01126_, _01466_);
  and (_01925_, _01130_, _01455_);
  or (_01926_, _01925_, _01924_);
  or (_01927_, _01926_, _01923_);
  and (_01928_, _01117_, _01445_);
  and (_01929_, _01155_, _01476_);
  and (_01930_, _01158_, _01478_);
  and (_01931_, _01162_, _01461_);
  or (_01932_, _01931_, _01930_);
  or (_01933_, _01932_, _01929_);
  or (_01934_, _01933_, _01928_);
  and (_01935_, _01152_, _01485_);
  and (_01936_, _01109_, _01457_);
  or (_01937_, _01936_, _01935_);
  or (_01938_, _01937_, _01934_);
  or (_01939_, _01938_, _01927_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01939_, _01914_);
  and (_01940_, _01117_, _01494_);
  and (_01941_, _01113_, _01490_);
  and (_01942_, _01109_, _01500_);
  or (_01943_, _01942_, _01941_);
  or (_01944_, _01943_, _01940_);
  and (_01945_, _01123_, _01513_);
  and (_01946_, _01143_, _01492_);
  and (_01947_, _01134_, _01498_);
  or (_01948_, _01947_, _01946_);
  and (_01949_, _01140_, _01521_);
  and (_01950_, _01137_, _01517_);
  or (_01951_, _01950_, _01949_);
  or (_01952_, _01951_, _01948_);
  or (_01953_, _01952_, _01945_);
  and (_01954_, _01126_, _01511_);
  and (_01955_, _01130_, _01502_);
  or (_01956_, _01955_, _01954_);
  or (_01957_, _01956_, _01953_);
  and (_01958_, _01167_, _41957_);
  and (_01959_, _01155_, _01519_);
  and (_01960_, _01162_, _01506_);
  and (_01961_, _01158_, _01523_);
  or (_01962_, _01961_, _01960_);
  or (_01963_, _01962_, _01959_);
  or (_01964_, _01963_, _01958_);
  and (_01965_, _01170_, _01528_);
  and (_01966_, _01152_, _01530_);
  or (_01967_, _01966_, _01965_);
  or (_01968_, _01967_, _01964_);
  or (_01969_, _01968_, _01957_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01969_, _01944_);
  and (_01970_, _01113_, _01535_);
  and (_01971_, _01170_, _01573_);
  and (_01972_, _01117_, _01539_);
  or (_01973_, _01972_, _01971_);
  or (_01974_, _01973_, _01970_);
  and (_01975_, _01123_, _01548_);
  and (_01976_, _01134_, _01543_);
  and (_01977_, _01137_, _01562_);
  or (_01978_, _01977_, _01976_);
  and (_01979_, _01143_, _01537_);
  and (_01980_, _01140_, _01566_);
  or (_01981_, _01980_, _01979_);
  or (_01982_, _01981_, _01978_);
  or (_01983_, _01982_, _01975_);
  and (_01984_, _01126_, _01545_);
  and (_01985_, _01130_, _01552_);
  or (_01986_, _01985_, _01984_);
  or (_01987_, _01986_, _01983_);
  and (_01988_, _01109_, _01550_);
  and (_01989_, _01155_, _01564_);
  and (_01990_, _01158_, _01568_);
  and (_01991_, _01162_, _01556_);
  or (_01992_, _01991_, _01990_);
  or (_01993_, _01992_, _01989_);
  or (_01994_, _01993_, _01988_);
  and (_01995_, _01167_, _41964_);
  and (_01996_, _01152_, _01575_);
  or (_01997_, _01996_, _01995_);
  or (_01998_, _01997_, _01994_);
  or (_01999_, _01998_, _01987_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _01999_, _01974_);
  and (_02000_, _01143_, _01269_);
  and (_02001_, _01162_, _01265_);
  and (_02002_, _01158_, _01267_);
  or (_02003_, _02002_, _02001_);
  or (_02004_, _02003_, _02000_);
  and (_02005_, _01167_, _01294_);
  and (_02006_, _01113_, _01280_);
  or (_02007_, _02006_, _02005_);
  or (_02008_, _02007_, _02004_);
  and (_02009_, _01117_, _01275_);
  and (_02010_, _01130_, _01305_);
  and (_02011_, _01123_, _01300_);
  and (_02012_, _01137_, _01303_);
  or (_02013_, _02012_, _02011_);
  or (_02014_, _02013_, _02010_);
  or (_02015_, _02014_, _02009_);
  or (_02016_, _02015_, _02008_);
  and (_02017_, _01155_, _01286_);
  and (_02018_, _01152_, _41922_);
  and (_02019_, _01170_, _01296_);
  or (_02020_, _02019_, _02018_);
  or (_02021_, _02020_, _02017_);
  and (_02022_, _01140_, _01292_);
  and (_02023_, _01109_, _01273_);
  and (_02024_, _01134_, _01278_);
  and (_02025_, _01126_, _01282_);
  or (_02026_, _02025_, _02024_);
  or (_02027_, _02026_, _02023_);
  or (_02028_, _02027_, _02022_);
  or (_02029_, _02028_, _02021_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02029_, _02016_);
  and (_02030_, _01170_, _01341_);
  and (_02031_, _01117_, _01318_);
  and (_02032_, _01109_, _01320_);
  or (_02033_, _02032_, _02031_);
  or (_02034_, _02033_, _02030_);
  and (_02035_, _01123_, _01345_);
  and (_02036_, _01140_, _01337_);
  and (_02037_, _01134_, _01323_);
  or (_02038_, _02037_, _02036_);
  and (_02039_, _01143_, _01314_);
  and (_02040_, _01137_, _01348_);
  or (_02041_, _02040_, _02039_);
  or (_02042_, _02041_, _02038_);
  or (_02043_, _02042_, _02035_);
  and (_02044_, _01130_, _01350_);
  and (_02045_, _01126_, _01327_);
  or (_02046_, _02045_, _02044_);
  or (_02047_, _02046_, _02043_);
  and (_02048_, _01113_, _01325_);
  and (_02049_, _01162_, _01310_);
  and (_02050_, _01155_, _01331_);
  and (_02051_, _01158_, _01312_);
  or (_02052_, _02051_, _02050_);
  or (_02053_, _02052_, _02049_);
  or (_02054_, _02053_, _02048_);
  and (_02055_, _01152_, _41929_);
  and (_02056_, _01167_, _01339_);
  or (_02057_, _02056_, _02055_);
  or (_02058_, _02057_, _02054_);
  or (_02059_, _02058_, _02047_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02059_, _02034_);
  and (_02060_, _01167_, _01384_);
  and (_02061_, _01109_, _01365_);
  and (_02062_, _01113_, _01370_);
  or (_02063_, _02062_, _02061_);
  or (_02064_, _02063_, _02060_);
  and (_02065_, _01130_, _01395_);
  and (_02066_, _01123_, _01390_);
  or (_02067_, _02066_, _02065_);
  and (_02068_, _01126_, _01372_);
  and (_02069_, _01137_, _01393_);
  and (_02070_, _01134_, _01368_);
  or (_02071_, _02070_, _02069_);
  and (_02072_, _01143_, _01359_);
  and (_02073_, _01140_, _01382_);
  or (_02074_, _02073_, _02072_);
  or (_02075_, _02074_, _02071_);
  or (_02076_, _02075_, _02068_);
  or (_02077_, _02076_, _02067_);
  and (_02078_, _01152_, _41936_);
  and (_02079_, _01162_, _01355_);
  and (_02080_, _01158_, _01357_);
  and (_02081_, _01155_, _01376_);
  or (_02082_, _02081_, _02080_);
  or (_02083_, _02082_, _02079_);
  or (_02084_, _02083_, _02078_);
  and (_02085_, _01117_, _01363_);
  and (_02086_, _01170_, _01386_);
  or (_02087_, _02086_, _02085_);
  or (_02088_, _02087_, _02084_);
  or (_02089_, _02088_, _02077_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02089_, _02064_);
  and (_02090_, _01113_, _01415_);
  and (_02091_, _01158_, _01402_);
  and (_02092_, _01162_, _01404_);
  or (_02093_, _02092_, _02091_);
  or (_02094_, _02093_, _02090_);
  and (_02095_, _01143_, _01400_);
  and (_02096_, _01155_, _01421_);
  or (_02097_, _02096_, _02095_);
  or (_02098_, _02097_, _02094_);
  and (_02099_, _01117_, _01408_);
  and (_02100_, _01130_, _01440_);
  and (_02101_, _01123_, _01427_);
  and (_02102_, _01137_, _01438_);
  or (_02103_, _02102_, _02101_);
  or (_02104_, _02103_, _02100_);
  or (_02105_, _02104_, _02099_);
  or (_02106_, _02105_, _02098_);
  and (_02107_, _01152_, _41943_);
  and (_02108_, _01167_, _01431_);
  and (_02109_, _01170_, _01433_);
  or (_02110_, _02109_, _02108_);
  or (_02111_, _02110_, _02107_);
  and (_02112_, _01140_, _01429_);
  and (_02113_, _01109_, _01410_);
  and (_02114_, _01134_, _01413_);
  and (_02115_, _01126_, _01417_);
  or (_02116_, _02115_, _02114_);
  or (_02117_, _02116_, _02113_);
  or (_02118_, _02117_, _02112_);
  or (_02119_, _02118_, _02111_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02119_, _02106_);
  and (_02120_, _01109_, _01466_);
  and (_02121_, _01152_, _41950_);
  and (_02122_, _01113_, _01457_);
  or (_02123_, _02122_, _02121_);
  or (_02124_, _02123_, _02120_);
  and (_02125_, _01130_, _01485_);
  and (_02126_, _01140_, _01478_);
  and (_02127_, _01137_, _01483_);
  or (_02128_, _02127_, _02126_);
  and (_02129_, _01143_, _01445_);
  and (_02130_, _01134_, _01468_);
  or (_02131_, _02130_, _02129_);
  or (_02132_, _02131_, _02128_);
  or (_02133_, _02132_, _02125_);
  and (_02134_, _01123_, _01447_);
  and (_02135_, _01126_, _01455_);
  or (_02136_, _02135_, _02134_);
  or (_02137_, _02136_, _02133_);
  and (_02138_, _01170_, _01474_);
  and (_02139_, _01162_, _01449_);
  and (_02140_, _01155_, _01461_);
  and (_02141_, _01158_, _01472_);
  or (_02142_, _02141_, _02140_);
  or (_02143_, _02142_, _02139_);
  or (_02144_, _02143_, _02138_);
  and (_02145_, _01167_, _01476_);
  and (_02146_, _01117_, _01453_);
  or (_02147_, _02146_, _02145_);
  or (_02148_, _02147_, _02144_);
  or (_02149_, _02148_, _02137_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02149_, _02124_);
  and (_02150_, _01113_, _01500_);
  and (_02151_, _01152_, _41957_);
  and (_02152_, _01109_, _01511_);
  or (_02153_, _02152_, _02151_);
  or (_02154_, _02153_, _02150_);
  and (_02155_, _01123_, _01517_);
  and (_02156_, _01137_, _01528_);
  and (_02157_, _01143_, _01494_);
  or (_02158_, _02157_, _02156_);
  and (_02159_, _01134_, _01513_);
  and (_02160_, _01140_, _01523_);
  or (_02161_, _02160_, _02159_);
  or (_02162_, _02161_, _02158_);
  or (_02163_, _02162_, _02155_);
  and (_02164_, _01130_, _01530_);
  and (_02165_, _01126_, _01502_);
  or (_02166_, _02165_, _02164_);
  or (_02167_, _02166_, _02163_);
  and (_02168_, _01170_, _01521_);
  and (_02169_, _01162_, _01490_);
  and (_02170_, _01158_, _01492_);
  and (_02171_, _01155_, _01506_);
  or (_02172_, _02171_, _02170_);
  or (_02173_, _02172_, _02169_);
  or (_02174_, _02173_, _02168_);
  and (_02175_, _01117_, _01498_);
  and (_02176_, _01167_, _01519_);
  or (_02177_, _02176_, _02175_);
  or (_02178_, _02177_, _02174_);
  or (_02179_, _02178_, _02167_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02179_, _02154_);
  and (_02180_, _01113_, _01550_);
  and (_02181_, _01167_, _01564_);
  and (_02182_, _01109_, _01545_);
  or (_02183_, _02182_, _02181_);
  or (_02184_, _02183_, _02180_);
  and (_02185_, _01123_, _01562_);
  and (_02186_, _01140_, _01568_);
  and (_02187_, _01134_, _01548_);
  or (_02188_, _02187_, _02186_);
  and (_02189_, _01143_, _01539_);
  and (_02190_, _01137_, _01573_);
  or (_02191_, _02190_, _02189_);
  or (_02192_, _02191_, _02188_);
  or (_02193_, _02192_, _02185_);
  and (_02194_, _01130_, _01575_);
  and (_02195_, _01126_, _01552_);
  or (_02196_, _02195_, _02194_);
  or (_02197_, _02196_, _02193_);
  and (_02198_, _01152_, _41964_);
  and (_02199_, _01170_, _01566_);
  or (_02200_, _02199_, _02198_);
  and (_02201_, _01117_, _01543_);
  and (_02202_, _01158_, _01537_);
  and (_02203_, _01155_, _01556_);
  and (_02204_, _01162_, _01535_);
  or (_02205_, _02204_, _02203_);
  or (_02206_, _02205_, _02202_);
  or (_02207_, _02206_, _02201_);
  or (_02208_, _02207_, _02200_);
  or (_02209_, _02208_, _02197_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02209_, _02184_);
  nand (_02210_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02211_, \oc8051_golden_model_1.PC [3]);
  or (_02212_, \oc8051_golden_model_1.PC [2], _02211_);
  or (_02213_, _02212_, _02210_);
  or (_02214_, _02213_, _41737_);
  not (_02215_, \oc8051_golden_model_1.PC [1]);
  or (_02216_, _02215_, \oc8051_golden_model_1.PC [0]);
  or (_02217_, _02216_, _02212_);
  or (_02218_, _02217_, _41683_);
  and (_02219_, _02218_, _02214_);
  not (_02220_, \oc8051_golden_model_1.PC [2]);
  or (_02221_, _02220_, \oc8051_golden_model_1.PC [3]);
  or (_02222_, _02221_, _02210_);
  or (_02223_, _02222_, _41555_);
  or (_02224_, _02221_, _02216_);
  or (_02225_, _02224_, _41514_);
  and (_02226_, _02225_, _02223_);
  and (_02227_, _02226_, _02219_);
  and (_02228_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_02229_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_02230_, _02229_, _02228_);
  nand (_02231_, _02230_, _41964_);
  nand (_02232_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02233_, _02232_, _02216_);
  or (_02234_, _02233_, _41907_);
  and (_02235_, _02234_, _02231_);
  or (_02236_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02237_, _02236_, _02210_);
  or (_02238_, _02237_, _41389_);
  or (_02239_, _02236_, _02216_);
  or (_02240_, _02239_, _41348_);
  and (_02241_, _02240_, _02238_);
  and (_02242_, _02241_, _02235_);
  and (_02243_, _02242_, _02227_);
  not (_02244_, \oc8051_golden_model_1.PC [0]);
  or (_02245_, \oc8051_golden_model_1.PC [1], _02244_);
  or (_02246_, _02245_, _02232_);
  or (_02247_, _02246_, _41850_);
  or (_02248_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02249_, _02248_, _02232_);
  or (_02250_, _02249_, _41793_);
  and (_02251_, _02250_, _02247_);
  or (_02252_, _02236_, _02248_);
  or (_02253_, _02252_, _41238_);
  or (_02254_, _02236_, _02245_);
  or (_02255_, _02254_, _41279_);
  and (_02256_, _02255_, _02253_);
  and (_02257_, _02256_, _02251_);
  or (_02258_, _02245_, _02212_);
  or (_02259_, _02258_, _41637_);
  or (_02260_, _02248_, _02212_);
  or (_02261_, _02260_, _41596_);
  and (_02262_, _02261_, _02259_);
  or (_02263_, _02245_, _02221_);
  or (_02264_, _02263_, _41473_);
  or (_02265_, _02248_, _02221_);
  or (_02266_, _02265_, _41432_);
  and (_02267_, _02266_, _02264_);
  and (_02268_, _02267_, _02262_);
  and (_02269_, _02268_, _02257_);
  and (_02270_, _02269_, _02243_);
  or (_02271_, _02213_, _41690_);
  or (_02272_, _02217_, _41643_);
  and (_02273_, _02272_, _02271_);
  or (_02274_, _02222_, _41520_);
  or (_02275_, _02224_, _41479_);
  and (_02276_, _02275_, _02274_);
  and (_02277_, _02276_, _02273_);
  nand (_02278_, _02230_, _41915_);
  or (_02279_, _02233_, _41859_);
  and (_02280_, _02279_, _02278_);
  or (_02281_, _02237_, _41354_);
  or (_02282_, _02239_, _41289_);
  and (_02283_, _02282_, _02281_);
  and (_02284_, _02283_, _02280_);
  and (_02285_, _02284_, _02277_);
  or (_02286_, _02246_, _41801_);
  or (_02287_, _02249_, _41745_);
  and (_02288_, _02287_, _02286_);
  or (_02289_, _02252_, _41203_);
  or (_02290_, _02254_, _41244_);
  and (_02291_, _02290_, _02289_);
  and (_02292_, _02291_, _02288_);
  or (_02293_, _02258_, _41602_);
  or (_02294_, _02260_, _41561_);
  and (_02295_, _02294_, _02293_);
  or (_02296_, _02263_, _41438_);
  or (_02297_, _02265_, _41395_);
  and (_02298_, _02297_, _02296_);
  and (_02299_, _02298_, _02295_);
  and (_02300_, _02299_, _02292_);
  and (_02301_, _02300_, _02285_);
  and (_02302_, _02301_, _02270_);
  or (_02303_, _02213_, _41724_);
  or (_02304_, _02217_, _41670_);
  and (_02305_, _02304_, _02303_);
  or (_02306_, _02222_, _41545_);
  or (_02307_, _02224_, _41504_);
  and (_02308_, _02307_, _02306_);
  and (_02309_, _02308_, _02305_);
  nand (_02310_, _02230_, _41950_);
  or (_02311_, _02233_, _41894_);
  and (_02312_, _02311_, _02310_);
  or (_02313_, _02237_, _41379_);
  or (_02314_, _02239_, _41338_);
  and (_02315_, _02314_, _02313_);
  and (_02316_, _02315_, _02312_);
  and (_02317_, _02316_, _02309_);
  or (_02318_, _02246_, _41836_);
  or (_02319_, _02249_, _41780_);
  and (_02320_, _02319_, _02318_);
  or (_02321_, _02252_, _41228_);
  or (_02322_, _02254_, _41269_);
  and (_02323_, _02322_, _02321_);
  and (_02324_, _02323_, _02320_);
  or (_02325_, _02258_, _41627_);
  or (_02326_, _02260_, _41586_);
  and (_02327_, _02326_, _02325_);
  or (_02328_, _02263_, _41463_);
  or (_02329_, _02265_, _41422_);
  and (_02330_, _02329_, _02328_);
  and (_02331_, _02330_, _02327_);
  and (_02332_, _02331_, _02324_);
  and (_02333_, _02332_, _02317_);
  or (_02334_, _02213_, _41730_);
  or (_02335_, _02217_, _41677_);
  and (_02336_, _02335_, _02334_);
  or (_02337_, _02222_, _41550_);
  or (_02338_, _02224_, _41509_);
  and (_02339_, _02338_, _02337_);
  and (_02340_, _02339_, _02336_);
  nand (_02341_, _02230_, _41957_);
  or (_02342_, _02233_, _41901_);
  and (_02343_, _02342_, _02341_);
  or (_02344_, _02237_, _41384_);
  or (_02345_, _02239_, _41343_);
  and (_02346_, _02345_, _02344_);
  and (_02347_, _02346_, _02343_);
  and (_02348_, _02347_, _02340_);
  or (_02349_, _02246_, _41844_);
  or (_02350_, _02249_, _41787_);
  and (_02351_, _02350_, _02349_);
  or (_02352_, _02252_, _41233_);
  or (_02353_, _02254_, _41274_);
  and (_02354_, _02353_, _02352_);
  and (_02355_, _02354_, _02351_);
  or (_02356_, _02258_, _41632_);
  or (_02357_, _02260_, _41591_);
  and (_02358_, _02357_, _02356_);
  or (_02359_, _02263_, _41468_);
  or (_02360_, _02265_, _41427_);
  and (_02361_, _02360_, _02359_);
  and (_02362_, _02361_, _02358_);
  and (_02363_, _02362_, _02355_);
  nand (_02364_, _02363_, _02348_);
  or (_02365_, _02364_, _02333_);
  not (_02366_, _02365_);
  and (_02367_, _02366_, _02302_);
  or (_02368_, _02213_, _41710_);
  or (_02369_, _02217_, _41658_);
  and (_02370_, _02369_, _02368_);
  or (_02371_, _02222_, _41535_);
  or (_02372_, _02224_, _41494_);
  and (_02373_, _02372_, _02371_);
  and (_02374_, _02373_, _02370_);
  nand (_02375_, _02230_, _41936_);
  or (_02376_, _02233_, _41880_);
  and (_02377_, _02376_, _02375_);
  or (_02378_, _02237_, _41369_);
  or (_02379_, _02239_, _41322_);
  and (_02380_, _02379_, _02378_);
  and (_02381_, _02380_, _02377_);
  and (_02382_, _02381_, _02374_);
  or (_02383_, _02246_, _41822_);
  or (_02384_, _02249_, _41766_);
  and (_02385_, _02384_, _02383_);
  or (_02386_, _02252_, _41218_);
  or (_02387_, _02254_, _41259_);
  and (_02388_, _02387_, _02386_);
  and (_02389_, _02388_, _02385_);
  or (_02390_, _02258_, _41617_);
  or (_02391_, _02260_, _41576_);
  and (_02392_, _02391_, _02390_);
  or (_02393_, _02263_, _41453_);
  or (_02394_, _02265_, _41411_);
  and (_02395_, _02394_, _02393_);
  and (_02396_, _02395_, _02392_);
  and (_02397_, _02396_, _02389_);
  nand (_02398_, _02397_, _02382_);
  or (_02399_, _02213_, _41717_);
  or (_02400_, _02217_, _41664_);
  and (_02401_, _02400_, _02399_);
  or (_02402_, _02222_, _41540_);
  or (_02403_, _02224_, _41499_);
  and (_02404_, _02403_, _02402_);
  and (_02405_, _02404_, _02401_);
  nand (_02406_, _02230_, _41943_);
  or (_02407_, _02233_, _41887_);
  and (_02408_, _02407_, _02406_);
  or (_02409_, _02237_, _41374_);
  or (_02410_, _02239_, _41333_);
  and (_02411_, _02410_, _02409_);
  and (_02412_, _02411_, _02408_);
  and (_02413_, _02412_, _02405_);
  or (_02414_, _02246_, _41829_);
  or (_02415_, _02249_, _41773_);
  and (_02416_, _02415_, _02414_);
  or (_02417_, _02252_, _41223_);
  or (_02418_, _02254_, _41264_);
  and (_02419_, _02418_, _02417_);
  and (_02420_, _02419_, _02416_);
  or (_02421_, _02258_, _41622_);
  or (_02422_, _02260_, _41581_);
  and (_02423_, _02422_, _02421_);
  or (_02424_, _02263_, _41458_);
  or (_02425_, _02265_, _41416_);
  and (_02426_, _02425_, _02424_);
  and (_02427_, _02426_, _02423_);
  and (_02428_, _02427_, _02420_);
  nand (_02429_, _02428_, _02413_);
  or (_02430_, _02429_, _02398_);
  not (_02431_, _02430_);
  or (_02432_, _02213_, _41697_);
  or (_02433_, _02217_, _41648_);
  and (_02434_, _02433_, _02432_);
  or (_02435_, _02222_, _41525_);
  or (_02436_, _02224_, _41484_);
  and (_02437_, _02436_, _02435_);
  and (_02438_, _02437_, _02434_);
  nand (_02439_, _02230_, _41922_);
  or (_02440_, _02233_, _41866_);
  and (_02441_, _02440_, _02439_);
  or (_02442_, _02237_, _41359_);
  or (_02443_, _02239_, _41300_);
  and (_02444_, _02443_, _02442_);
  and (_02445_, _02444_, _02441_);
  and (_02446_, _02445_, _02438_);
  or (_02447_, _02246_, _41808_);
  or (_02448_, _02249_, _41752_);
  and (_02449_, _02448_, _02447_);
  or (_02450_, _02252_, _41208_);
  or (_02451_, _02254_, _41249_);
  and (_02452_, _02451_, _02450_);
  and (_02453_, _02452_, _02449_);
  or (_02454_, _02258_, _41607_);
  or (_02455_, _02260_, _41566_);
  and (_02456_, _02455_, _02454_);
  or (_02457_, _02263_, _41443_);
  or (_02458_, _02265_, _41400_);
  and (_02459_, _02458_, _02457_);
  and (_02460_, _02459_, _02456_);
  and (_02461_, _02460_, _02453_);
  and (_02462_, _02461_, _02446_);
  or (_02463_, _02213_, _41703_);
  or (_02464_, _02217_, _41653_);
  and (_02465_, _02464_, _02463_);
  or (_02466_, _02222_, _41530_);
  or (_02467_, _02224_, _41489_);
  and (_02468_, _02467_, _02466_);
  and (_02469_, _02468_, _02465_);
  nand (_02470_, _02230_, _41929_);
  or (_02471_, _02233_, _41873_);
  and (_02472_, _02471_, _02470_);
  or (_02473_, _02237_, _41364_);
  or (_02474_, _02239_, _41311_);
  and (_02475_, _02474_, _02473_);
  and (_02476_, _02475_, _02472_);
  and (_02477_, _02476_, _02469_);
  or (_02478_, _02246_, _41816_);
  or (_02479_, _02249_, _41759_);
  and (_02480_, _02479_, _02478_);
  or (_02481_, _02252_, _41213_);
  or (_02482_, _02254_, _41254_);
  and (_02483_, _02482_, _02481_);
  and (_02484_, _02483_, _02480_);
  or (_02485_, _02258_, _41612_);
  or (_02486_, _02260_, _41571_);
  and (_02487_, _02486_, _02485_);
  or (_02488_, _02263_, _41448_);
  or (_02489_, _02265_, _41405_);
  and (_02490_, _02489_, _02488_);
  and (_02491_, _02490_, _02487_);
  and (_02492_, _02491_, _02484_);
  nand (_02493_, _02492_, _02477_);
  not (_02494_, _02493_);
  and (_02495_, _02494_, _02462_);
  and (_02496_, _02495_, _02431_);
  and (_02497_, _02496_, _02367_);
  not (_02498_, _02497_);
  or (_02499_, _02493_, _02462_);
  or (_02500_, _02499_, _02430_);
  not (_02501_, _02500_);
  nand (_02502_, _02332_, _02317_);
  and (_02503_, _02363_, _02348_);
  or (_02504_, _02503_, _02502_);
  not (_02505_, _02504_);
  nand (_02506_, _02269_, _02243_);
  and (_02507_, _02301_, _02506_);
  and (_02508_, _02507_, _02505_);
  and (_02509_, _02508_, _02501_);
  not (_02510_, _02509_);
  or (_02511_, _02503_, _02333_);
  not (_02512_, _02511_);
  and (_02513_, _02512_, _02507_);
  and (_02514_, _02513_, _02501_);
  or (_02515_, _02364_, _02502_);
  or (_02516_, _02301_, _02506_);
  nor (_02517_, _02516_, _02515_);
  and (_02518_, _02517_, _02501_);
  nor (_02519_, _02518_, _02514_);
  and (_02520_, _02519_, _02510_);
  not (_02521_, _02515_);
  and (_02522_, _02302_, _02521_);
  and (_02523_, _02522_, _02501_);
  not (_02524_, _02523_);
  and (_02525_, _02367_, _02501_);
  not (_02526_, _02525_);
  not (_02527_, _02302_);
  or (_02528_, _02527_, _02511_);
  or (_02529_, _02528_, _02500_);
  not (_02530_, _02507_);
  or (_02531_, _02365_, _02530_);
  or (_02532_, _02531_, _02500_);
  and (_02533_, _02532_, _02529_);
  or (_02534_, _02515_, _02530_);
  or (_02535_, _02534_, _02500_);
  or (_02536_, _02527_, _02504_);
  or (_02537_, _02536_, _02500_);
  and (_02538_, _02537_, _02535_);
  and (_02539_, _02538_, _02533_);
  and (_02540_, _02539_, _02526_);
  and (_02541_, _02540_, _02524_);
  and (_02542_, _02541_, _02520_);
  not (_02543_, _02462_);
  and (_02544_, _02493_, _02543_);
  and (_02545_, _02544_, _02431_);
  and (_02546_, _02545_, _02517_);
  and (_02547_, _02228_, \oc8051_golden_model_1.PC [2]);
  and (_02548_, _02210_, _02220_);
  nor (_02549_, _02548_, _02547_);
  and (_02550_, _02549_, \oc8051_golden_model_1.ACC [2]);
  not (_02551_, \oc8051_golden_model_1.ACC [1]);
  and (_02552_, _02245_, _02216_);
  nor (_02553_, _02552_, _02551_);
  and (_02554_, \oc8051_golden_model_1.ACC [0], _02244_);
  and (_02555_, _02552_, _02551_);
  nor (_02556_, _02555_, _02553_);
  and (_02557_, _02556_, _02554_);
  nor (_02558_, _02557_, _02553_);
  nor (_02559_, _02549_, \oc8051_golden_model_1.ACC [2]);
  nor (_02560_, _02559_, _02550_);
  not (_02561_, _02560_);
  nor (_02562_, _02561_, _02558_);
  nor (_02563_, _02562_, _02550_);
  not (_02564_, \oc8051_golden_model_1.ACC [3]);
  not (_02565_, _02222_);
  nor (_02566_, _02547_, _02211_);
  nor (_02567_, _02566_, _02565_);
  nor (_02568_, _02567_, _02564_);
  and (_02569_, _02567_, _02564_);
  nor (_02570_, _02569_, _02568_);
  nor (_02571_, _02570_, _02563_);
  and (_02572_, _02570_, _02563_);
  or (_02573_, _02572_, _02571_);
  and (_02574_, _02573_, _02546_);
  not (_02575_, _02499_);
  not (_02576_, _02429_);
  and (_02577_, _02576_, _02398_);
  and (_02578_, _02577_, _02575_);
  and (_02579_, _02578_, _02517_);
  nor (_02580_, _02365_, _02516_);
  and (_02581_, _02580_, _02501_);
  nor (_02582_, _02581_, _02579_);
  and (_02583_, _02580_, _02545_);
  and (_02584_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  and (_02585_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_02586_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02587_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02588_, _02587_, _02585_);
  and (_02589_, _02588_, _02586_);
  nor (_02590_, _02589_, _02585_);
  nor (_02591_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02592_, _02591_, _02584_);
  not (_02593_, _02592_);
  nor (_02594_, _02593_, _02590_);
  nor (_02595_, _02594_, _02584_);
  and (_02596_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02597_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02598_, _02597_, _02596_);
  not (_02599_, _02598_);
  nor (_02600_, _02599_, _02595_);
  and (_02601_, _02599_, _02595_);
  nor (_02602_, _02601_, _02600_);
  nand (_02603_, _02602_, _02583_);
  and (_02604_, _02603_, _02582_);
  not (_02605_, _02583_);
  not (_02606_, _02567_);
  or (_02607_, _02301_, _02270_);
  or (_02608_, _02607_, _02365_);
  or (_02609_, _02608_, _02500_);
  or (_02610_, _02607_, _02511_);
  or (_02611_, _02610_, _02500_);
  and (_02612_, _02611_, _02609_);
  or (_02613_, _02516_, _02511_);
  or (_02614_, _02613_, _02500_);
  or (_02615_, _02607_, _02504_);
  or (_02616_, _02615_, _02500_);
  and (_02617_, _02616_, _02614_);
  or (_02618_, _02516_, _02504_);
  or (_02619_, _02618_, _02500_);
  or (_02620_, _02607_, _02515_);
  or (_02621_, _02620_, _02500_);
  and (_02622_, _02621_, _02619_);
  and (_02623_, _02622_, _02617_);
  nand (_02624_, _02623_, _02612_);
  or (_02625_, _02624_, _02606_);
  and (_02626_, _02229_, \oc8051_golden_model_1.PC [1]);
  and (_02627_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02628_, _02627_, \oc8051_golden_model_1.PC [3]);
  nor (_02629_, _02628_, _02626_);
  and (_02630_, _02623_, _02612_);
  or (_02631_, _02630_, _02629_);
  and (_02632_, _02631_, _02625_);
  nand (_02633_, _02632_, _02605_);
  nand (_02634_, _02633_, _02604_);
  not (_02635_, _02546_);
  or (_02636_, _02582_, _02629_);
  and (_02637_, _02636_, _02635_);
  and (_02638_, _02637_, _02634_);
  or (_02639_, _02638_, _02574_);
  and (_02640_, _02639_, _02542_);
  not (_02641_, _02629_);
  nor (_02642_, _02641_, _02542_);
  nor (_02643_, _02642_, _02640_);
  and (_02644_, _02561_, _02558_);
  nor (_02645_, _02644_, _02562_);
  and (_02646_, _02645_, _02546_);
  nor (_02647_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02648_, _02647_, _02627_);
  or (_02649_, _02648_, _02630_);
  or (_02650_, _02648_, _02582_);
  and (_02651_, _02650_, _02635_);
  and (_02652_, _02593_, _02590_);
  nor (_02653_, _02652_, _02594_);
  nand (_02654_, _02653_, _02583_);
  and (_02655_, _02654_, _02582_);
  or (_02656_, _02624_, _02549_);
  nand (_02657_, _02656_, _02605_);
  nand (_02658_, _02657_, _02655_);
  nand (_02659_, _02658_, _02651_);
  nand (_02660_, _02659_, _02542_);
  and (_02661_, _02660_, _02649_);
  or (_02662_, _02661_, _02646_);
  or (_02663_, _02648_, _02542_);
  nand (_02664_, _02663_, _02662_);
  or (_02665_, _02664_, _02643_);
  or (_02666_, _02542_, \oc8051_golden_model_1.PC [0]);
  not (_02667_, \oc8051_golden_model_1.ACC [0]);
  and (_02668_, _02667_, \oc8051_golden_model_1.PC [0]);
  nor (_02669_, _02668_, _02554_);
  and (_02670_, _02669_, _02546_);
  and (_02671_, _02630_, _02582_);
  or (_02672_, _02671_, \oc8051_golden_model_1.PC [0]);
  not (_02673_, _02542_);
  or (_02674_, _02624_, _02244_);
  and (_02675_, _02674_, _02605_);
  nor (_02676_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02677_, _02676_, _02586_);
  nand (_02678_, _02677_, _02583_);
  nand (_02679_, _02678_, _02582_);
  or (_02680_, _02679_, _02675_);
  and (_02681_, _02680_, _02635_);
  or (_02682_, _02681_, _02673_);
  and (_02683_, _02682_, _02672_);
  or (_02684_, _02683_, _02670_);
  nand (_02685_, _02684_, _02666_);
  or (_02686_, _02630_, \oc8051_golden_model_1.PC [1]);
  or (_02687_, _02624_, _02552_);
  nand (_02689_, _02687_, _02686_);
  nand (_02690_, _02689_, _02605_);
  nor (_02691_, _02588_, _02586_);
  nor (_02692_, _02691_, _02589_);
  nand (_02693_, _02692_, _02583_);
  and (_02694_, _02693_, _02582_);
  nand (_02695_, _02694_, _02690_);
  or (_02696_, _02582_, _02215_);
  and (_02697_, _02696_, _02635_);
  and (_02698_, _02697_, _02695_);
  nor (_02699_, _02556_, _02554_);
  nor (_02700_, _02699_, _02557_);
  and (_02701_, _02700_, _02546_);
  or (_02702_, _02701_, _02698_);
  and (_02703_, _02702_, _02542_);
  nor (_02704_, _02542_, \oc8051_golden_model_1.PC [1]);
  nor (_02705_, _02704_, _02703_);
  or (_02706_, _02705_, _02685_);
  nor (_02707_, _02706_, _02665_);
  nand (_02708_, _02707_, _41915_);
  or (_02709_, _02704_, _02703_);
  or (_02710_, _02709_, _02685_);
  or (_02711_, _02642_, _02640_);
  and (_02712_, _02663_, _02662_);
  or (_02713_, _02712_, _02711_);
  or (_02714_, _02713_, _02710_);
  or (_02715_, _02714_, _41244_);
  and (_02716_, _02715_, _02708_);
  or (_02717_, _02712_, _02643_);
  or (_02718_, _02717_, _02706_);
  or (_02719_, _02718_, _41690_);
  and (_02720_, _02684_, _02666_);
  or (_02721_, _02709_, _02720_);
  or (_02722_, _02713_, _02721_);
  or (_02723_, _02722_, _41203_);
  and (_02724_, _02723_, _02719_);
  and (_02725_, _02724_, _02716_);
  or (_02726_, _02717_, _02710_);
  or (_02727_, _02726_, _41602_);
  or (_02728_, _02705_, _02720_);
  or (_02729_, _02713_, _02728_);
  or (_02730_, _02729_, _41289_);
  and (_02731_, _02730_, _02727_);
  or (_02732_, _02664_, _02711_);
  or (_02733_, _02732_, _02706_);
  or (_02734_, _02733_, _41520_);
  or (_02735_, _02732_, _02710_);
  or (_02736_, _02735_, _41438_);
  and (_02737_, _02736_, _02734_);
  and (_02738_, _02737_, _02731_);
  and (_02739_, _02738_, _02725_);
  or (_02740_, _02713_, _02706_);
  or (_02741_, _02740_, _41354_);
  or (_02742_, _02732_, _02721_);
  or (_02743_, _02742_, _41395_);
  and (_02744_, _02743_, _02741_);
  or (_02745_, _02728_, _02665_);
  or (_02746_, _02745_, _41859_);
  or (_02747_, _02717_, _02728_);
  or (_02748_, _02747_, _41643_);
  and (_02749_, _02748_, _02746_);
  and (_02750_, _02749_, _02744_);
  or (_02751_, _02721_, _02665_);
  or (_02752_, _02751_, _41745_);
  or (_02753_, _02717_, _02721_);
  or (_02754_, _02753_, _41561_);
  and (_02755_, _02754_, _02752_);
  or (_02756_, _02710_, _02665_);
  or (_02757_, _02756_, _41801_);
  or (_02758_, _02732_, _02728_);
  or (_02759_, _02758_, _41479_);
  and (_02760_, _02759_, _02757_);
  and (_02761_, _02760_, _02755_);
  and (_02762_, _02761_, _02750_);
  nand (_02763_, _02762_, _02739_);
  or (_02764_, _02751_, _41773_);
  or (_02765_, _02718_, _41717_);
  and (_02766_, _02765_, _02764_);
  nand (_02767_, _02707_, _41943_);
  or (_02768_, _02745_, _41887_);
  and (_02769_, _02768_, _02767_);
  and (_02770_, _02769_, _02766_);
  or (_02771_, _02742_, _41416_);
  or (_02772_, _02729_, _41333_);
  and (_02773_, _02772_, _02771_);
  or (_02774_, _02733_, _41540_);
  or (_02775_, _02735_, _41458_);
  and (_02776_, _02775_, _02774_);
  and (_02777_, _02776_, _02773_);
  and (_02778_, _02777_, _02770_);
  or (_02779_, _02726_, _41622_);
  or (_02780_, _02714_, _41264_);
  and (_02781_, _02780_, _02779_);
  or (_02782_, _02753_, _41581_);
  or (_02783_, _02740_, _41374_);
  and (_02784_, _02783_, _02782_);
  and (_02785_, _02784_, _02781_);
  or (_02786_, _02756_, _41829_);
  or (_02787_, _02722_, _41223_);
  and (_02788_, _02787_, _02786_);
  or (_02789_, _02747_, _41664_);
  or (_02790_, _02758_, _41499_);
  and (_02791_, _02790_, _02789_);
  and (_02792_, _02791_, _02788_);
  and (_02793_, _02792_, _02785_);
  and (_02794_, _02793_, _02778_);
  or (_02795_, _02794_, _02763_);
  nor (_02796_, _02795_, _02498_);
  nor (_02797_, _02498_, _02763_);
  not (_02798_, _02797_);
  and (_02799_, _02462_, _02429_);
  and (_02800_, _02799_, _02367_);
  nor (_02801_, _02529_, \oc8051_golden_model_1.SP [0]);
  and (_02802_, _02578_, _02513_);
  not (_02803_, _02802_);
  nor (_02804_, _02803_, _02763_);
  or (_02805_, _02718_, _41697_);
  or (_02806_, _02747_, _41648_);
  and (_02807_, _02806_, _02805_);
  or (_02808_, _02733_, _41525_);
  or (_02809_, _02758_, _41484_);
  and (_02810_, _02809_, _02808_);
  and (_02811_, _02810_, _02807_);
  nand (_02812_, _02707_, _41922_);
  or (_02813_, _02745_, _41866_);
  and (_02814_, _02813_, _02812_);
  or (_02815_, _02740_, _41359_);
  or (_02816_, _02729_, _41300_);
  and (_02817_, _02816_, _02815_);
  and (_02818_, _02817_, _02814_);
  and (_02819_, _02818_, _02811_);
  or (_02820_, _02756_, _41808_);
  or (_02821_, _02751_, _41752_);
  and (_02822_, _02821_, _02820_);
  or (_02823_, _02722_, _41208_);
  or (_02824_, _02714_, _41249_);
  and (_02825_, _02824_, _02823_);
  and (_02826_, _02825_, _02822_);
  or (_02827_, _02726_, _41607_);
  or (_02828_, _02753_, _41566_);
  and (_02829_, _02828_, _02827_);
  or (_02830_, _02735_, _41443_);
  or (_02831_, _02742_, _41400_);
  and (_02832_, _02831_, _02830_);
  and (_02833_, _02832_, _02829_);
  and (_02834_, _02833_, _02826_);
  nand (_02835_, _02834_, _02819_);
  and (_02836_, _02835_, _02804_);
  and (_02837_, _02834_, _02819_);
  not (_02838_, _02579_);
  and (_02839_, _02429_, _02398_);
  and (_02840_, _02839_, _02495_);
  and (_02841_, _02840_, _02517_);
  not (_02842_, _02841_);
  not (_02843_, _02398_);
  and (_02844_, _02429_, _02843_);
  and (_02845_, _02844_, _02493_);
  and (_02846_, _02839_, _02575_);
  and (_02847_, _02839_, _02493_);
  or (_02848_, _02847_, _02846_);
  or (_02849_, _02848_, _02845_);
  nand (_02850_, _02849_, _02517_);
  and (_02851_, _02850_, _02842_);
  and (_02852_, _02577_, _02493_);
  and (_02853_, _02852_, _02517_);
  and (_02854_, _02844_, _02494_);
  and (_02855_, _02854_, _02517_);
  nor (_02856_, _02855_, _02853_);
  and (_02857_, _02856_, _02851_);
  and (_02858_, _02857_, _02838_);
  nor (_02859_, _02858_, _02763_);
  and (_02860_, _02859_, _02837_);
  and (_02861_, _02493_, _02462_);
  and (_02862_, _02861_, _02431_);
  and (_02863_, _02862_, _02580_);
  not (_02864_, _02863_);
  nor (_02865_, _02795_, _02864_);
  not (_02866_, \oc8051_golden_model_1.SP [0]);
  nor (_02867_, _02614_, _02866_);
  not (_02868_, _02613_);
  and (_02869_, _02862_, _02868_);
  not (_02870_, _02869_);
  nor (_02871_, _02795_, _02870_);
  nor (_02872_, _02870_, _02763_);
  not (_02873_, _02872_);
  not (_02874_, _02620_);
  and (_02875_, _02496_, _02874_);
  and (_02876_, _02862_, _02874_);
  not (_02877_, _02876_);
  nor (_02878_, _02795_, _02877_);
  not (_02879_, _02608_);
  and (_02880_, _02862_, _02879_);
  not (_02881_, _02880_);
  or (_02882_, _02795_, _02881_);
  nor (_02883_, _02881_, _02763_);
  not (_02884_, _02610_);
  and (_02885_, _02852_, _02884_);
  and (_02886_, _02852_, _02879_);
  nor (_02887_, _02886_, _02885_);
  and (_02888_, _02578_, _02522_);
  not (_02890_, _02888_);
  not (_02891_, _02536_);
  and (_02892_, _02862_, _02891_);
  not (_02893_, _02892_);
  and (_02894_, _02578_, _02891_);
  and (_02895_, _02794_, _02894_);
  not (_02896_, _02894_);
  and (_02897_, _02707_, _41964_);
  nor (_02898_, _02718_, _41737_);
  nor (_02899_, _02898_, _02897_);
  nor (_02900_, _02733_, _41555_);
  nor (_02901_, _02722_, _41238_);
  nor (_02902_, _02901_, _02900_);
  and (_02903_, _02902_, _02899_);
  nor (_02904_, _02745_, _41907_);
  nor (_02905_, _02756_, _41850_);
  nor (_02906_, _02905_, _02904_);
  nor (_02907_, _02747_, _41683_);
  nor (_02908_, _02726_, _41637_);
  nor (_02909_, _02908_, _02907_);
  and (_02910_, _02909_, _02906_);
  and (_02911_, _02910_, _02903_);
  nor (_02912_, _02742_, _41432_);
  nor (_02913_, _02740_, _41389_);
  nor (_02914_, _02913_, _02912_);
  nor (_02915_, _02758_, _41514_);
  nor (_02916_, _02735_, _41473_);
  nor (_02917_, _02916_, _02915_);
  and (_02918_, _02917_, _02914_);
  nor (_02919_, _02729_, _41348_);
  nor (_02920_, _02714_, _41279_);
  nor (_02921_, _02920_, _02919_);
  nor (_02922_, _02751_, _41793_);
  nor (_02923_, _02753_, _41596_);
  nor (_02924_, _02923_, _02922_);
  and (_02925_, _02924_, _02921_);
  and (_02926_, _02925_, _02918_);
  and (_02927_, _02926_, _02911_);
  nor (_02928_, _02927_, _02763_);
  not (_02929_, _02794_);
  and (_02930_, _02929_, _02763_);
  nor (_02931_, _02930_, _02928_);
  and (_02932_, _02862_, _02513_);
  and (_02933_, _02862_, _02517_);
  nor (_02934_, _02933_, _02932_);
  not (_02935_, _02934_);
  and (_02936_, _02935_, _02931_);
  and (_02937_, _02862_, _02522_);
  nor (_02938_, _02937_, _02497_);
  and (_02939_, _02862_, _02367_);
  and (_02940_, _02496_, _02891_);
  nor (_02941_, _02940_, _02939_);
  and (_02942_, _02941_, _02938_);
  or (_02943_, _02613_, _02543_);
  and (_02944_, _02839_, _02494_);
  nor (_02945_, _02944_, _02845_);
  nor (_02946_, _02945_, _02943_);
  and (_02947_, _02844_, _02544_);
  and (_02948_, _02947_, _02868_);
  nor (_02949_, _02948_, _02946_);
  and (_02950_, _02868_, _02578_);
  and (_02951_, _02495_, _02577_);
  and (_02952_, _02951_, _02868_);
  nor (_02953_, _02952_, _02950_);
  and (_02954_, _02854_, _02868_);
  not (_02955_, _02954_);
  and (_02956_, _02955_, _02953_);
  and (_02957_, _02956_, _02949_);
  and (_02958_, _02957_, _02942_);
  and (_02959_, _02846_, _02868_);
  and (_02960_, _02839_, _02861_);
  and (_02961_, _02960_, _02868_);
  or (_02962_, _02961_, _02959_);
  not (_02963_, _02962_);
  not (_02964_, _02534_);
  and (_02965_, _02545_, _02964_);
  nor (_02966_, _02965_, _02802_);
  not (_02967_, _02528_);
  and (_02968_, _02496_, _02967_);
  not (_02969_, _02531_);
  and (_02970_, _02545_, _02969_);
  nor (_02971_, _02970_, _02968_);
  and (_02972_, _02971_, _02966_);
  and (_02973_, _02972_, _02963_);
  and (_02974_, _02879_, _02578_);
  and (_02975_, _02839_, _02544_);
  and (_02976_, _02975_, _02868_);
  nor (_02977_, _02976_, _02974_);
  and (_02978_, _02852_, _02868_);
  not (_02979_, _02978_);
  and (_02980_, _02545_, _02508_);
  and (_02981_, _02496_, _02580_);
  nor (_02982_, _02981_, _02980_);
  and (_02983_, _02982_, _02979_);
  and (_02984_, _02983_, _02977_);
  and (_02985_, _02984_, _02973_);
  and (_02986_, _02985_, _02958_);
  nand (_02987_, _02986_, _02244_);
  and (_02988_, _02987_, _02215_);
  nor (_02989_, _02987_, _02215_);
  nor (_02990_, _02989_, _02988_);
  or (_02991_, _02986_, _02244_);
  nand (_02992_, _02991_, _02987_);
  nor (_02993_, _02992_, _02990_);
  nor (_02994_, _02986_, _02648_);
  not (_02995_, _02549_);
  and (_02996_, _02986_, _02995_);
  nor (_02997_, _02996_, _02994_);
  nor (_02998_, _02986_, _02641_);
  and (_02999_, _02986_, _02606_);
  nor (_03000_, _02999_, _02998_);
  and (_03001_, _03000_, _02997_);
  and (_03002_, _03001_, _02993_);
  and (_03003_, _03002_, _01408_);
  and (_03004_, _02992_, _02990_);
  and (_03005_, _03004_, _03001_);
  and (_03006_, _03005_, _01410_);
  nor (_03007_, _03006_, _03003_);
  not (_03008_, _03000_);
  and (_03009_, _03008_, _02997_);
  not (_03010_, _02990_);
  and (_03011_, _02992_, _03010_);
  and (_03012_, _03011_, _03009_);
  and (_03013_, _03012_, _41943_);
  nor (_03014_, _03000_, _02997_);
  and (_03015_, _03014_, _03011_);
  and (_03016_, _03015_, _01421_);
  nor (_03017_, _03016_, _03013_);
  and (_03018_, _03017_, _03007_);
  and (_03019_, _03009_, _02993_);
  and (_03020_, _03019_, _01433_);
  and (_03021_, _03009_, _03004_);
  and (_03022_, _03021_, _01431_);
  nor (_03023_, _03022_, _03020_);
  and (_03024_, _03014_, _02993_);
  and (_03025_, _03024_, _01402_);
  and (_03026_, _03014_, _03004_);
  and (_03027_, _03026_, _01404_);
  nor (_03028_, _03027_, _03025_);
  and (_03029_, _03028_, _03023_);
  and (_03030_, _03029_, _03018_);
  nor (_03031_, _02992_, _03010_);
  nor (_03032_, _03008_, _02997_);
  and (_03033_, _03032_, _03031_);
  and (_03034_, _03033_, _01438_);
  and (_03035_, _03032_, _02993_);
  and (_03036_, _03035_, _01427_);
  nor (_03037_, _03036_, _03034_);
  and (_03038_, _03011_, _03001_);
  and (_03039_, _03038_, _01415_);
  and (_03040_, _03031_, _03001_);
  and (_03041_, _03040_, _01413_);
  nor (_03042_, _03041_, _03039_);
  and (_03043_, _03042_, _03037_);
  and (_03044_, _03031_, _03009_);
  and (_03045_, _03044_, _01429_);
  and (_03046_, _03031_, _03014_);
  and (_03047_, _03046_, _01400_);
  nor (_03048_, _03047_, _03045_);
  and (_03049_, _03032_, _03011_);
  and (_03051_, _03049_, _01417_);
  and (_03052_, _03032_, _03004_);
  and (_03053_, _03052_, _01440_);
  nor (_03054_, _03053_, _03051_);
  and (_03055_, _03054_, _03048_);
  and (_03056_, _03055_, _03043_);
  and (_03057_, _03056_, _03030_);
  nor (_03058_, _03057_, _02838_);
  nor (_03059_, _02618_, _02576_);
  and (_03060_, _03059_, _02794_);
  and (_03062_, _02496_, _02868_);
  or (_03063_, _03062_, _02869_);
  not (_03064_, _03063_);
  nor (_03065_, _03064_, _02931_);
  nor (_03066_, _02877_, _02931_);
  and (_03067_, _02931_, _02880_);
  not (_03068_, \oc8051_golden_model_1.SP [3]);
  and (_03069_, _02496_, _02879_);
  and (_03070_, _03069_, _03068_);
  not (_03071_, _02615_);
  and (_03072_, _03071_, _02578_);
  nor (_03073_, _03072_, _02974_);
  or (_03074_, _03073_, _02794_);
  and (_03075_, _02874_, _02578_);
  nor (_03076_, _03069_, _02880_);
  nand (_03077_, _03073_, \oc8051_golden_model_1.PSW [3]);
  and (_03078_, _03077_, _03076_);
  or (_03079_, _03078_, _03075_);
  and (_03080_, _03079_, _03074_);
  or (_03081_, _03080_, _03070_);
  nor (_03083_, _03081_, _03067_);
  not (_03084_, _03075_);
  nor (_03085_, _03084_, _02794_);
  nor (_03086_, _03085_, _03083_);
  nor (_03087_, _03086_, _02876_);
  nor (_03088_, _02950_, _02875_);
  not (_03089_, _03088_);
  or (_03090_, _03089_, _03087_);
  nor (_03091_, _03090_, _03066_);
  and (_03092_, _03089_, _02794_);
  or (_03094_, _03063_, _03092_);
  nor (_03095_, _03094_, _03091_);
  or (_03096_, _03095_, _03059_);
  nor (_03097_, _03096_, _03065_);
  nor (_03098_, _03097_, _03060_);
  not (_03099_, _02618_);
  and (_03100_, _02496_, _03099_);
  and (_03101_, _02862_, _03099_);
  nor (_03102_, _03101_, _03100_);
  not (_03103_, _03102_);
  nor (_03105_, _03103_, _03098_);
  and (_03106_, _02580_, _02578_);
  and (_03107_, _03103_, _02931_);
  nor (_03108_, _03107_, _03106_);
  not (_03109_, _03108_);
  nor (_03110_, _03109_, _03105_);
  not (_03111_, _03106_);
  nor (_03112_, _03111_, _02794_);
  or (_03113_, _03112_, _03110_);
  and (_03114_, _03113_, _02864_);
  nor (_03115_, _02864_, _02931_);
  or (_03116_, _03115_, _03114_);
  and (_03117_, _03116_, _02838_);
  or (_03118_, _03117_, _02935_);
  nor (_03119_, _03118_, _03058_);
  nor (_03120_, _03119_, _02936_);
  and (_03121_, _02578_, _02964_);
  not (_03122_, _03121_);
  and (_03123_, _02862_, _02964_);
  nor (_03124_, _03123_, _02965_);
  and (_03126_, _03124_, _03122_);
  and (_03127_, _02862_, _02508_);
  not (_03128_, _03127_);
  and (_03129_, _02578_, _02508_);
  nor (_03130_, _03129_, _02980_);
  and (_03131_, _03130_, _03128_);
  and (_03132_, _03131_, _03126_);
  and (_03133_, _02578_, _02967_);
  not (_03134_, _03133_);
  and (_03135_, _02862_, _02969_);
  not (_03137_, _03135_);
  and (_03138_, _02578_, _02969_);
  nor (_03139_, _03138_, _02970_);
  and (_03140_, _03139_, _03137_);
  and (_03141_, _03140_, _03134_);
  and (_03142_, _03141_, _03132_);
  not (_03143_, _03142_);
  nor (_03144_, _03143_, _03120_);
  and (_03145_, _02862_, _02967_);
  and (_03146_, _03143_, _02794_);
  nor (_03148_, _03146_, _03145_);
  not (_03149_, _03148_);
  nor (_03150_, _03149_, _03144_);
  and (_03151_, _03145_, \oc8051_golden_model_1.SP [3]);
  or (_03152_, _03151_, _02968_);
  nor (_03153_, _03152_, _03150_);
  and (_03154_, _02931_, _02968_);
  or (_03155_, _03154_, _03153_);
  and (_03156_, _03155_, _02896_);
  or (_03157_, _03156_, _02895_);
  nand (_03159_, _03157_, _02893_);
  and (_03160_, _02892_, _03068_);
  nor (_03161_, _03160_, _02940_);
  nand (_03162_, _03161_, _03159_);
  and (_03163_, _02578_, _02367_);
  not (_03164_, _02940_);
  nor (_03165_, _03164_, _02931_);
  nor (_03166_, _03165_, _03163_);
  nand (_03167_, _03166_, _03162_);
  and (_03168_, _03163_, _02794_);
  nor (_03170_, _03168_, _02497_);
  and (_03171_, _03170_, _03167_);
  nor (_03172_, _02931_, _02498_);
  or (_03173_, _03172_, _03171_);
  nand (_03174_, _03173_, _02890_);
  nor (_03175_, _02794_, _02890_);
  not (_03176_, _03175_);
  and (_03177_, _03176_, _03174_);
  nor (_03178_, _02733_, _41550_);
  nor (_03179_, _02714_, _41274_);
  nor (_03181_, _03179_, _03178_);
  nor (_03182_, _02726_, _41632_);
  nor (_03183_, _02729_, _41343_);
  nor (_03184_, _03183_, _03182_);
  and (_03185_, _03184_, _03181_);
  nor (_03186_, _02756_, _41844_);
  nor (_03187_, _02751_, _41787_);
  nor (_03188_, _03187_, _03186_);
  nor (_03189_, _02735_, _41468_);
  nor (_03190_, _02742_, _41427_);
  nor (_03192_, _03190_, _03189_);
  and (_03193_, _03192_, _03188_);
  and (_03194_, _03193_, _03185_);
  nor (_03195_, _02745_, _41901_);
  nor (_03196_, _02718_, _41730_);
  nor (_03197_, _03196_, _03195_);
  nor (_03198_, _02740_, _41384_);
  nor (_03199_, _02722_, _41233_);
  nor (_03200_, _03199_, _03198_);
  and (_03201_, _03200_, _03197_);
  and (_03203_, _02707_, _41957_);
  nor (_03204_, _02758_, _41509_);
  nor (_03205_, _03204_, _03203_);
  nor (_03206_, _02747_, _41677_);
  nor (_03207_, _02753_, _41591_);
  nor (_03208_, _03207_, _03206_);
  and (_03209_, _03208_, _03205_);
  and (_03210_, _03209_, _03201_);
  and (_03211_, _03210_, _03194_);
  nor (_03212_, _03211_, _02763_);
  and (_03214_, _03212_, _02880_);
  not (_03215_, _03214_);
  nor (_03216_, _02940_, _02968_);
  and (_03217_, _03216_, _02864_);
  and (_03218_, _03102_, _03064_);
  nor (_03219_, _02876_, _02497_);
  and (_03220_, _03219_, _02934_);
  and (_03221_, _03220_, _03218_);
  and (_03222_, _03221_, _03217_);
  not (_03223_, _03222_);
  and (_03224_, _03223_, _03212_);
  not (_03225_, _03224_);
  nor (_03226_, _02733_, _41535_);
  nor (_03227_, _02714_, _41259_);
  nor (_03228_, _03227_, _03226_);
  nor (_03229_, _02726_, _41617_);
  nor (_03230_, _02740_, _41369_);
  nor (_03231_, _03230_, _03229_);
  and (_03232_, _03231_, _03228_);
  nor (_03233_, _02718_, _41710_);
  nor (_03234_, _02722_, _41218_);
  nor (_03235_, _03234_, _03233_);
  and (_03236_, _02707_, _41936_);
  nor (_03237_, _02756_, _41822_);
  nor (_03238_, _03237_, _03236_);
  and (_03239_, _03238_, _03235_);
  and (_03240_, _03239_, _03232_);
  nor (_03241_, _02745_, _41880_);
  nor (_03242_, _02729_, _41322_);
  nor (_03243_, _03242_, _03241_);
  nor (_03244_, _02753_, _41576_);
  nor (_03245_, _02758_, _41494_);
  nor (_03246_, _03245_, _03244_);
  and (_03247_, _03246_, _03243_);
  nor (_03248_, _02747_, _41658_);
  nor (_03249_, _02742_, _41411_);
  nor (_03250_, _03249_, _03248_);
  nor (_03251_, _02751_, _41766_);
  nor (_03252_, _02735_, _41453_);
  nor (_03253_, _03252_, _03251_);
  and (_03254_, _03253_, _03250_);
  and (_03255_, _03254_, _03247_);
  and (_03256_, _03255_, _03240_);
  nor (_03257_, _03106_, _03059_);
  nor (_03258_, _03163_, _03075_);
  and (_03259_, _03258_, _03257_);
  nor (_03260_, _02894_, _02888_);
  and (_03261_, _03260_, _03088_);
  and (_03262_, _03261_, _03073_);
  and (_03263_, _03262_, _03259_);
  and (_03264_, _03263_, _03142_);
  nor (_03265_, _03264_, _03256_);
  not (_03266_, _03265_);
  and (_03267_, _03012_, _41936_);
  and (_03268_, _03015_, _01376_);
  nor (_03269_, _03268_, _03267_);
  and (_03270_, _03005_, _01365_);
  and (_03271_, _03035_, _01390_);
  nor (_03272_, _03271_, _03270_);
  and (_03273_, _03272_, _03269_);
  and (_03274_, _03019_, _01386_);
  and (_03275_, _03021_, _01384_);
  nor (_03276_, _03275_, _03274_);
  and (_03277_, _03024_, _01357_);
  and (_03278_, _03026_, _01355_);
  nor (_03279_, _03278_, _03277_);
  and (_03280_, _03279_, _03276_);
  and (_03281_, _03280_, _03273_);
  and (_03282_, _03040_, _01368_);
  and (_03283_, _03049_, _01372_);
  nor (_03284_, _03283_, _03282_);
  and (_03285_, _03038_, _01370_);
  and (_03286_, _03033_, _01393_);
  nor (_03287_, _03286_, _03285_);
  and (_03288_, _03287_, _03284_);
  and (_03289_, _03044_, _01382_);
  and (_03290_, _03046_, _01359_);
  nor (_03291_, _03290_, _03289_);
  and (_03292_, _03002_, _01363_);
  and (_03293_, _03052_, _01395_);
  nor (_03294_, _03293_, _03292_);
  and (_03295_, _03294_, _03291_);
  and (_03296_, _03295_, _03288_);
  and (_03297_, _03296_, _03281_);
  nor (_03298_, _03297_, _02838_);
  not (_03299_, _02847_);
  nor (_03300_, _03299_, _02531_);
  not (_03301_, _03300_);
  and (_03302_, _02839_, _02522_);
  and (_03303_, _02944_, _02367_);
  nor (_03305_, _03303_, _03302_);
  and (_03306_, _03305_, _03301_);
  not (_03307_, _02944_);
  nor (_03308_, _03307_, _02534_);
  not (_03309_, _02839_);
  nor (_03310_, _03309_, _02615_);
  nor (_03311_, _03310_, _03308_);
  nor (_03312_, _03299_, _02528_);
  nor (_03313_, _03307_, _02531_);
  nor (_03314_, _03313_, _03312_);
  and (_03315_, _03314_, _03311_);
  and (_03316_, _03315_, _03306_);
  and (_03317_, _02847_, _02367_);
  and (_03318_, _02847_, _02874_);
  nor (_03319_, _03318_, _03317_);
  nor (_03320_, _02516_, _02333_);
  or (_03321_, _03320_, _02879_);
  and (_03322_, _03321_, _02847_);
  nor (_03323_, _03299_, _02534_);
  nor (_03324_, _03323_, _03322_);
  and (_03325_, _03324_, _03319_);
  and (_03326_, _03325_, _03316_);
  and (_03327_, _02608_, _02528_);
  nor (_03328_, _02868_, _02508_);
  nor (_03329_, _02516_, _02364_);
  nor (_03330_, _03329_, _02874_);
  and (_03331_, _03330_, _03328_);
  and (_03332_, _03331_, _03327_);
  nor (_03333_, _03332_, _03307_);
  not (_03334_, _03333_);
  not (_03335_, \oc8051_golden_model_1.SP [2]);
  not (_03336_, _03069_);
  nor (_03337_, _03145_, _02892_);
  and (_03338_, _03337_, _03336_);
  nor (_03339_, _03338_, _03335_);
  nor (_03340_, _03309_, _02536_);
  nor (_03341_, _02517_, _02508_);
  nor (_03342_, _03341_, _03299_);
  nor (_03343_, _03342_, _03340_);
  not (_03344_, _03343_);
  nor (_03345_, _03344_, _03339_);
  and (_03346_, _03345_, _03334_);
  and (_03347_, _03346_, _03326_);
  not (_03348_, _03347_);
  nor (_03349_, _03348_, _03298_);
  and (_03350_, _03349_, _03266_);
  and (_03351_, _03350_, _03225_);
  and (_03352_, _03351_, _03215_);
  not (_03353_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_03354_, _02835_, _02888_);
  not (_03355_, _03354_);
  and (_03356_, _02835_, _03106_);
  and (_03357_, _02835_, _02950_);
  or (_03358_, _02837_, _03084_);
  and (_03359_, _02835_, _02974_);
  and (_03360_, _02845_, _03071_);
  not (_03361_, _03360_);
  not (_03362_, _02885_);
  and (_03363_, _02852_, _03071_);
  nor (_03364_, _03363_, _03310_);
  and (_03365_, _03364_, _03362_);
  and (_03366_, _03365_, _03361_);
  nor (_03367_, _03366_, _02543_);
  and (_03368_, _02844_, _02495_);
  and (_03369_, _03368_, _03071_);
  and (_03370_, _02862_, _02884_);
  nor (_03371_, _03370_, _03369_);
  not (_03372_, _03371_);
  nor (_03373_, _03372_, _03367_);
  and (_03374_, _02944_, _02879_);
  or (_03375_, _03374_, _02886_);
  and (_03376_, _03375_, _02462_);
  and (_03377_, _02960_, _02879_);
  and (_03378_, _02844_, _02462_);
  and (_03379_, _03378_, _02879_);
  and (_03380_, _02862_, _03071_);
  or (_03381_, _03380_, _02974_);
  or (_03382_, _03381_, _03379_);
  or (_03383_, _03382_, _03377_);
  nor (_03384_, _03383_, _03376_);
  and (_03385_, _03384_, _03373_);
  or (_03386_, _03385_, _03359_);
  not (_03387_, _03072_);
  or (_03388_, _02835_, _03387_);
  and (_03389_, _03388_, _02881_);
  nand (_03390_, _03389_, _03386_);
  nand (_03391_, _02882_, _03390_);
  and (_03392_, _02845_, _02874_);
  nor (_03393_, _03392_, _03318_);
  nor (_03394_, _03393_, _02543_);
  and (_03395_, _03069_, _02866_);
  nor (_03396_, _03395_, _03075_);
  and (_03397_, _02840_, _02874_);
  and (_03398_, _03368_, _02874_);
  and (_03399_, _02852_, _02874_);
  and (_03400_, _03399_, _02462_);
  or (_03401_, _03400_, _03398_);
  nor (_03402_, _03401_, _03397_);
  nand (_03403_, _03402_, _03396_);
  nor (_03404_, _03403_, _03394_);
  nand (_03405_, _03404_, _03391_);
  nand (_03406_, _03405_, _03358_);
  and (_03407_, _03406_, _02877_);
  or (_03408_, _02878_, _03407_);
  and (_03409_, _02837_, _02875_);
  not (_03410_, _03368_);
  and (_03411_, _02861_, _02577_);
  nor (_03412_, _03411_, _02578_);
  and (_03413_, _03412_, _03410_);
  or (_03414_, _03413_, _02613_);
  nor (_03415_, _02961_, _02946_);
  and (_03416_, _03415_, _03414_);
  not (_03417_, _03416_);
  nor (_03418_, _03417_, _03409_);
  and (_03419_, _03418_, _03408_);
  or (_03420_, _03419_, _03357_);
  nand (_03421_, _03420_, _03064_);
  nor (_03422_, _02795_, _03064_);
  nor (_03423_, _03422_, _03059_);
  nand (_03424_, _03423_, _03421_);
  and (_03425_, _02837_, _03059_);
  and (_03426_, _03411_, _03099_);
  nor (_03427_, _03426_, _03103_);
  not (_03428_, _03427_);
  nor (_03429_, _03428_, _03425_);
  and (_03430_, _03429_, _03424_);
  nor (_03431_, _02795_, _03102_);
  or (_03432_, _03431_, _03430_);
  and (_03433_, _02854_, _02580_);
  and (_03434_, _02852_, _02580_);
  nor (_03435_, _03434_, _03433_);
  nor (_03436_, _03435_, _02543_);
  not (_03437_, _03436_);
  and (_03438_, _02840_, _02580_);
  not (_03439_, _03438_);
  and (_03440_, _02861_, _02429_);
  and (_03441_, _03440_, _02580_);
  nor (_03442_, _03441_, _03106_);
  and (_03443_, _03442_, _03439_);
  and (_03444_, _03443_, _03437_);
  and (_03445_, _03444_, _03432_);
  or (_03446_, _03445_, _03356_);
  and (_03447_, _03446_, _02864_);
  or (_03448_, _02865_, _03447_);
  and (_03449_, _03411_, _02517_);
  and (_03450_, _03368_, _02517_);
  nor (_03451_, _03450_, _03449_);
  and (_03452_, _03440_, _02517_);
  nor (_03453_, _03452_, _02841_);
  and (_03454_, _03453_, _03451_);
  and (_03455_, _03454_, _03448_);
  and (_03456_, _03015_, _01286_);
  and (_03457_, _03038_, _01280_);
  nor (_03458_, _03457_, _03456_);
  and (_03459_, _03002_, _01275_);
  and (_03460_, _03033_, _01303_);
  nor (_03461_, _03460_, _03459_);
  and (_03462_, _03461_, _03458_);
  and (_03463_, _03012_, _41922_);
  and (_03464_, _03049_, _01282_);
  nor (_03465_, _03464_, _03463_);
  and (_03466_, _03019_, _01296_);
  and (_03467_, _03046_, _01269_);
  nor (_03468_, _03467_, _03466_);
  and (_03469_, _03468_, _03465_);
  and (_03470_, _03469_, _03462_);
  and (_03471_, _03005_, _01273_);
  and (_03472_, _03040_, _01278_);
  nor (_03473_, _03472_, _03471_);
  and (_03474_, _03024_, _01267_);
  and (_03475_, _03052_, _01305_);
  nor (_03476_, _03475_, _03474_);
  and (_03477_, _03476_, _03473_);
  and (_03478_, _03044_, _01292_);
  and (_03479_, _03035_, _01300_);
  nor (_03480_, _03479_, _03478_);
  and (_03481_, _03021_, _01294_);
  and (_03482_, _03026_, _01265_);
  nor (_03483_, _03482_, _03481_);
  and (_03484_, _03483_, _03480_);
  and (_03485_, _03484_, _03477_);
  and (_03486_, _03485_, _03470_);
  and (_03487_, _03486_, _02579_);
  nor (_03488_, _03487_, _02933_);
  and (_03489_, _03488_, _03455_);
  not (_03490_, _02933_);
  nor (_03491_, _02795_, _03490_);
  or (_03492_, _03491_, _03489_);
  and (_03493_, _03411_, _02513_);
  nor (_03494_, _03493_, _02932_);
  and (_03495_, _03494_, _03492_);
  not (_03496_, _02932_);
  nor (_03497_, _02795_, _03496_);
  or (_03498_, _03497_, _03495_);
  and (_03499_, _03368_, _02508_);
  not (_03500_, _03499_);
  and (_03501_, _02960_, _02508_);
  not (_03502_, _03501_);
  and (_03503_, _02840_, _02508_);
  and (_03504_, _03411_, _02508_);
  nor (_03506_, _03504_, _03503_);
  and (_03507_, _03506_, _03502_);
  and (_03508_, _02844_, _02861_);
  and (_03509_, _03508_, _02508_);
  not (_03510_, _03509_);
  and (_03511_, _03510_, _03507_);
  and (_03512_, _03511_, _03500_);
  and (_03513_, _03512_, _03498_);
  nor (_03514_, _02835_, _03131_);
  and (_03515_, _02840_, _02969_);
  not (_03516_, _03515_);
  and (_03517_, _03411_, _02969_);
  and (_03518_, _03368_, _02969_);
  nor (_03519_, _03518_, _03517_);
  and (_03520_, _02960_, _02969_);
  and (_03521_, _03508_, _02969_);
  nor (_03522_, _03521_, _03520_);
  and (_03523_, _03522_, _03519_);
  and (_03524_, _03523_, _03516_);
  not (_03525_, _03524_);
  nor (_03526_, _03525_, _03514_);
  and (_03527_, _03526_, _03513_);
  and (_03528_, _03368_, _02964_);
  not (_03529_, _03528_);
  nor (_03530_, _02835_, _03140_);
  and (_03531_, _03411_, _02964_);
  and (_03532_, _02960_, _02964_);
  not (_03533_, _03532_);
  and (_03534_, _02840_, _02964_);
  and (_03535_, _03508_, _02964_);
  nor (_03536_, _03535_, _03534_);
  nand (_03537_, _03536_, _03533_);
  or (_03538_, _03537_, _03531_);
  nor (_03539_, _03538_, _03530_);
  and (_03540_, _03539_, _03529_);
  and (_03541_, _03540_, _03527_);
  nor (_03542_, _02835_, _03126_);
  and (_03543_, _03508_, _02967_);
  nor (_03544_, _03543_, _03133_);
  and (_03545_, _02960_, _02967_);
  and (_03546_, _03368_, _02967_);
  nor (_03547_, _03546_, _03545_);
  and (_03548_, _02840_, _02967_);
  and (_03549_, _03411_, _02967_);
  nor (_03550_, _03549_, _03548_);
  and (_03551_, _03550_, _03547_);
  and (_03552_, _03551_, _03544_);
  not (_03553_, _03552_);
  nor (_03554_, _03553_, _03542_);
  and (_03555_, _03554_, _03541_);
  and (_03556_, _02835_, _03133_);
  or (_03557_, _03556_, _03555_);
  and (_03558_, _03145_, _02866_);
  nor (_03559_, _03558_, _02968_);
  and (_03560_, _03559_, _03557_);
  not (_03561_, _02968_);
  nor (_03562_, _02795_, _03561_);
  nor (_03563_, _03562_, _03560_);
  not (_03564_, _02799_);
  and (_03565_, _03564_, _03412_);
  nor (_03566_, _03565_, _02536_);
  nor (_03567_, _03566_, _03563_);
  and (_03568_, _02835_, _02894_);
  or (_03569_, _03568_, _03567_);
  and (_03570_, _02892_, _02866_);
  nor (_03571_, _03570_, _02940_);
  and (_03572_, _03571_, _03569_);
  nor (_03573_, _02795_, _03164_);
  or (_03574_, _03573_, _03572_);
  and (_03575_, _02852_, _02367_);
  and (_03576_, _03575_, _02462_);
  not (_03577_, _03576_);
  nor (_03578_, _02800_, _03163_);
  and (_03579_, _03578_, _03577_);
  and (_03580_, _03579_, _03574_);
  and (_03581_, _02835_, _03163_);
  or (_03582_, _03581_, _03580_);
  and (_03583_, _03582_, _02498_);
  or (_03584_, _02796_, _03583_);
  and (_03585_, _03411_, _02522_);
  and (_03586_, _03368_, _02522_);
  nor (_03587_, _03586_, _03585_);
  and (_03588_, _02960_, _02522_);
  not (_03589_, _03588_);
  and (_03590_, _02840_, _02522_);
  and (_03591_, _03508_, _02522_);
  nor (_03592_, _03591_, _03590_);
  and (_03593_, _03592_, _03589_);
  and (_03594_, _03593_, _02890_);
  and (_03595_, _03594_, _03587_);
  nand (_03596_, _03595_, _03584_);
  nand (_03597_, _03596_, _03355_);
  or (_03598_, _03597_, _03353_);
  and (_03599_, _02707_, _41950_);
  nor (_03600_, _02714_, _41269_);
  nor (_03601_, _03600_, _03599_);
  nor (_03602_, _02747_, _41670_);
  nor (_03603_, _02722_, _41228_);
  nor (_03604_, _03603_, _03602_);
  and (_03605_, _03604_, _03601_);
  nor (_03606_, _02753_, _41586_);
  nor (_03607_, _02729_, _41338_);
  nor (_03608_, _03607_, _03606_);
  nor (_03609_, _02733_, _41545_);
  nor (_03610_, _02735_, _41463_);
  nor (_03611_, _03610_, _03609_);
  and (_03612_, _03611_, _03608_);
  and (_03613_, _03612_, _03605_);
  nor (_03614_, _02740_, _41379_);
  nor (_03615_, _02742_, _41422_);
  nor (_03616_, _03615_, _03614_);
  nor (_03617_, _02745_, _41894_);
  nor (_03618_, _02718_, _41724_);
  nor (_03619_, _03618_, _03617_);
  and (_03620_, _03619_, _03616_);
  nor (_03621_, _02751_, _41780_);
  nor (_03622_, _02726_, _41627_);
  nor (_03623_, _03622_, _03621_);
  nor (_03624_, _02756_, _41836_);
  nor (_03625_, _02758_, _41504_);
  nor (_03626_, _03625_, _03624_);
  and (_03627_, _03626_, _03623_);
  and (_03628_, _03627_, _03620_);
  and (_03629_, _03628_, _03613_);
  nor (_03630_, _03629_, _02763_);
  and (_03631_, _03223_, _03630_);
  not (_03632_, _03631_);
  and (_03633_, _02880_, _03630_);
  not (_03634_, _03633_);
  nor (_03635_, _02745_, _41873_);
  nor (_03636_, _02756_, _41816_);
  nor (_03637_, _03636_, _03635_);
  nor (_03638_, _02733_, _41530_);
  nor (_03639_, _02740_, _41364_);
  nor (_03640_, _03639_, _03638_);
  and (_03641_, _03640_, _03637_);
  nor (_03642_, _02729_, _41311_);
  nor (_03643_, _02714_, _41254_);
  nor (_03644_, _03643_, _03642_);
  nor (_03645_, _02758_, _41489_);
  nor (_03646_, _02742_, _41405_);
  nor (_03647_, _03646_, _03645_);
  and (_03648_, _03647_, _03644_);
  and (_03649_, _03648_, _03641_);
  nor (_03650_, _02747_, _41653_);
  nor (_03651_, _02753_, _41571_);
  nor (_03652_, _03651_, _03650_);
  and (_03653_, _02707_, _41929_);
  nor (_03654_, _02751_, _41759_);
  nor (_03655_, _03654_, _03653_);
  and (_03656_, _03655_, _03652_);
  nor (_03657_, _02735_, _41448_);
  nor (_03658_, _02722_, _41213_);
  nor (_03659_, _03658_, _03657_);
  nor (_03660_, _02718_, _41703_);
  nor (_03661_, _02726_, _41612_);
  nor (_03662_, _03661_, _03660_);
  and (_03663_, _03662_, _03659_);
  and (_03664_, _03663_, _03656_);
  and (_03665_, _03664_, _03649_);
  nor (_03666_, _03264_, _03665_);
  not (_03667_, _03666_);
  and (_03668_, _03038_, _01325_);
  and (_03669_, _03049_, _01327_);
  nor (_03670_, _03669_, _03668_);
  and (_03671_, _03012_, _41929_);
  and (_03672_, _03046_, _01314_);
  nor (_03673_, _03672_, _03671_);
  and (_03674_, _03673_, _03670_);
  and (_03675_, _03035_, _01345_);
  and (_03676_, _03052_, _01350_);
  nor (_03677_, _03676_, _03675_);
  and (_03678_, _03002_, _01318_);
  and (_03679_, _03040_, _01323_);
  nor (_03680_, _03679_, _03678_);
  and (_03681_, _03680_, _03677_);
  and (_03682_, _03681_, _03674_);
  and (_03683_, _03021_, _01339_);
  and (_03684_, _03015_, _01331_);
  nor (_03685_, _03684_, _03683_);
  and (_03686_, _03019_, _01341_);
  and (_03687_, _03044_, _01337_);
  nor (_03688_, _03687_, _03686_);
  and (_03689_, _03688_, _03685_);
  and (_03690_, _03024_, _01312_);
  and (_03691_, _03026_, _01310_);
  nor (_03692_, _03691_, _03690_);
  and (_03693_, _03005_, _01320_);
  and (_03694_, _03033_, _01348_);
  nor (_03695_, _03694_, _03693_);
  and (_03696_, _03695_, _03692_);
  and (_03697_, _03696_, _03689_);
  and (_03698_, _03697_, _03682_);
  nor (_03699_, _03698_, _02838_);
  not (_03700_, \oc8051_golden_model_1.SP [1]);
  nor (_03701_, _03338_, _03700_);
  not (_03702_, _03701_);
  and (_03703_, _02947_, _02517_);
  not (_03704_, _03703_);
  nor (_03705_, _03543_, _03360_);
  and (_03707_, _03705_, _03704_);
  and (_03708_, _03508_, _02517_);
  and (_03709_, _02947_, _02580_);
  nor (_03710_, _03709_, _03708_);
  and (_03711_, _03508_, _02580_);
  and (_03712_, _02847_, _03071_);
  nor (_03713_, _03712_, _03711_);
  and (_03714_, _03713_, _03710_);
  and (_03715_, _03714_, _03707_);
  and (_03716_, _03715_, _03702_);
  and (_03717_, _02847_, _02522_);
  and (_03718_, _02845_, _02367_);
  nor (_03719_, _03718_, _03717_);
  and (_03720_, _03719_, _03325_);
  nor (_03721_, _03299_, _02536_);
  not (_03722_, _03721_);
  and (_03723_, _02845_, _02868_);
  nor (_03724_, _03312_, _03723_);
  and (_03725_, _03724_, _03722_);
  and (_03726_, _02947_, _02967_);
  nor (_03727_, _03726_, _03342_);
  and (_03728_, _03727_, _03725_);
  and (_03729_, _02845_, _02879_);
  and (_03730_, _02845_, _02891_);
  nor (_03731_, _03730_, _03729_);
  and (_03732_, _02845_, _02964_);
  nor (_03733_, _03732_, _03392_);
  and (_03734_, _03733_, _03731_);
  and (_03735_, _02845_, _02508_);
  nor (_03736_, _03735_, _03300_);
  and (_03737_, _02845_, _02522_);
  and (_03738_, _02845_, _02969_);
  nor (_03739_, _03738_, _03737_);
  and (_03740_, _03739_, _03736_);
  and (_03741_, _03740_, _03734_);
  and (_03742_, _03741_, _03728_);
  and (_03743_, _03742_, _03720_);
  and (_03744_, _03743_, _03716_);
  not (_03745_, _03744_);
  nor (_03746_, _03745_, _03699_);
  and (_03747_, _03746_, _03667_);
  and (_03748_, _03747_, _03634_);
  and (_03749_, _03748_, _03632_);
  not (_03750_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_03751_, _03596_, _03355_);
  or (_03752_, _03751_, _03750_);
  and (_03753_, _03752_, _03749_);
  nand (_03754_, _03753_, _03598_);
  not (_03755_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_03756_, _03751_, _03755_);
  not (_03757_, _03749_);
  not (_03758_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_03759_, _03597_, _03758_);
  and (_03760_, _03759_, _03757_);
  nand (_03761_, _03760_, _03756_);
  nand (_03762_, _03761_, _03754_);
  nand (_03763_, _03762_, _03352_);
  not (_03764_, _03352_);
  not (_03765_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_03766_, _03751_, _03765_);
  not (_03767_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_03768_, _03597_, _03767_);
  and (_03769_, _03768_, _03757_);
  nand (_03770_, _03769_, _03766_);
  not (_03771_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_03772_, _03597_, _03771_);
  not (_03773_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_03774_, _03751_, _03773_);
  and (_03775_, _03774_, _03749_);
  nand (_03776_, _03775_, _03772_);
  nand (_03777_, _03776_, _03770_);
  nand (_03778_, _03777_, _03764_);
  nand (_03779_, _03778_, _03763_);
  nand (_03780_, _03779_, _03177_);
  not (_03781_, _03177_);
  not (_03782_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03783_, _03751_, _03782_);
  nand (_03784_, _03751_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03785_, _03784_, _03757_);
  nand (_03786_, _03785_, _03783_);
  not (_03787_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03788_, _03597_, _03787_);
  nand (_03789_, _03597_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03790_, _03789_, _03749_);
  nand (_03791_, _03790_, _03788_);
  nand (_03792_, _03791_, _03786_);
  nand (_03793_, _03792_, _03352_);
  not (_03794_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03795_, _03751_, _03794_);
  nand (_03796_, _03751_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03797_, _03796_, _03757_);
  nand (_03798_, _03797_, _03795_);
  not (_03799_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03800_, _03597_, _03799_);
  nand (_03801_, _03597_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_03802_, _03801_, _03749_);
  nand (_03803_, _03802_, _03800_);
  nand (_03804_, _03803_, _03798_);
  nand (_03805_, _03804_, _03764_);
  nand (_03806_, _03805_, _03793_);
  nand (_03807_, _03806_, _03781_);
  and (_03808_, _03807_, _03780_);
  or (_03809_, _03808_, _02887_);
  not (_03810_, _02974_);
  nor (_03811_, _03810_, _02763_);
  not (_03812_, _03811_);
  and (_03813_, _02884_, _02578_);
  not (_03814_, _03813_);
  nor (_03815_, _03814_, _02763_);
  nor (_03816_, _03564_, _02610_);
  nor (_03817_, _03816_, _03815_);
  not (_03818_, _02611_);
  and (_03819_, _03815_, _02835_);
  or (_03820_, _03819_, _03818_);
  or (_03821_, _03820_, _03817_);
  nor (_03822_, _02611_, _02866_);
  nor (_03823_, _03564_, _02608_);
  nor (_03824_, _03823_, _03822_);
  and (_03825_, _03824_, _03821_);
  and (_03826_, _03825_, _03812_);
  and (_03827_, _03826_, _03809_);
  and (_03828_, _02835_, _03811_);
  nor (_03829_, _03828_, _03827_);
  nor (_03830_, _03829_, _02883_);
  not (_03831_, _03830_);
  and (_03832_, _03831_, _02882_);
  nor (_03833_, _02609_, _02866_);
  nor (_03834_, _03833_, _03832_);
  nor (_03835_, _03564_, _02620_);
  nor (_03836_, _03336_, _02763_);
  and (_03837_, _03836_, _02837_);
  nor (_03838_, _03837_, _03835_);
  and (_03839_, _03838_, _03834_);
  not (_03840_, _03399_);
  nor (_03841_, _03808_, _03840_);
  not (_03842_, _03841_);
  and (_03843_, _03842_, _03839_);
  nor (_03844_, _02877_, _02763_);
  nor (_03845_, _03084_, _02763_);
  and (_03846_, _03845_, _02837_);
  nor (_03847_, _03846_, _03844_);
  and (_03848_, _03847_, _03843_);
  nor (_03849_, _03848_, _02878_);
  nor (_03850_, _03849_, _02875_);
  and (_03851_, _02875_, _02866_);
  or (_03852_, _03851_, _03850_);
  and (_03853_, _03852_, _02873_);
  nor (_03854_, _03853_, _02871_);
  and (_03855_, _03059_, _02462_);
  or (_03856_, _03855_, _03854_);
  nor (_03857_, _03856_, _02867_);
  nor (_03858_, _02864_, _02763_);
  and (_03859_, _02852_, _03099_);
  not (_03860_, _03859_);
  nor (_03861_, _03808_, _03860_);
  nor (_03862_, _03861_, _03858_);
  and (_03863_, _03862_, _03857_);
  nor (_03864_, _03863_, _02865_);
  nor (_03865_, _03864_, _02581_);
  and (_03866_, _02581_, _02866_);
  nor (_03867_, _03866_, _03865_);
  and (_03868_, _02799_, _02513_);
  or (_03869_, _03868_, _03867_);
  nor (_03870_, _03869_, _02860_);
  and (_03871_, _02852_, _02513_);
  not (_03872_, _03808_);
  and (_03873_, _03872_, _03871_);
  nor (_03874_, _03873_, _02804_);
  and (_03875_, _03874_, _03870_);
  nor (_03876_, _03875_, _02836_);
  nor (_03877_, _03876_, _02514_);
  and (_03878_, _02514_, _02866_);
  nor (_03879_, _03878_, _03877_);
  not (_03880_, _02532_);
  nor (_03881_, _03137_, _02763_);
  not (_03882_, _03881_);
  not (_03883_, _02970_);
  nor (_03884_, _03883_, _02763_);
  not (_03885_, _03884_);
  nor (_03886_, _03128_, _02763_);
  not (_03887_, _02980_);
  nor (_03888_, _03887_, _02763_);
  nor (_03889_, _03888_, _03886_);
  and (_03890_, _03889_, _03885_);
  and (_03891_, _03890_, _03882_);
  nor (_03892_, _03891_, _02835_);
  nor (_03893_, _03892_, _03880_);
  not (_03894_, _03893_);
  nor (_03895_, _03894_, _03879_);
  nor (_03896_, _02532_, \oc8051_golden_model_1.SP [0]);
  nor (_03897_, _03896_, _03895_);
  not (_03898_, _02529_);
  nor (_03899_, _03124_, _02763_);
  and (_03900_, _03899_, _02837_);
  nor (_03901_, _03900_, _03898_);
  not (_03902_, _03901_);
  nor (_03903_, _03902_, _03897_);
  nor (_03904_, _03903_, _02801_);
  nor (_03905_, _03904_, _02800_);
  not (_03906_, _03163_);
  nor (_03908_, _03906_, _02763_);
  not (_03909_, _03575_);
  nor (_03910_, _03808_, _03909_);
  nor (_03911_, _03910_, _03908_);
  and (_03912_, _03911_, _03905_);
  and (_03913_, _03908_, _02835_);
  nor (_03914_, _03913_, _03912_);
  nor (_03915_, _02939_, _02525_);
  nor (_03916_, _03915_, _02866_);
  nor (_03917_, _03916_, _03914_);
  and (_03918_, _03917_, _02798_);
  nor (_03919_, _03918_, _02796_);
  and (_03920_, _02852_, _02522_);
  not (_03921_, _03920_);
  nor (_03922_, _03808_, _03921_);
  nor (_03923_, _02890_, _02763_);
  and (_03924_, _02799_, _02522_);
  or (_03925_, _03924_, _03923_);
  or (_03926_, _03925_, _03922_);
  nor (_03927_, _03926_, _03919_);
  and (_03928_, _03923_, _02835_);
  nor (_03929_, _03928_, _03927_);
  not (_03930_, _03929_);
  and (_03931_, _03630_, _02497_);
  and (_03932_, _03700_, \oc8051_golden_model_1.SP [0]);
  and (_03933_, \oc8051_golden_model_1.SP [1], _02866_);
  nor (_03934_, _03933_, _03932_);
  nor (_03935_, _03934_, _02529_);
  not (_03936_, _03665_);
  and (_03937_, _02804_, _03936_);
  and (_03938_, _02863_, _03630_);
  not (_03939_, _03934_);
  and (_03940_, _02875_, _03939_);
  not (_03941_, _02875_);
  and (_03942_, _03811_, _03936_);
  not (_03943_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03944_, _03597_, _03943_);
  not (_03945_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_03946_, _03751_, _03945_);
  and (_03947_, _03946_, _03749_);
  nand (_03948_, _03947_, _03944_);
  not (_03949_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03950_, _03751_, _03949_);
  not (_03951_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03952_, _03597_, _03951_);
  and (_03953_, _03952_, _03757_);
  nand (_03954_, _03953_, _03950_);
  nand (_03955_, _03954_, _03948_);
  nand (_03956_, _03955_, _03352_);
  not (_03957_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03958_, _03751_, _03957_);
  not (_03959_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03960_, _03597_, _03959_);
  and (_03961_, _03960_, _03757_);
  nand (_03962_, _03961_, _03958_);
  not (_03963_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03964_, _03597_, _03963_);
  not (_03965_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03966_, _03751_, _03965_);
  and (_03967_, _03966_, _03749_);
  nand (_03968_, _03967_, _03964_);
  nand (_03969_, _03968_, _03962_);
  nand (_03970_, _03969_, _03764_);
  nand (_03971_, _03970_, _03956_);
  nand (_03972_, _03971_, _03177_);
  not (_03973_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03974_, _03751_, _03973_);
  nand (_03975_, _03751_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03976_, _03975_, _03757_);
  nand (_03977_, _03976_, _03974_);
  not (_03978_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_03979_, _03597_, _03978_);
  nand (_03980_, _03597_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03981_, _03980_, _03749_);
  nand (_03982_, _03981_, _03979_);
  nand (_03983_, _03982_, _03977_);
  nand (_03984_, _03983_, _03352_);
  not (_03985_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_03986_, _03751_, _03985_);
  nand (_03987_, _03751_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_03988_, _03987_, _03757_);
  nand (_03989_, _03988_, _03986_);
  not (_03990_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03991_, _03597_, _03990_);
  not (_03992_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_03993_, _03751_, _03992_);
  and (_03994_, _03993_, _03749_);
  nand (_03995_, _03994_, _03991_);
  nand (_03996_, _03995_, _03989_);
  nand (_03997_, _03996_, _03764_);
  nand (_03998_, _03997_, _03984_);
  nand (_03999_, _03998_, _03781_);
  and (_04000_, _03999_, _03972_);
  or (_04001_, _04000_, _02887_);
  and (_04002_, _02494_, _02429_);
  and (_04003_, _04002_, _02884_);
  nor (_04004_, _04003_, _03815_);
  and (_04005_, _03815_, _03936_);
  or (_04006_, _04005_, _03818_);
  or (_04007_, _04006_, _04004_);
  and (_04008_, _03368_, _02879_);
  and (_04009_, _02844_, _02575_);
  and (_04010_, _04009_, _02879_);
  nor (_04011_, _04010_, _04008_);
  nor (_04012_, _03939_, _02611_);
  nor (_04013_, _04012_, _03374_);
  and (_04014_, _04013_, _04011_);
  and (_04015_, _04014_, _04007_);
  and (_04016_, _04015_, _03812_);
  and (_04017_, _04016_, _04001_);
  nor (_04018_, _04017_, _03942_);
  nor (_04019_, _04018_, _02883_);
  nor (_04020_, _04019_, _03633_);
  nor (_04021_, _03939_, _02609_);
  nor (_04022_, _04021_, _04020_);
  and (_04023_, _03836_, _03665_);
  and (_04024_, _04002_, _02874_);
  nor (_04025_, _04024_, _04023_);
  and (_04026_, _04025_, _04022_);
  nor (_04027_, _04000_, _03840_);
  nor (_04028_, _04027_, _03845_);
  and (_04029_, _04028_, _04026_);
  and (_04030_, _03845_, _03936_);
  nor (_04031_, _04030_, _04029_);
  and (_04032_, _03844_, _03629_);
  nor (_04033_, _04032_, _04031_);
  and (_04034_, _04033_, _03941_);
  nor (_04035_, _04034_, _03940_);
  and (_04036_, _02872_, _03629_);
  or (_04037_, _04036_, _04035_);
  and (_04038_, _04002_, _03099_);
  nor (_04039_, _03939_, _02614_);
  nor (_04040_, _04039_, _04038_);
  not (_04041_, _04040_);
  nor (_04042_, _04041_, _04037_);
  nor (_04043_, _04000_, _03860_);
  nor (_04044_, _04043_, _03858_);
  and (_04045_, _04044_, _04042_);
  nor (_04046_, _04045_, _03938_);
  nor (_04047_, _04046_, _02581_);
  and (_04048_, _03939_, _02581_);
  nor (_04049_, _04048_, _04047_);
  and (_04050_, _02859_, _03665_);
  and (_04051_, _04002_, _02513_);
  nor (_04052_, _04051_, _04050_);
  not (_04053_, _04052_);
  nor (_04054_, _04053_, _04049_);
  not (_04055_, _04000_);
  and (_04056_, _04055_, _03871_);
  nor (_04057_, _04056_, _02804_);
  and (_04058_, _04057_, _04054_);
  nor (_04059_, _04058_, _03937_);
  nor (_04060_, _04059_, _02514_);
  and (_04061_, _03939_, _02514_);
  nor (_04062_, _04061_, _04060_);
  nor (_04063_, _03891_, _03936_);
  nor (_04064_, _04063_, _03880_);
  not (_04065_, _04064_);
  nor (_04066_, _04065_, _04062_);
  nor (_04067_, _03934_, _02532_);
  nor (_04068_, _04067_, _04066_);
  and (_04069_, _03899_, _03665_);
  nor (_04070_, _04069_, _03898_);
  not (_04071_, _04070_);
  nor (_04072_, _04071_, _04068_);
  nor (_04073_, _04072_, _03935_);
  and (_04074_, _04002_, _02367_);
  nor (_04075_, _04074_, _04073_);
  nor (_04076_, _04000_, _03909_);
  nor (_04077_, _04076_, _03908_);
  and (_04078_, _04077_, _04075_);
  and (_04079_, _03908_, _03936_);
  nor (_04080_, _04079_, _04078_);
  nor (_04081_, _03915_, _03939_);
  nor (_04082_, _04081_, _02797_);
  not (_04083_, _04082_);
  nor (_04084_, _04083_, _04080_);
  nor (_04085_, _04084_, _03931_);
  and (_04086_, _04002_, _02522_);
  nor (_04087_, _04086_, _04085_);
  nor (_04088_, _04000_, _03921_);
  nor (_04089_, _04088_, _03923_);
  and (_04090_, _04089_, _04087_);
  and (_04091_, _03923_, _03936_);
  nor (_04092_, _04091_, _04090_);
  not (_04093_, _02514_);
  and (_04094_, _02533_, _04093_);
  not (_04095_, _02614_);
  nor (_04096_, _04095_, _02581_);
  and (_04097_, _04096_, _02612_);
  and (_04098_, _04097_, _04094_);
  and (_04099_, _02944_, _02522_);
  not (_04100_, _04099_);
  and (_04101_, _02844_, _02513_);
  and (_04102_, _04101_, _02575_);
  and (_04103_, _03059_, _02398_);
  nor (_04104_, _04103_, _04102_);
  and (_04105_, _04104_, _04100_);
  nor (_04106_, _03575_, _03871_);
  and (_04107_, _04106_, _03915_);
  and (_04109_, _04101_, _02495_);
  nor (_04110_, _04109_, _03398_);
  and (_04111_, _04110_, _04107_);
  and (_04112_, _04111_, _04105_);
  and (_04113_, _04112_, _04098_);
  and (_04114_, _02844_, _03099_);
  and (_04115_, _04114_, _02493_);
  not (_04116_, _04115_);
  nor (_04117_, _03586_, _03920_);
  not (_04118_, _04117_);
  and (_04119_, _02854_, _02522_);
  and (_04120_, _04119_, _02543_);
  nor (_04121_, _04120_, _04118_);
  and (_04122_, _04121_, _04116_);
  and (_04123_, _04011_, _03719_);
  and (_04124_, _02947_, _02513_);
  not (_04125_, _04124_);
  and (_04126_, _02840_, _02513_);
  and (_04127_, _03508_, _02513_);
  nor (_04128_, _04127_, _04126_);
  and (_04129_, _04128_, _04125_);
  and (_04130_, _02854_, _03099_);
  not (_04131_, _04130_);
  and (_04132_, _04131_, _04129_);
  and (_04133_, _04132_, _04123_);
  nor (_04134_, _03317_, _03303_);
  nor (_04135_, _03737_, _03729_);
  and (_04136_, _04135_, _04134_);
  nor (_04137_, _03859_, _02875_);
  nor (_04138_, _03309_, _02620_);
  nor (_04139_, _03399_, _04138_);
  and (_04140_, _04139_, _04137_);
  and (_04141_, _04140_, _04136_);
  and (_04142_, _02844_, _02884_);
  nor (_04143_, _03309_, _02608_);
  nor (_04144_, _04143_, _04142_);
  and (_04145_, _02846_, _02513_);
  and (_04146_, _02847_, _02513_);
  or (_04147_, _04146_, _04145_);
  not (_04148_, _02844_);
  nor (_04149_, _04148_, _02495_);
  and (_04150_, _04149_, _02874_);
  nor (_04151_, _04150_, _04147_);
  and (_04152_, _04151_, _04144_);
  and (_04153_, _02854_, _02367_);
  nor (_04154_, _03309_, _02610_);
  nor (_04155_, _04154_, _04153_);
  and (_04156_, _04155_, _02887_);
  and (_04157_, _04156_, _04152_);
  and (_04158_, _04157_, _04141_);
  and (_04159_, _04158_, _04133_);
  and (_04160_, _04159_, _04122_);
  and (_04161_, _04160_, _04113_);
  and (_04162_, _04161_, _02798_);
  nor (_04163_, _03844_, _02872_);
  nor (_04164_, _03899_, _02804_);
  and (_04165_, _04164_, _04163_);
  and (_04166_, _04165_, _04162_);
  nor (_04167_, _03845_, _03858_);
  nor (_04168_, _03908_, _03881_);
  and (_04169_, _04168_, _04167_);
  nor (_04170_, _03836_, _02883_);
  nor (_04171_, _03815_, _03811_);
  and (_04172_, _04171_, _04170_);
  and (_04173_, _04172_, _04169_);
  nor (_04174_, _02857_, _02763_);
  not (_04175_, _04174_);
  nor (_04176_, _02763_, _02838_);
  nor (_04177_, _03923_, _04176_);
  and (_04178_, _04177_, _04175_);
  and (_04179_, _04178_, _03890_);
  and (_04180_, _04179_, _04173_);
  and (_04181_, _04180_, _04166_);
  and (_04182_, _43220_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_04183_, _04182_);
  nor (_04184_, _04183_, _04181_);
  not (_04185_, _04184_);
  nor (_04186_, _04185_, _04092_);
  and (_04187_, _04186_, _03930_);
  not (_04188_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04189_, _03597_, _04188_);
  not (_04190_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_04191_, _03751_, _04190_);
  and (_04192_, _04191_, _03749_);
  nand (_04193_, _04192_, _04189_);
  not (_04194_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_04195_, _03751_, _04194_);
  not (_04196_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04197_, _03597_, _04196_);
  and (_04198_, _04197_, _03757_);
  nand (_04199_, _04198_, _04195_);
  nand (_04200_, _04199_, _04193_);
  nand (_04201_, _04200_, _03352_);
  not (_04202_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04203_, _03751_, _04202_);
  not (_04204_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04205_, _03597_, _04204_);
  and (_04206_, _04205_, _03757_);
  nand (_04207_, _04206_, _04203_);
  not (_04208_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04209_, _03597_, _04208_);
  not (_04210_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04211_, _03751_, _04210_);
  and (_04212_, _04211_, _03749_);
  nand (_04213_, _04212_, _04209_);
  nand (_04214_, _04213_, _04207_);
  nand (_04215_, _04214_, _03764_);
  nand (_04216_, _04215_, _04201_);
  nand (_04217_, _04216_, _03177_);
  nand (_04218_, _03597_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04219_, _03751_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04220_, _04219_, _03757_);
  nand (_04221_, _04220_, _04218_);
  nand (_04222_, _03751_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04223_, _03597_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04224_, _04223_, _03749_);
  nand (_04225_, _04224_, _04222_);
  nand (_04226_, _04225_, _04221_);
  nand (_04227_, _04226_, _03352_);
  nand (_04228_, _03597_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04229_, _03751_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04230_, _04229_, _03757_);
  nand (_04231_, _04230_, _04228_);
  nand (_04232_, _03751_, \oc8051_golden_model_1.IRAM[12] [3]);
  not (_04233_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_04234_, _03751_, _04233_);
  and (_04235_, _04234_, _03749_);
  nand (_04236_, _04235_, _04232_);
  nand (_04237_, _04236_, _04231_);
  nand (_04238_, _04237_, _03764_);
  nand (_04239_, _04238_, _04227_);
  nand (_04240_, _04239_, _03781_);
  and (_04241_, _04240_, _04217_);
  nor (_04242_, _04241_, _03921_);
  and (_04243_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04244_, _04243_, \oc8051_golden_model_1.SP [2]);
  or (_04245_, _04244_, \oc8051_golden_model_1.SP [3]);
  and (_04246_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04247_, _04246_, \oc8051_golden_model_1.SP [3]);
  nand (_04248_, _04247_, \oc8051_golden_model_1.SP [0]);
  and (_04249_, _04248_, _04245_);
  and (_04250_, _04249_, _02581_);
  not (_04251_, _02581_);
  not (_04252_, _02609_);
  nand (_04253_, _02927_, _02883_);
  or (_04254_, _02885_, \oc8051_golden_model_1.PSW [3]);
  or (_04255_, _04241_, _03362_);
  and (_04256_, _04255_, _04254_);
  or (_04257_, _04256_, _03815_);
  nand (_04258_, _03815_, _02794_);
  and (_04259_, _04258_, _02611_);
  and (_04260_, _04259_, _04257_);
  not (_04261_, _04249_);
  nor (_04262_, _04261_, _02611_);
  or (_04263_, _04262_, _02886_);
  or (_04264_, _04263_, _04260_);
  not (_04265_, _02886_);
  or (_04266_, _04241_, _04265_);
  and (_04267_, _04266_, _03812_);
  and (_04268_, _04267_, _04264_);
  nor (_04269_, _02795_, _03810_);
  or (_04270_, _04269_, _02883_);
  or (_04271_, _04270_, _04268_);
  and (_04272_, _04271_, _04253_);
  or (_04273_, _04272_, _04252_);
  nor (_04274_, _04249_, _02609_);
  nor (_04275_, _04274_, _03836_);
  and (_04276_, _04275_, _04273_);
  and (_04277_, _03836_, _02929_);
  or (_04278_, _04277_, _03399_);
  or (_04279_, _04278_, _04276_);
  nor (_04280_, _04241_, _03840_);
  nor (_04281_, _04280_, _03845_);
  and (_04282_, _04281_, _04279_);
  nor (_04283_, _02795_, _03084_);
  or (_04284_, _04283_, _03844_);
  or (_04285_, _04284_, _04282_);
  nand (_04286_, _03844_, _02927_);
  and (_04287_, _04286_, _03941_);
  and (_04288_, _04287_, _04285_);
  and (_04289_, _04249_, _02875_);
  or (_04290_, _04289_, _02872_);
  or (_04291_, _04290_, _04288_);
  nand (_04292_, _02927_, _02872_);
  and (_04293_, _04292_, _02614_);
  and (_04294_, _04293_, _04291_);
  nor (_04295_, _04261_, _02614_);
  or (_04296_, _04295_, _03859_);
  or (_04297_, _04296_, _04294_);
  not (_04298_, _03858_);
  or (_04299_, _04241_, _03860_);
  and (_04300_, _04299_, _04298_);
  and (_04301_, _04300_, _04297_);
  nor (_04302_, _04298_, _02931_);
  or (_04303_, _04302_, _04301_);
  and (_04304_, _04303_, _04251_);
  nor (_04305_, _04304_, _04250_);
  nor (_04306_, _04305_, _02859_);
  and (_04307_, _02859_, _02929_);
  or (_04308_, _04307_, _03871_);
  or (_04310_, _04308_, _04306_);
  not (_04311_, _04241_);
  and (_04312_, _04311_, _03871_);
  nor (_04313_, _04312_, _02804_);
  and (_04314_, _04313_, _04310_);
  and (_04315_, _02929_, _02804_);
  or (_04316_, _04315_, _04314_);
  and (_04317_, _04316_, _04093_);
  nand (_04318_, _04249_, _02514_);
  nand (_04319_, _04318_, _03891_);
  or (_04320_, _04319_, _04317_);
  or (_04321_, _03891_, _02929_);
  and (_04322_, _04321_, _02532_);
  and (_04323_, _04322_, _04320_);
  nor (_04324_, _04261_, _02532_);
  or (_04325_, _04324_, _03899_);
  or (_04326_, _04325_, _04323_);
  nand (_04327_, _03899_, _02794_);
  and (_04328_, _04327_, _02529_);
  and (_04329_, _04328_, _04326_);
  nor (_04330_, _04261_, _02529_);
  or (_04331_, _04330_, _03575_);
  or (_04332_, _04331_, _04329_);
  not (_04333_, _03908_);
  or (_04334_, _04241_, _03909_);
  and (_04335_, _04334_, _04333_);
  and (_04336_, _04335_, _04332_);
  not (_04337_, _03915_);
  and (_04338_, _03908_, _02929_);
  or (_04339_, _04338_, _04337_);
  or (_04340_, _04339_, _04336_);
  nor (_04341_, _04249_, _03915_);
  nor (_04342_, _04341_, _02797_);
  and (_04343_, _04342_, _04340_);
  not (_04344_, _02927_);
  and (_04345_, _04344_, _02797_);
  or (_04346_, _04345_, _03920_);
  nor (_04347_, _04346_, _04343_);
  or (_04348_, _04347_, _03923_);
  nor (_04349_, _04348_, _04242_);
  and (_04350_, _03923_, _02929_);
  nor (_04351_, _04350_, _04349_);
  not (_04352_, _04351_);
  and (_04353_, _02844_, _02522_);
  and (_04354_, _03212_, _02497_);
  nor (_04355_, _04243_, \oc8051_golden_model_1.SP [2]);
  nor (_04356_, _04355_, _04244_);
  not (_04358_, _04356_);
  nor (_04359_, _04358_, _02529_);
  not (_04361_, _03256_);
  and (_04362_, _04361_, _02804_);
  and (_04364_, _03212_, _02863_);
  and (_04365_, _04356_, _02875_);
  and (_04367_, _04361_, _03811_);
  not (_04368_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_04370_, _03597_, _04368_);
  not (_04371_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_04373_, _03751_, _04371_);
  and (_04374_, _04373_, _03749_);
  nand (_04376_, _04374_, _04370_);
  not (_04377_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_04379_, _03751_, _04377_);
  not (_04380_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04382_, _03597_, _04380_);
  and (_04383_, _04382_, _03757_);
  nand (_04385_, _04383_, _04379_);
  nand (_04386_, _04385_, _04376_);
  nand (_04388_, _04386_, _03352_);
  not (_04389_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_04391_, _03751_, _04389_);
  not (_04392_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04394_, _03597_, _04392_);
  and (_04395_, _04394_, _03757_);
  nand (_04396_, _04395_, _04391_);
  not (_04397_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04398_, _03597_, _04397_);
  not (_04399_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_04400_, _03751_, _04399_);
  and (_04401_, _04400_, _03749_);
  nand (_04402_, _04401_, _04398_);
  nand (_04403_, _04402_, _04396_);
  nand (_04404_, _04403_, _03764_);
  nand (_04405_, _04404_, _04388_);
  nand (_04406_, _04405_, _03177_);
  not (_04407_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_04408_, _03751_, _04407_);
  not (_04409_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04410_, _03597_, _04409_);
  and (_04411_, _04410_, _03757_);
  nand (_04412_, _04411_, _04408_);
  nand (_04413_, _03751_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_04414_, _03597_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04415_, _04414_, _03749_);
  nand (_04416_, _04415_, _04413_);
  nand (_04417_, _04416_, _04412_);
  nand (_04418_, _04417_, _03352_);
  not (_04419_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_04420_, _03751_, _04419_);
  not (_04421_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04422_, _03597_, _04421_);
  and (_04424_, _04422_, _03757_);
  nand (_04425_, _04424_, _04420_);
  nand (_04426_, _03751_, \oc8051_golden_model_1.IRAM[12] [2]);
  not (_04427_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_04428_, _03751_, _04427_);
  and (_04429_, _04428_, _03749_);
  nand (_04430_, _04429_, _04426_);
  nand (_04431_, _04430_, _04425_);
  nand (_04432_, _04431_, _03764_);
  nand (_04433_, _04432_, _04418_);
  nand (_04434_, _04433_, _03781_);
  and (_04435_, _04434_, _04406_);
  or (_04436_, _04435_, _02887_);
  nor (_04437_, _04142_, _03815_);
  and (_04438_, _03815_, _04361_);
  or (_04439_, _04438_, _03818_);
  or (_04440_, _04439_, _04437_);
  nor (_04441_, _04356_, _02611_);
  and (_04442_, _02844_, _02879_);
  nor (_04443_, _04442_, _04441_);
  and (_04444_, _04443_, _04440_);
  and (_04445_, _04444_, _03812_);
  and (_04446_, _04445_, _04436_);
  nor (_04447_, _04446_, _04367_);
  nor (_04448_, _04447_, _02883_);
  nor (_04449_, _04448_, _03214_);
  nor (_04450_, _04356_, _02609_);
  nor (_04451_, _04450_, _04449_);
  and (_04452_, _03836_, _03256_);
  and (_04454_, _02844_, _02874_);
  nor (_04456_, _04454_, _04452_);
  and (_04457_, _04456_, _04451_);
  nor (_04459_, _04435_, _03840_);
  nor (_04460_, _04459_, _03845_);
  and (_04462_, _04460_, _04457_);
  and (_04463_, _03845_, _04361_);
  nor (_04465_, _04463_, _04462_);
  and (_04466_, _03844_, _03211_);
  nor (_04468_, _04466_, _04465_);
  and (_04469_, _04468_, _03941_);
  nor (_04471_, _04469_, _04365_);
  and (_04472_, _03211_, _02872_);
  or (_04474_, _04472_, _04471_);
  nor (_04475_, _04356_, _02614_);
  nor (_04477_, _04475_, _04114_);
  not (_04478_, _04477_);
  nor (_04480_, _04478_, _04474_);
  nor (_04481_, _04435_, _03860_);
  nor (_04483_, _04481_, _03858_);
  and (_04484_, _04483_, _04480_);
  nor (_04486_, _04484_, _04364_);
  nor (_04487_, _04486_, _02581_);
  and (_04488_, _04356_, _02581_);
  nor (_04489_, _04488_, _04487_);
  and (_04490_, _02859_, _03256_);
  nor (_04491_, _04490_, _04101_);
  not (_04492_, _04491_);
  nor (_04493_, _04492_, _04489_);
  not (_04494_, _04435_);
  and (_04495_, _04494_, _03871_);
  nor (_04496_, _04495_, _02804_);
  and (_04497_, _04496_, _04493_);
  nor (_04498_, _04497_, _04362_);
  nor (_04499_, _04498_, _02514_);
  and (_04500_, _04356_, _02514_);
  nor (_04501_, _04500_, _04499_);
  nor (_04502_, _03891_, _04361_);
  nor (_04503_, _04502_, _03880_);
  not (_04504_, _04503_);
  nor (_04505_, _04504_, _04501_);
  nor (_04506_, _04358_, _02532_);
  nor (_04507_, _04506_, _04505_);
  and (_04508_, _03899_, _03256_);
  nor (_04509_, _04508_, _03898_);
  not (_04510_, _04509_);
  nor (_04511_, _04510_, _04507_);
  nor (_04512_, _04511_, _04359_);
  nor (_04513_, _04153_, _03718_);
  not (_04514_, _04513_);
  nor (_04515_, _04514_, _04512_);
  nor (_04516_, _04435_, _03909_);
  nor (_04517_, _04516_, _03908_);
  and (_04518_, _04517_, _04515_);
  and (_04519_, _03908_, _04361_);
  nor (_04520_, _04519_, _04518_);
  nor (_04521_, _04356_, _03915_);
  nor (_04522_, _04521_, _02797_);
  not (_04523_, _04522_);
  nor (_04524_, _04523_, _04520_);
  nor (_04525_, _04524_, _04354_);
  nor (_04526_, _04525_, _04353_);
  nor (_04527_, _04435_, _03921_);
  nor (_04528_, _04527_, _03923_);
  and (_04529_, _04528_, _04526_);
  and (_04530_, _03923_, _04361_);
  nor (_04531_, _04530_, _04529_);
  nor (_04532_, _04185_, _04531_);
  and (_04533_, _04532_, _04352_);
  and (_04534_, _04533_, _04187_);
  or (_04535_, _04534_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04537_, _04246_, _02866_);
  nor (_04538_, _04356_, _03933_);
  nor (_04539_, _04538_, _04537_);
  and (_04540_, _04247_, _02866_);
  nor (_04541_, _04537_, _04249_);
  nor (_04542_, _04541_, _04540_);
  and (_04543_, _04098_, _03915_);
  nor (_04544_, _04543_, _04183_);
  and (_04545_, _04544_, _04542_);
  and (_04546_, _04545_, _04539_);
  and (_04547_, _04546_, _03932_);
  not (_04548_, _04547_);
  and (_04549_, _04548_, _04535_);
  not (_04550_, _04534_);
  not (_04551_, _02763_);
  nand (_04552_, _03751_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand (_04553_, _03597_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_04554_, _04553_, _03749_);
  nand (_04555_, _04554_, _04552_);
  not (_04556_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_04557_, _03751_, _04556_);
  not (_04558_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_04559_, _03597_, _04558_);
  and (_04560_, _04559_, _03757_);
  nand (_04561_, _04560_, _04557_);
  nand (_04562_, _04561_, _04555_);
  nand (_04563_, _04562_, _03352_);
  not (_04564_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_04565_, _03751_, _04564_);
  not (_04566_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04567_, _03597_, _04566_);
  and (_04568_, _04567_, _03757_);
  nand (_04569_, _04568_, _04565_);
  nand (_04570_, _03751_, \oc8051_golden_model_1.IRAM[4] [7]);
  nand (_04571_, _03597_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_04572_, _04571_, _03749_);
  nand (_04573_, _04572_, _04570_);
  nand (_04574_, _04573_, _04569_);
  nand (_04575_, _04574_, _03764_);
  nand (_04576_, _04575_, _04563_);
  nand (_04577_, _04576_, _03177_);
  not (_04578_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_04579_, _03751_, _04578_);
  not (_04580_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04581_, _03597_, _04580_);
  and (_04582_, _04581_, _03757_);
  nand (_04583_, _04582_, _04579_);
  nand (_04584_, _03751_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_04585_, _03597_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_04586_, _04585_, _03749_);
  nand (_04587_, _04586_, _04584_);
  nand (_04588_, _04587_, _04583_);
  nand (_04589_, _04588_, _03352_);
  not (_04590_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_04591_, _03751_, _04590_);
  not (_04592_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04593_, _03597_, _04592_);
  and (_04594_, _04593_, _03757_);
  nand (_04595_, _04594_, _04591_);
  nand (_04596_, _03751_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_04597_, _03597_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_04598_, _04597_, _03749_);
  nand (_04599_, _04598_, _04596_);
  nand (_04600_, _04599_, _04595_);
  nand (_04601_, _04600_, _03764_);
  nand (_04602_, _04601_, _04589_);
  nand (_04603_, _04602_, _03781_);
  and (_04604_, _04603_, _04577_);
  nand (_04605_, _04604_, _04551_);
  and (_04606_, _02927_, _02763_);
  and (_04607_, _04606_, _03211_);
  and (_04608_, _04607_, _03629_);
  and (_04609_, _04608_, _02794_);
  nor (_04610_, _02835_, _03665_);
  and (_04611_, _04610_, _03256_);
  and (_04612_, _04611_, _04609_);
  and (_04613_, _04612_, \oc8051_golden_model_1.DPL [7]);
  not (_04614_, _04613_);
  and (_04615_, _02835_, _03665_);
  and (_04616_, _04615_, _03256_);
  and (_04617_, _04616_, _04609_);
  and (_04618_, _04617_, \oc8051_golden_model_1.SP [7]);
  and (_04619_, _02837_, _03665_);
  and (_04620_, _04619_, _03256_);
  and (_04621_, _04620_, _02929_);
  and (_04622_, _04621_, _04608_);
  and (_04623_, _04622_, \oc8051_golden_model_1.TCON [7]);
  nor (_04624_, _04623_, _04618_);
  and (_04625_, _04624_, _04614_);
  and (_04626_, _03256_, _02794_);
  and (_04627_, _04619_, _04626_);
  and (_04628_, _04627_, _04608_);
  and (_04629_, _04628_, \oc8051_golden_model_1.P0 [7]);
  not (_04630_, _04629_);
  not (_04631_, _03629_);
  and (_04632_, _03211_, _04631_);
  and (_04633_, _04632_, _04606_);
  and (_04634_, _04633_, _04627_);
  and (_04635_, _04634_, \oc8051_golden_model_1.P1 [7]);
  not (_04636_, _04635_);
  not (_04638_, _03211_);
  and (_04639_, _04638_, _03629_);
  and (_04640_, _04639_, _04606_);
  and (_04641_, _04640_, _04627_);
  and (_04642_, _04641_, \oc8051_golden_model_1.P2 [7]);
  nor (_04643_, _03211_, _03629_);
  and (_04644_, _04643_, _04606_);
  and (_04645_, _04644_, _04627_);
  and (_04646_, _04645_, \oc8051_golden_model_1.P3 [7]);
  nor (_04647_, _04646_, _04642_);
  and (_04648_, _04647_, _04636_);
  and (_04649_, _04648_, _04630_);
  and (_04650_, _04649_, _04625_);
  not (_04651_, _04608_);
  nand (_04652_, _03256_, _02929_);
  nor (_04653_, _02837_, _03665_);
  not (_04654_, _04653_);
  or (_04655_, _04654_, _04652_);
  nor (_04656_, _04655_, _04651_);
  and (_04657_, _04656_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04658_, _03256_, _02794_);
  nand (_04659_, _04658_, _04615_);
  nor (_04660_, _04659_, _04651_);
  and (_04661_, _04660_, \oc8051_golden_model_1.TH1 [7]);
  nor (_04662_, _04661_, _04657_);
  and (_04663_, _04616_, _02929_);
  and (_04664_, _04663_, _04608_);
  and (_04665_, _04664_, \oc8051_golden_model_1.TMOD [7]);
  and (_04666_, _04633_, _04621_);
  and (_04667_, _04666_, \oc8051_golden_model_1.SCON [7]);
  nor (_04668_, _04667_, _04665_);
  and (_04669_, _04668_, _04662_);
  and (_04670_, _04653_, _03256_);
  and (_04671_, _04670_, _04609_);
  and (_04672_, _04671_, \oc8051_golden_model_1.DPH [7]);
  not (_04673_, _04672_);
  not (_04674_, _04610_);
  or (_04675_, _04652_, _04674_);
  nor (_04676_, _04675_, _04651_);
  and (_04677_, _04676_, \oc8051_golden_model_1.TL0 [7]);
  nand (_04678_, _04658_, _04619_);
  nor (_04679_, _04678_, _04651_);
  and (_04680_, _04679_, \oc8051_golden_model_1.TH0 [7]);
  nor (_04681_, _04680_, _04677_);
  and (_04682_, _04681_, _04673_);
  and (_04683_, _04682_, _04669_);
  and (_04684_, _04653_, _04361_);
  and (_04685_, _04684_, _04609_);
  and (_04686_, _04685_, \oc8051_golden_model_1.PCON [7]);
  not (_04687_, _04686_);
  nor (_04688_, _02927_, _04551_);
  and (_04689_, _04688_, _04632_);
  and (_04690_, _04689_, _04627_);
  and (_04691_, _04690_, \oc8051_golden_model_1.PSW [7]);
  not (_04692_, _04691_);
  and (_04693_, _04644_, _04621_);
  and (_04694_, _04693_, \oc8051_golden_model_1.IP [7]);
  and (_04695_, _04688_, _04643_);
  and (_04696_, _04695_, _04627_);
  and (_04697_, _04696_, \oc8051_golden_model_1.B [7]);
  nor (_04698_, _04697_, _04694_);
  and (_04699_, _04698_, _04692_);
  and (_04700_, _04663_, _04633_);
  and (_04701_, _04700_, \oc8051_golden_model_1.SBUF [7]);
  not (_04702_, _04701_);
  and (_04703_, _04640_, _04621_);
  and (_04704_, _04703_, \oc8051_golden_model_1.IE [7]);
  and (_04705_, _04688_, _04639_);
  and (_04706_, _04705_, _04627_);
  and (_04707_, _04706_, \oc8051_golden_model_1.ACC [7]);
  nor (_04708_, _04707_, _04704_);
  and (_04709_, _04708_, _04702_);
  and (_04710_, _04709_, _04699_);
  and (_04711_, _04710_, _04687_);
  and (_04712_, _04711_, _04683_);
  and (_04713_, _04712_, _04650_);
  and (_04714_, _04713_, _04605_);
  not (_04715_, _04714_);
  not (_04716_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_04717_, _03597_, _04716_);
  not (_04718_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_04719_, _03751_, _04718_);
  and (_04720_, _04719_, _03749_);
  nand (_04721_, _04720_, _04717_);
  not (_04722_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_04723_, _03751_, _04722_);
  not (_04724_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_04725_, _03597_, _04724_);
  and (_04726_, _04725_, _03757_);
  nand (_04727_, _04726_, _04723_);
  nand (_04728_, _04727_, _04721_);
  nand (_04729_, _04728_, _03352_);
  not (_04730_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_04731_, _03751_, _04730_);
  not (_04732_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_04733_, _03597_, _04732_);
  and (_04734_, _04733_, _03757_);
  nand (_04735_, _04734_, _04731_);
  not (_04736_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04737_, _03597_, _04736_);
  not (_04739_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_04740_, _03751_, _04739_);
  and (_04741_, _04740_, _03749_);
  nand (_04742_, _04741_, _04737_);
  nand (_04743_, _04742_, _04735_);
  nand (_04744_, _04743_, _03764_);
  nand (_04745_, _04744_, _04729_);
  nand (_04746_, _04745_, _03177_);
  nand (_04747_, _03597_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04748_, _03751_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04749_, _04748_, _03757_);
  nand (_04750_, _04749_, _04747_);
  nand (_04751_, _03751_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04752_, _03597_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04753_, _04752_, _03749_);
  nand (_04754_, _04753_, _04751_);
  nand (_04755_, _04754_, _04750_);
  nand (_04756_, _04755_, _03352_);
  nand (_04757_, _03597_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04758_, _03751_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04759_, _04758_, _03757_);
  nand (_04760_, _04759_, _04757_);
  nand (_04761_, _03751_, \oc8051_golden_model_1.IRAM[12] [6]);
  not (_04762_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_04763_, _03751_, _04762_);
  and (_04764_, _04763_, _03749_);
  nand (_04765_, _04764_, _04761_);
  nand (_04766_, _04765_, _04760_);
  nand (_04767_, _04766_, _03764_);
  nand (_04768_, _04767_, _04756_);
  nand (_04769_, _04768_, _03781_);
  and (_04770_, _04769_, _04746_);
  nand (_04771_, _04770_, _04551_);
  and (_04772_, _04693_, \oc8051_golden_model_1.IP [6]);
  not (_04773_, _04772_);
  and (_04774_, _04690_, \oc8051_golden_model_1.PSW [6]);
  not (_04775_, _04774_);
  and (_04776_, _04706_, \oc8051_golden_model_1.ACC [6]);
  and (_04777_, _04696_, \oc8051_golden_model_1.B [6]);
  nor (_04778_, _04777_, _04776_);
  and (_04779_, _04778_, _04775_);
  and (_04780_, _04779_, _04773_);
  and (_04781_, _04628_, \oc8051_golden_model_1.P0 [6]);
  and (_04782_, _04653_, _04626_);
  and (_04783_, _04782_, _04608_);
  and (_04784_, _04783_, \oc8051_golden_model_1.DPH [6]);
  nor (_04785_, _04784_, _04781_);
  and (_04786_, _04641_, \oc8051_golden_model_1.P2 [6]);
  and (_04787_, _04645_, \oc8051_golden_model_1.P3 [6]);
  nor (_04788_, _04787_, _04786_);
  and (_04789_, _04685_, \oc8051_golden_model_1.PCON [6]);
  not (_04790_, _04789_);
  and (_04791_, _04700_, \oc8051_golden_model_1.SBUF [6]);
  and (_04792_, _04703_, \oc8051_golden_model_1.IE [6]);
  nor (_04793_, _04792_, _04791_);
  and (_04794_, _04793_, _04790_);
  and (_04795_, _04794_, _04788_);
  and (_04796_, _04622_, \oc8051_golden_model_1.TCON [6]);
  and (_04797_, _04679_, \oc8051_golden_model_1.TH0 [6]);
  nor (_04798_, _04797_, _04796_);
  and (_04799_, _04634_, \oc8051_golden_model_1.P1 [6]);
  and (_04800_, _04656_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04798_);
  and (_04803_, _04660_, \oc8051_golden_model_1.TH1 [6]);
  and (_04804_, _04666_, \oc8051_golden_model_1.SCON [6]);
  nor (_04805_, _04804_, _04803_);
  and (_04806_, _04664_, \oc8051_golden_model_1.TMOD [6]);
  and (_04807_, _04676_, \oc8051_golden_model_1.TL0 [6]);
  nor (_04808_, _04807_, _04806_);
  and (_04809_, _04808_, _04805_);
  and (_04810_, _04809_, _04802_);
  and (_04811_, _04612_, \oc8051_golden_model_1.DPL [6]);
  and (_04812_, _04617_, \oc8051_golden_model_1.SP [6]);
  nor (_04813_, _04812_, _04811_);
  and (_04814_, _04813_, _04810_);
  and (_04815_, _04814_, _04795_);
  and (_04816_, _04815_, _04785_);
  and (_04817_, _04816_, _04780_);
  and (_04818_, _04817_, _04771_);
  not (_04819_, _04818_);
  not (_04820_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_04821_, _03597_, _04820_);
  not (_04822_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_04823_, _03751_, _04822_);
  and (_04824_, _04823_, _03749_);
  nand (_04825_, _04824_, _04821_);
  not (_04826_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_04827_, _03751_, _04826_);
  not (_04828_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_04829_, _03597_, _04828_);
  and (_04830_, _04829_, _03757_);
  nand (_04831_, _04830_, _04827_);
  nand (_04832_, _04831_, _04825_);
  nand (_04833_, _04832_, _03352_);
  not (_04834_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_04835_, _03751_, _04834_);
  not (_04836_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_04837_, _03597_, _04836_);
  and (_04838_, _04837_, _03757_);
  nand (_04840_, _04838_, _04835_);
  not (_04841_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_04842_, _03597_, _04841_);
  not (_04843_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_04844_, _03751_, _04843_);
  and (_04845_, _04844_, _03749_);
  nand (_04846_, _04845_, _04842_);
  nand (_04847_, _04846_, _04840_);
  nand (_04848_, _04847_, _03764_);
  nand (_04849_, _04848_, _04833_);
  nand (_04850_, _04849_, _03177_);
  nand (_04851_, _03597_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_04852_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_04853_, _03597_, _04852_);
  and (_04854_, _04853_, _03757_);
  nand (_04855_, _04854_, _04851_);
  nand (_04856_, _03751_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_04857_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_04858_, _03751_, _04857_);
  and (_04859_, _04858_, _03749_);
  nand (_04860_, _04859_, _04856_);
  nand (_04861_, _04860_, _04855_);
  nand (_04862_, _04861_, _03352_);
  nand (_04863_, _03597_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_04864_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_04865_, _03597_, _04864_);
  and (_04866_, _04865_, _03757_);
  nand (_04867_, _04866_, _04863_);
  nand (_04868_, _03751_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_04869_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_04870_, _03751_, _04869_);
  and (_04871_, _04870_, _03749_);
  nand (_04872_, _04871_, _04868_);
  nand (_04873_, _04872_, _04867_);
  nand (_04874_, _04873_, _03764_);
  nand (_04875_, _04874_, _04862_);
  nand (_04876_, _04875_, _03781_);
  and (_04877_, _04876_, _04850_);
  nand (_04878_, _04877_, _04551_);
  and (_04879_, _04700_, \oc8051_golden_model_1.SBUF [5]);
  and (_04880_, _04703_, \oc8051_golden_model_1.IE [5]);
  nor (_04881_, _04880_, _04879_);
  and (_04882_, _04645_, \oc8051_golden_model_1.P3 [5]);
  not (_04883_, _04882_);
  and (_04884_, _04641_, \oc8051_golden_model_1.P2 [5]);
  and (_04885_, _04685_, \oc8051_golden_model_1.PCON [5]);
  nor (_04886_, _04885_, _04884_);
  and (_04887_, _04886_, _04883_);
  and (_04888_, _04887_, _04881_);
  and (_04889_, _04690_, \oc8051_golden_model_1.PSW [5]);
  and (_04890_, _04706_, \oc8051_golden_model_1.ACC [5]);
  nor (_04891_, _04890_, _04889_);
  and (_04892_, _04693_, \oc8051_golden_model_1.IP [5]);
  and (_04893_, _04696_, \oc8051_golden_model_1.B [5]);
  nor (_04894_, _04893_, _04892_);
  and (_04895_, _04894_, _04891_);
  and (_04896_, _04622_, \oc8051_golden_model_1.TCON [5]);
  and (_04897_, _04679_, \oc8051_golden_model_1.TH0 [5]);
  nor (_04898_, _04897_, _04896_);
  and (_04899_, _04634_, \oc8051_golden_model_1.P1 [5]);
  and (_04900_, _04656_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04901_, _04900_, _04899_);
  and (_04902_, _04901_, _04898_);
  and (_04903_, _04660_, \oc8051_golden_model_1.TH1 [5]);
  and (_04904_, _04666_, \oc8051_golden_model_1.SCON [5]);
  nor (_04905_, _04904_, _04903_);
  and (_04906_, _04676_, \oc8051_golden_model_1.TL0 [5]);
  and (_04907_, _04664_, \oc8051_golden_model_1.TMOD [5]);
  nor (_04908_, _04907_, _04906_);
  and (_04909_, _04908_, _04905_);
  and (_04910_, _04909_, _04902_);
  and (_04911_, _04910_, _04895_);
  and (_04912_, _04911_, _04888_);
  and (_04913_, _04628_, \oc8051_golden_model_1.P0 [5]);
  not (_04914_, _04913_);
  and (_04915_, _04783_, \oc8051_golden_model_1.DPH [5]);
  not (_04916_, _04915_);
  and (_04917_, _04612_, \oc8051_golden_model_1.DPL [5]);
  and (_04918_, _04617_, \oc8051_golden_model_1.SP [5]);
  nor (_04919_, _04918_, _04917_);
  and (_04920_, _04919_, _04916_);
  and (_04921_, _04920_, _04914_);
  and (_04922_, _04921_, _04912_);
  and (_04923_, _04922_, _04878_);
  not (_04924_, _04923_);
  not (_04925_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_04926_, _03597_, _04925_);
  not (_04927_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_04928_, _03751_, _04927_);
  and (_04929_, _04928_, _03749_);
  nand (_04930_, _04929_, _04926_);
  not (_04931_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_04932_, _03751_, _04931_);
  not (_04933_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_04934_, _03597_, _04933_);
  and (_04935_, _04934_, _03757_);
  nand (_04936_, _04935_, _04932_);
  nand (_04937_, _04936_, _04930_);
  nand (_04938_, _04937_, _03352_);
  not (_04939_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_04941_, _03751_, _04939_);
  not (_04942_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_04943_, _03597_, _04942_);
  and (_04944_, _04943_, _03757_);
  nand (_04945_, _04944_, _04941_);
  not (_04946_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_04947_, _03597_, _04946_);
  not (_04948_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_04949_, _03751_, _04948_);
  and (_04950_, _04949_, _03749_);
  nand (_04951_, _04950_, _04947_);
  nand (_04952_, _04951_, _04945_);
  nand (_04953_, _04952_, _03764_);
  nand (_04954_, _04953_, _04938_);
  nand (_04955_, _04954_, _03177_);
  nand (_04956_, _03597_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_04957_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_04958_, _03597_, _04957_);
  and (_04959_, _04958_, _03757_);
  nand (_04960_, _04959_, _04956_);
  nand (_04961_, _03751_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_04962_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_04963_, _03751_, _04962_);
  and (_04964_, _04963_, _03749_);
  nand (_04965_, _04964_, _04961_);
  nand (_04966_, _04965_, _04960_);
  nand (_04967_, _04966_, _03352_);
  nand (_04968_, _03597_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_04969_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_04970_, _03597_, _04969_);
  and (_04971_, _04970_, _03757_);
  nand (_04972_, _04971_, _04968_);
  nand (_04973_, _03751_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_04974_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_04975_, _03751_, _04974_);
  and (_04976_, _04975_, _03749_);
  nand (_04977_, _04976_, _04973_);
  nand (_04978_, _04977_, _04972_);
  nand (_04979_, _04978_, _03764_);
  nand (_04980_, _04979_, _04967_);
  nand (_04981_, _04980_, _03781_);
  and (_04982_, _04981_, _04955_);
  nand (_04983_, _04982_, _04551_);
  and (_04984_, _04671_, \oc8051_golden_model_1.DPH [4]);
  not (_04985_, _04984_);
  and (_04986_, _04679_, \oc8051_golden_model_1.TH0 [4]);
  and (_04987_, _04656_, \oc8051_golden_model_1.TL1 [4]);
  nor (_04988_, _04987_, _04986_);
  and (_04989_, _04988_, _04985_);
  and (_04990_, _04617_, \oc8051_golden_model_1.SP [4]);
  and (_04991_, _04612_, \oc8051_golden_model_1.DPL [4]);
  nor (_04992_, _04991_, _04990_);
  and (_04993_, _04685_, \oc8051_golden_model_1.PCON [4]);
  not (_04994_, _04993_);
  and (_04995_, _04700_, \oc8051_golden_model_1.SBUF [4]);
  and (_04996_, _04703_, \oc8051_golden_model_1.IE [4]);
  nor (_04997_, _04996_, _04995_);
  and (_04998_, _04997_, _04994_);
  and (_04999_, _04998_, _04992_);
  and (_05000_, _04999_, _04989_);
  and (_05001_, _04664_, \oc8051_golden_model_1.TMOD [4]);
  and (_05002_, _04666_, \oc8051_golden_model_1.SCON [4]);
  nor (_05003_, _05002_, _05001_);
  and (_05004_, _04676_, \oc8051_golden_model_1.TL0 [4]);
  not (_05005_, _05004_);
  and (_05006_, _04622_, \oc8051_golden_model_1.TCON [4]);
  and (_05007_, _04660_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05008_, _05007_, _05006_);
  and (_05009_, _05008_, _05005_);
  and (_05010_, _05009_, _05003_);
  and (_05011_, _04690_, \oc8051_golden_model_1.PSW [4]);
  and (_05012_, _04696_, \oc8051_golden_model_1.B [4]);
  nor (_05013_, _05012_, _05011_);
  and (_05014_, _04693_, \oc8051_golden_model_1.IP [4]);
  and (_05015_, _04706_, \oc8051_golden_model_1.ACC [4]);
  nor (_05016_, _05015_, _05014_);
  and (_05017_, _05016_, _05013_);
  and (_05018_, _04628_, \oc8051_golden_model_1.P0 [4]);
  not (_05019_, _05018_);
  and (_05020_, _04634_, \oc8051_golden_model_1.P1 [4]);
  not (_05021_, _05020_);
  and (_05022_, _04641_, \oc8051_golden_model_1.P2 [4]);
  and (_05023_, _04645_, \oc8051_golden_model_1.P3 [4]);
  nor (_05024_, _05023_, _05022_);
  and (_05025_, _05024_, _05021_);
  and (_05026_, _05025_, _05019_);
  and (_05027_, _05026_, _05017_);
  and (_05028_, _05027_, _05010_);
  and (_05029_, _05028_, _05000_);
  and (_05030_, _05029_, _04983_);
  not (_05031_, _05030_);
  nand (_05032_, _04241_, _04551_);
  and (_05033_, _04685_, \oc8051_golden_model_1.PCON [3]);
  not (_05034_, _05033_);
  and (_05035_, _04700_, \oc8051_golden_model_1.SBUF [3]);
  and (_05036_, _04703_, \oc8051_golden_model_1.IE [3]);
  nor (_05037_, _05036_, _05035_);
  and (_05038_, _05037_, _05034_);
  and (_05039_, _04641_, \oc8051_golden_model_1.P2 [3]);
  and (_05040_, _04645_, \oc8051_golden_model_1.P3 [3]);
  nor (_05042_, _05040_, _05039_);
  and (_05043_, _05042_, _05038_);
  and (_05044_, _04693_, \oc8051_golden_model_1.IP [3]);
  and (_05045_, _04706_, \oc8051_golden_model_1.ACC [3]);
  nor (_05046_, _05045_, _05044_);
  and (_05047_, _04690_, \oc8051_golden_model_1.PSW [3]);
  and (_05048_, _04696_, \oc8051_golden_model_1.B [3]);
  nor (_05049_, _05048_, _05047_);
  and (_05050_, _05049_, _05046_);
  and (_05051_, _04622_, \oc8051_golden_model_1.TCON [3]);
  and (_05052_, _04679_, \oc8051_golden_model_1.TH0 [3]);
  nor (_05053_, _05052_, _05051_);
  and (_05054_, _04634_, \oc8051_golden_model_1.P1 [3]);
  and (_05055_, _04656_, \oc8051_golden_model_1.TL1 [3]);
  nor (_05056_, _05055_, _05054_);
  and (_05057_, _05056_, _05053_);
  and (_05058_, _04666_, \oc8051_golden_model_1.SCON [3]);
  and (_05059_, _04660_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05060_, _05059_, _05058_);
  and (_05061_, _04664_, \oc8051_golden_model_1.TMOD [3]);
  and (_05062_, _04676_, \oc8051_golden_model_1.TL0 [3]);
  nor (_05063_, _05062_, _05061_);
  and (_05064_, _05063_, _05060_);
  and (_05065_, _05064_, _05057_);
  and (_05066_, _05065_, _05050_);
  and (_05067_, _05066_, _05043_);
  and (_05068_, _04628_, \oc8051_golden_model_1.P0 [3]);
  not (_05069_, _05068_);
  and (_05070_, _04617_, \oc8051_golden_model_1.SP [3]);
  and (_05071_, _04612_, \oc8051_golden_model_1.DPL [3]);
  nor (_05072_, _05071_, _05070_);
  and (_05073_, _04783_, \oc8051_golden_model_1.DPH [3]);
  not (_05074_, _05073_);
  and (_05075_, _05074_, _05072_);
  and (_05076_, _05075_, _05069_);
  and (_05077_, _05076_, _05067_);
  and (_05078_, _05077_, _05032_);
  not (_05079_, _05078_);
  nand (_05080_, _04435_, _04551_);
  and (_05081_, _04612_, \oc8051_golden_model_1.DPL [2]);
  not (_05082_, _05081_);
  and (_05083_, _04617_, \oc8051_golden_model_1.SP [2]);
  and (_05084_, _04622_, \oc8051_golden_model_1.TCON [2]);
  nor (_05085_, _05084_, _05083_);
  and (_05086_, _05085_, _05082_);
  and (_05087_, _04628_, \oc8051_golden_model_1.P0 [2]);
  not (_05088_, _05087_);
  and (_05089_, _04634_, \oc8051_golden_model_1.P1 [2]);
  not (_05090_, _05089_);
  and (_05091_, _04641_, \oc8051_golden_model_1.P2 [2]);
  and (_05092_, _04645_, \oc8051_golden_model_1.P3 [2]);
  nor (_05093_, _05092_, _05091_);
  and (_05094_, _05093_, _05090_);
  and (_05095_, _05094_, _05088_);
  and (_05096_, _05095_, _05086_);
  and (_05097_, _04656_, \oc8051_golden_model_1.TL1 [2]);
  and (_05098_, _04660_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05099_, _05098_, _05097_);
  and (_05100_, _04664_, \oc8051_golden_model_1.TMOD [2]);
  and (_05101_, _04666_, \oc8051_golden_model_1.SCON [2]);
  nor (_05102_, _05101_, _05100_);
  and (_05103_, _05102_, _05099_);
  and (_05104_, _04671_, \oc8051_golden_model_1.DPH [2]);
  not (_05105_, _05104_);
  and (_05106_, _04676_, \oc8051_golden_model_1.TL0 [2]);
  and (_05107_, _04679_, \oc8051_golden_model_1.TH0 [2]);
  nor (_05108_, _05107_, _05106_);
  and (_05109_, _05108_, _05105_);
  and (_05110_, _05109_, _05103_);
  and (_05111_, _04685_, \oc8051_golden_model_1.PCON [2]);
  not (_05112_, _05111_);
  and (_05113_, _04690_, \oc8051_golden_model_1.PSW [2]);
  not (_05114_, _05113_);
  and (_05115_, _04693_, \oc8051_golden_model_1.IP [2]);
  and (_05116_, _04696_, \oc8051_golden_model_1.B [2]);
  nor (_05117_, _05116_, _05115_);
  and (_05118_, _05117_, _05114_);
  and (_05119_, _04700_, \oc8051_golden_model_1.SBUF [2]);
  not (_05120_, _05119_);
  and (_05121_, _04703_, \oc8051_golden_model_1.IE [2]);
  and (_05122_, _04706_, \oc8051_golden_model_1.ACC [2]);
  nor (_05123_, _05122_, _05121_);
  and (_05124_, _05123_, _05120_);
  and (_05125_, _05124_, _05118_);
  and (_05126_, _05125_, _05112_);
  and (_05127_, _05126_, _05110_);
  and (_05128_, _05127_, _05096_);
  and (_05129_, _05128_, _05080_);
  not (_05130_, _05129_);
  nand (_05131_, _04000_, _04551_);
  and (_05132_, _04671_, \oc8051_golden_model_1.DPH [1]);
  not (_05133_, _05132_);
  and (_05134_, _04679_, \oc8051_golden_model_1.TH0 [1]);
  and (_05135_, _04656_, \oc8051_golden_model_1.TL1 [1]);
  nor (_05136_, _05135_, _05134_);
  and (_05137_, _05136_, _05133_);
  and (_05138_, _04617_, \oc8051_golden_model_1.SP [1]);
  and (_05139_, _04612_, \oc8051_golden_model_1.DPL [1]);
  nor (_05140_, _05139_, _05138_);
  and (_05141_, _04685_, \oc8051_golden_model_1.PCON [1]);
  not (_05142_, _05141_);
  and (_05143_, _04700_, \oc8051_golden_model_1.SBUF [1]);
  and (_05144_, _04703_, \oc8051_golden_model_1.IE [1]);
  nor (_05145_, _05144_, _05143_);
  and (_05146_, _05145_, _05142_);
  and (_05147_, _05146_, _05140_);
  and (_05148_, _05147_, _05137_);
  and (_05149_, _04664_, \oc8051_golden_model_1.TMOD [1]);
  and (_05150_, _04666_, \oc8051_golden_model_1.SCON [1]);
  nor (_05151_, _05150_, _05149_);
  and (_05152_, _04676_, \oc8051_golden_model_1.TL0 [1]);
  not (_05153_, _05152_);
  and (_05154_, _04622_, \oc8051_golden_model_1.TCON [1]);
  and (_05155_, _04660_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05156_, _05155_, _05154_);
  and (_05157_, _05156_, _05153_);
  and (_05158_, _05157_, _05151_);
  and (_05159_, _04628_, \oc8051_golden_model_1.P0 [1]);
  not (_05160_, _05159_);
  and (_05161_, _04690_, \oc8051_golden_model_1.PSW [1]);
  and (_05162_, _04706_, \oc8051_golden_model_1.ACC [1]);
  nor (_05163_, _05162_, _05161_);
  and (_05164_, _04693_, \oc8051_golden_model_1.IP [1]);
  and (_05165_, _04696_, \oc8051_golden_model_1.B [1]);
  nor (_05166_, _05165_, _05164_);
  and (_05167_, _05166_, _05163_);
  and (_05168_, _04634_, \oc8051_golden_model_1.P1 [1]);
  not (_05169_, _05168_);
  and (_05170_, _04641_, \oc8051_golden_model_1.P2 [1]);
  and (_05171_, _04645_, \oc8051_golden_model_1.P3 [1]);
  nor (_05172_, _05171_, _05170_);
  and (_05173_, _05172_, _05169_);
  and (_05174_, _05173_, _05167_);
  and (_05175_, _05174_, _05160_);
  and (_05176_, _05175_, _05158_);
  and (_05177_, _05176_, _05148_);
  and (_05178_, _05177_, _05131_);
  nand (_05179_, _03808_, _04551_);
  and (_05180_, _04671_, \oc8051_golden_model_1.DPH [0]);
  not (_05181_, _05180_);
  and (_05182_, _04679_, \oc8051_golden_model_1.TH0 [0]);
  and (_05183_, _04656_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05184_, _05183_, _05182_);
  and (_05185_, _05184_, _05181_);
  and (_05186_, _04617_, \oc8051_golden_model_1.SP [0]);
  and (_05187_, _04612_, \oc8051_golden_model_1.DPL [0]);
  nor (_05188_, _05187_, _05186_);
  and (_05189_, _04685_, \oc8051_golden_model_1.PCON [0]);
  not (_05190_, _05189_);
  and (_05191_, _04700_, \oc8051_golden_model_1.SBUF [0]);
  and (_05192_, _04703_, \oc8051_golden_model_1.IE [0]);
  nor (_05193_, _05192_, _05191_);
  and (_05194_, _05193_, _05190_);
  and (_05195_, _05194_, _05188_);
  and (_05196_, _05195_, _05185_);
  and (_05197_, _04676_, \oc8051_golden_model_1.TL0 [0]);
  and (_05198_, _04666_, \oc8051_golden_model_1.SCON [0]);
  nor (_05199_, _05198_, _05197_);
  and (_05200_, _04660_, \oc8051_golden_model_1.TH1 [0]);
  not (_05201_, _05200_);
  and (_05202_, _04622_, \oc8051_golden_model_1.TCON [0]);
  and (_05203_, _04664_, \oc8051_golden_model_1.TMOD [0]);
  nor (_05204_, _05203_, _05202_);
  and (_05205_, _05204_, _05201_);
  and (_05206_, _05205_, _05199_);
  and (_05207_, _04628_, \oc8051_golden_model_1.P0 [0]);
  not (_05208_, _05207_);
  and (_05209_, _04693_, \oc8051_golden_model_1.IP [0]);
  and (_05210_, _04706_, \oc8051_golden_model_1.ACC [0]);
  nor (_05211_, _05210_, _05209_);
  and (_05212_, _04690_, \oc8051_golden_model_1.PSW [0]);
  and (_05213_, _04696_, \oc8051_golden_model_1.B [0]);
  nor (_05214_, _05213_, _05212_);
  and (_05215_, _05214_, _05211_);
  and (_05216_, _04634_, \oc8051_golden_model_1.P1 [0]);
  not (_05217_, _05216_);
  and (_05218_, _04641_, \oc8051_golden_model_1.P2 [0]);
  and (_05219_, _04645_, \oc8051_golden_model_1.P3 [0]);
  nor (_05220_, _05219_, _05218_);
  and (_05221_, _05220_, _05217_);
  and (_05222_, _05221_, _05215_);
  and (_05223_, _05222_, _05208_);
  and (_05224_, _05223_, _05206_);
  and (_05225_, _05224_, _05196_);
  and (_05226_, _05225_, _05179_);
  nor (_05227_, _05226_, _05178_);
  and (_05228_, _05227_, _05130_);
  and (_05229_, _05228_, _05079_);
  and (_05230_, _05229_, _05031_);
  and (_05231_, _05230_, _04924_);
  and (_05232_, _05231_, _04819_);
  nor (_05233_, _05232_, _04715_);
  and (_05234_, _05232_, _04715_);
  nor (_05235_, _05234_, _05233_);
  and (_05236_, _05235_, _03923_);
  nand (_05237_, _02522_, _02429_);
  not (_05238_, _04119_);
  and (_05239_, _03808_, _04000_);
  and (_05240_, _04241_, _04435_);
  and (_05241_, _05240_, _05239_);
  and (_05242_, _05241_, _04982_);
  and (_05243_, _05242_, _04877_);
  nor (_05244_, _04770_, _04604_);
  and (_05245_, _04770_, _04604_);
  nor (_05246_, _05245_, _05244_);
  and (_05247_, _05246_, _05243_);
  not (_05248_, _04604_);
  nor (_05249_, _05248_, _05243_);
  or (_05250_, _05249_, _05247_);
  and (_05251_, _05250_, _05238_);
  or (_05252_, _05251_, _05237_);
  and (_05253_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05254_, _05253_, \oc8051_golden_model_1.PC [6]);
  and (_05255_, _02248_, _02229_);
  and (_05256_, _05255_, _05254_);
  and (_05257_, _05256_, \oc8051_golden_model_1.PC [7]);
  nor (_05258_, _05256_, \oc8051_golden_model_1.PC [7]);
  nor (_05259_, _05258_, _05257_);
  not (_05260_, _05259_);
  nand (_05261_, _05260_, _02939_);
  not (_05262_, _04153_);
  and (_05263_, _02846_, _02367_);
  or (_05264_, _05263_, _03317_);
  not (_05265_, _05264_);
  and (_05266_, _02840_, _02367_);
  nor (_05267_, _03718_, _05266_);
  and (_05268_, _05267_, _05265_);
  not (_05269_, _04770_);
  nor (_05270_, _04982_, _04877_);
  nor (_05271_, _03808_, _04000_);
  nor (_05272_, _04241_, _04435_);
  and (_05273_, _05272_, _05271_);
  and (_05274_, _05273_, _05270_);
  and (_05275_, _05274_, _05269_);
  or (_05276_, _05275_, _04604_);
  nand (_05277_, _05275_, _04604_);
  and (_05278_, _05277_, _05276_);
  or (_05279_, _05278_, _05268_);
  and (_05280_, _05279_, _05262_);
  and (_05281_, _03012_, _41915_);
  and (_05282_, _03049_, _01136_);
  nor (_05283_, _05282_, _05281_);
  and (_05284_, _03021_, _01157_);
  and (_05285_, _03046_, _01083_);
  nor (_05286_, _05285_, _05284_);
  and (_05287_, _05286_, _05283_);
  and (_05288_, _03015_, _01142_);
  and (_05289_, _03038_, _01132_);
  nor (_05290_, _05289_, _05288_);
  and (_05291_, _03002_, _01125_);
  and (_05292_, _03033_, _01166_);
  nor (_05293_, _05292_, _05291_);
  and (_05294_, _05293_, _05290_);
  and (_05295_, _05294_, _05287_);
  and (_05296_, _03019_, _01154_);
  and (_05297_, _03044_, _01161_);
  nor (_05298_, _05297_, _05296_);
  and (_05299_, _03026_, _01115_);
  and (_05300_, _03035_, _01149_);
  nor (_05301_, _05300_, _05299_);
  and (_05302_, _05301_, _05298_);
  and (_05303_, _03024_, _01111_);
  and (_05304_, _03040_, _01129_);
  nor (_05305_, _05304_, _05303_);
  and (_05306_, _03005_, _01121_);
  and (_05307_, _03052_, _01169_);
  nor (_05308_, _05307_, _05306_);
  and (_05309_, _05308_, _05305_);
  and (_05310_, _05309_, _05302_);
  and (_05311_, _05310_, _05295_);
  nor (_05312_, _05311_, _04714_);
  and (_05313_, _05312_, _03884_);
  nand (_05314_, _05311_, _02804_);
  not (_05315_, _03844_);
  not (_05316_, _02795_);
  nor (_05317_, _05316_, _03630_);
  nor (_05318_, _03212_, _02931_);
  and (_05319_, _05318_, _05317_);
  and (_05320_, _05319_, _04608_);
  and (_05321_, _05320_, \oc8051_golden_model_1.TCON [7]);
  not (_05322_, _03212_);
  and (_05323_, _05322_, _02931_);
  and (_05324_, _05323_, _05317_);
  and (_05325_, _04705_, _05324_);
  and (_05326_, _05325_, \oc8051_golden_model_1.ACC [7]);
  nor (_05327_, _05326_, _05321_);
  and (_05328_, _05319_, _04644_);
  and (_05329_, _05328_, \oc8051_golden_model_1.IP [7]);
  not (_05330_, _05329_);
  and (_05331_, _04689_, _05324_);
  and (_05332_, _05331_, \oc8051_golden_model_1.PSW [7]);
  and (_05333_, _04695_, _05324_);
  and (_05334_, _05333_, \oc8051_golden_model_1.B [7]);
  nor (_05335_, _05334_, _05332_);
  and (_05336_, _05335_, _05330_);
  and (_05337_, _05336_, _05327_);
  and (_05338_, _05319_, _04633_);
  and (_05339_, _05338_, \oc8051_golden_model_1.SCON [7]);
  and (_05340_, _05319_, _04640_);
  and (_05341_, _05340_, \oc8051_golden_model_1.IE [7]);
  nor (_05342_, _05341_, _05339_);
  and (_05343_, _04609_, \oc8051_golden_model_1.P0 [7]);
  and (_05344_, _04633_, _05324_);
  and (_05345_, _05344_, \oc8051_golden_model_1.P1 [7]);
  nor (_05346_, _05345_, _05343_);
  and (_05347_, _04640_, _05324_);
  and (_05348_, _05347_, \oc8051_golden_model_1.P2 [7]);
  and (_05349_, _04644_, _05324_);
  and (_05350_, _05349_, \oc8051_golden_model_1.P3 [7]);
  nor (_05351_, _05350_, _05348_);
  and (_05352_, _05351_, _05346_);
  and (_05353_, _05352_, _05342_);
  and (_05354_, _05353_, _05337_);
  and (_05355_, _05354_, _04605_);
  nor (_05356_, _05355_, _04684_);
  or (_05357_, _05356_, _05315_);
  not (_05358_, _02883_);
  not (_05359_, _04684_);
  nand (_05360_, _05355_, _05359_);
  or (_05361_, _05360_, _05358_);
  nor (_05362_, _04442_, _04143_);
  not (_05363_, _05362_);
  and (_05364_, _05363_, _05278_);
  and (_05365_, _05254_, _02626_);
  and (_05366_, _05365_, \oc8051_golden_model_1.PC [7]);
  nor (_05367_, _05365_, \oc8051_golden_model_1.PC [7]);
  nor (_05368_, _05367_, _05366_);
  not (_05369_, _05368_);
  nor (_05370_, _05369_, _02611_);
  and (_05371_, _02611_, \oc8051_golden_model_1.ACC [7]);
  or (_05372_, _05371_, _05370_);
  and (_05373_, _05372_, _05362_);
  or (_05374_, _05373_, _02886_);
  or (_05375_, _05374_, _05364_);
  nor (_05376_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05377_, _05376_, _03335_);
  nor (_05378_, _05377_, _03068_);
  nor (_05379_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05380_, _05379_, _03068_);
  and (_05381_, _05380_, _02866_);
  nor (_05382_, _05381_, _05378_);
  nor (_05383_, _05382_, _03337_);
  not (_05384_, _05383_);
  or (_05385_, _04241_, _03859_);
  not (_05386_, _03337_);
  and (_05387_, _03859_, _02794_);
  nor (_05388_, _05387_, _05386_);
  nand (_05389_, _05388_, _05385_);
  and (_05390_, _05389_, _05384_);
  not (_05391_, _05390_);
  nor (_05392_, _05376_, _03335_);
  nor (_05393_, _05392_, _05377_);
  nor (_05394_, _05393_, _03337_);
  not (_05395_, _05394_);
  or (_05396_, _04435_, _03859_);
  and (_05397_, _03859_, _03256_);
  nor (_05398_, _05397_, _05386_);
  nand (_05399_, _05398_, _05396_);
  and (_05400_, _05399_, _05395_);
  not (_05401_, _05400_);
  nor (_05402_, _03337_, _03934_);
  not (_05403_, _05402_);
  and (_05404_, _04000_, _03860_);
  nor (_05405_, _03860_, _03665_);
  or (_05406_, _05405_, _05386_);
  or (_05407_, _05406_, _05404_);
  nand (_05408_, _05407_, _05403_);
  or (_05409_, _03808_, _03859_);
  and (_05410_, _03859_, _02837_);
  nor (_05411_, _05410_, _05386_);
  nand (_05412_, _05411_, _05409_);
  nor (_05413_, _03337_, \oc8051_golden_model_1.SP [0]);
  not (_05414_, _05413_);
  and (_05415_, _05414_, _05412_);
  and (_05416_, _05415_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand (_05417_, _05414_, _05412_);
  and (_05418_, _05417_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05419_, _05418_, _05416_);
  and (_05420_, _05419_, _05408_);
  and (_05421_, _05407_, _05403_);
  and (_05422_, _05415_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_05423_, _05417_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05424_, _05423_, _05422_);
  and (_05425_, _05424_, _05421_);
  or (_05426_, _05425_, _05420_);
  nor (_05427_, _05426_, _05401_);
  and (_05428_, _05415_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_05429_, _05417_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05430_, _05429_, _05428_);
  and (_05431_, _05430_, _05408_);
  and (_05432_, _05415_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_05433_, _05417_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05434_, _05433_, _05432_);
  and (_05435_, _05434_, _05421_);
  or (_05436_, _05435_, _05431_);
  nor (_05437_, _05436_, _05400_);
  nor (_05438_, _05437_, _05427_);
  nor (_05439_, _05438_, _05391_);
  and (_05440_, _05415_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_05441_, _05417_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_05442_, _05441_, _05440_);
  and (_05443_, _05442_, _05408_);
  and (_05444_, _05415_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_05445_, _05417_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_05446_, _05445_, _05444_);
  and (_05447_, _05446_, _05421_);
  or (_05448_, _05447_, _05443_);
  nor (_05449_, _05448_, _05401_);
  and (_05450_, _05415_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_05451_, _05417_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05452_, _05451_, _05450_);
  and (_05453_, _05452_, _05408_);
  and (_05454_, _05415_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_05455_, _05417_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_05456_, _05455_, _05454_);
  and (_05457_, _05456_, _05421_);
  or (_05458_, _05457_, _05453_);
  nor (_05459_, _05458_, _05400_);
  nor (_05460_, _05459_, _05449_);
  nor (_05461_, _05460_, _05390_);
  nor (_05462_, _05461_, _05439_);
  or (_05463_, _05462_, _04265_);
  and (_05464_, _05463_, _05375_);
  or (_05465_, _05464_, _03811_);
  and (_05466_, _05030_, _04923_);
  and (_05467_, _05226_, _05178_);
  and (_05468_, _05129_, _05078_);
  and (_05469_, _05468_, _05467_);
  and (_05470_, _05469_, _05466_);
  and (_05471_, _05470_, _04818_);
  nor (_05472_, _05471_, _04715_);
  and (_05473_, _05471_, _04715_);
  nor (_05474_, _05473_, _05472_);
  or (_05475_, _05474_, _03812_);
  and (_05476_, _05475_, _05465_);
  or (_05477_, _05476_, _02883_);
  and (_05478_, _05477_, _05361_);
  or (_05479_, _05478_, _04252_);
  nor (_05480_, _05368_, _02609_);
  nor (_05481_, _05480_, _03836_);
  and (_05482_, _05481_, _05479_);
  and (_05483_, _04604_, _03836_);
  or (_05484_, _05483_, _03844_);
  or (_05485_, _05484_, _05482_);
  and (_05486_, _05485_, _05357_);
  or (_05487_, _05486_, _02875_);
  and (_05488_, _04641_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05489_, _04645_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05490_, _05489_, _05488_);
  and (_05491_, _04628_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05492_, _04634_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_05493_, _05492_, _05491_);
  and (_05494_, _05493_, _05490_);
  and (_05495_, _05494_, _04625_);
  and (_05496_, _05495_, _04712_);
  and (_05497_, _05496_, _04605_);
  nand (_05498_, _05497_, _02875_);
  and (_05499_, _05498_, _02873_);
  and (_05500_, _05499_, _05487_);
  nor (_05501_, _05355_, _05359_);
  not (_05502_, _05501_);
  and (_05503_, _05502_, _05360_);
  and (_05504_, _05503_, _02872_);
  or (_05505_, _05504_, _05500_);
  and (_05506_, _05505_, _02614_);
  nor (_05507_, _05369_, _02614_);
  or (_05508_, _05507_, _03059_);
  or (_05509_, _05508_, _05506_);
  nand (_05510_, _05497_, _03059_);
  and (_05511_, _05510_, _05509_);
  or (_05512_, _05511_, _03859_);
  and (_05513_, _05462_, _04551_);
  nand (_05514_, _05496_, _03859_);
  or (_05515_, _05514_, _05513_);
  and (_05516_, _05515_, _04298_);
  and (_05517_, _05516_, _05512_);
  and (_05518_, _04609_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05519_, _05347_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05520_, _05519_, _05518_);
  and (_05521_, _05344_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05522_, _05349_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05523_, _05522_, _05521_);
  and (_05524_, _05523_, _05520_);
  and (_05525_, _05524_, _05342_);
  and (_05526_, _05525_, _05337_);
  and (_05527_, _05526_, _04605_);
  nor (_05528_, _05527_, _04684_);
  and (_05529_, _04684_, \oc8051_golden_model_1.PSW [7]);
  nor (_05530_, _05529_, _05528_);
  nor (_05531_, _05530_, _04298_);
  or (_05532_, _05531_, _02581_);
  or (_05533_, _05532_, _05517_);
  not (_05534_, _02855_);
  and (_05535_, _02851_, _05534_);
  nor (_05536_, _05535_, _02763_);
  and (_05537_, _05369_, _02581_);
  nor (_05538_, _05537_, _05536_);
  and (_05539_, _05538_, _05533_);
  not (_05540_, _02853_);
  nor (_05541_, _05540_, _02763_);
  and (_05542_, _04604_, _05536_);
  or (_05543_, _05542_, _05541_);
  or (_05544_, _05543_, _05539_);
  not (_05545_, _04176_);
  not (_05546_, _05541_);
  or (_05547_, _05462_, _05546_);
  and (_05548_, _05547_, _05545_);
  and (_05549_, _05548_, _05544_);
  and (_05550_, _05311_, _04604_);
  not (_05551_, _05550_);
  and (_05552_, _03012_, _41950_);
  and (_05553_, _03052_, _01485_);
  nor (_05554_, _05553_, _05552_);
  and (_05555_, _03024_, _01472_);
  and (_05556_, _03033_, _01483_);
  nor (_05557_, _05556_, _05555_);
  and (_05558_, _05557_, _05554_);
  and (_05559_, _03046_, _01445_);
  and (_05560_, _03035_, _01447_);
  nor (_05561_, _05560_, _05559_);
  and (_05562_, _03038_, _01457_);
  and (_05563_, _03040_, _01468_);
  nor (_05564_, _05563_, _05562_);
  and (_05565_, _05564_, _05561_);
  and (_05566_, _05565_, _05558_);
  and (_05567_, _03005_, _01466_);
  and (_05568_, _03049_, _01455_);
  nor (_05569_, _05568_, _05567_);
  and (_05570_, _03021_, _01476_);
  and (_05571_, _03015_, _01461_);
  nor (_05572_, _05571_, _05570_);
  and (_05573_, _05572_, _05569_);
  and (_05574_, _03019_, _01474_);
  and (_05575_, _03026_, _01449_);
  nor (_05576_, _05575_, _05574_);
  and (_05577_, _03044_, _01478_);
  and (_05578_, _03002_, _01453_);
  nor (_05579_, _05578_, _05577_);
  and (_05580_, _05579_, _05576_);
  and (_05581_, _05580_, _05573_);
  and (_05582_, _05581_, _05566_);
  and (_05583_, _03019_, _01521_);
  and (_05584_, _03021_, _01519_);
  nor (_05585_, _05584_, _05583_);
  and (_05586_, _03005_, _01511_);
  and (_05587_, _03049_, _01502_);
  nor (_05588_, _05587_, _05586_);
  and (_05589_, _05588_, _05585_);
  and (_05590_, _03035_, _01517_);
  and (_05591_, _03052_, _01530_);
  nor (_05592_, _05591_, _05590_);
  and (_05593_, _03002_, _01498_);
  and (_05594_, _03040_, _01513_);
  nor (_05595_, _05594_, _05593_);
  and (_05596_, _05595_, _05592_);
  and (_05597_, _05596_, _05589_);
  and (_05598_, _03024_, _01492_);
  and (_05599_, _03046_, _01494_);
  nor (_05600_, _05599_, _05598_);
  and (_05601_, _03012_, _41957_);
  and (_05602_, _03044_, _01523_);
  nor (_05603_, _05602_, _05601_);
  and (_05604_, _05603_, _05600_);
  and (_05605_, _03038_, _01500_);
  and (_05606_, _03033_, _01528_);
  nor (_05607_, _05606_, _05605_);
  and (_05608_, _03015_, _01506_);
  and (_05609_, _03026_, _01490_);
  nor (_05610_, _05609_, _05608_);
  and (_05611_, _05610_, _05607_);
  and (_05612_, _05611_, _05604_);
  and (_05613_, _05612_, _05597_);
  not (_05614_, _05613_);
  and (_05615_, _05614_, _05582_);
  and (_05616_, _03698_, _03486_);
  and (_05617_, _03297_, _03057_);
  and (_05618_, _05617_, _05616_);
  and (_05619_, _03038_, _01550_);
  and (_05620_, _03033_, _01573_);
  nor (_05621_, _05620_, _05619_);
  and (_05622_, _03019_, _01566_);
  and (_05623_, _03049_, _01552_);
  nor (_05624_, _05623_, _05622_);
  and (_05625_, _05624_, _05621_);
  and (_05626_, _03021_, _01564_);
  and (_05627_, _03044_, _01568_);
  nor (_05628_, _05627_, _05626_);
  and (_05629_, _03005_, _01545_);
  and (_05630_, _03040_, _01548_);
  nor (_05631_, _05630_, _05629_);
  and (_05632_, _05631_, _05628_);
  and (_05633_, _05632_, _05625_);
  and (_05634_, _03035_, _01562_);
  and (_05635_, _03052_, _01575_);
  nor (_05636_, _05635_, _05634_);
  and (_05637_, _03024_, _01537_);
  and (_05638_, _03046_, _01539_);
  nor (_05639_, _05638_, _05637_);
  and (_05640_, _05639_, _05636_);
  and (_05641_, _03012_, _41964_);
  and (_05642_, _03002_, _01543_);
  nor (_05643_, _05642_, _05641_);
  and (_05644_, _03015_, _01556_);
  and (_05645_, _03026_, _01535_);
  nor (_05646_, _05645_, _05644_);
  and (_05647_, _05646_, _05643_);
  and (_05648_, _05647_, _05640_);
  and (_05649_, _05648_, _05633_);
  nor (_05650_, _05649_, _05311_);
  and (_05651_, _05650_, _05618_);
  and (_05652_, _05651_, _05615_);
  and (_05653_, _05652_, \oc8051_golden_model_1.ACC [7]);
  nor (_05654_, _05613_, _05582_);
  and (_05655_, _05654_, _05651_);
  and (_05656_, _05655_, \oc8051_golden_model_1.B [7]);
  nor (_05657_, _05656_, _05653_);
  not (_05658_, _03057_);
  and (_05659_, _03297_, _05658_);
  and (_05660_, _05659_, _05616_);
  not (_05661_, _05311_);
  and (_05662_, _05649_, _05661_);
  and (_05663_, _05662_, _05654_);
  and (_05664_, _05663_, _05660_);
  and (_05665_, _05664_, \oc8051_golden_model_1.IP [7]);
  not (_05666_, _05582_);
  and (_05667_, _05613_, _05666_);
  and (_05668_, _05667_, _05651_);
  and (_05669_, _05668_, \oc8051_golden_model_1.PSW [7]);
  nor (_05670_, _05669_, _05665_);
  and (_05671_, _05670_, _05657_);
  not (_05672_, _03486_);
  and (_05673_, _03698_, _05672_);
  and (_05674_, _05613_, _05582_);
  and (_05675_, _05674_, _05662_);
  nor (_05676_, _03297_, _03057_);
  and (_05677_, _05676_, _05675_);
  and (_05678_, _05677_, _05673_);
  and (_05679_, _05678_, \oc8051_golden_model_1.TH1 [7]);
  not (_05680_, _05679_);
  and (_05681_, _05675_, _05617_);
  and (_05682_, _05681_, _05673_);
  and (_05683_, _05682_, \oc8051_golden_model_1.SP [7]);
  not (_05684_, _03698_);
  and (_05685_, _05684_, _03486_);
  and (_05686_, _05675_, _05659_);
  and (_05687_, _05686_, _05685_);
  and (_05688_, _05687_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05689_, _05688_, _05683_);
  and (_05690_, _05689_, _05680_);
  and (_05691_, _05690_, _05671_);
  and (_05692_, _05677_, _05616_);
  and (_05693_, _05692_, \oc8051_golden_model_1.TH0 [7]);
  nor (_05694_, _03698_, _03486_);
  and (_05695_, _05694_, _05675_);
  and (_05696_, _05695_, _05659_);
  and (_05697_, _05696_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05698_, _05697_, _05693_);
  and (_05699_, _05675_, _05660_);
  and (_05700_, _05699_, \oc8051_golden_model_1.TCON [7]);
  not (_05701_, _03297_);
  and (_05702_, _05701_, _03057_);
  and (_05703_, _05695_, _05702_);
  and (_05704_, _05703_, \oc8051_golden_model_1.PCON [7]);
  nor (_05705_, _05704_, _05700_);
  and (_05706_, _05705_, _05698_);
  and (_05707_, _05685_, _05681_);
  and (_05708_, _05707_, \oc8051_golden_model_1.DPL [7]);
  not (_05709_, _05708_);
  and (_05710_, _05675_, _05618_);
  and (_05711_, _05710_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05712_, _05711_);
  and (_05713_, _05654_, _05618_);
  and (_05714_, _05662_, _05713_);
  nand (_05715_, _05714_, \oc8051_golden_model_1.P3INREG [7]);
  and (_05716_, _05667_, _05662_);
  and (_05717_, _05716_, _05618_);
  and (_05718_, _05717_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05719_, _05662_, _05615_);
  and (_05720_, _05719_, _05618_);
  and (_05721_, _05720_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05722_, _05721_, _05718_);
  and (_05723_, _05722_, _05715_);
  and (_05724_, _05723_, _05712_);
  and (_05725_, _05724_, _05709_);
  and (_05726_, _05719_, _05660_);
  and (_05727_, _05726_, \oc8051_golden_model_1.IE [7]);
  and (_05728_, _05673_, _05659_);
  and (_05729_, _05728_, _05716_);
  and (_05730_, _05729_, \oc8051_golden_model_1.SBUF [7]);
  and (_05731_, _05716_, _05660_);
  and (_05732_, _05731_, \oc8051_golden_model_1.SCON [7]);
  or (_05733_, _05732_, _05730_);
  nor (_05734_, _05733_, _05727_);
  and (_05735_, _05686_, _05673_);
  and (_05736_, _05735_, \oc8051_golden_model_1.TMOD [7]);
  and (_05737_, _05695_, _05617_);
  and (_05738_, _05737_, \oc8051_golden_model_1.DPH [7]);
  nor (_05739_, _05738_, _05736_);
  and (_05740_, _05739_, _05734_);
  and (_05741_, _05740_, _05725_);
  and (_05742_, _05741_, _05706_);
  and (_05743_, _05742_, _05691_);
  and (_05744_, _05743_, _05551_);
  nor (_05745_, _05744_, _05545_);
  not (_05746_, _02513_);
  and (_05747_, _02577_, _02544_);
  nor (_05748_, _03368_, _05747_);
  nor (_05749_, _05748_, _05746_);
  nor (_05750_, _05749_, _03493_);
  nor (_05751_, _04147_, _04102_);
  and (_05752_, _05751_, _04129_);
  and (_05753_, _05752_, _05750_);
  not (_05754_, _05753_);
  or (_05755_, _05754_, _05745_);
  or (_05756_, _05755_, _05549_);
  or (_05757_, _05753_, _02763_);
  and (_05758_, _05757_, _05756_);
  or (_05759_, _05758_, _02804_);
  and (_05760_, _05759_, _05314_);
  or (_05761_, _05760_, _02514_);
  and (_05762_, _05369_, _02514_);
  nor (_05763_, _05762_, _03888_);
  and (_05764_, _05763_, _05761_);
  and (_05765_, _05311_, _04714_);
  nor (_05766_, _05765_, _05312_);
  nor (_05767_, _05766_, _03886_);
  nor (_05768_, _05767_, _03889_);
  or (_05769_, _05768_, _05764_);
  not (_05770_, _03886_);
  not (_05771_, \oc8051_golden_model_1.ACC [7]);
  nor (_05772_, _04714_, _05771_);
  and (_05773_, _04714_, _05771_);
  nor (_05774_, _05773_, _05772_);
  or (_05775_, _05774_, _05770_);
  and (_05776_, _05775_, _03885_);
  and (_05777_, _05776_, _05769_);
  or (_05778_, _05777_, _05313_);
  and (_05779_, _05778_, _03882_);
  and (_05780_, _05772_, _03881_);
  or (_05781_, _05780_, _03880_);
  or (_05782_, _05781_, _05779_);
  not (_05783_, _02965_);
  nor (_05784_, _05783_, _02763_);
  nor (_05785_, _05368_, _02532_);
  nor (_05786_, _05785_, _05784_);
  and (_05787_, _05786_, _05782_);
  not (_05788_, _03123_);
  nor (_05789_, _05788_, _02763_);
  not (_05790_, _05784_);
  nor (_05791_, _05765_, _05790_);
  or (_05792_, _05791_, _05789_);
  or (_05793_, _05792_, _05787_);
  nand (_05794_, _05773_, _05789_);
  and (_05795_, _05794_, _02529_);
  and (_05796_, _05795_, _05793_);
  or (_05797_, _05369_, _02529_);
  nand (_05798_, _05797_, _05268_);
  or (_05799_, _05798_, _05796_);
  and (_05800_, _05799_, _05280_);
  and (_05801_, _05278_, _04153_);
  or (_05802_, _05801_, _03575_);
  or (_05803_, _05802_, _05800_);
  not (_05804_, _05462_);
  or (_05805_, _05417_, _04716_);
  or (_05806_, _05415_, _04718_);
  and (_05807_, _05806_, _05408_);
  nand (_05808_, _05807_, _05805_);
  or (_05809_, _05417_, _04724_);
  or (_05810_, _05415_, _04722_);
  and (_05811_, _05810_, _05421_);
  nand (_05812_, _05811_, _05809_);
  nand (_05813_, _05812_, _05808_);
  nand (_05814_, _05813_, _05400_);
  or (_05815_, _05417_, _04736_);
  or (_05816_, _05415_, _04739_);
  and (_05817_, _05816_, _05408_);
  nand (_05818_, _05817_, _05815_);
  or (_05819_, _05417_, _04732_);
  or (_05820_, _05415_, _04730_);
  and (_05821_, _05820_, _05421_);
  nand (_05822_, _05821_, _05819_);
  nand (_05823_, _05822_, _05818_);
  nand (_05824_, _05823_, _05401_);
  and (_05825_, _05824_, _05390_);
  and (_05826_, _05825_, _05814_);
  or (_05827_, _05417_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05828_, _05415_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05829_, _05828_, _05827_);
  nand (_05830_, _05829_, _05421_);
  or (_05831_, _05417_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_05832_, _05415_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_05833_, _05832_, _05831_);
  nand (_05834_, _05833_, _05408_);
  nand (_05835_, _05834_, _05830_);
  nand (_05836_, _05835_, _05400_);
  or (_05837_, _05417_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05838_, _05415_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05839_, _05838_, _05837_);
  nand (_05840_, _05839_, _05421_);
  or (_05841_, _05417_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_05842_, _05415_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_05843_, _05842_, _05841_);
  nand (_05844_, _05843_, _05408_);
  nand (_05845_, _05844_, _05840_);
  nand (_05846_, _05845_, _05401_);
  and (_05847_, _05846_, _05391_);
  and (_05848_, _05847_, _05836_);
  or (_05849_, _05848_, _05826_);
  not (_05850_, _05849_);
  or (_05851_, _05417_, _03943_);
  or (_05852_, _05415_, _03945_);
  and (_05853_, _05852_, _05408_);
  nand (_05854_, _05853_, _05851_);
  or (_05855_, _05417_, _03951_);
  or (_05856_, _05415_, _03949_);
  and (_05857_, _05856_, _05421_);
  nand (_05858_, _05857_, _05855_);
  nand (_05859_, _05858_, _05854_);
  nand (_05860_, _05859_, _05400_);
  or (_05861_, _05417_, _03963_);
  or (_05862_, _05415_, _03965_);
  and (_05863_, _05862_, _05408_);
  nand (_05864_, _05863_, _05861_);
  or (_05865_, _05417_, _03959_);
  or (_05866_, _05415_, _03957_);
  and (_05867_, _05866_, _05421_);
  nand (_05868_, _05867_, _05865_);
  nand (_05869_, _05868_, _05864_);
  nand (_05870_, _05869_, _05401_);
  and (_05871_, _05870_, _05390_);
  and (_05872_, _05871_, _05860_);
  or (_05873_, _05417_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_05874_, _05415_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_05875_, _05874_, _05873_);
  nand (_05876_, _05875_, _05421_);
  or (_05877_, _05417_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_05878_, _05415_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_05879_, _05878_, _05877_);
  nand (_05880_, _05879_, _05408_);
  nand (_05881_, _05880_, _05876_);
  nand (_05882_, _05881_, _05400_);
  or (_05883_, _05417_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_05884_, _05415_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_05885_, _05884_, _05883_);
  nand (_05886_, _05885_, _05421_);
  or (_05887_, _05417_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_05888_, _05415_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_05889_, _05888_, _05887_);
  nand (_05890_, _05889_, _05408_);
  nand (_05891_, _05890_, _05886_);
  nand (_05892_, _05891_, _05401_);
  and (_05893_, _05892_, _05391_);
  and (_05894_, _05893_, _05882_);
  nor (_05895_, _05894_, _05872_);
  or (_05896_, _05417_, _03353_);
  or (_05897_, _05415_, _03750_);
  and (_05898_, _05897_, _05408_);
  nand (_05899_, _05898_, _05896_);
  or (_05900_, _05417_, _03758_);
  or (_05901_, _05415_, _03755_);
  and (_05902_, _05901_, _05421_);
  nand (_05903_, _05902_, _05900_);
  nand (_05904_, _05903_, _05899_);
  nand (_05905_, _05904_, _05400_);
  or (_05906_, _05417_, _03771_);
  or (_05907_, _05415_, _03773_);
  and (_05908_, _05907_, _05408_);
  nand (_05909_, _05908_, _05906_);
  or (_05910_, _05417_, _03767_);
  or (_05911_, _05415_, _03765_);
  and (_05912_, _05911_, _05421_);
  nand (_05913_, _05912_, _05910_);
  nand (_05914_, _05913_, _05909_);
  nand (_05915_, _05914_, _05401_);
  and (_05916_, _05915_, _05390_);
  and (_05917_, _05916_, _05905_);
  or (_05918_, _05417_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_05919_, _05415_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_05920_, _05919_, _05918_);
  nand (_05921_, _05920_, _05421_);
  or (_05922_, _05417_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_05923_, _05415_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_05924_, _05923_, _05922_);
  nand (_05925_, _05924_, _05408_);
  nand (_05926_, _05925_, _05921_);
  nand (_05927_, _05926_, _05400_);
  or (_05928_, _05417_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_05929_, _05415_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_05930_, _05929_, _05928_);
  nand (_05931_, _05930_, _05421_);
  or (_05932_, _05417_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_05933_, _05415_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_05934_, _05933_, _05932_);
  nand (_05935_, _05934_, _05408_);
  nand (_05936_, _05935_, _05931_);
  nand (_05937_, _05936_, _05401_);
  and (_05938_, _05937_, _05391_);
  and (_05939_, _05938_, _05927_);
  nor (_05940_, _05939_, _05917_);
  and (_05941_, _05940_, _05895_);
  or (_05942_, _05417_, _04188_);
  or (_05943_, _05415_, _04190_);
  and (_05944_, _05943_, _05408_);
  nand (_05945_, _05944_, _05942_);
  or (_05946_, _05417_, _04196_);
  or (_05947_, _05415_, _04194_);
  and (_05948_, _05947_, _05421_);
  nand (_05949_, _05948_, _05946_);
  nand (_05950_, _05949_, _05945_);
  nand (_05951_, _05950_, _05400_);
  or (_05952_, _05417_, _04208_);
  or (_05953_, _05415_, _04210_);
  and (_05954_, _05953_, _05408_);
  nand (_05955_, _05954_, _05952_);
  or (_05956_, _05417_, _04204_);
  or (_05957_, _05415_, _04202_);
  and (_05958_, _05957_, _05421_);
  nand (_05959_, _05958_, _05956_);
  nand (_05960_, _05959_, _05955_);
  nand (_05961_, _05960_, _05401_);
  and (_05962_, _05961_, _05390_);
  and (_05963_, _05962_, _05951_);
  or (_05964_, _05417_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05965_, _05415_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_05966_, _05965_, _05964_);
  nand (_05967_, _05966_, _05421_);
  or (_05968_, _05417_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_05969_, _05415_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_05970_, _05969_, _05968_);
  nand (_05971_, _05970_, _05408_);
  nand (_05972_, _05971_, _05967_);
  nand (_05973_, _05972_, _05400_);
  or (_05974_, _05417_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05975_, _05415_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_05976_, _05975_, _05974_);
  nand (_05977_, _05976_, _05421_);
  or (_05978_, _05417_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_05979_, _05415_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_05980_, _05979_, _05978_);
  nand (_05981_, _05980_, _05408_);
  nand (_05982_, _05981_, _05977_);
  nand (_05983_, _05982_, _05401_);
  and (_05984_, _05983_, _05391_);
  and (_05985_, _05984_, _05973_);
  nor (_05986_, _05985_, _05963_);
  or (_05987_, _05417_, _04368_);
  or (_05988_, _05415_, _04371_);
  and (_05989_, _05988_, _05408_);
  nand (_05990_, _05989_, _05987_);
  or (_05991_, _05417_, _04380_);
  or (_05992_, _05415_, _04377_);
  and (_05993_, _05992_, _05421_);
  nand (_05994_, _05993_, _05991_);
  nand (_05995_, _05994_, _05990_);
  nand (_05996_, _05995_, _05400_);
  or (_05997_, _05417_, _04397_);
  or (_05998_, _05415_, _04399_);
  and (_05999_, _05998_, _05408_);
  nand (_06000_, _05999_, _05997_);
  or (_06001_, _05417_, _04392_);
  or (_06002_, _05415_, _04389_);
  and (_06003_, _06002_, _05421_);
  nand (_06004_, _06003_, _06001_);
  nand (_06005_, _06004_, _06000_);
  nand (_06006_, _06005_, _05401_);
  and (_06007_, _06006_, _05390_);
  and (_06008_, _06007_, _05996_);
  or (_06009_, _05417_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06010_, _05415_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_06011_, _06010_, _06009_);
  nand (_06012_, _06011_, _05421_);
  or (_06013_, _05417_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_06014_, _05415_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_06015_, _06014_, _06013_);
  nand (_06016_, _06015_, _05408_);
  nand (_06017_, _06016_, _06012_);
  nand (_06018_, _06017_, _05400_);
  or (_06019_, _05417_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06020_, _05415_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_06021_, _06020_, _06019_);
  nand (_06022_, _06021_, _05421_);
  or (_06023_, _05417_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_06024_, _05415_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_06025_, _06024_, _06023_);
  nand (_06026_, _06025_, _05408_);
  nand (_06027_, _06026_, _06022_);
  nand (_06028_, _06027_, _05401_);
  and (_06029_, _06028_, _05391_);
  and (_06030_, _06029_, _06018_);
  nor (_06031_, _06030_, _06008_);
  and (_06032_, _06031_, _05986_);
  and (_06033_, _06032_, _05941_);
  or (_06034_, _05417_, _04820_);
  or (_06035_, _05415_, _04822_);
  and (_06036_, _06035_, _05408_);
  nand (_06037_, _06036_, _06034_);
  or (_06038_, _05417_, _04828_);
  or (_06039_, _05415_, _04826_);
  and (_06040_, _06039_, _05421_);
  nand (_06041_, _06040_, _06038_);
  nand (_06042_, _06041_, _06037_);
  nand (_06043_, _06042_, _05400_);
  or (_06044_, _05417_, _04841_);
  or (_06045_, _05415_, _04843_);
  and (_06046_, _06045_, _05408_);
  nand (_06047_, _06046_, _06044_);
  or (_06048_, _05417_, _04836_);
  or (_06049_, _05415_, _04834_);
  and (_06050_, _06049_, _05421_);
  nand (_06051_, _06050_, _06048_);
  nand (_06052_, _06051_, _06047_);
  nand (_06053_, _06052_, _05401_);
  and (_06054_, _06053_, _05390_);
  and (_06055_, _06054_, _06043_);
  or (_06056_, _05417_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06057_, _05415_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_06058_, _06057_, _06056_);
  nand (_06059_, _06058_, _05421_);
  or (_06060_, _05417_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_06061_, _05415_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_06062_, _06061_, _06060_);
  nand (_06063_, _06062_, _05408_);
  nand (_06064_, _06063_, _06059_);
  nand (_06065_, _06064_, _05400_);
  or (_06066_, _05417_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06067_, _05415_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_06068_, _06067_, _06066_);
  nand (_06069_, _06068_, _05421_);
  or (_06070_, _05417_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_06071_, _05415_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_06072_, _06071_, _06070_);
  nand (_06073_, _06072_, _05408_);
  nand (_06074_, _06073_, _06069_);
  nand (_06075_, _06074_, _05401_);
  and (_06076_, _06075_, _05391_);
  and (_06077_, _06076_, _06065_);
  nor (_06078_, _06077_, _06055_);
  or (_06079_, _05417_, _04925_);
  or (_06080_, _05415_, _04927_);
  and (_06081_, _06080_, _05408_);
  nand (_06082_, _06081_, _06079_);
  or (_06083_, _05417_, _04933_);
  or (_06084_, _05415_, _04931_);
  and (_06085_, _06084_, _05421_);
  nand (_06086_, _06085_, _06083_);
  nand (_06087_, _06086_, _06082_);
  nand (_06088_, _06087_, _05400_);
  or (_06089_, _05417_, _04946_);
  or (_06090_, _05415_, _04948_);
  and (_06091_, _06090_, _05408_);
  nand (_06092_, _06091_, _06089_);
  or (_06093_, _05417_, _04942_);
  or (_06094_, _05415_, _04939_);
  and (_06095_, _06094_, _05421_);
  nand (_06096_, _06095_, _06093_);
  nand (_06097_, _06096_, _06092_);
  nand (_06098_, _06097_, _05401_);
  and (_06099_, _06098_, _05390_);
  and (_06100_, _06099_, _06088_);
  or (_06101_, _05417_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06102_, _05415_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_06103_, _06102_, _06101_);
  nand (_06104_, _06103_, _05421_);
  or (_06105_, _05417_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_06106_, _05415_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_06107_, _06106_, _06105_);
  nand (_06108_, _06107_, _05408_);
  nand (_06109_, _06108_, _06104_);
  nand (_06110_, _06109_, _05400_);
  or (_06111_, _05417_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06112_, _05415_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_06113_, _06112_, _06111_);
  nand (_06114_, _06113_, _05421_);
  or (_06115_, _05417_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_06116_, _05415_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_06117_, _06116_, _06115_);
  nand (_06118_, _06117_, _05408_);
  nand (_06119_, _06118_, _06114_);
  nand (_06120_, _06119_, _05401_);
  and (_06121_, _06120_, _05391_);
  and (_06122_, _06121_, _06110_);
  nor (_06123_, _06122_, _06100_);
  and (_06124_, _06123_, _06078_);
  and (_06125_, _06124_, _06033_);
  and (_06126_, _06125_, _05850_);
  nor (_06127_, _06126_, _05804_);
  and (_06128_, _06126_, _05804_);
  or (_06129_, _06128_, _06127_);
  or (_06130_, _06129_, _03909_);
  and (_06131_, _06130_, _04333_);
  and (_06132_, _06131_, _05803_);
  and (_06133_, _05474_, _03908_);
  or (_06134_, _06133_, _02939_);
  or (_06135_, _06134_, _06132_);
  and (_06136_, _06135_, _05261_);
  or (_06137_, _06136_, _02525_);
  and (_06138_, _05369_, _02525_);
  nor (_06139_, _06138_, _02797_);
  and (_06140_, _06139_, _06137_);
  nor (_06141_, _03737_, _03302_);
  not (_06142_, _06141_);
  and (_06143_, _05528_, _02797_);
  or (_06144_, _06143_, _06142_);
  or (_06145_, _06144_, _06140_);
  and (_06146_, _06145_, _05252_);
  and (_06147_, _05250_, _04119_);
  or (_06148_, _06147_, _03920_);
  or (_06149_, _06148_, _06146_);
  not (_06150_, _03923_);
  or (_06151_, _05894_, _05872_);
  or (_06152_, _05939_, _05917_);
  and (_06153_, _06152_, _06151_);
  or (_06154_, _05985_, _05963_);
  or (_06155_, _06030_, _06008_);
  and (_06156_, _06155_, _06154_);
  and (_06157_, _06156_, _06153_);
  or (_06158_, _06077_, _06055_);
  or (_06159_, _06122_, _06100_);
  and (_06160_, _06159_, _06158_);
  and (_06161_, _06160_, _06157_);
  and (_06162_, _06161_, _05849_);
  nor (_06163_, _06162_, _05804_);
  and (_06164_, _06162_, _05804_);
  or (_06165_, _06164_, _06163_);
  or (_06166_, _06165_, _03921_);
  and (_06167_, _06166_, _06150_);
  and (_06168_, _06167_, _06149_);
  or (_06169_, _06168_, _05236_);
  and (_06170_, _06169_, _04184_);
  or (_06171_, _06170_, _04550_);
  and (_06172_, _06171_, _04549_);
  not (_06173_, _02939_);
  and (_06174_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06175_, _06174_, \oc8051_golden_model_1.PC [10]);
  and (_06176_, _06175_, _05257_);
  and (_06177_, _06176_, \oc8051_golden_model_1.PC [11]);
  and (_06178_, _06177_, \oc8051_golden_model_1.PC [12]);
  and (_06179_, _06178_, \oc8051_golden_model_1.PC [13]);
  and (_06180_, _06179_, \oc8051_golden_model_1.PC [14]);
  nor (_06181_, _06180_, \oc8051_golden_model_1.PC [15]);
  and (_06182_, _06174_, _05257_);
  and (_06183_, _06182_, \oc8051_golden_model_1.PC [10]);
  and (_06184_, _06183_, \oc8051_golden_model_1.PC [11]);
  and (_06185_, _06184_, \oc8051_golden_model_1.PC [12]);
  and (_06186_, _06185_, \oc8051_golden_model_1.PC [13]);
  and (_06187_, _06186_, \oc8051_golden_model_1.PC [14]);
  and (_06188_, _06187_, \oc8051_golden_model_1.PC [15]);
  nor (_06189_, _06188_, _06181_);
  or (_06190_, _06189_, _06173_);
  and (_06191_, _06175_, _05366_);
  and (_06192_, _06191_, \oc8051_golden_model_1.PC [11]);
  and (_06193_, _06192_, \oc8051_golden_model_1.PC [12]);
  and (_06194_, _06193_, \oc8051_golden_model_1.PC [13]);
  and (_06195_, _06194_, \oc8051_golden_model_1.PC [14]);
  nor (_06196_, _06195_, \oc8051_golden_model_1.PC [15]);
  and (_06197_, _05366_, \oc8051_golden_model_1.PC [8]);
  and (_06198_, _06197_, \oc8051_golden_model_1.PC [9]);
  and (_06199_, _06198_, \oc8051_golden_model_1.PC [10]);
  and (_06200_, _06199_, \oc8051_golden_model_1.PC [11]);
  and (_06201_, _06200_, \oc8051_golden_model_1.PC [12]);
  and (_06202_, _06201_, \oc8051_golden_model_1.PC [13]);
  and (_06203_, _06202_, \oc8051_golden_model_1.PC [14]);
  and (_06204_, _06203_, \oc8051_golden_model_1.PC [15]);
  nor (_06205_, _06204_, _06196_);
  or (_06206_, _06205_, _02939_);
  and (_06207_, _06206_, _06190_);
  and (_06208_, _06207_, _04544_);
  and (_06209_, _06208_, _04547_);
  or (_40484_, _06209_, _06172_);
  not (_06210_, \oc8051_golden_model_1.B [7]);
  nor (_06211_, _42668_, _06210_);
  nor (_06212_, _04696_, _06210_);
  and (_06213_, _05774_, _04696_);
  or (_06214_, _06213_, _06212_);
  and (_06215_, _06214_, _03127_);
  and (_06216_, _04696_, _04604_);
  or (_06217_, _06216_, _06212_);
  or (_06218_, _06217_, _05535_);
  nor (_06219_, _05333_, _06210_);
  and (_06220_, _05356_, _05333_);
  or (_06221_, _06220_, _06219_);
  and (_06222_, _06221_, _02876_);
  and (_06223_, _05474_, _04696_);
  or (_06224_, _06223_, _06212_);
  or (_06225_, _06224_, _03810_);
  and (_06226_, _04696_, \oc8051_golden_model_1.ACC [7]);
  or (_06227_, _06226_, _06212_);
  and (_06228_, _06227_, _03813_);
  nor (_06229_, _03813_, _06210_);
  or (_06230_, _06229_, _02974_);
  or (_06231_, _06230_, _06228_);
  and (_06232_, _06231_, _02881_);
  and (_06233_, _06232_, _06225_);
  and (_06234_, _05360_, _05333_);
  or (_06235_, _06234_, _06219_);
  and (_06236_, _06235_, _02880_);
  or (_06237_, _06236_, _03069_);
  or (_06238_, _06237_, _06233_);
  or (_06239_, _06217_, _03336_);
  and (_06240_, _06239_, _06238_);
  or (_06241_, _06240_, _03075_);
  or (_06242_, _06227_, _03084_);
  and (_06243_, _06242_, _02877_);
  and (_06244_, _06243_, _06241_);
  or (_06245_, _06244_, _06222_);
  and (_06246_, _06245_, _02870_);
  and (_06247_, _02951_, _03099_);
  or (_06248_, _06219_, _05502_);
  and (_06249_, _06248_, _02869_);
  and (_06250_, _06249_, _06235_);
  or (_06251_, _06250_, _06247_);
  or (_06252_, _06251_, _06246_);
  not (_06253_, _06247_);
  and (_06254_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06255_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06256_, _06255_, _06254_);
  and (_06257_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06258_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_06259_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_06260_, _06259_, _06258_);
  nor (_06261_, _06260_, _06256_);
  and (_06262_, _06261_, _06257_);
  nor (_06263_, _06262_, _06256_);
  and (_06264_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06265_, _06264_, _06258_);
  and (_06266_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06267_, _06266_, _06254_);
  nor (_06268_, _06267_, _06265_);
  not (_06269_, _06268_);
  nor (_06270_, _06269_, _06263_);
  and (_06271_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06272_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06273_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06274_, _06273_, _06272_);
  nor (_06275_, _06273_, _06272_);
  nor (_06276_, _06275_, _06274_);
  and (_06277_, _06276_, _06271_);
  nor (_06278_, _06276_, _06271_);
  nor (_06279_, _06278_, _06277_);
  and (_06280_, _06269_, _06263_);
  nor (_06281_, _06280_, _06270_);
  and (_06282_, _06281_, _06279_);
  nor (_06283_, _06282_, _06270_);
  not (_06284_, _06258_);
  and (_06285_, _06264_, _06284_);
  and (_06286_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06287_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06288_, _06287_, _06272_);
  and (_06289_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06290_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06291_, _06290_, _06289_);
  nor (_06292_, _06291_, _06288_);
  and (_06293_, _06292_, _06286_);
  nor (_06294_, _06292_, _06286_);
  nor (_06295_, _06294_, _06293_);
  and (_06296_, _06295_, _06285_);
  nor (_06297_, _06295_, _06285_);
  nor (_06298_, _06297_, _06296_);
  not (_06299_, _06298_);
  nor (_06300_, _06299_, _06283_);
  and (_06301_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06302_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06303_, _06302_, _06301_);
  nor (_06304_, _06277_, _06274_);
  and (_06305_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06306_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06307_, _06306_, _06305_);
  nor (_06308_, _06306_, _06305_);
  nor (_06309_, _06308_, _06307_);
  not (_06310_, _06309_);
  nor (_06311_, _06310_, _06304_);
  and (_06312_, _06310_, _06304_);
  nor (_06313_, _06312_, _06311_);
  and (_06314_, _06313_, _06303_);
  nor (_06315_, _06313_, _06303_);
  nor (_06316_, _06315_, _06314_);
  and (_06317_, _06299_, _06283_);
  nor (_06318_, _06317_, _06300_);
  and (_06319_, _06318_, _06316_);
  nor (_06320_, _06319_, _06300_);
  nor (_06321_, _06293_, _06288_);
  and (_06322_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06323_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06324_, _06323_, _06322_);
  nor (_06325_, _06323_, _06322_);
  nor (_06326_, _06325_, _06324_);
  not (_06327_, _06326_);
  nor (_06328_, _06327_, _06321_);
  and (_06329_, _06327_, _06321_);
  nor (_06330_, _06329_, _06328_);
  and (_06331_, _06330_, _06307_);
  nor (_06332_, _06330_, _06307_);
  nor (_06333_, _06332_, _06331_);
  nor (_06334_, _06296_, _06265_);
  and (_06335_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_06336_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_06337_, _06336_, _06287_);
  nor (_06338_, _06336_, _06287_);
  nor (_06339_, _06338_, _06337_);
  and (_06340_, _06339_, _06335_);
  nor (_06341_, _06339_, _06335_);
  nor (_06342_, _06341_, _06340_);
  not (_06343_, _06342_);
  nor (_06344_, _06343_, _06334_);
  and (_06345_, _06343_, _06334_);
  nor (_06346_, _06345_, _06344_);
  and (_06347_, _06346_, _06333_);
  nor (_06348_, _06346_, _06333_);
  nor (_06349_, _06348_, _06347_);
  not (_06350_, _06349_);
  nor (_06351_, _06350_, _06320_);
  nor (_06352_, _06314_, _06311_);
  not (_06353_, _06352_);
  and (_06354_, _06350_, _06320_);
  nor (_06355_, _06354_, _06351_);
  and (_06356_, _06355_, _06353_);
  nor (_06357_, _06356_, _06351_);
  nor (_06358_, _06331_, _06328_);
  not (_06359_, _06358_);
  nor (_06360_, _06347_, _06344_);
  not (_06361_, _06360_);
  and (_06362_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_06363_, _06362_, _06287_);
  and (_06364_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_06365_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_06366_, _06365_, _06364_);
  nor (_06367_, _06366_, _06363_);
  nor (_06368_, _06340_, _06337_);
  and (_06369_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_06370_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_06371_, _06370_, _06369_);
  nor (_06372_, _06370_, _06369_);
  nor (_06373_, _06372_, _06371_);
  not (_06374_, _06373_);
  nor (_06375_, _06374_, _06368_);
  and (_06376_, _06374_, _06368_);
  nor (_06377_, _06376_, _06375_);
  and (_06378_, _06377_, _06324_);
  nor (_06379_, _06377_, _06324_);
  nor (_06380_, _06379_, _06378_);
  and (_06381_, _06380_, _06367_);
  nor (_06382_, _06380_, _06367_);
  nor (_06383_, _06382_, _06381_);
  and (_06384_, _06383_, _06361_);
  nor (_06385_, _06383_, _06361_);
  nor (_06386_, _06385_, _06384_);
  and (_06387_, _06386_, _06359_);
  nor (_06388_, _06386_, _06359_);
  nor (_06389_, _06388_, _06387_);
  not (_06390_, _06389_);
  nor (_06391_, _06390_, _06357_);
  nor (_06392_, _06387_, _06384_);
  nor (_06393_, _06378_, _06375_);
  not (_06394_, _06393_);
  and (_06395_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_06396_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_06397_, _06396_, _06395_);
  nor (_06398_, _06396_, _06395_);
  nor (_06399_, _06398_, _06397_);
  and (_06400_, _06399_, _06363_);
  nor (_06401_, _06399_, _06363_);
  nor (_06402_, _06401_, _06400_);
  and (_06403_, _06402_, _06371_);
  nor (_06404_, _06402_, _06371_);
  nor (_06405_, _06404_, _06403_);
  and (_06406_, _06405_, _06362_);
  nor (_06407_, _06405_, _06362_);
  nor (_06408_, _06407_, _06406_);
  and (_06409_, _06408_, _06381_);
  nor (_06410_, _06408_, _06381_);
  nor (_06411_, _06410_, _06409_);
  and (_06412_, _06411_, _06394_);
  nor (_06413_, _06411_, _06394_);
  nor (_06414_, _06413_, _06412_);
  not (_06415_, _06414_);
  nor (_06416_, _06415_, _06392_);
  and (_06417_, _06415_, _06392_);
  nor (_06418_, _06417_, _06416_);
  and (_06419_, _06418_, _06391_);
  nor (_06420_, _06412_, _06409_);
  nor (_06421_, _06403_, _06400_);
  not (_06422_, _06421_);
  and (_06423_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_06424_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_06425_, _06424_, _06423_);
  nor (_06426_, _06424_, _06423_);
  nor (_06427_, _06426_, _06425_);
  and (_06428_, _06427_, _06397_);
  nor (_06429_, _06427_, _06397_);
  nor (_06430_, _06429_, _06428_);
  and (_06431_, _06430_, _06406_);
  nor (_06432_, _06430_, _06406_);
  nor (_06433_, _06432_, _06431_);
  and (_06434_, _06433_, _06422_);
  nor (_06435_, _06433_, _06422_);
  nor (_06436_, _06435_, _06434_);
  not (_06437_, _06436_);
  nor (_06438_, _06437_, _06420_);
  and (_06439_, _06437_, _06420_);
  nor (_06440_, _06439_, _06438_);
  and (_06441_, _06440_, _06416_);
  nor (_06442_, _06440_, _06416_);
  nor (_06443_, _06442_, _06441_);
  nor (_06444_, _06443_, _06419_);
  and (_06445_, _06443_, _06419_);
  not (_06446_, _06445_);
  and (_06447_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_06448_, _06447_, _06258_);
  and (_06449_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_06450_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_06451_, _06450_, _06255_);
  nor (_06452_, _06451_, _06448_);
  and (_06453_, _06452_, _06449_);
  nor (_06454_, _06453_, _06448_);
  not (_06455_, _06454_);
  nor (_06456_, _06261_, _06257_);
  nor (_06457_, _06456_, _06262_);
  and (_06458_, _06457_, _06455_);
  and (_06459_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_06460_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_06461_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_06462_, _06461_, _06460_);
  nor (_06463_, _06461_, _06460_);
  nor (_06464_, _06463_, _06462_);
  and (_06465_, _06464_, _06459_);
  nor (_06466_, _06464_, _06459_);
  nor (_06467_, _06466_, _06465_);
  nor (_06468_, _06457_, _06455_);
  nor (_06469_, _06468_, _06458_);
  and (_06470_, _06469_, _06467_);
  nor (_06471_, _06470_, _06458_);
  nor (_06472_, _06281_, _06279_);
  nor (_06473_, _06472_, _06282_);
  not (_06474_, _06473_);
  nor (_06475_, _06474_, _06471_);
  and (_06476_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_06477_, _06476_, _06302_);
  nor (_06478_, _06465_, _06462_);
  nor (_06479_, _06302_, _06301_);
  nor (_06480_, _06479_, _06303_);
  not (_06481_, _06480_);
  nor (_06482_, _06481_, _06478_);
  and (_06483_, _06481_, _06478_);
  nor (_06484_, _06483_, _06482_);
  and (_06485_, _06484_, _06477_);
  nor (_06486_, _06484_, _06477_);
  nor (_06487_, _06486_, _06485_);
  and (_06488_, _06474_, _06471_);
  nor (_06489_, _06488_, _06475_);
  and (_06490_, _06489_, _06487_);
  nor (_06491_, _06490_, _06475_);
  nor (_06492_, _06318_, _06316_);
  nor (_06493_, _06492_, _06319_);
  not (_06494_, _06493_);
  nor (_06495_, _06494_, _06491_);
  nor (_06496_, _06485_, _06482_);
  not (_06497_, _06496_);
  and (_06498_, _06494_, _06491_);
  nor (_06499_, _06498_, _06495_);
  and (_06500_, _06499_, _06497_);
  nor (_06501_, _06500_, _06495_);
  nor (_06502_, _06355_, _06353_);
  nor (_06503_, _06502_, _06356_);
  not (_06504_, _06503_);
  nor (_06505_, _06504_, _06501_);
  and (_06506_, _06390_, _06357_);
  nor (_06507_, _06506_, _06391_);
  and (_06508_, _06507_, _06505_);
  nor (_06509_, _06418_, _06391_);
  nor (_06510_, _06509_, _06419_);
  and (_06511_, _06510_, _06508_);
  and (_06512_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_06513_, _06512_, _06447_);
  and (_06514_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_06515_, _06512_, _06447_);
  nor (_06516_, _06515_, _06513_);
  and (_06517_, _06516_, _06514_);
  nor (_06518_, _06517_, _06513_);
  not (_06519_, _06518_);
  nor (_06520_, _06452_, _06449_);
  nor (_06521_, _06520_, _06453_);
  and (_06522_, _06521_, _06519_);
  and (_06523_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_06524_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_06525_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_06526_, _06525_, _06524_);
  nor (_06527_, _06525_, _06524_);
  nor (_06528_, _06527_, _06526_);
  and (_06529_, _06528_, _06523_);
  nor (_06530_, _06528_, _06523_);
  nor (_06531_, _06530_, _06529_);
  nor (_06532_, _06521_, _06519_);
  nor (_06533_, _06532_, _06522_);
  and (_06534_, _06533_, _06531_);
  nor (_06535_, _06534_, _06522_);
  not (_06536_, _06535_);
  nor (_06537_, _06469_, _06467_);
  nor (_06538_, _06537_, _06470_);
  and (_06539_, _06538_, _06536_);
  nor (_06540_, _06529_, _06526_);
  and (_06541_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_06542_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_06543_, _06542_, _06541_);
  nor (_06544_, _06543_, _06477_);
  not (_06545_, _06544_);
  nor (_06546_, _06545_, _06540_);
  and (_06547_, _06545_, _06540_);
  nor (_06548_, _06547_, _06546_);
  nor (_06549_, _06538_, _06536_);
  nor (_06550_, _06549_, _06539_);
  and (_06551_, _06550_, _06548_);
  nor (_06552_, _06551_, _06539_);
  nor (_06553_, _06489_, _06487_);
  nor (_06554_, _06553_, _06490_);
  not (_06555_, _06554_);
  nor (_06556_, _06555_, _06552_);
  and (_06557_, _06555_, _06552_);
  nor (_06558_, _06557_, _06556_);
  and (_06559_, _06558_, _06546_);
  nor (_06560_, _06559_, _06556_);
  nor (_06561_, _06499_, _06497_);
  nor (_06562_, _06561_, _06500_);
  not (_06563_, _06562_);
  nor (_06564_, _06563_, _06560_);
  and (_06565_, _06504_, _06501_);
  nor (_06566_, _06565_, _06505_);
  and (_06567_, _06566_, _06564_);
  nor (_06568_, _06507_, _06505_);
  nor (_06569_, _06568_, _06508_);
  and (_06570_, _06569_, _06567_);
  nor (_06571_, _06569_, _06567_);
  nor (_06572_, _06571_, _06570_);
  and (_06573_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_06574_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_06575_, _06574_, _06573_);
  and (_06576_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06577_, _06574_, _06573_);
  nor (_06578_, _06577_, _06575_);
  and (_06579_, _06578_, _06576_);
  nor (_06580_, _06579_, _06575_);
  not (_06581_, _06580_);
  nor (_06582_, _06516_, _06514_);
  nor (_06583_, _06582_, _06517_);
  and (_06584_, _06583_, _06581_);
  and (_06585_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_06586_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_06587_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_06588_, _06587_, _06586_);
  nor (_06589_, _06587_, _06586_);
  nor (_06590_, _06589_, _06588_);
  and (_06591_, _06590_, _06585_);
  nor (_06592_, _06590_, _06585_);
  nor (_06593_, _06592_, _06591_);
  nor (_06594_, _06583_, _06581_);
  nor (_06595_, _06594_, _06584_);
  and (_06596_, _06595_, _06593_);
  nor (_06597_, _06596_, _06584_);
  not (_06598_, _06597_);
  nor (_06599_, _06533_, _06531_);
  nor (_06600_, _06599_, _06534_);
  and (_06601_, _06600_, _06598_);
  not (_06602_, _06476_);
  nor (_06603_, _06591_, _06588_);
  nor (_06604_, _06603_, _06602_);
  and (_06605_, _06603_, _06602_);
  nor (_06606_, _06605_, _06604_);
  nor (_06607_, _06600_, _06598_);
  nor (_06608_, _06607_, _06601_);
  and (_06609_, _06608_, _06606_);
  nor (_06610_, _06609_, _06601_);
  not (_06611_, _06610_);
  nor (_06612_, _06550_, _06548_);
  nor (_06613_, _06612_, _06551_);
  and (_06614_, _06613_, _06611_);
  nor (_06615_, _06613_, _06611_);
  nor (_06616_, _06615_, _06614_);
  and (_06617_, _06616_, _06604_);
  nor (_06618_, _06617_, _06614_);
  nor (_06619_, _06558_, _06546_);
  nor (_06620_, _06619_, _06559_);
  not (_06621_, _06620_);
  nor (_06622_, _06621_, _06618_);
  and (_06623_, _06563_, _06560_);
  nor (_06624_, _06623_, _06564_);
  and (_06625_, _06624_, _06622_);
  nor (_06626_, _06566_, _06564_);
  nor (_06627_, _06626_, _06567_);
  and (_06628_, _06627_, _06625_);
  nor (_06629_, _06627_, _06625_);
  nor (_06630_, _06629_, _06628_);
  and (_06631_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_06632_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_06633_, _06632_, _06631_);
  and (_06634_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06635_, _06632_, _06631_);
  nor (_06636_, _06635_, _06633_);
  and (_06637_, _06636_, _06634_);
  nor (_06638_, _06637_, _06633_);
  not (_06639_, _06638_);
  nor (_06640_, _06578_, _06576_);
  nor (_06641_, _06640_, _06579_);
  and (_06642_, _06641_, _06639_);
  and (_06643_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_06644_, _06643_, _06587_);
  and (_06645_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_06646_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_06647_, _06646_, _06645_);
  nor (_06648_, _06647_, _06644_);
  nor (_06649_, _06641_, _06639_);
  nor (_06650_, _06649_, _06642_);
  and (_06651_, _06650_, _06648_);
  nor (_06652_, _06651_, _06642_);
  not (_06653_, _06652_);
  nor (_06654_, _06595_, _06593_);
  nor (_06655_, _06654_, _06596_);
  and (_06656_, _06655_, _06653_);
  nor (_06657_, _06655_, _06653_);
  nor (_06658_, _06657_, _06656_);
  and (_06659_, _06658_, _06644_);
  nor (_06660_, _06659_, _06656_);
  not (_06661_, _06660_);
  nor (_06662_, _06608_, _06606_);
  nor (_06663_, _06662_, _06609_);
  and (_06664_, _06663_, _06661_);
  nor (_06665_, _06616_, _06604_);
  nor (_06666_, _06665_, _06617_);
  and (_06667_, _06666_, _06664_);
  and (_06668_, _06621_, _06618_);
  nor (_06669_, _06668_, _06622_);
  and (_06670_, _06669_, _06667_);
  nor (_06671_, _06624_, _06622_);
  nor (_06672_, _06671_, _06625_);
  and (_06673_, _06672_, _06670_);
  nor (_06674_, _06672_, _06670_);
  nor (_06675_, _06674_, _06673_);
  and (_06676_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_06677_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_06678_, _06677_, _06676_);
  and (_06679_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_06680_, _06677_, _06676_);
  nor (_06681_, _06680_, _06678_);
  and (_06682_, _06681_, _06679_);
  nor (_06683_, _06682_, _06678_);
  not (_06684_, _06683_);
  nor (_06685_, _06636_, _06634_);
  nor (_06686_, _06685_, _06637_);
  and (_06687_, _06686_, _06684_);
  nor (_06688_, _06686_, _06684_);
  nor (_06689_, _06688_, _06687_);
  and (_06690_, _06689_, _06643_);
  nor (_06691_, _06690_, _06687_);
  not (_06692_, _06691_);
  nor (_06693_, _06650_, _06648_);
  nor (_06694_, _06693_, _06651_);
  and (_06695_, _06694_, _06692_);
  nor (_06696_, _06658_, _06644_);
  nor (_06697_, _06696_, _06659_);
  and (_06698_, _06697_, _06695_);
  nor (_06699_, _06663_, _06661_);
  nor (_06700_, _06699_, _06664_);
  and (_06701_, _06700_, _06698_);
  nor (_06702_, _06666_, _06664_);
  nor (_06703_, _06702_, _06667_);
  and (_06704_, _06703_, _06701_);
  nor (_06705_, _06669_, _06667_);
  nor (_06706_, _06705_, _06670_);
  and (_06707_, _06706_, _06704_);
  and (_06708_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_06709_, _06708_, _06677_);
  nor (_06710_, _06681_, _06679_);
  nor (_06711_, _06710_, _06682_);
  and (_06712_, _06711_, _06709_);
  nor (_06713_, _06689_, _06643_);
  nor (_06714_, _06713_, _06690_);
  and (_06715_, _06714_, _06712_);
  nor (_06716_, _06694_, _06692_);
  nor (_06717_, _06716_, _06695_);
  and (_06718_, _06717_, _06715_);
  nor (_06719_, _06697_, _06695_);
  nor (_06720_, _06719_, _06698_);
  and (_06721_, _06720_, _06718_);
  nor (_06722_, _06700_, _06698_);
  nor (_06723_, _06722_, _06701_);
  and (_06724_, _06723_, _06721_);
  nor (_06725_, _06703_, _06701_);
  nor (_06726_, _06725_, _06704_);
  and (_06727_, _06726_, _06724_);
  nor (_06728_, _06706_, _06704_);
  nor (_06729_, _06728_, _06707_);
  and (_06730_, _06729_, _06727_);
  nor (_06732_, _06730_, _06707_);
  not (_06733_, _06732_);
  and (_06734_, _06733_, _06675_);
  nor (_06735_, _06734_, _06673_);
  not (_06736_, _06735_);
  and (_06737_, _06736_, _06630_);
  nor (_06738_, _06737_, _06628_);
  not (_06739_, _06738_);
  and (_06740_, _06739_, _06572_);
  nor (_06741_, _06740_, _06570_);
  not (_06742_, _06741_);
  nor (_06743_, _06510_, _06508_);
  nor (_06744_, _06743_, _06511_);
  and (_06745_, _06744_, _06742_);
  nor (_06746_, _06745_, _06511_);
  and (_06747_, _06746_, _06446_);
  or (_06748_, _06747_, _06444_);
  not (_06749_, _06748_);
  and (_06750_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_06751_, _06750_);
  nor (_06752_, _06751_, _06396_);
  nor (_06753_, _06752_, _06428_);
  nor (_06754_, _06434_, _06431_);
  nor (_06755_, _06754_, _06753_);
  and (_06756_, _06754_, _06753_);
  nor (_06757_, _06756_, _06755_);
  not (_06758_, _06757_);
  nor (_06759_, _06441_, _06438_);
  nor (_06760_, _06759_, _06758_);
  and (_06761_, _06759_, _06758_);
  nor (_06762_, _06761_, _06760_);
  and (_06763_, _06762_, _06749_);
  or (_06764_, _06755_, _06425_);
  or (_06765_, _06764_, _06760_);
  or (_06766_, _06765_, _06763_);
  or (_06767_, _06766_, _06253_);
  and (_06768_, _06767_, _02864_);
  and (_06769_, _06768_, _06252_);
  not (_06770_, _05535_);
  not (_06771_, _05333_);
  nor (_06772_, _05530_, _06771_);
  or (_06773_, _06772_, _06219_);
  and (_06774_, _06773_, _02863_);
  or (_06775_, _06774_, _06770_);
  or (_06776_, _06775_, _06769_);
  and (_06777_, _06776_, _06218_);
  or (_06778_, _06777_, _02853_);
  and (_06779_, _04696_, _05462_);
  or (_06780_, _06212_, _05540_);
  or (_06781_, _06780_, _06779_);
  and (_06782_, _06781_, _02838_);
  and (_06783_, _06782_, _06778_);
  and (_06784_, _02951_, _02517_);
  not (_06785_, _04696_);
  nor (_06786_, _05744_, _06785_);
  or (_06787_, _06786_, _06212_);
  and (_06788_, _06787_, _02579_);
  or (_06789_, _06788_, _06784_);
  or (_06790_, _06789_, _06783_);
  not (_06791_, _06784_);
  nor (_06792_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_06793_, _06792_, _06259_);
  and (_06794_, \oc8051_golden_model_1.B [0], _05771_);
  not (_06795_, _06794_);
  not (_06796_, \oc8051_golden_model_1.B [1]);
  nor (_06797_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_06798_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_06799_, _06798_, _06797_);
  and (_06800_, _06799_, _06796_);
  nor (_06801_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_06802_, _06801_, _06800_);
  and (_06803_, _06802_, _06795_);
  and (_06804_, _06803_, _06793_);
  nor (_06805_, _06803_, _05771_);
  not (_06806_, \oc8051_golden_model_1.ACC [6]);
  and (_06807_, \oc8051_golden_model_1.B [0], _06806_);
  nor (_06808_, _06807_, _05771_);
  nor (_06809_, _06808_, _06796_);
  and (_06810_, _06801_, _06799_);
  not (_06811_, _06810_);
  nor (_06812_, _06811_, _06809_);
  not (_06813_, _06812_);
  and (_06814_, _06813_, _06805_);
  nor (_06815_, _06814_, _06804_);
  and (_06816_, _06812_, \oc8051_golden_model_1.B [0]);
  nor (_06817_, _06816_, _06806_);
  and (_06818_, _06817_, _06796_);
  nor (_06819_, _06817_, _06796_);
  nor (_06820_, _06819_, _06818_);
  nor (_06821_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06822_, _06821_, _06447_);
  nor (_06823_, _06822_, \oc8051_golden_model_1.ACC [4]);
  nor (_06824_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  not (_06825_, \oc8051_golden_model_1.B [0]);
  and (_06826_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06827_, _06826_, _06825_);
  nor (_06828_, _06827_, _06824_);
  nor (_06829_, _06828_, _06823_);
  not (_06830_, _06829_);
  and (_06831_, _06830_, _06820_);
  not (_06832_, _06831_);
  nor (_06833_, _06815_, \oc8051_golden_model_1.B [2]);
  nor (_06834_, _06833_, _06818_);
  and (_06835_, _06834_, _06832_);
  not (_06836_, \oc8051_golden_model_1.B [3]);
  nor (_06837_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06838_, _06837_, _06797_);
  and (_06839_, _06838_, _06836_);
  and (_06840_, \oc8051_golden_model_1.B [2], _05771_);
  not (_06841_, _06840_);
  and (_06842_, _06841_, _06839_);
  not (_06843_, _06842_);
  nor (_06844_, _06843_, _06835_);
  nor (_06845_, _06844_, _06815_);
  nor (_06846_, _06845_, _06804_);
  and (_06847_, _06838_, \oc8051_golden_model_1.ACC [7]);
  nor (_06848_, _06847_, _06839_);
  nor (_06849_, _06846_, \oc8051_golden_model_1.B [3]);
  not (_06850_, \oc8051_golden_model_1.B [2]);
  nor (_06851_, _06830_, _06820_);
  nor (_06852_, _06851_, _06831_);
  not (_06853_, _06852_);
  and (_06854_, _06853_, _06844_);
  nor (_06855_, _06844_, _06817_);
  nor (_06856_, _06855_, _06854_);
  and (_06857_, _06856_, _06850_);
  nor (_06858_, _06856_, _06850_);
  nor (_06859_, _06858_, _06857_);
  not (_06860_, _06859_);
  not (_06861_, \oc8051_golden_model_1.ACC [5]);
  nor (_06862_, _06844_, _06861_);
  and (_06863_, _06844_, _06822_);
  or (_06864_, _06863_, _06862_);
  and (_06865_, _06864_, _06796_);
  nor (_06866_, _06864_, _06796_);
  not (_06867_, \oc8051_golden_model_1.ACC [4]);
  and (_06868_, \oc8051_golden_model_1.B [0], _06867_);
  nor (_06869_, _06868_, _06866_);
  nor (_06870_, _06869_, _06865_);
  nor (_06871_, _06870_, _06860_);
  or (_06872_, _06871_, _06857_);
  nor (_06873_, _06872_, _06849_);
  nor (_06874_, _06873_, _06848_);
  nor (_06875_, _06874_, _06846_);
  nor (_06876_, _06875_, _06804_);
  not (_06877_, _06874_);
  and (_06878_, _06870_, _06860_);
  nor (_06879_, _06878_, _06871_);
  nor (_06880_, _06879_, _06877_);
  nor (_06881_, _06874_, _06856_);
  nor (_06882_, _06881_, _06880_);
  and (_06883_, _06882_, _06836_);
  nor (_06884_, _06882_, _06836_);
  nor (_06885_, _06884_, _06883_);
  not (_06886_, _06885_);
  nor (_06887_, _06874_, _06864_);
  nor (_06888_, _06866_, _06865_);
  and (_06889_, _06888_, _06868_);
  nor (_06890_, _06888_, _06868_);
  nor (_06891_, _06890_, _06889_);
  and (_06892_, _06891_, _06874_);
  or (_06893_, _06892_, _06887_);
  nor (_06894_, _06893_, \oc8051_golden_model_1.B [2]);
  and (_06895_, _06893_, \oc8051_golden_model_1.B [2]);
  nor (_06896_, _06874_, _06867_);
  nor (_06897_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06898_, _06897_, _06573_);
  and (_06899_, _06874_, _06898_);
  or (_06900_, _06899_, _06896_);
  and (_06901_, _06900_, _06796_);
  nor (_06902_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06903_, _06902_, _06631_);
  nor (_06904_, _06903_, \oc8051_golden_model_1.ACC [2]);
  nor (_06905_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06906_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06907_, _06906_, _06825_);
  nor (_06908_, _06907_, _06905_);
  nor (_06909_, _06908_, _06904_);
  not (_06910_, _06909_);
  nor (_06911_, _06900_, _06796_);
  nor (_06912_, _06911_, _06901_);
  and (_06913_, _06912_, _06910_);
  nor (_06914_, _06913_, _06901_);
  nor (_06915_, _06914_, _06895_);
  nor (_06916_, _06915_, _06894_);
  nor (_06917_, _06916_, _06886_);
  nor (_06918_, _06876_, \oc8051_golden_model_1.B [4]);
  nor (_06919_, _06918_, _06883_);
  not (_06920_, _06919_);
  nor (_06921_, _06920_, _06917_);
  not (_06922_, \oc8051_golden_model_1.B [5]);
  and (_06923_, _06837_, _06922_);
  and (_06924_, \oc8051_golden_model_1.B [4], _05771_);
  not (_06925_, _06924_);
  and (_06926_, _06925_, _06923_);
  not (_06927_, _06926_);
  nor (_06928_, _06927_, _06921_);
  nor (_06929_, _06928_, _06876_);
  nor (_06930_, _06929_, _06804_);
  not (_06931_, \oc8051_golden_model_1.B [4]);
  and (_06932_, _06916_, _06886_);
  nor (_06933_, _06932_, _06917_);
  not (_06934_, _06933_);
  and (_06935_, _06934_, _06928_);
  nor (_06936_, _06928_, _06882_);
  nor (_06937_, _06936_, _06935_);
  and (_06938_, _06937_, _06931_);
  nor (_06939_, _06937_, _06931_);
  nor (_06940_, _06939_, _06938_);
  not (_06941_, _06940_);
  nor (_06942_, _06928_, _06893_);
  nor (_06943_, _06895_, _06894_);
  and (_06944_, _06943_, _06914_);
  nor (_06945_, _06943_, _06914_);
  nor (_06946_, _06945_, _06944_);
  not (_06947_, _06946_);
  and (_06948_, _06947_, _06928_);
  nor (_06949_, _06948_, _06942_);
  nor (_06950_, _06949_, \oc8051_golden_model_1.B [3]);
  and (_06951_, _06949_, \oc8051_golden_model_1.B [3]);
  nor (_06952_, _06912_, _06910_);
  nor (_06953_, _06952_, _06913_);
  not (_06954_, _06953_);
  and (_06955_, _06954_, _06928_);
  nor (_06956_, _06928_, _06900_);
  nor (_06957_, _06956_, _06955_);
  and (_06958_, _06957_, _06850_);
  nor (_06959_, _06928_, _02564_);
  and (_06960_, _06928_, _06903_);
  or (_06961_, _06960_, _06959_);
  and (_06962_, _06961_, _06796_);
  nor (_06963_, _06961_, _06796_);
  not (_06964_, \oc8051_golden_model_1.ACC [2]);
  and (_06965_, \oc8051_golden_model_1.B [0], _06964_);
  nor (_06966_, _06965_, _06963_);
  nor (_06967_, _06966_, _06962_);
  nor (_06968_, _06957_, _06850_);
  nor (_06969_, _06968_, _06958_);
  not (_06970_, _06969_);
  nor (_06971_, _06970_, _06967_);
  nor (_06972_, _06971_, _06958_);
  nor (_06973_, _06972_, _06951_);
  nor (_06974_, _06973_, _06950_);
  nor (_06975_, _06974_, _06941_);
  nor (_06976_, _06930_, \oc8051_golden_model_1.B [5]);
  nor (_06977_, _06976_, _06938_);
  not (_06978_, _06977_);
  nor (_06979_, _06978_, _06975_);
  not (_06980_, _06979_);
  not (_06981_, _06837_);
  and (_06982_, \oc8051_golden_model_1.B [5], _05771_);
  nor (_06983_, _06982_, _06981_);
  and (_06984_, _06983_, _06980_);
  nor (_06985_, _06984_, _06930_);
  not (_06986_, _06984_);
  and (_06987_, _06974_, _06941_);
  nor (_06988_, _06987_, _06975_);
  nor (_06989_, _06988_, _06986_);
  nor (_06990_, _06984_, _06937_);
  nor (_06991_, _06990_, _06989_);
  and (_06992_, _06991_, _06922_);
  nor (_06993_, _06991_, _06922_);
  nor (_06994_, _06993_, _06992_);
  not (_06995_, _06994_);
  nor (_06996_, _06984_, _06949_);
  nor (_06997_, _06951_, _06950_);
  nor (_06998_, _06997_, _06972_);
  and (_06999_, _06997_, _06972_);
  or (_07000_, _06999_, _06998_);
  and (_07001_, _07000_, _06984_);
  or (_07002_, _07001_, _06996_);
  and (_07003_, _07002_, _06931_);
  nor (_07004_, _07002_, _06931_);
  and (_07005_, _06970_, _06967_);
  nor (_07006_, _07005_, _06971_);
  nor (_07007_, _07006_, _06986_);
  nor (_07008_, _06984_, _06957_);
  nor (_07009_, _07008_, _07007_);
  and (_07010_, _07009_, _06836_);
  nor (_07011_, _06963_, _06962_);
  nor (_07012_, _07011_, _06965_);
  and (_07013_, _07011_, _06965_);
  or (_07014_, _07013_, _07012_);
  nor (_07015_, _07014_, _06986_);
  nor (_07016_, _06984_, _06961_);
  nor (_07017_, _07016_, _07015_);
  and (_07018_, _07017_, _06850_);
  nor (_07019_, _07017_, _06850_);
  nor (_07020_, _06984_, _06964_);
  nor (_07021_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07022_, _07021_, _06676_);
  and (_07023_, _06984_, _07022_);
  or (_07024_, _07023_, _07020_);
  and (_07025_, _07024_, _06796_);
  and (_07026_, \oc8051_golden_model_1.B [0], _02551_);
  not (_07027_, _07026_);
  nor (_07028_, _07024_, _06796_);
  nor (_07029_, _07028_, _07025_);
  and (_07030_, _07029_, _07027_);
  nor (_07031_, _07030_, _07025_);
  nor (_07032_, _07031_, _07019_);
  nor (_07033_, _07032_, _07018_);
  nor (_07034_, _07009_, _06836_);
  nor (_07035_, _07034_, _07010_);
  not (_07036_, _07035_);
  nor (_07037_, _07036_, _07033_);
  nor (_07038_, _07037_, _07010_);
  nor (_07039_, _07038_, _07004_);
  nor (_07040_, _07039_, _07003_);
  nor (_07041_, _07040_, _06995_);
  nor (_07042_, _07041_, _06992_);
  and (_07043_, _06210_, \oc8051_golden_model_1.ACC [7]);
  nor (_07044_, _07043_, _06837_);
  nor (_07045_, _07044_, _07042_);
  nor (_07046_, _06985_, _06804_);
  nor (_07047_, _07046_, _06981_);
  nor (_07048_, _07047_, _07045_);
  and (_07049_, _07048_, _06985_);
  nor (_07050_, _07049_, _06804_);
  and (_07051_, _07050_, \oc8051_golden_model_1.B [7]);
  and (_07052_, _07050_, _06210_);
  nor (_07053_, _07052_, _06750_);
  not (_07054_, _07053_);
  not (_07055_, \oc8051_golden_model_1.B [6]);
  and (_07056_, _07040_, _06995_);
  nor (_07057_, _07056_, _07041_);
  nor (_07058_, _07057_, _07048_);
  not (_07059_, _07048_);
  nor (_07060_, _07059_, _06991_);
  nor (_07061_, _07060_, _07058_);
  nor (_07062_, _07061_, _07055_);
  and (_07063_, _07061_, _07055_);
  nor (_07064_, _07004_, _07003_);
  nor (_07065_, _07064_, _07038_);
  and (_07066_, _07064_, _07038_);
  or (_07067_, _07066_, _07065_);
  nor (_07068_, _07067_, _07048_);
  nor (_07069_, _07059_, _07002_);
  nor (_07070_, _07069_, _07068_);
  nor (_07071_, _07070_, _06922_);
  and (_07072_, _07070_, _06922_);
  not (_07073_, _07072_);
  and (_07074_, _07036_, _07033_);
  nor (_07075_, _07074_, _07037_);
  nor (_07076_, _07075_, _07048_);
  nor (_07077_, _07059_, _07009_);
  nor (_07078_, _07077_, _07076_);
  nor (_07079_, _07078_, _06931_);
  and (_07080_, _07048_, _07017_);
  nor (_07081_, _07019_, _07018_);
  and (_07082_, _07081_, _07031_);
  nor (_07083_, _07081_, _07031_);
  nor (_07084_, _07083_, _07082_);
  nor (_07085_, _07084_, _07048_);
  or (_07086_, _07085_, _07080_);
  nor (_07087_, _07086_, _06836_);
  and (_07088_, _07086_, _06836_);
  nor (_07089_, _07088_, _07087_);
  nor (_07090_, _07029_, _07027_);
  nor (_07091_, _07090_, _07030_);
  nor (_07092_, _07091_, _07048_);
  nor (_07093_, _07059_, _07024_);
  nor (_07094_, _07093_, _07092_);
  nor (_07095_, _07094_, _06850_);
  and (_07096_, _07094_, _06850_);
  nor (_07097_, _07096_, _07095_);
  and (_07098_, _07097_, _07089_);
  and (_07099_, _07048_, _02551_);
  and (_07100_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07101_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07102_, _07101_, _07100_);
  nor (_07103_, _07048_, _07102_);
  nor (_07104_, _07103_, _07099_);
  and (_07105_, _07104_, _06796_);
  nor (_07106_, _07104_, _06796_);
  and (_07107_, _06825_, \oc8051_golden_model_1.ACC [0]);
  not (_07108_, _07107_);
  nor (_07109_, _07108_, _07106_);
  nor (_07110_, _07109_, _07105_);
  and (_07111_, _07110_, _07098_);
  and (_07112_, _07095_, _07089_);
  nor (_07113_, _07112_, _07087_);
  not (_07114_, _07113_);
  nor (_07115_, _07114_, _07111_);
  and (_07116_, _07078_, _06931_);
  nor (_07117_, _07116_, _07115_);
  or (_07118_, _07117_, _07079_);
  and (_07119_, _07118_, _07073_);
  nor (_07120_, _07119_, _07071_);
  nor (_07121_, _07120_, _07063_);
  or (_07122_, _07121_, _07062_);
  and (_07123_, _07122_, _07054_);
  nor (_07124_, _07123_, _07051_);
  nor (_07125_, _07063_, _07062_);
  and (_07126_, _07125_, _07054_);
  nor (_07127_, _07116_, _07079_);
  nor (_07128_, _07072_, _07071_);
  and (_07129_, _07128_, _07127_);
  and (_07130_, _07129_, _07126_);
  and (_07131_, \oc8051_golden_model_1.B [0], _02667_);
  not (_07132_, _07131_);
  nor (_07133_, _07106_, _07105_);
  and (_07134_, _07133_, _07132_);
  and (_07135_, _07134_, _07108_);
  and (_07136_, _07135_, _07098_);
  and (_07137_, _07136_, _07130_);
  nor (_07138_, _07137_, _07124_);
  and (_07139_, _07138_, _07049_);
  or (_07140_, _07139_, _06804_);
  or (_07141_, _07140_, _06791_);
  and (_07142_, _07141_, _02803_);
  and (_07143_, _07142_, _06790_);
  and (_07144_, _05661_, _04696_);
  or (_07145_, _07144_, _06212_);
  and (_07146_, _07145_, _02802_);
  or (_07147_, _07146_, _02980_);
  or (_07148_, _07147_, _07143_);
  and (_07149_, _05766_, _04696_);
  or (_07150_, _06212_, _03887_);
  or (_07151_, _07150_, _07149_);
  and (_07152_, _07151_, _03128_);
  and (_07153_, _07152_, _07148_);
  or (_07154_, _07153_, _06215_);
  and (_07155_, _07154_, _03883_);
  or (_07156_, _06212_, _04715_);
  and (_07157_, _07145_, _02970_);
  and (_07158_, _07157_, _07156_);
  or (_07159_, _07158_, _07155_);
  and (_07160_, _07159_, _03137_);
  and (_07161_, _06227_, _03135_);
  and (_07162_, _07161_, _07156_);
  or (_07163_, _07162_, _02965_);
  or (_07164_, _07163_, _07160_);
  nor (_07165_, _05765_, _06785_);
  or (_07166_, _06212_, _05783_);
  or (_07167_, _07166_, _07165_);
  and (_07168_, _07167_, _05788_);
  and (_07169_, _07168_, _07164_);
  nor (_07170_, _05773_, _06785_);
  or (_07171_, _07170_, _06212_);
  and (_07172_, _07171_, _03123_);
  or (_07173_, _07172_, _03163_);
  or (_07174_, _07173_, _07169_);
  or (_07175_, _06224_, _03906_);
  and (_07176_, _07175_, _02498_);
  and (_07177_, _07176_, _07174_);
  and (_07178_, _06221_, _02497_);
  or (_07179_, _07178_, _02888_);
  or (_07180_, _07179_, _07177_);
  and (_07181_, _05235_, _04696_);
  or (_07182_, _06212_, _02890_);
  or (_07183_, _07182_, _07181_);
  and (_07184_, _07183_, _42668_);
  and (_07185_, _07184_, _07180_);
  or (_07186_, _07185_, _06211_);
  and (_40486_, _07186_, _43998_);
  nor (_07187_, _42668_, _05771_);
  and (_07188_, _02852_, _02891_);
  nor (_07189_, _04604_, \oc8051_golden_model_1.ACC [7]);
  and (_07190_, _04604_, \oc8051_golden_model_1.ACC [7]);
  nor (_07191_, _07190_, _07189_);
  and (_07192_, _04770_, \oc8051_golden_model_1.ACC [6]);
  nor (_07193_, _04770_, \oc8051_golden_model_1.ACC [6]);
  nor (_07194_, _07193_, _07192_);
  and (_07195_, _04877_, \oc8051_golden_model_1.ACC [5]);
  nor (_07196_, _04877_, \oc8051_golden_model_1.ACC [5]);
  nor (_07197_, _07196_, _07195_);
  not (_07198_, _07197_);
  and (_07199_, _04982_, \oc8051_golden_model_1.ACC [4]);
  nor (_07200_, _04982_, \oc8051_golden_model_1.ACC [4]);
  nor (_07201_, _07200_, _07199_);
  nor (_07202_, _04241_, \oc8051_golden_model_1.ACC [3]);
  not (_07203_, _07202_);
  and (_07204_, _04241_, \oc8051_golden_model_1.ACC [3]);
  not (_07205_, _07204_);
  and (_07206_, _04435_, \oc8051_golden_model_1.ACC [2]);
  nor (_07207_, _04435_, \oc8051_golden_model_1.ACC [2]);
  nor (_07208_, _07207_, _07206_);
  not (_07209_, _07208_);
  and (_07210_, _04000_, \oc8051_golden_model_1.ACC [1]);
  nor (_07211_, _04000_, \oc8051_golden_model_1.ACC [1]);
  nor (_07212_, _07211_, _07210_);
  and (_07213_, _03808_, \oc8051_golden_model_1.ACC [0]);
  and (_07214_, _07213_, _07212_);
  nor (_07215_, _07214_, _07210_);
  nor (_07216_, _07215_, _07209_);
  nor (_07217_, _07216_, _07206_);
  nand (_07218_, _07217_, _07205_);
  and (_07219_, _07218_, _07203_);
  and (_07220_, _07219_, _07201_);
  nor (_07221_, _07220_, _07199_);
  nor (_07222_, _07221_, _07198_);
  or (_07223_, _07222_, _07195_);
  and (_07224_, _07223_, _07194_);
  nor (_07225_, _07224_, _07192_);
  nor (_07226_, _07225_, _07191_);
  and (_07227_, _07225_, _07191_);
  or (_07228_, _07227_, _07226_);
  and (_07229_, _03368_, _02891_);
  not (_07230_, _07229_);
  or (_07231_, _02839_, _02947_);
  and (_07232_, _07231_, _02891_);
  not (_07233_, _07232_);
  and (_07234_, _03508_, _02891_);
  and (_07235_, _04009_, _02891_);
  nor (_07236_, _07235_, _07234_);
  and (_07237_, _07236_, _07233_);
  and (_07238_, _07237_, _07230_);
  or (_07239_, _07238_, _07228_);
  and (_07240_, _02852_, _02967_);
  not (_07241_, _07240_);
  and (_07242_, _06162_, \oc8051_golden_model_1.PSW [7]);
  nor (_07243_, _07242_, _05804_);
  and (_07244_, _07242_, _05804_);
  nor (_07245_, _07244_, _07243_);
  and (_07246_, _07245_, \oc8051_golden_model_1.ACC [7]);
  nor (_07247_, _07245_, \oc8051_golden_model_1.ACC [7]);
  nor (_07248_, _07247_, _07246_);
  and (_07249_, _06161_, \oc8051_golden_model_1.PSW [7]);
  nor (_07250_, _07249_, _05849_);
  nor (_07251_, _07250_, _07242_);
  and (_07252_, _07251_, \oc8051_golden_model_1.ACC [6]);
  nor (_07253_, _07251_, _06806_);
  and (_07254_, _07251_, _06806_);
  nor (_07255_, _07254_, _07253_);
  and (_07256_, _06159_, _06157_);
  and (_07257_, _07256_, \oc8051_golden_model_1.PSW [7]);
  nor (_07258_, _07257_, _06158_);
  nor (_07259_, _07258_, _07249_);
  and (_07260_, _07259_, \oc8051_golden_model_1.ACC [5]);
  nor (_07261_, _07259_, _06861_);
  and (_07262_, _07259_, _06861_);
  nor (_07263_, _07262_, _07261_);
  and (_07264_, _06153_, \oc8051_golden_model_1.PSW [7]);
  and (_07265_, _07264_, _06156_);
  nor (_07266_, _07265_, _06159_);
  nor (_07267_, _07266_, _07257_);
  and (_07268_, _07267_, \oc8051_golden_model_1.ACC [4]);
  nor (_07269_, _07267_, _06867_);
  and (_07270_, _07267_, _06867_);
  nor (_07271_, _07270_, _07269_);
  and (_07272_, _06155_, _06153_);
  and (_07273_, _07272_, \oc8051_golden_model_1.PSW [7]);
  nor (_07274_, _07273_, _06154_);
  nor (_07275_, _07274_, _07265_);
  and (_07276_, _07275_, \oc8051_golden_model_1.ACC [3]);
  nor (_07277_, _07275_, _02564_);
  and (_07278_, _07275_, _02564_);
  nor (_07279_, _07278_, _07277_);
  nor (_07280_, _07264_, _06155_);
  nor (_07281_, _07280_, _07273_);
  and (_07282_, _07281_, \oc8051_golden_model_1.ACC [2]);
  nor (_07283_, _07281_, _06964_);
  and (_07284_, _07281_, _06964_);
  nor (_07285_, _07284_, _07283_);
  and (_07286_, _06152_, \oc8051_golden_model_1.PSW [7]);
  nor (_07287_, _07286_, _06151_);
  nor (_07288_, _07287_, _07264_);
  and (_07289_, _07288_, \oc8051_golden_model_1.ACC [1]);
  and (_07290_, _07288_, _02551_);
  nor (_07291_, _07288_, _02551_);
  nor (_07292_, _07291_, _07290_);
  not (_07293_, \oc8051_golden_model_1.PSW [7]);
  and (_07294_, _05940_, _07293_);
  nor (_07295_, _07294_, _07286_);
  and (_07296_, _07295_, \oc8051_golden_model_1.ACC [0]);
  not (_07297_, _07296_);
  nor (_07298_, _07297_, _07292_);
  nor (_07299_, _07298_, _07289_);
  nor (_07300_, _07299_, _07285_);
  nor (_07301_, _07300_, _07282_);
  nor (_07302_, _07301_, _07279_);
  nor (_07303_, _07302_, _07276_);
  nor (_07304_, _07303_, _07271_);
  nor (_07305_, _07304_, _07268_);
  nor (_07306_, _07305_, _07263_);
  nor (_07307_, _07306_, _07260_);
  nor (_07308_, _07307_, _07255_);
  nor (_07309_, _07308_, _07252_);
  nor (_07310_, _07309_, _07248_);
  and (_07311_, _07309_, _07248_);
  nor (_07312_, _07311_, _07310_);
  or (_07313_, _07312_, _07241_);
  and (_07314_, _07313_, _03134_);
  and (_07315_, _02854_, _02967_);
  not (_07316_, _07315_);
  not (_07317_, _03543_);
  not (_07318_, _03726_);
  or (_07319_, _03309_, _02528_);
  and (_07320_, _07319_, _07318_);
  and (_07321_, _07320_, _07317_);
  and (_07322_, _07321_, _07316_);
  and (_07323_, _05243_, \oc8051_golden_model_1.PSW [7]);
  and (_07324_, _07323_, _04770_);
  nor (_07325_, _07324_, _05248_);
  and (_07326_, _07324_, _05248_);
  nor (_07327_, _07326_, _07325_);
  and (_07328_, _07327_, \oc8051_golden_model_1.ACC [7]);
  nor (_07329_, _07327_, \oc8051_golden_model_1.ACC [7]);
  nor (_07330_, _07329_, _07328_);
  nor (_07331_, _07323_, _04770_);
  nor (_07332_, _07331_, _07324_);
  and (_07333_, _07332_, \oc8051_golden_model_1.ACC [6]);
  nor (_07334_, _07332_, _06806_);
  and (_07335_, _07332_, _06806_);
  nor (_07336_, _07335_, _07334_);
  and (_07337_, _05242_, \oc8051_golden_model_1.PSW [7]);
  nor (_07338_, _07337_, _04877_);
  nor (_07339_, _07338_, _07323_);
  and (_07340_, _07339_, \oc8051_golden_model_1.ACC [5]);
  nor (_07341_, _07339_, _06861_);
  and (_07342_, _07339_, _06861_);
  nor (_07343_, _07342_, _07341_);
  and (_07344_, _05239_, \oc8051_golden_model_1.PSW [7]);
  and (_07345_, _07344_, _05240_);
  nor (_07346_, _07345_, _04982_);
  nor (_07347_, _07346_, _07337_);
  and (_07348_, _07347_, \oc8051_golden_model_1.ACC [4]);
  nor (_07349_, _07347_, _06867_);
  and (_07350_, _07347_, _06867_);
  nor (_07351_, _07350_, _07349_);
  and (_07352_, _05239_, _04435_);
  and (_07353_, _07352_, \oc8051_golden_model_1.PSW [7]);
  nor (_07354_, _07353_, _04241_);
  nor (_07355_, _07354_, _07345_);
  and (_07356_, _07355_, \oc8051_golden_model_1.ACC [3]);
  nor (_07357_, _07355_, _02564_);
  and (_07358_, _07355_, _02564_);
  nor (_07359_, _07358_, _07357_);
  nor (_07360_, _07344_, _04435_);
  nor (_07361_, _07360_, _07353_);
  and (_07362_, _07361_, \oc8051_golden_model_1.ACC [2]);
  nor (_07363_, _07361_, _06964_);
  and (_07364_, _07361_, _06964_);
  nor (_07365_, _07364_, _07363_);
  and (_07366_, _03808_, \oc8051_golden_model_1.PSW [7]);
  nor (_07367_, _07366_, _04000_);
  nor (_07368_, _07367_, _07344_);
  and (_07369_, _07368_, \oc8051_golden_model_1.ACC [1]);
  and (_07370_, _07368_, _02551_);
  nor (_07371_, _07368_, _02551_);
  nor (_07372_, _07371_, _07370_);
  nor (_07373_, _03808_, \oc8051_golden_model_1.PSW [7]);
  nor (_07374_, _07373_, _07366_);
  and (_07375_, _07374_, \oc8051_golden_model_1.ACC [0]);
  not (_07376_, _07375_);
  nor (_07377_, _07376_, _07372_);
  nor (_07378_, _07377_, _07369_);
  nor (_07379_, _07378_, _07365_);
  nor (_07380_, _07379_, _07362_);
  nor (_07381_, _07380_, _07359_);
  nor (_07382_, _07381_, _07356_);
  nor (_07383_, _07382_, _07351_);
  nor (_07384_, _07383_, _07348_);
  nor (_07385_, _07384_, _07343_);
  nor (_07386_, _07385_, _07340_);
  nor (_07387_, _07386_, _07336_);
  nor (_07388_, _07387_, _07333_);
  nor (_07389_, _07388_, _07330_);
  and (_07390_, _07388_, _07330_);
  nor (_07391_, _07390_, _07389_);
  and (_07392_, _07391_, _07316_);
  or (_07393_, _07392_, _07322_);
  and (_07394_, _02951_, _02969_);
  not (_07395_, _07394_);
  not (_07396_, _03138_);
  or (_07397_, _05772_, _07396_);
  and (_07398_, _07397_, _07395_);
  and (_07399_, _02951_, _02508_);
  nor (_07400_, _04706_, _05771_);
  and (_07401_, _04706_, _04604_);
  nor (_07402_, _07401_, _07400_);
  nand (_07403_, _07402_, _06770_);
  and (_07404_, _02951_, _02580_);
  not (_07405_, _07404_);
  not (_07406_, _04796_);
  not (_07407_, _04784_);
  and (_07408_, _04813_, _07407_);
  and (_07409_, _07408_, _07406_);
  and (_07410_, _04641_, \oc8051_golden_model_1.P2INREG [6]);
  and (_07411_, _04645_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_07412_, _07411_, _07410_);
  and (_07413_, _04628_, \oc8051_golden_model_1.P0INREG [6]);
  and (_07414_, _04634_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_07415_, _07414_, _07413_);
  and (_07416_, _07415_, _07412_);
  nor (_07417_, _04797_, _04800_);
  and (_07418_, _07417_, _04808_);
  and (_07419_, _07418_, _07416_);
  and (_07420_, _07419_, _07409_);
  and (_07421_, _04805_, _04794_);
  and (_07422_, _07421_, _04780_);
  and (_07423_, _07422_, _07420_);
  and (_07424_, _07423_, _04771_);
  not (_07425_, _07424_);
  not (_07426_, _05051_);
  nor (_07427_, _05055_, _05052_);
  and (_07428_, _07427_, _05063_);
  and (_07429_, _07428_, _07426_);
  and (_07430_, _07429_, _05075_);
  and (_07431_, _05060_, _05038_);
  and (_07432_, _04641_, \oc8051_golden_model_1.P2INREG [3]);
  and (_07433_, _04645_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_07434_, _07433_, _07432_);
  and (_07435_, _04634_, \oc8051_golden_model_1.P1INREG [3]);
  and (_07436_, _04628_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_07437_, _07436_, _07435_);
  and (_07438_, _07437_, _07434_);
  and (_07439_, _07438_, _05050_);
  and (_07440_, _07439_, _07431_);
  and (_07441_, _07440_, _07430_);
  and (_07442_, _07441_, _05032_);
  not (_07443_, _07442_);
  and (_07444_, _04641_, \oc8051_golden_model_1.P2INREG [2]);
  and (_07445_, _04645_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_07446_, _07445_, _07444_);
  and (_07447_, _04628_, \oc8051_golden_model_1.P0INREG [2]);
  and (_07448_, _04634_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_07449_, _07448_, _07447_);
  and (_07450_, _07449_, _07446_);
  and (_07451_, _07450_, _05086_);
  and (_07452_, _07451_, _05127_);
  and (_07453_, _07452_, _05080_);
  not (_07454_, _07453_);
  and (_07455_, _04628_, \oc8051_golden_model_1.P0INREG [1]);
  not (_07456_, _07455_);
  and (_07457_, _04634_, \oc8051_golden_model_1.P1INREG [1]);
  not (_07458_, _07457_);
  and (_07459_, _04641_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07460_, _04645_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_07461_, _07460_, _07459_);
  and (_07462_, _07461_, _07458_);
  and (_07463_, _07462_, _05167_);
  and (_07464_, _07463_, _07456_);
  and (_07465_, _07464_, _05158_);
  and (_07466_, _07465_, _05148_);
  and (_07467_, _07466_, _05131_);
  not (_07468_, _07467_);
  and (_07469_, _04628_, \oc8051_golden_model_1.P0INREG [0]);
  not (_07470_, _07469_);
  and (_07471_, _04634_, \oc8051_golden_model_1.P1INREG [0]);
  not (_07472_, _07471_);
  and (_07473_, _04641_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07474_, _04645_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07475_, _07474_, _07473_);
  and (_07476_, _07475_, _07472_);
  and (_07477_, _07476_, _05215_);
  and (_07478_, _07477_, _07470_);
  and (_07479_, _07478_, _05206_);
  and (_07480_, _07479_, _05196_);
  and (_07481_, _07480_, _05179_);
  nor (_07482_, _07481_, _07293_);
  and (_07483_, _07482_, _07468_);
  and (_07484_, _07483_, _07454_);
  and (_07485_, _07484_, _07443_);
  not (_07486_, _04896_);
  nor (_07487_, _04900_, _04897_);
  and (_07488_, _04908_, _07487_);
  and (_07489_, _07488_, _07486_);
  and (_07490_, _07489_, _04920_);
  not (_07491_, _04885_);
  and (_07492_, _07491_, _04905_);
  and (_07493_, _07492_, _04881_);
  and (_07494_, _04641_, \oc8051_golden_model_1.P2INREG [5]);
  and (_07495_, _04645_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_07496_, _07495_, _07494_);
  and (_07497_, _04634_, \oc8051_golden_model_1.P1INREG [5]);
  and (_07498_, _04628_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_07499_, _07498_, _07497_);
  and (_07500_, _07499_, _07496_);
  and (_07501_, _07500_, _04895_);
  and (_07502_, _07501_, _07493_);
  and (_07503_, _07502_, _07490_);
  and (_07504_, _07503_, _04878_);
  and (_07505_, _04628_, \oc8051_golden_model_1.P0INREG [4]);
  not (_07506_, _07505_);
  and (_07507_, _04634_, \oc8051_golden_model_1.P1INREG [4]);
  not (_07508_, _07507_);
  and (_07509_, _04641_, \oc8051_golden_model_1.P2INREG [4]);
  and (_07510_, _04645_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_07511_, _07510_, _07509_);
  and (_07512_, _07511_, _07508_);
  and (_07513_, _07512_, _05017_);
  and (_07514_, _07513_, _07506_);
  and (_07515_, _07514_, _05010_);
  and (_07516_, _07515_, _05000_);
  and (_07517_, _07516_, _04983_);
  nor (_07518_, _07517_, _07504_);
  and (_07519_, _07518_, _07485_);
  and (_07520_, _07519_, _07425_);
  nor (_07521_, _07520_, _05497_);
  and (_07522_, _07520_, _05497_);
  nor (_07523_, _07522_, _07521_);
  and (_07524_, _07523_, \oc8051_golden_model_1.ACC [7]);
  nor (_07525_, _07523_, \oc8051_golden_model_1.ACC [7]);
  nor (_07526_, _07525_, _07524_);
  not (_07527_, _07526_);
  nor (_07528_, _07519_, _07425_);
  nor (_07529_, _07528_, _07520_);
  nor (_07530_, _07529_, _06806_);
  and (_07531_, _07529_, _06806_);
  not (_07532_, _07504_);
  not (_07533_, _07517_);
  and (_07534_, _07485_, _07533_);
  nor (_07535_, _07534_, _07532_);
  nor (_07536_, _07535_, _07519_);
  nor (_07537_, _07536_, _06861_);
  and (_07538_, _07536_, _06861_);
  nor (_07539_, _07538_, _07537_);
  nor (_07540_, _07485_, _07533_);
  nor (_07541_, _07540_, _07534_);
  nor (_07542_, _07541_, _06867_);
  and (_07543_, _07541_, _06867_);
  nor (_07544_, _07543_, _07542_);
  and (_07545_, _07544_, _07539_);
  not (_07546_, _07545_);
  nor (_07547_, _07484_, _07443_);
  nor (_07548_, _07547_, _07485_);
  nor (_07549_, _07548_, _02564_);
  and (_07550_, _07548_, _02564_);
  nor (_07551_, _07550_, _07549_);
  nor (_07552_, _07483_, _07454_);
  nor (_07553_, _07552_, _07484_);
  nor (_07554_, _07553_, _06964_);
  and (_07555_, _07553_, _06964_);
  nor (_07556_, _07555_, _07554_);
  and (_07557_, _07556_, _07551_);
  not (_07558_, _07557_);
  nor (_07559_, _07482_, _07468_);
  nor (_07560_, _07559_, _07483_);
  and (_07561_, _07560_, _02551_);
  nor (_07562_, _07560_, _02551_);
  and (_07563_, _07481_, _07293_);
  nor (_07564_, _07563_, _07482_);
  nor (_07565_, _07564_, _02667_);
  nor (_07566_, _07565_, _07562_);
  nor (_07567_, _07566_, _07561_);
  nor (_07568_, _07567_, _07558_);
  nor (_07569_, _07555_, _07550_);
  nor (_07570_, _07569_, _07549_);
  nor (_07571_, _07570_, _07568_);
  and (_07572_, _07564_, _02667_);
  nor (_07573_, _07565_, _07572_);
  nor (_07574_, _07467_, \oc8051_golden_model_1.ACC [1]);
  and (_07575_, _07467_, \oc8051_golden_model_1.ACC [1]);
  nor (_07576_, _07575_, _07574_);
  and (_07577_, \oc8051_golden_model_1.PSW [7], _02667_);
  and (_07578_, _07293_, \oc8051_golden_model_1.ACC [0]);
  nor (_07579_, _07578_, _07481_);
  nor (_07580_, _07579_, _07577_);
  and (_07581_, _07580_, _07576_);
  nor (_07582_, _07580_, _07576_);
  or (_07583_, _07582_, _07581_);
  nand (_07584_, _07583_, _07573_);
  nor (_07585_, _07584_, _07558_);
  nor (_07586_, _07585_, _07571_);
  nor (_07587_, _07586_, _07546_);
  not (_07588_, _07587_);
  nor (_07589_, _07542_, _07537_);
  or (_07590_, _07589_, _07538_);
  and (_07591_, _07590_, _07588_);
  nor (_07592_, _07591_, _07531_);
  or (_07593_, _07592_, _07530_);
  and (_07594_, _07593_, _07527_);
  nor (_07595_, _07593_, _07527_);
  nor (_07596_, _07595_, _07594_);
  nand (_07597_, _07596_, _03106_);
  and (_07598_, _07597_, _07405_);
  not (_07599_, _07248_);
  nor (_07600_, _07269_, _07261_);
  nor (_07601_, _07600_, _07262_);
  and (_07602_, _07271_, _07263_);
  not (_07603_, _07602_);
  and (_07604_, _07285_, _07279_);
  nor (_07605_, _07295_, _02667_);
  nor (_07606_, _07605_, _07291_);
  or (_07607_, _07606_, _07290_);
  and (_07608_, _07607_, _07604_);
  not (_07609_, _07608_);
  and (_07610_, _07284_, _07279_);
  nor (_07611_, _07610_, _07278_);
  and (_07612_, _07611_, _07609_);
  and (_07613_, _07295_, _02667_);
  nor (_07614_, _07605_, _07613_);
  and (_07615_, _07614_, _07292_);
  and (_07616_, _07615_, _07604_);
  nor (_07617_, _07616_, _07612_);
  nor (_07618_, _07617_, _07603_);
  nor (_07619_, _07618_, _07601_);
  nor (_07620_, _07619_, _07254_);
  or (_07621_, _07620_, _07253_);
  and (_07622_, _07621_, _07599_);
  nor (_07623_, _07621_, _07599_);
  or (_07624_, _07623_, _07622_);
  and (_07625_, _07624_, _03434_);
  not (_07626_, _03434_);
  not (_07627_, _04024_);
  and (_07628_, _07627_, _03393_);
  or (_07629_, _07628_, _04604_);
  nor (_07630_, _05497_, _03387_);
  not (_07631_, _03363_);
  or (_07632_, _05462_, _07631_);
  nor (_07633_, _02615_, _02576_);
  and (_07634_, _07633_, _04604_);
  not (_07635_, _07633_);
  and (_07636_, _02951_, _02884_);
  and (_07637_, _07636_, _05771_);
  nor (_07638_, _07636_, _05771_);
  or (_07639_, _07638_, _07637_);
  and (_07640_, _07639_, _07635_);
  or (_07641_, _07640_, _03363_);
  or (_07642_, _07641_, _07634_);
  and (_07643_, _07642_, _03387_);
  and (_07644_, _07643_, _07632_);
  or (_07645_, _07644_, _07630_);
  and (_07646_, _02951_, _03071_);
  nor (_07647_, _07646_, _02974_);
  and (_07648_, _07647_, _07645_);
  and (_07649_, _02951_, _02879_);
  and (_07650_, _05474_, _04706_);
  nor (_07651_, _07650_, _07400_);
  nor (_07652_, _07651_, _03810_);
  or (_07653_, _07652_, _07649_);
  or (_07654_, _07653_, _07648_);
  nor (_07655_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07656_, _07655_, _02564_);
  and (_07657_, _07656_, _06826_);
  and (_07658_, _07657_, \oc8051_golden_model_1.ACC [6]);
  and (_07659_, _07658_, \oc8051_golden_model_1.ACC [7]);
  nor (_07660_, _07658_, \oc8051_golden_model_1.ACC [7]);
  nor (_07661_, _07660_, _07659_);
  and (_07662_, _07656_, \oc8051_golden_model_1.ACC [4]);
  nor (_07663_, _07662_, \oc8051_golden_model_1.ACC [5]);
  nor (_07664_, _07663_, _07657_);
  nor (_07665_, _07657_, \oc8051_golden_model_1.ACC [6]);
  nor (_07666_, _07665_, _07658_);
  nor (_07667_, _07666_, _07664_);
  not (_07668_, _07667_);
  and (_07669_, _07668_, _07661_);
  nor (_07670_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_07671_, _07670_, _07667_);
  nor (_07672_, _07671_, _07661_);
  nor (_07673_, _07672_, _07669_);
  not (_07674_, _07673_);
  nand (_07675_, _07674_, _07649_);
  and (_07676_, _07675_, _03076_);
  and (_07677_, _07676_, _07654_);
  nor (_07678_, _05325_, _05771_);
  and (_07679_, _05360_, _05325_);
  nor (_07680_, _07679_, _07678_);
  nor (_07681_, _07680_, _02881_);
  not (_07682_, _07628_);
  nor (_07683_, _07402_, _03336_);
  or (_07684_, _07683_, _07682_);
  or (_07685_, _07684_, _07681_);
  or (_07686_, _07685_, _07677_);
  and (_07687_, _07686_, _07629_);
  or (_07688_, _07687_, _03399_);
  or (_07689_, _05462_, _03840_);
  and (_07690_, _07689_, _03084_);
  and (_07691_, _07690_, _07688_);
  and (_07692_, _02951_, _02874_);
  nor (_07693_, _05497_, _03084_);
  or (_07694_, _07693_, _07692_);
  or (_07695_, _07694_, _07691_);
  nand (_07696_, _07692_, _02564_);
  and (_07697_, _07696_, _07695_);
  or (_07698_, _07697_, _02876_);
  and (_07699_, _05356_, _05325_);
  nor (_07700_, _07699_, _07678_);
  nand (_07701_, _07700_, _02876_);
  and (_07702_, _07701_, _02870_);
  and (_07703_, _07702_, _07698_);
  and (_07704_, _07679_, _05502_);
  nor (_07705_, _07704_, _07678_);
  nor (_07706_, _07705_, _02870_);
  or (_07707_, _07706_, _06247_);
  or (_07708_, _07707_, _07703_);
  nor (_07709_, _06726_, _06724_);
  nor (_07710_, _07709_, _06727_);
  or (_07711_, _07710_, _06253_);
  not (_07712_, _03433_);
  and (_07713_, _02848_, _02580_);
  not (_07714_, _07713_);
  nor (_07715_, _03709_, _03438_);
  nand (_07716_, _07715_, _07714_);
  nor (_07717_, _07716_, _03711_);
  and (_07718_, _07717_, _07712_);
  and (_07719_, _07718_, _07711_);
  and (_07720_, _07719_, _07708_);
  not (_07721_, _07330_);
  nor (_07722_, _07349_, _07341_);
  nor (_07723_, _07722_, _07342_);
  and (_07724_, _07351_, _07343_);
  not (_07725_, _07724_);
  and (_07726_, _07365_, _07359_);
  nor (_07727_, _07374_, _02667_);
  nor (_07728_, _07727_, _07371_);
  nor (_07729_, _07728_, _07370_);
  not (_07730_, _07729_);
  and (_07731_, _07730_, _07726_);
  not (_07732_, _07731_);
  and (_07733_, _07364_, _07359_);
  nor (_07734_, _07733_, _07358_);
  and (_07735_, _07734_, _07732_);
  and (_07736_, _07374_, _02667_);
  nor (_07737_, _07727_, _07736_);
  and (_07738_, _07737_, _07372_);
  and (_07739_, _07738_, _07726_);
  nor (_07740_, _07739_, _07735_);
  nor (_07741_, _07740_, _07725_);
  nor (_07742_, _07741_, _07723_);
  nor (_07743_, _07742_, _07335_);
  or (_07744_, _07743_, _07334_);
  and (_07745_, _07744_, _07721_);
  nor (_07746_, _07744_, _07721_);
  nor (_07747_, _07746_, _07745_);
  nor (_07748_, _07747_, _07718_);
  or (_07749_, _07748_, _07720_);
  and (_07750_, _07749_, _07626_);
  or (_07751_, _07750_, _03106_);
  or (_07752_, _07751_, _07625_);
  and (_07753_, _07752_, _07598_);
  and (_07754_, _04653_, \oc8051_golden_model_1.PSW [7]);
  and (_07755_, _07754_, _04658_);
  and (_07756_, _07755_, _04643_);
  and (_07757_, _07756_, _04344_);
  nor (_07758_, _07757_, _04551_);
  and (_07759_, _07756_, _02928_);
  nor (_07760_, _07759_, _07758_);
  and (_07761_, _07760_, \oc8051_golden_model_1.ACC [7]);
  nor (_07762_, _07760_, \oc8051_golden_model_1.ACC [7]);
  nor (_07763_, _07762_, _07761_);
  not (_07764_, _07763_);
  nor (_07765_, _07756_, _04344_);
  nor (_07766_, _07765_, _07757_);
  nor (_07767_, _07766_, _06806_);
  and (_07768_, _07766_, _06806_);
  nor (_07769_, _07767_, _07768_);
  and (_07770_, _07755_, _04631_);
  nor (_07771_, _07770_, _04638_);
  nor (_07772_, _07771_, _07756_);
  nor (_07773_, _07772_, _06861_);
  and (_07774_, _07772_, _06861_);
  nor (_07775_, _07774_, _07773_);
  nor (_07776_, _07755_, _04631_);
  nor (_07777_, _07776_, _07770_);
  nor (_07778_, _07777_, _06867_);
  and (_07779_, _07777_, _06867_);
  nor (_07780_, _07779_, _07778_);
  and (_07781_, _07780_, _07775_);
  nor (_07782_, _05529_, _02929_);
  nor (_07783_, _07782_, _07755_);
  nor (_07784_, _07783_, _02564_);
  and (_07785_, _07783_, _02564_);
  nor (_07786_, _07785_, _07784_);
  nor (_07787_, _07754_, _04361_);
  nor (_07788_, _07787_, _05529_);
  nor (_07789_, _07788_, _06964_);
  and (_07790_, _07788_, _06964_);
  nor (_07791_, _07790_, _07789_);
  and (_07792_, _07791_, _07786_);
  and (_07793_, _02835_, \oc8051_golden_model_1.PSW [7]);
  nor (_07794_, _07793_, _03936_);
  nor (_07795_, _07794_, _07754_);
  and (_07796_, _07795_, _02551_);
  nor (_07797_, _07795_, _02551_);
  nor (_07798_, _07797_, _07796_);
  and (_07799_, _02835_, _07293_);
  and (_07800_, _02837_, \oc8051_golden_model_1.PSW [7]);
  nor (_07801_, _07800_, _07799_);
  nor (_07802_, _07801_, _02667_);
  and (_07803_, _07801_, _02667_);
  or (_07804_, _07803_, _07802_);
  and (_07805_, _07804_, _07798_);
  and (_07806_, _07805_, _07792_);
  and (_07807_, _07801_, \oc8051_golden_model_1.ACC [0]);
  not (_07808_, _07807_);
  nor (_07809_, _07808_, _07796_);
  nor (_07810_, _07809_, _07797_);
  and (_07811_, _07810_, _07792_);
  not (_07812_, _07811_);
  and (_07813_, _07790_, _07786_);
  nor (_07814_, _07813_, _07785_);
  and (_07815_, _07814_, _07812_);
  nor (_07816_, _07815_, _07806_);
  not (_07817_, _07816_);
  and (_07818_, _07817_, _07781_);
  nor (_07819_, _07778_, _07773_);
  nor (_07820_, _07819_, _07774_);
  or (_07821_, _07820_, _07818_);
  and (_07822_, _07821_, _07769_);
  or (_07823_, _07822_, _07767_);
  and (_07824_, _07823_, _07764_);
  nor (_07825_, _07823_, _07764_);
  or (_07826_, _07825_, _07824_);
  and (_07827_, _07826_, _07404_);
  or (_07828_, _07827_, _02583_);
  or (_07829_, _07828_, _07753_);
  or (_07830_, _02763_, _02605_);
  and (_07831_, _07830_, _02864_);
  and (_07832_, _07831_, _07829_);
  not (_07833_, _05325_);
  nor (_07834_, _05530_, _07833_);
  nor (_07835_, _07834_, _07678_);
  nor (_07836_, _07835_, _02864_);
  or (_07837_, _07836_, _06770_);
  or (_07838_, _07837_, _07832_);
  and (_07839_, _07838_, _07403_);
  or (_07840_, _07839_, _02853_);
  and (_07841_, _04706_, _05462_);
  or (_07842_, _07841_, _07400_);
  or (_07843_, _07842_, _05540_);
  and (_07844_, _07843_, _02838_);
  and (_07845_, _07844_, _07840_);
  not (_07846_, _04706_);
  nor (_07847_, _05744_, _07846_);
  nor (_07848_, _07847_, _07400_);
  nor (_07849_, _07848_, _02838_);
  or (_07850_, _07849_, _06784_);
  or (_07851_, _07850_, _07845_);
  not (_07852_, _06803_);
  nand (_07853_, _07852_, _06784_);
  and (_07854_, _07853_, _07851_);
  and (_07855_, _07854_, _02635_);
  and (_07856_, _02763_, _02546_);
  or (_07857_, _07856_, _02802_);
  or (_07858_, _07857_, _07855_);
  and (_07859_, _02951_, _02513_);
  not (_07860_, _07859_);
  and (_07861_, _05661_, _04706_);
  nor (_07862_, _07861_, _07400_);
  nand (_07863_, _07862_, _02802_);
  and (_07864_, _07863_, _07860_);
  and (_07865_, _07864_, _07858_);
  and (_07866_, _07859_, _02763_);
  and (_07867_, _02947_, _02508_);
  nor (_07868_, _07867_, _03503_);
  and (_07869_, _02848_, _02508_);
  not (_07870_, _07869_);
  and (_07871_, _07870_, _07868_);
  and (_07872_, _04009_, _02508_);
  nor (_07873_, _07872_, _03509_);
  and (_07874_, _07873_, _03500_);
  and (_07875_, _07874_, _07871_);
  not (_07876_, _07875_);
  or (_07877_, _07876_, _07866_);
  or (_07878_, _07877_, _07865_);
  and (_07879_, _02852_, _02508_);
  not (_07880_, _07879_);
  or (_07881_, _07875_, _07191_);
  and (_07882_, _07881_, _07880_);
  and (_07883_, _07882_, _07878_);
  nor (_07884_, _05462_, \oc8051_golden_model_1.ACC [7]);
  and (_07885_, _05462_, \oc8051_golden_model_1.ACC [7]);
  nor (_07886_, _07885_, _07884_);
  and (_07887_, _07886_, _07879_);
  or (_07888_, _07887_, _03129_);
  or (_07889_, _07888_, _07883_);
  not (_07890_, _03129_);
  or (_07891_, _05774_, _07890_);
  and (_07892_, _07891_, _07889_);
  or (_07893_, _07892_, _07399_);
  nor (_07894_, _02763_, \oc8051_golden_model_1.ACC [7]);
  and (_07895_, _02763_, \oc8051_golden_model_1.ACC [7]);
  nor (_07896_, _07895_, _07894_);
  not (_07897_, _07399_);
  or (_07898_, _07897_, _07896_);
  and (_07899_, _07898_, _07893_);
  or (_07900_, _07899_, _02980_);
  and (_07901_, _05766_, _04706_);
  nor (_07902_, _07901_, _07400_);
  nand (_07903_, _07902_, _02980_);
  and (_07904_, _07903_, _03128_);
  and (_07905_, _07904_, _07900_);
  and (_07906_, _07400_, _03127_);
  or (_07907_, _02531_, _02576_);
  not (_07908_, _07907_);
  or (_07909_, _07908_, _07906_);
  or (_07910_, _07909_, _07905_);
  and (_07911_, _02852_, _02969_);
  not (_07912_, _07911_);
  or (_07913_, _07907_, _07190_);
  and (_07914_, _07913_, _07912_);
  and (_07915_, _07914_, _07910_);
  and (_07916_, _07885_, _07911_);
  or (_07917_, _07916_, _03138_);
  or (_07918_, _07917_, _07915_);
  and (_07919_, _07918_, _07398_);
  and (_07920_, _07895_, _07394_);
  or (_07921_, _07920_, _07919_);
  and (_07922_, _07921_, _03883_);
  or (_07923_, _07862_, _05773_);
  nor (_07924_, _07923_, _03883_);
  nor (_07925_, _03309_, _02534_);
  nor (_07926_, _07925_, _03732_);
  not (_07927_, _07926_);
  or (_07928_, _07927_, _07924_);
  or (_07929_, _07928_, _07922_);
  and (_07930_, _02854_, _02964_);
  not (_07931_, _07930_);
  nand (_07932_, _07927_, _07189_);
  and (_07933_, _07932_, _07931_);
  and (_07934_, _07933_, _07929_);
  and (_07935_, _02852_, _02964_);
  nor (_07936_, _07189_, _07931_);
  or (_07937_, _07936_, _07935_);
  or (_07938_, _07937_, _07934_);
  nand (_07939_, _07884_, _07935_);
  and (_07940_, _07939_, _03122_);
  and (_07941_, _07940_, _07938_);
  and (_07942_, _02951_, _02964_);
  nor (_07943_, _07942_, _03121_);
  not (_07944_, _07943_);
  not (_07945_, _07942_);
  nand (_07946_, _07945_, _05773_);
  and (_07947_, _07946_, _07944_);
  or (_07948_, _07947_, _07941_);
  nand (_07949_, _07942_, _07894_);
  and (_07950_, _07949_, _05783_);
  and (_07951_, _07950_, _07948_);
  nor (_07952_, _05765_, _07846_);
  nor (_07953_, _07952_, _07400_);
  or (_07954_, _07953_, _05783_);
  nand (_07955_, _07954_, _07321_);
  or (_07956_, _07955_, _07951_);
  and (_07957_, _07956_, _07393_);
  and (_07958_, _07391_, _07315_);
  or (_07959_, _07958_, _07240_);
  or (_07960_, _07959_, _07957_);
  and (_07961_, _07960_, _07314_);
  and (_07962_, _02951_, _02967_);
  and (_07963_, _07529_, \oc8051_golden_model_1.ACC [6]);
  nor (_07964_, _07530_, _07531_);
  and (_07965_, _07536_, \oc8051_golden_model_1.ACC [5]);
  and (_07966_, _07541_, \oc8051_golden_model_1.ACC [4]);
  and (_07967_, _07548_, \oc8051_golden_model_1.ACC [3]);
  and (_07968_, _07553_, \oc8051_golden_model_1.ACC [2]);
  and (_07969_, _07560_, \oc8051_golden_model_1.ACC [1]);
  nor (_07970_, _07562_, _07561_);
  and (_07971_, _07564_, \oc8051_golden_model_1.ACC [0]);
  not (_07972_, _07971_);
  nor (_07973_, _07972_, _07970_);
  nor (_07974_, _07973_, _07969_);
  nor (_07975_, _07974_, _07556_);
  nor (_07976_, _07975_, _07968_);
  nor (_07977_, _07976_, _07551_);
  nor (_07978_, _07977_, _07967_);
  nor (_07979_, _07978_, _07544_);
  nor (_07980_, _07979_, _07966_);
  nor (_07981_, _07980_, _07539_);
  nor (_07982_, _07981_, _07965_);
  nor (_07983_, _07982_, _07964_);
  nor (_07984_, _07983_, _07963_);
  nor (_07985_, _07984_, _07526_);
  and (_07986_, _07984_, _07526_);
  nor (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _03133_);
  or (_07989_, _07988_, _07962_);
  or (_07990_, _07989_, _07961_);
  and (_07991_, _02545_, _02967_);
  not (_07992_, _07991_);
  not (_07993_, _07962_);
  and (_07994_, _07766_, \oc8051_golden_model_1.ACC [6]);
  and (_07995_, _07772_, \oc8051_golden_model_1.ACC [5]);
  and (_07996_, _07777_, \oc8051_golden_model_1.ACC [4]);
  and (_07997_, _07783_, \oc8051_golden_model_1.ACC [3]);
  and (_07998_, _07788_, \oc8051_golden_model_1.ACC [2]);
  and (_07999_, _07795_, \oc8051_golden_model_1.ACC [1]);
  not (_08000_, _07802_);
  nor (_08001_, _08000_, _07798_);
  nor (_08002_, _08001_, _07999_);
  nor (_08003_, _08002_, _07791_);
  nor (_08004_, _08003_, _07998_);
  nor (_08005_, _08004_, _07786_);
  nor (_08006_, _08005_, _07997_);
  nor (_08007_, _08006_, _07780_);
  nor (_08008_, _08007_, _07996_);
  nor (_08009_, _08008_, _07775_);
  nor (_08010_, _08009_, _07995_);
  nor (_08011_, _08010_, _07769_);
  nor (_08012_, _08011_, _07994_);
  nor (_08013_, _08012_, _07763_);
  and (_08014_, _08012_, _07763_);
  nor (_08015_, _08014_, _08013_);
  or (_08016_, _08015_, _07993_);
  and (_08017_, _08016_, _07992_);
  and (_08018_, _08017_, _07990_);
  nand (_08019_, _07991_, \oc8051_golden_model_1.ACC [6]);
  nand (_08020_, _08019_, _07238_);
  or (_08021_, _08020_, _08018_);
  and (_08022_, _08021_, _07239_);
  or (_08023_, _08022_, _07188_);
  not (_08024_, _07188_);
  and (_08025_, _05849_, \oc8051_golden_model_1.ACC [6]);
  nor (_08026_, _05849_, \oc8051_golden_model_1.ACC [6]);
  nor (_08027_, _08025_, _08026_);
  and (_08028_, _06158_, \oc8051_golden_model_1.ACC [5]);
  and (_08029_, _06078_, _06861_);
  nor (_08030_, _08029_, _08028_);
  not (_08031_, _08030_);
  and (_08032_, _06159_, \oc8051_golden_model_1.ACC [4]);
  and (_08033_, _06123_, _06867_);
  nor (_08034_, _08032_, _08033_);
  and (_08035_, _05986_, _02564_);
  not (_08036_, _08035_);
  and (_08037_, _06154_, \oc8051_golden_model_1.ACC [3]);
  not (_08038_, _08037_);
  and (_08039_, _06155_, \oc8051_golden_model_1.ACC [2]);
  and (_08040_, _06031_, _06964_);
  nor (_08041_, _08039_, _08040_);
  not (_08042_, _08041_);
  and (_08043_, _06151_, \oc8051_golden_model_1.ACC [1]);
  and (_08044_, _05895_, _02551_);
  nor (_08045_, _08043_, _08044_);
  and (_08046_, _06152_, \oc8051_golden_model_1.ACC [0]);
  and (_08047_, _08046_, _08045_);
  nor (_08048_, _08047_, _08043_);
  nor (_08049_, _08048_, _08042_);
  nor (_08050_, _08049_, _08039_);
  nand (_08051_, _08050_, _08038_);
  and (_08052_, _08051_, _08036_);
  and (_08053_, _08052_, _08034_);
  nor (_08054_, _08053_, _08032_);
  nor (_08055_, _08054_, _08031_);
  or (_08056_, _08055_, _08028_);
  and (_08057_, _08056_, _08027_);
  nor (_08058_, _08057_, _08025_);
  nor (_08059_, _08058_, _07886_);
  and (_08060_, _08058_, _07886_);
  or (_08061_, _08060_, _08059_);
  or (_08062_, _08061_, _08024_);
  and (_08063_, _08062_, _02896_);
  and (_08064_, _08063_, _08023_);
  and (_08065_, _02951_, _02891_);
  nor (_08066_, _08065_, _02894_);
  not (_08067_, _08066_);
  and (_08068_, _05497_, _05771_);
  nor (_08069_, _05497_, _05771_);
  nor (_08070_, _08069_, _08068_);
  nor (_08071_, _07424_, _06806_);
  and (_08072_, _07424_, \oc8051_golden_model_1.ACC [6]);
  nor (_08073_, _07424_, \oc8051_golden_model_1.ACC [6]);
  nor (_08074_, _08073_, _08072_);
  nor (_08075_, _07504_, _06861_);
  nor (_08076_, _07504_, \oc8051_golden_model_1.ACC [5]);
  and (_08077_, _07504_, \oc8051_golden_model_1.ACC [5]);
  nor (_08078_, _08077_, _08076_);
  nor (_08079_, _07517_, _06867_);
  and (_08080_, _07517_, \oc8051_golden_model_1.ACC [4]);
  nor (_08081_, _07517_, \oc8051_golden_model_1.ACC [4]);
  nor (_08082_, _08081_, _08080_);
  not (_08083_, _08082_);
  nor (_08084_, _07453_, _06964_);
  and (_08085_, _07453_, \oc8051_golden_model_1.ACC [2]);
  nor (_08086_, _07453_, \oc8051_golden_model_1.ACC [2]);
  nor (_08087_, _08086_, _08085_);
  nor (_08088_, _07467_, _02551_);
  nor (_08089_, _07481_, _02667_);
  not (_08090_, _08089_);
  nor (_08091_, _08090_, _07576_);
  nor (_08092_, _08091_, _08088_);
  nor (_08093_, _08092_, _08087_);
  nor (_08094_, _08093_, _08084_);
  nor (_08095_, _08094_, _07442_);
  or (_08096_, _08095_, \oc8051_golden_model_1.ACC [3]);
  nand (_08097_, _08094_, _07442_);
  and (_08098_, _08097_, _08096_);
  and (_08099_, _08098_, _08083_);
  nor (_08100_, _08099_, _08079_);
  nor (_08101_, _08100_, _08078_);
  nor (_08102_, _08101_, _08075_);
  nor (_08103_, _08102_, _08074_);
  nor (_08104_, _08103_, _08071_);
  nor (_08105_, _08104_, _08070_);
  and (_08106_, _08104_, _08070_);
  or (_08107_, _08106_, _08105_);
  or (_08108_, _08107_, _08065_);
  and (_08109_, _08108_, _08067_);
  or (_08110_, _08109_, _08064_);
  and (_08111_, _02545_, _02891_);
  not (_08112_, _08111_);
  not (_08113_, _08065_);
  nor (_08114_, _02927_, _06806_);
  and (_08115_, _02927_, _06806_);
  nor (_08116_, _08115_, _08114_);
  nor (_08117_, _03211_, _06861_);
  and (_08118_, _03211_, _06861_);
  nor (_08119_, _08118_, _08117_);
  not (_08120_, _08119_);
  nor (_08121_, _03629_, _06867_);
  and (_08122_, _03629_, _06867_);
  nor (_08123_, _08122_, _08121_);
  nor (_08124_, _02794_, _02564_);
  and (_08125_, _02794_, _02564_);
  nor (_08126_, _03256_, _06964_);
  and (_08127_, _03256_, _06964_);
  or (_08128_, _08127_, _08126_);
  nor (_08129_, _03665_, _02551_);
  and (_08130_, _03665_, _02551_);
  nor (_08131_, _08130_, _08129_);
  and (_08132_, _02835_, \oc8051_golden_model_1.ACC [0]);
  and (_08133_, _08132_, _08131_);
  nor (_08134_, _08133_, _08129_);
  nor (_08135_, _08134_, _08128_);
  nor (_08136_, _08135_, _08126_);
  nor (_08137_, _08136_, _08125_);
  or (_08138_, _08137_, _08124_);
  and (_08139_, _08138_, _08123_);
  nor (_08140_, _08139_, _08121_);
  nor (_08141_, _08140_, _08120_);
  or (_08142_, _08141_, _08117_);
  and (_08143_, _08142_, _08116_);
  nor (_08144_, _08143_, _08114_);
  nor (_08145_, _08144_, _07896_);
  and (_08146_, _08144_, _07896_);
  or (_08147_, _08146_, _08145_);
  or (_08148_, _08147_, _08113_);
  and (_08149_, _08148_, _08112_);
  and (_08150_, _08149_, _08110_);
  and (_08151_, _08111_, \oc8051_golden_model_1.ACC [6]);
  or (_08152_, _08151_, _03163_);
  or (_08153_, _08152_, _08150_);
  and (_08154_, _02951_, _02367_);
  not (_08155_, _08154_);
  nand (_08156_, _07651_, _03163_);
  and (_08157_, _08156_, _08155_);
  and (_08158_, _08157_, _08153_);
  and (_08159_, _02545_, _02367_);
  nor (_08160_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08161_, _08160_, _06905_);
  and (_08162_, _08161_, _06824_);
  and (_08163_, _08162_, _06806_);
  nor (_08164_, _08163_, _05771_);
  and (_08165_, _08163_, _05771_);
  nor (_08166_, _08165_, _08164_);
  nor (_08167_, _08166_, _08155_);
  or (_08168_, _08167_, _08159_);
  or (_08169_, _08168_, _08158_);
  nand (_08170_, _08159_, _07293_);
  and (_08171_, _08170_, _02498_);
  and (_08172_, _08171_, _08169_);
  nor (_08173_, _07700_, _02498_);
  or (_08174_, _08173_, _02888_);
  or (_08175_, _08174_, _08172_);
  and (_08176_, _02951_, _02522_);
  not (_08177_, _08176_);
  and (_08178_, _05235_, _04706_);
  nor (_08179_, _08178_, _07400_);
  nand (_08180_, _08179_, _02888_);
  and (_08181_, _08180_, _08177_);
  and (_08182_, _08181_, _08175_);
  and (_08183_, _02545_, _02522_);
  and (_08184_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08185_, _08184_, _06906_);
  nor (_08186_, _08185_, _06867_);
  and (_08187_, _08186_, \oc8051_golden_model_1.ACC [5]);
  and (_08188_, _08187_, \oc8051_golden_model_1.ACC [6]);
  nor (_08189_, _08188_, \oc8051_golden_model_1.ACC [7]);
  and (_08190_, _08188_, \oc8051_golden_model_1.ACC [7]);
  nor (_08191_, _08190_, _08189_);
  and (_08192_, _08191_, _08176_);
  or (_08193_, _08192_, _08183_);
  or (_08194_, _08193_, _08182_);
  nand (_08195_, _08183_, _02667_);
  and (_08196_, _08195_, _42668_);
  and (_08197_, _08196_, _08194_);
  or (_08198_, _08197_, _07187_);
  and (_40487_, _08198_, _43998_);
  or (_08199_, _42668_, \oc8051_golden_model_1.DPL [7]);
  and (_08200_, _08199_, _43998_);
  not (_08201_, \oc8051_golden_model_1.DPL [7]);
  nor (_08202_, _04612_, _08201_);
  and (_08203_, _05774_, _04612_);
  or (_08204_, _08203_, _08202_);
  and (_08205_, _08204_, _03127_);
  and (_08206_, _04612_, _04604_);
  or (_08207_, _08206_, _08202_);
  or (_08208_, _08207_, _05535_);
  not (_08209_, _02981_);
  and (_08210_, _05474_, _04612_);
  or (_08211_, _08210_, _08202_);
  or (_08212_, _08211_, _03810_);
  and (_08213_, _04612_, \oc8051_golden_model_1.ACC [7]);
  or (_08214_, _08213_, _08202_);
  and (_08215_, _08214_, _03813_);
  nor (_08216_, _03813_, _08201_);
  or (_08217_, _08216_, _02974_);
  or (_08218_, _08217_, _08215_);
  and (_08219_, _08218_, _03336_);
  and (_08220_, _08219_, _08212_);
  and (_08221_, _08207_, _03069_);
  or (_08222_, _08221_, _03075_);
  or (_08223_, _08222_, _08220_);
  and (_08224_, _03099_, _02545_);
  not (_08225_, _08224_);
  or (_08226_, _08214_, _03084_);
  and (_08227_, _08226_, _08225_);
  and (_08228_, _08227_, _08223_);
  and (_08229_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08230_, _08229_, \oc8051_golden_model_1.DPL [2]);
  and (_08231_, _08230_, \oc8051_golden_model_1.DPL [3]);
  and (_08232_, _08231_, \oc8051_golden_model_1.DPL [4]);
  and (_08233_, _08232_, \oc8051_golden_model_1.DPL [5]);
  and (_08234_, _08233_, \oc8051_golden_model_1.DPL [6]);
  nor (_08235_, _08234_, \oc8051_golden_model_1.DPL [7]);
  and (_08236_, _08234_, \oc8051_golden_model_1.DPL [7]);
  nor (_08237_, _08236_, _08235_);
  and (_08238_, _08237_, _08224_);
  or (_08239_, _08238_, _08228_);
  and (_08240_, _08239_, _08209_);
  nor (_08241_, _05311_, _08209_);
  or (_08242_, _08241_, _06770_);
  or (_08243_, _08242_, _08240_);
  and (_08244_, _08243_, _08208_);
  or (_08245_, _08244_, _02853_);
  and (_08246_, _04612_, _05462_);
  or (_08247_, _08202_, _05540_);
  or (_08248_, _08247_, _08246_);
  and (_08249_, _08248_, _02838_);
  and (_08250_, _08249_, _08245_);
  not (_08251_, _04612_);
  nor (_08252_, _05744_, _08251_);
  or (_08253_, _08252_, _08202_);
  and (_08254_, _08253_, _02579_);
  or (_08255_, _08254_, _02802_);
  or (_08256_, _08255_, _08250_);
  and (_08257_, _05661_, _04612_);
  or (_08258_, _08257_, _08202_);
  or (_08259_, _08258_, _02803_);
  and (_08260_, _08259_, _08256_);
  or (_08261_, _08260_, _02980_);
  and (_08262_, _05766_, _04612_);
  or (_08263_, _08202_, _03887_);
  or (_08264_, _08263_, _08262_);
  and (_08265_, _08264_, _03128_);
  and (_08266_, _08265_, _08261_);
  or (_08267_, _08266_, _08205_);
  and (_08268_, _08267_, _03883_);
  or (_08269_, _08202_, _04715_);
  and (_08270_, _08258_, _02970_);
  and (_08271_, _08270_, _08269_);
  or (_08272_, _08271_, _08268_);
  and (_08273_, _08272_, _03137_);
  and (_08274_, _08214_, _03135_);
  and (_08275_, _08274_, _08269_);
  or (_08276_, _08275_, _02965_);
  or (_08277_, _08276_, _08273_);
  nor (_08278_, _05765_, _08251_);
  or (_08279_, _08202_, _05783_);
  or (_08280_, _08279_, _08278_);
  and (_08281_, _08280_, _05788_);
  and (_08282_, _08281_, _08277_);
  nor (_08283_, _05773_, _08251_);
  or (_08284_, _08283_, _08202_);
  and (_08285_, _08284_, _03123_);
  or (_08286_, _08285_, _03163_);
  or (_08287_, _08286_, _08282_);
  or (_08288_, _08211_, _03906_);
  and (_08289_, _08288_, _02890_);
  and (_08290_, _08289_, _08287_);
  and (_08291_, _05235_, _04612_);
  or (_08292_, _08291_, _08202_);
  and (_08293_, _08292_, _02888_);
  or (_08294_, _08293_, _42672_);
  or (_08295_, _08294_, _08290_);
  and (_40488_, _08295_, _08200_);
  or (_08296_, _42668_, \oc8051_golden_model_1.DPH [7]);
  and (_08297_, _08296_, _43998_);
  not (_08298_, \oc8051_golden_model_1.DPH [7]);
  nor (_08299_, _04783_, _08298_);
  and (_08300_, _05774_, _04671_);
  or (_08301_, _08300_, _08299_);
  and (_08302_, _08301_, _03127_);
  and (_08303_, _04671_, _04604_);
  or (_08304_, _08303_, _08299_);
  or (_08305_, _08304_, _05535_);
  and (_08306_, _05474_, _04671_);
  or (_08307_, _08306_, _08299_);
  or (_08308_, _08307_, _03810_);
  and (_08309_, _04783_, \oc8051_golden_model_1.ACC [7]);
  or (_08310_, _08309_, _08299_);
  and (_08311_, _08310_, _03813_);
  nor (_08312_, _03813_, _08298_);
  or (_08313_, _08312_, _02974_);
  or (_08314_, _08313_, _08311_);
  and (_08315_, _08314_, _03336_);
  and (_08316_, _08315_, _08308_);
  and (_08317_, _08304_, _03069_);
  or (_08318_, _08317_, _03075_);
  or (_08319_, _08318_, _08316_);
  or (_08320_, _08310_, _03084_);
  and (_08321_, _08320_, _08225_);
  and (_08322_, _08321_, _08319_);
  and (_08323_, _08236_, \oc8051_golden_model_1.DPH [0]);
  and (_08324_, _08323_, \oc8051_golden_model_1.DPH [1]);
  and (_08325_, _08324_, \oc8051_golden_model_1.DPH [2]);
  and (_08326_, _08325_, \oc8051_golden_model_1.DPH [3]);
  and (_08327_, _08326_, \oc8051_golden_model_1.DPH [4]);
  and (_08328_, _08327_, \oc8051_golden_model_1.DPH [5]);
  and (_08329_, _08328_, \oc8051_golden_model_1.DPH [6]);
  nand (_08330_, _08329_, \oc8051_golden_model_1.DPH [7]);
  or (_08331_, _08329_, \oc8051_golden_model_1.DPH [7]);
  and (_08332_, _08331_, _08224_);
  and (_08333_, _08332_, _08330_);
  or (_08334_, _08333_, _08322_);
  and (_08335_, _08334_, _08209_);
  and (_08336_, _02981_, _02763_);
  or (_08337_, _08336_, _06770_);
  or (_08338_, _08337_, _08335_);
  and (_08339_, _08338_, _08305_);
  or (_08340_, _08339_, _02853_);
  or (_08341_, _08299_, _05540_);
  and (_08342_, _04783_, _05462_);
  or (_08343_, _08342_, _08341_);
  and (_08344_, _08343_, _02838_);
  and (_08345_, _08344_, _08340_);
  not (_08346_, _04783_);
  nor (_08347_, _05744_, _08346_);
  or (_08348_, _08347_, _08299_);
  and (_08349_, _08348_, _02579_);
  or (_08350_, _08349_, _02802_);
  or (_08351_, _08350_, _08345_);
  and (_08352_, _05661_, _04783_);
  or (_08353_, _08352_, _08299_);
  or (_08354_, _08353_, _02803_);
  and (_08355_, _08354_, _08351_);
  or (_08356_, _08355_, _02980_);
  and (_08357_, _05766_, _04671_);
  or (_08358_, _08299_, _03887_);
  or (_08359_, _08358_, _08357_);
  and (_08360_, _08359_, _03128_);
  and (_08361_, _08360_, _08356_);
  or (_08362_, _08361_, _08302_);
  and (_08363_, _08362_, _03883_);
  or (_08364_, _08299_, _04715_);
  and (_08365_, _08353_, _02970_);
  and (_08366_, _08365_, _08364_);
  or (_08367_, _08366_, _08363_);
  and (_08368_, _08367_, _03137_);
  and (_08369_, _08310_, _03135_);
  and (_08370_, _08369_, _08364_);
  or (_08371_, _08370_, _02965_);
  or (_08372_, _08371_, _08368_);
  not (_08373_, _04671_);
  nor (_08374_, _05765_, _08373_);
  or (_08375_, _08299_, _05783_);
  or (_08376_, _08375_, _08374_);
  and (_08377_, _08376_, _05788_);
  and (_08378_, _08377_, _08372_);
  nor (_08379_, _05773_, _08373_);
  or (_08380_, _08379_, _08299_);
  and (_08381_, _08380_, _03123_);
  or (_08382_, _08381_, _03163_);
  or (_08383_, _08382_, _08378_);
  or (_08384_, _08307_, _03906_);
  and (_08385_, _08384_, _02890_);
  and (_08386_, _08385_, _08383_);
  and (_08387_, _05235_, _04671_);
  or (_08388_, _08387_, _08299_);
  and (_08389_, _08388_, _02888_);
  or (_08390_, _08389_, _42672_);
  or (_08391_, _08390_, _08386_);
  and (_40489_, _08391_, _08297_);
  not (_08392_, \oc8051_golden_model_1.IE [7]);
  nor (_08393_, _04703_, _08392_);
  and (_08394_, _05774_, _04703_);
  nor (_08395_, _08394_, _08393_);
  nor (_08396_, _08395_, _03128_);
  and (_08397_, _04703_, _04604_);
  nor (_08398_, _08397_, _08393_);
  and (_08399_, _08398_, _06770_);
  nor (_08400_, _05340_, _08392_);
  and (_08401_, _05356_, _05340_);
  nor (_08402_, _08401_, _08400_);
  nor (_08403_, _08402_, _02877_);
  and (_08404_, _04703_, \oc8051_golden_model_1.ACC [7]);
  nor (_08405_, _08404_, _08393_);
  nor (_08406_, _08405_, _03814_);
  nor (_08407_, _03813_, _08392_);
  or (_08408_, _08407_, _08406_);
  and (_08409_, _08408_, _03810_);
  and (_08410_, _05474_, _04703_);
  nor (_08411_, _08410_, _08393_);
  nor (_08412_, _08411_, _03810_);
  or (_08413_, _08412_, _08409_);
  and (_08414_, _08413_, _02881_);
  and (_08415_, _05360_, _05340_);
  nor (_08416_, _08415_, _08400_);
  nor (_08417_, _08416_, _02881_);
  or (_08418_, _08417_, _03069_);
  or (_08419_, _08418_, _08414_);
  nand (_08420_, _08398_, _03069_);
  and (_08421_, _08420_, _08419_);
  and (_08422_, _08421_, _03084_);
  nor (_08423_, _08405_, _03084_);
  or (_08424_, _08423_, _08422_);
  and (_08425_, _08424_, _02877_);
  nor (_08426_, _08425_, _08403_);
  nor (_08427_, _08426_, _02869_);
  and (_08428_, _05503_, _05340_);
  nor (_08429_, _08428_, _08400_);
  nor (_08430_, _08429_, _02870_);
  nor (_08431_, _08430_, _08427_);
  nor (_08432_, _08431_, _02863_);
  not (_08433_, _05340_);
  nor (_08434_, _05530_, _08433_);
  nor (_08435_, _08434_, _08400_);
  nor (_08436_, _08435_, _02864_);
  nor (_08437_, _08436_, _06770_);
  not (_08438_, _08437_);
  nor (_08439_, _08438_, _08432_);
  nor (_08440_, _08439_, _08399_);
  nor (_08441_, _08440_, _02853_);
  and (_08442_, _04703_, _05462_);
  nor (_08443_, _08393_, _05540_);
  not (_08444_, _08443_);
  nor (_08445_, _08444_, _08442_);
  nor (_08446_, _08445_, _02579_);
  not (_08447_, _08446_);
  nor (_08448_, _08447_, _08441_);
  not (_08449_, _04703_);
  nor (_08450_, _05744_, _08449_);
  nor (_08451_, _08450_, _08393_);
  nor (_08452_, _08451_, _02838_);
  or (_08453_, _08452_, _02802_);
  or (_08454_, _08453_, _08448_);
  and (_08455_, _05661_, _04703_);
  nor (_08456_, _08455_, _08393_);
  nand (_08457_, _08456_, _02802_);
  and (_08458_, _08457_, _08454_);
  and (_08459_, _08458_, _03887_);
  and (_08460_, _05766_, _04703_);
  nor (_08461_, _08460_, _08393_);
  nor (_08462_, _08461_, _03887_);
  or (_08463_, _08462_, _08459_);
  and (_08464_, _08463_, _03128_);
  nor (_08465_, _08464_, _08396_);
  nor (_08466_, _08465_, _02970_);
  nor (_08467_, _08393_, _04715_);
  not (_08468_, _08467_);
  nor (_08469_, _08456_, _03883_);
  and (_08470_, _08469_, _08468_);
  nor (_08471_, _08470_, _08466_);
  nor (_08472_, _08471_, _03135_);
  nor (_08473_, _08405_, _03137_);
  and (_08474_, _08473_, _08468_);
  nor (_08475_, _08474_, _02965_);
  not (_08476_, _08475_);
  nor (_08477_, _08476_, _08472_);
  nor (_08478_, _05765_, _08449_);
  or (_08479_, _08393_, _05783_);
  nor (_08480_, _08479_, _08478_);
  or (_08481_, _08480_, _03123_);
  nor (_08482_, _08481_, _08477_);
  nor (_08483_, _05773_, _08449_);
  nor (_08484_, _08483_, _08393_);
  nor (_08485_, _08484_, _05788_);
  or (_08486_, _08485_, _08482_);
  and (_08487_, _08486_, _03906_);
  nor (_08488_, _08411_, _03906_);
  or (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _02498_);
  nor (_08491_, _08402_, _02498_);
  or (_08492_, _08491_, _08490_);
  and (_08493_, _08492_, _02890_);
  and (_08494_, _05235_, _04703_);
  nor (_08495_, _08494_, _08393_);
  nor (_08496_, _08495_, _02890_);
  or (_08497_, _08496_, _08493_);
  or (_08498_, _08497_, _42672_);
  or (_08499_, _42668_, \oc8051_golden_model_1.IE [7]);
  and (_08500_, _08499_, _43998_);
  and (_40490_, _08500_, _08498_);
  not (_08501_, \oc8051_golden_model_1.IP [7]);
  nor (_08502_, _04693_, _08501_);
  and (_08503_, _05774_, _04693_);
  nor (_08504_, _08503_, _08502_);
  nor (_08505_, _08504_, _03128_);
  and (_08506_, _04693_, _04604_);
  nor (_08507_, _08506_, _08502_);
  and (_08508_, _08507_, _06770_);
  nor (_08509_, _05328_, _08501_);
  and (_08510_, _05356_, _05328_);
  nor (_08511_, _08510_, _08509_);
  nor (_08512_, _08511_, _02877_);
  and (_08513_, _04693_, \oc8051_golden_model_1.ACC [7]);
  nor (_08514_, _08513_, _08502_);
  nor (_08515_, _08514_, _03814_);
  nor (_08516_, _03813_, _08501_);
  or (_08517_, _08516_, _08515_);
  and (_08518_, _08517_, _03810_);
  and (_08519_, _05474_, _04693_);
  nor (_08520_, _08519_, _08502_);
  nor (_08521_, _08520_, _03810_);
  or (_08522_, _08521_, _08518_);
  and (_08523_, _08522_, _02881_);
  and (_08524_, _05360_, _05328_);
  nor (_08525_, _08524_, _08509_);
  nor (_08526_, _08525_, _02881_);
  or (_08527_, _08526_, _03069_);
  or (_08528_, _08527_, _08523_);
  nand (_08529_, _08507_, _03069_);
  and (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _03084_);
  nor (_08532_, _08514_, _03084_);
  or (_08533_, _08532_, _08531_);
  and (_08534_, _08533_, _02877_);
  nor (_08535_, _08534_, _08512_);
  nor (_08536_, _08535_, _02869_);
  and (_08537_, _05503_, _05328_);
  nor (_08538_, _08537_, _08509_);
  nor (_08539_, _08538_, _02870_);
  nor (_08540_, _08539_, _08536_);
  nor (_08541_, _08540_, _02863_);
  not (_08542_, _05328_);
  nor (_08543_, _05530_, _08542_);
  nor (_08544_, _08543_, _08509_);
  nor (_08545_, _08544_, _02864_);
  nor (_08546_, _08545_, _06770_);
  not (_08547_, _08546_);
  nor (_08548_, _08547_, _08541_);
  nor (_08549_, _08548_, _08508_);
  nor (_08550_, _08549_, _02853_);
  and (_08551_, _04693_, _05462_);
  nor (_08552_, _08502_, _05540_);
  not (_08553_, _08552_);
  nor (_08554_, _08553_, _08551_);
  nor (_08555_, _08554_, _02579_);
  not (_08556_, _08555_);
  nor (_08557_, _08556_, _08550_);
  not (_08558_, _04693_);
  nor (_08559_, _05744_, _08558_);
  nor (_08560_, _08559_, _08502_);
  nor (_08561_, _08560_, _02838_);
  or (_08562_, _08561_, _02802_);
  or (_08563_, _08562_, _08557_);
  and (_08564_, _05661_, _04693_);
  nor (_08565_, _08564_, _08502_);
  nand (_08566_, _08565_, _02802_);
  and (_08567_, _08566_, _08563_);
  and (_08568_, _08567_, _03887_);
  and (_08569_, _05766_, _04693_);
  nor (_08570_, _08569_, _08502_);
  nor (_08571_, _08570_, _03887_);
  or (_08572_, _08571_, _08568_);
  and (_08573_, _08572_, _03128_);
  nor (_08574_, _08573_, _08505_);
  nor (_08575_, _08574_, _02970_);
  nor (_08576_, _08502_, _04715_);
  not (_08577_, _08576_);
  nor (_08578_, _08565_, _03883_);
  and (_08579_, _08578_, _08577_);
  nor (_08580_, _08579_, _08575_);
  nor (_08581_, _08580_, _03135_);
  nor (_08582_, _08514_, _03137_);
  and (_08583_, _08582_, _08577_);
  nor (_08584_, _08583_, _02965_);
  not (_08585_, _08584_);
  nor (_08586_, _08585_, _08581_);
  nor (_08587_, _05765_, _08558_);
  or (_08588_, _08502_, _05783_);
  nor (_08589_, _08588_, _08587_);
  or (_08590_, _08589_, _03123_);
  nor (_08591_, _08590_, _08586_);
  nor (_08592_, _05773_, _08558_);
  nor (_08593_, _08592_, _08502_);
  nor (_08594_, _08593_, _05788_);
  or (_08595_, _08594_, _08591_);
  and (_08596_, _08595_, _03906_);
  nor (_08597_, _08520_, _03906_);
  or (_08598_, _08597_, _08596_);
  and (_08599_, _08598_, _02498_);
  nor (_08600_, _08511_, _02498_);
  or (_08601_, _08600_, _08599_);
  and (_08602_, _08601_, _02890_);
  and (_08603_, _05235_, _04693_);
  nor (_08604_, _08603_, _08502_);
  nor (_08605_, _08604_, _02890_);
  or (_08606_, _08605_, _08602_);
  or (_08607_, _08606_, _42672_);
  or (_08608_, _42668_, \oc8051_golden_model_1.IP [7]);
  and (_08609_, _08608_, _43998_);
  and (_40491_, _08609_, _08607_);
  not (_08610_, \oc8051_golden_model_1.P0 [7]);
  nor (_08611_, _42668_, _08610_);
  or (_08612_, _08611_, rst);
  nor (_08613_, _04628_, _08610_);
  and (_08614_, _05774_, _04628_);
  or (_08615_, _08614_, _08613_);
  and (_08616_, _08615_, _03127_);
  and (_08617_, _04628_, _04604_);
  or (_08618_, _08617_, _08613_);
  or (_08619_, _08618_, _05535_);
  nor (_08620_, _04609_, _08610_);
  and (_08621_, _05356_, _04609_);
  or (_08622_, _08621_, _08620_);
  and (_08623_, _08622_, _02876_);
  and (_08624_, _05474_, _04628_);
  or (_08625_, _08624_, _08613_);
  or (_08626_, _08625_, _03810_);
  and (_08627_, _04628_, \oc8051_golden_model_1.ACC [7]);
  or (_08628_, _08627_, _08613_);
  and (_08629_, _08628_, _03813_);
  nor (_08630_, _03813_, _08610_);
  or (_08631_, _08630_, _02974_);
  or (_08632_, _08631_, _08629_);
  and (_08633_, _08632_, _02881_);
  and (_08634_, _08633_, _08626_);
  and (_08635_, _05360_, _04609_);
  or (_08636_, _08635_, _08620_);
  and (_08637_, _08636_, _02880_);
  or (_08638_, _08637_, _03069_);
  or (_08639_, _08638_, _08634_);
  or (_08640_, _08618_, _03336_);
  and (_08641_, _08640_, _08639_);
  or (_08642_, _08641_, _03075_);
  or (_08643_, _08628_, _03084_);
  and (_08644_, _08643_, _02877_);
  and (_08645_, _08644_, _08642_);
  or (_08646_, _08645_, _08623_);
  and (_08647_, _08646_, _02870_);
  or (_08648_, _08620_, _05502_);
  and (_08649_, _08648_, _02869_);
  and (_08650_, _08649_, _08636_);
  or (_08651_, _08650_, _08647_);
  and (_08652_, _08651_, _02864_);
  or (_08653_, _05529_, _05356_);
  and (_08654_, _08653_, _04609_);
  or (_08655_, _08654_, _08620_);
  and (_08656_, _08655_, _02863_);
  or (_08657_, _08656_, _06770_);
  or (_08658_, _08657_, _08652_);
  and (_08659_, _08658_, _08619_);
  or (_08660_, _08659_, _02853_);
  and (_08661_, _04628_, _05462_);
  or (_08662_, _08613_, _05540_);
  or (_08663_, _08662_, _08661_);
  and (_08664_, _08663_, _02838_);
  and (_08665_, _08664_, _08660_);
  and (_08666_, _05717_, \oc8051_golden_model_1.P1 [7]);
  and (_08667_, _05710_, \oc8051_golden_model_1.P0 [7]);
  and (_08668_, _05720_, \oc8051_golden_model_1.P2 [7]);
  and (_08669_, _05663_, _05618_);
  and (_08670_, _08669_, \oc8051_golden_model_1.P3 [7]);
  or (_08671_, _08670_, _08668_);
  or (_08672_, _08671_, _08667_);
  or (_08673_, _08672_, _08666_);
  nor (_08674_, _08673_, _05708_);
  and (_08675_, _08674_, _05740_);
  and (_08676_, _08675_, _05706_);
  nand (_08677_, _08676_, _05691_);
  or (_08678_, _08677_, _05550_);
  and (_08679_, _08678_, _04628_);
  or (_08680_, _08679_, _08613_);
  and (_08681_, _08680_, _02579_);
  or (_08682_, _08681_, _02802_);
  or (_08683_, _08682_, _08665_);
  and (_08684_, _05661_, _04628_);
  or (_08685_, _08684_, _08613_);
  or (_08686_, _08685_, _02803_);
  and (_08687_, _08686_, _08683_);
  or (_08688_, _08687_, _02980_);
  and (_08689_, _05766_, _04628_);
  or (_08690_, _08613_, _03887_);
  or (_08691_, _08690_, _08689_);
  and (_08692_, _08691_, _03128_);
  and (_08693_, _08692_, _08688_);
  or (_08694_, _08693_, _08616_);
  and (_08695_, _08694_, _03883_);
  or (_08696_, _08613_, _04715_);
  and (_08697_, _08685_, _02970_);
  and (_08698_, _08697_, _08696_);
  or (_08699_, _08698_, _08695_);
  and (_08700_, _08699_, _03137_);
  and (_08701_, _08628_, _03135_);
  and (_08702_, _08701_, _08696_);
  or (_08703_, _08702_, _02965_);
  or (_08704_, _08703_, _08700_);
  not (_08705_, _04628_);
  nor (_08706_, _05765_, _08705_);
  or (_08707_, _08613_, _05783_);
  or (_08708_, _08707_, _08706_);
  and (_08709_, _08708_, _05788_);
  and (_08710_, _08709_, _08704_);
  nor (_08711_, _05773_, _08705_);
  or (_08712_, _08711_, _08613_);
  and (_08713_, _08712_, _03123_);
  or (_08714_, _08713_, _03163_);
  or (_08715_, _08714_, _08710_);
  or (_08716_, _08625_, _03906_);
  and (_08717_, _08716_, _02498_);
  and (_08718_, _08717_, _08715_);
  and (_08719_, _08622_, _02497_);
  or (_08720_, _08719_, _02888_);
  or (_08721_, _08720_, _08718_);
  and (_08722_, _05235_, _04628_);
  or (_08723_, _08613_, _02890_);
  or (_08724_, _08723_, _08722_);
  and (_08725_, _08724_, _42668_);
  and (_08726_, _08725_, _08721_);
  or (_40492_, _08726_, _08612_);
  not (_08727_, \oc8051_golden_model_1.P1 [7]);
  nor (_08728_, _42668_, _08727_);
  or (_08729_, _08728_, rst);
  nor (_08730_, _04634_, _08727_);
  and (_08731_, _05774_, _04634_);
  or (_08732_, _08731_, _08730_);
  and (_08733_, _08732_, _03127_);
  and (_08734_, _04634_, _04604_);
  or (_08735_, _08734_, _08730_);
  or (_08736_, _08735_, _05535_);
  nor (_08737_, _05344_, _08727_);
  and (_08738_, _05356_, _05344_);
  or (_08739_, _08738_, _08737_);
  and (_08740_, _08739_, _02876_);
  and (_08741_, _05474_, _04634_);
  or (_08742_, _08741_, _08730_);
  or (_08743_, _08742_, _03810_);
  and (_08744_, _04634_, \oc8051_golden_model_1.ACC [7]);
  or (_08745_, _08744_, _08730_);
  and (_08746_, _08745_, _03813_);
  nor (_08747_, _03813_, _08727_);
  or (_08748_, _08747_, _02974_);
  or (_08749_, _08748_, _08746_);
  and (_08750_, _08749_, _02881_);
  and (_08751_, _08750_, _08743_);
  and (_08752_, _05360_, _05344_);
  or (_08753_, _08752_, _08737_);
  and (_08754_, _08753_, _02880_);
  or (_08755_, _08754_, _03069_);
  or (_08756_, _08755_, _08751_);
  or (_08757_, _08735_, _03336_);
  and (_08758_, _08757_, _08756_);
  or (_08759_, _08758_, _03075_);
  or (_08760_, _08745_, _03084_);
  and (_08761_, _08760_, _02877_);
  and (_08762_, _08761_, _08759_);
  or (_08763_, _08762_, _08740_);
  and (_08764_, _08763_, _02870_);
  and (_08765_, _05503_, _05344_);
  or (_08766_, _08765_, _08737_);
  and (_08767_, _08766_, _02869_);
  or (_08768_, _08767_, _08764_);
  and (_08769_, _08768_, _02864_);
  and (_08770_, _08653_, _05344_);
  or (_08771_, _08770_, _08737_);
  and (_08772_, _08771_, _02863_);
  or (_08773_, _08772_, _06770_);
  or (_08774_, _08773_, _08769_);
  and (_08775_, _08774_, _08736_);
  or (_08776_, _08775_, _02853_);
  and (_08777_, _04634_, _05462_);
  or (_08778_, _08730_, _05540_);
  or (_08779_, _08778_, _08777_);
  and (_08780_, _08779_, _02838_);
  and (_08781_, _08780_, _08776_);
  and (_08782_, _08678_, _04634_);
  or (_08783_, _08782_, _08730_);
  and (_08784_, _08783_, _02579_);
  or (_08785_, _08784_, _02802_);
  or (_08786_, _08785_, _08781_);
  and (_08787_, _05661_, _04634_);
  or (_08788_, _08787_, _08730_);
  or (_08789_, _08788_, _02803_);
  and (_08790_, _08789_, _08786_);
  or (_08791_, _08790_, _02980_);
  and (_08792_, _05766_, _04634_);
  or (_08793_, _08730_, _03887_);
  or (_08794_, _08793_, _08792_);
  and (_08795_, _08794_, _03128_);
  and (_08796_, _08795_, _08791_);
  or (_08797_, _08796_, _08733_);
  and (_08798_, _08797_, _03883_);
  or (_08799_, _08730_, _04715_);
  and (_08800_, _08788_, _02970_);
  and (_08801_, _08800_, _08799_);
  or (_08802_, _08801_, _08798_);
  and (_08803_, _08802_, _03137_);
  and (_08804_, _08745_, _03135_);
  and (_08805_, _08804_, _08799_);
  or (_08806_, _08805_, _02965_);
  or (_08807_, _08806_, _08803_);
  not (_08808_, _04634_);
  nor (_08809_, _05765_, _08808_);
  or (_08810_, _08730_, _05783_);
  or (_08811_, _08810_, _08809_);
  and (_08812_, _08811_, _05788_);
  and (_08813_, _08812_, _08807_);
  nor (_08814_, _05773_, _08808_);
  or (_08815_, _08814_, _08730_);
  and (_08816_, _08815_, _03123_);
  or (_08817_, _08816_, _03163_);
  or (_08818_, _08817_, _08813_);
  or (_08819_, _08742_, _03906_);
  and (_08820_, _08819_, _02498_);
  and (_08821_, _08820_, _08818_);
  and (_08822_, _08739_, _02497_);
  or (_08823_, _08822_, _02888_);
  or (_08824_, _08823_, _08821_);
  and (_08825_, _05235_, _04634_);
  or (_08826_, _08730_, _02890_);
  or (_08827_, _08826_, _08825_);
  and (_08828_, _08827_, _42668_);
  and (_08829_, _08828_, _08824_);
  or (_40493_, _08829_, _08729_);
  not (_08830_, \oc8051_golden_model_1.P2 [7]);
  nor (_08831_, _42668_, _08830_);
  or (_08832_, _08831_, rst);
  nor (_08833_, _04641_, _08830_);
  and (_08834_, _05774_, _04641_);
  or (_08835_, _08834_, _08833_);
  and (_08836_, _08835_, _03127_);
  and (_08837_, _04641_, _04604_);
  or (_08838_, _08837_, _08833_);
  or (_08839_, _08838_, _05535_);
  nor (_08840_, _05347_, _08830_);
  and (_08841_, _05356_, _05347_);
  or (_08842_, _08841_, _08840_);
  and (_08843_, _08842_, _02876_);
  and (_08844_, _05474_, _04641_);
  or (_08845_, _08844_, _08833_);
  or (_08846_, _08845_, _03810_);
  and (_08847_, _04641_, \oc8051_golden_model_1.ACC [7]);
  or (_08848_, _08847_, _08833_);
  and (_08849_, _08848_, _03813_);
  nor (_08850_, _03813_, _08830_);
  or (_08851_, _08850_, _02974_);
  or (_08852_, _08851_, _08849_);
  and (_08853_, _08852_, _02881_);
  and (_08854_, _08853_, _08846_);
  and (_08855_, _05360_, _05347_);
  or (_08856_, _08855_, _08840_);
  and (_08857_, _08856_, _02880_);
  or (_08858_, _08857_, _03069_);
  or (_08859_, _08858_, _08854_);
  or (_08860_, _08838_, _03336_);
  and (_08861_, _08860_, _08859_);
  or (_08862_, _08861_, _03075_);
  or (_08863_, _08848_, _03084_);
  and (_08864_, _08863_, _02877_);
  and (_08865_, _08864_, _08862_);
  or (_08866_, _08865_, _08843_);
  and (_08867_, _08866_, _02870_);
  or (_08868_, _08840_, _05502_);
  and (_08869_, _08868_, _02869_);
  and (_08870_, _08869_, _08856_);
  or (_08871_, _08870_, _08867_);
  and (_08872_, _08871_, _02864_);
  and (_08873_, _08653_, _05347_);
  or (_08874_, _08873_, _08840_);
  and (_08875_, _08874_, _02863_);
  or (_08876_, _08875_, _06770_);
  or (_08877_, _08876_, _08872_);
  and (_08878_, _08877_, _08839_);
  or (_08879_, _08878_, _02853_);
  and (_08880_, _04641_, _05462_);
  or (_08881_, _08833_, _05540_);
  or (_08882_, _08881_, _08880_);
  and (_08883_, _08882_, _02838_);
  and (_08884_, _08883_, _08879_);
  and (_08885_, _08678_, _04641_);
  or (_08886_, _08885_, _08833_);
  and (_08887_, _08886_, _02579_);
  or (_08888_, _08887_, _02802_);
  or (_08889_, _08888_, _08884_);
  and (_08890_, _05661_, _04641_);
  or (_08891_, _08890_, _08833_);
  or (_08892_, _08891_, _02803_);
  and (_08893_, _08892_, _08889_);
  or (_08894_, _08893_, _02980_);
  and (_08895_, _05766_, _04641_);
  or (_08896_, _08833_, _03887_);
  or (_08897_, _08896_, _08895_);
  and (_08898_, _08897_, _03128_);
  and (_08899_, _08898_, _08894_);
  or (_08900_, _08899_, _08836_);
  and (_08901_, _08900_, _03883_);
  or (_08902_, _08833_, _04715_);
  and (_08903_, _08891_, _02970_);
  and (_08904_, _08903_, _08902_);
  or (_08905_, _08904_, _08901_);
  and (_08906_, _08905_, _03137_);
  and (_08907_, _08848_, _03135_);
  and (_08908_, _08907_, _08902_);
  or (_08909_, _08908_, _02965_);
  or (_08910_, _08909_, _08906_);
  not (_08911_, _04641_);
  nor (_08912_, _05765_, _08911_);
  or (_08913_, _08833_, _05783_);
  or (_08914_, _08913_, _08912_);
  and (_08915_, _08914_, _05788_);
  and (_08916_, _08915_, _08910_);
  nor (_08917_, _05773_, _08911_);
  or (_08918_, _08917_, _08833_);
  and (_08919_, _08918_, _03123_);
  or (_08920_, _08919_, _03163_);
  or (_08921_, _08920_, _08916_);
  or (_08922_, _08845_, _03906_);
  and (_08923_, _08922_, _02498_);
  and (_08924_, _08923_, _08921_);
  and (_08925_, _08842_, _02497_);
  or (_08926_, _08925_, _02888_);
  or (_08927_, _08926_, _08924_);
  and (_08928_, _05235_, _04641_);
  or (_08929_, _08833_, _02890_);
  or (_08930_, _08929_, _08928_);
  and (_08931_, _08930_, _42668_);
  and (_08932_, _08931_, _08927_);
  or (_40494_, _08932_, _08832_);
  not (_08933_, \oc8051_golden_model_1.P3 [7]);
  nor (_08934_, _42668_, _08933_);
  or (_08935_, _08934_, rst);
  nor (_08936_, _04645_, _08933_);
  and (_08937_, _05774_, _04645_);
  or (_08938_, _08937_, _08936_);
  and (_08939_, _08938_, _03127_);
  and (_08940_, _04645_, _04604_);
  or (_08941_, _08940_, _08936_);
  or (_08942_, _08941_, _05535_);
  nor (_08943_, _05349_, _08933_);
  and (_08944_, _05356_, _05349_);
  or (_08945_, _08944_, _08943_);
  and (_08946_, _08945_, _02876_);
  and (_08947_, _05474_, _04645_);
  or (_08948_, _08947_, _08936_);
  or (_08949_, _08948_, _03810_);
  and (_08950_, _04645_, \oc8051_golden_model_1.ACC [7]);
  or (_08951_, _08950_, _08936_);
  and (_08952_, _08951_, _03813_);
  nor (_08953_, _03813_, _08933_);
  or (_08954_, _08953_, _02974_);
  or (_08955_, _08954_, _08952_);
  and (_08956_, _08955_, _02881_);
  and (_08957_, _08956_, _08949_);
  and (_08958_, _05360_, _05349_);
  or (_08959_, _08958_, _08943_);
  and (_08960_, _08959_, _02880_);
  or (_08961_, _08960_, _03069_);
  or (_08962_, _08961_, _08957_);
  or (_08964_, _08941_, _03336_);
  and (_08965_, _08964_, _08962_);
  or (_08966_, _08965_, _03075_);
  or (_08967_, _08951_, _03084_);
  and (_08968_, _08967_, _02877_);
  and (_08969_, _08968_, _08966_);
  or (_08970_, _08969_, _08946_);
  and (_08971_, _08970_, _02870_);
  and (_08972_, _05503_, _05349_);
  or (_08973_, _08972_, _08943_);
  and (_08975_, _08973_, _02869_);
  or (_08976_, _08975_, _08971_);
  and (_08977_, _08976_, _02864_);
  and (_08978_, _08653_, _05349_);
  or (_08979_, _08978_, _08943_);
  and (_08980_, _08979_, _02863_);
  or (_08981_, _08980_, _06770_);
  or (_08982_, _08981_, _08977_);
  and (_08983_, _08982_, _08942_);
  or (_08984_, _08983_, _02853_);
  and (_08986_, _04645_, _05462_);
  or (_08987_, _08936_, _05540_);
  or (_08988_, _08987_, _08986_);
  and (_08989_, _08988_, _02838_);
  and (_08990_, _08989_, _08984_);
  and (_08991_, _08678_, _04645_);
  or (_08992_, _08991_, _08936_);
  and (_08993_, _08992_, _02579_);
  or (_08994_, _08993_, _02802_);
  or (_08995_, _08994_, _08990_);
  and (_08997_, _05661_, _04645_);
  or (_08998_, _08997_, _08936_);
  or (_08999_, _08998_, _02803_);
  and (_09000_, _08999_, _08995_);
  or (_09001_, _09000_, _02980_);
  and (_09002_, _05766_, _04645_);
  or (_09003_, _08936_, _03887_);
  or (_09004_, _09003_, _09002_);
  and (_09005_, _09004_, _03128_);
  and (_09006_, _09005_, _09001_);
  or (_09008_, _09006_, _08939_);
  and (_09009_, _09008_, _03883_);
  or (_09010_, _08936_, _04715_);
  and (_09011_, _08998_, _02970_);
  and (_09012_, _09011_, _09010_);
  or (_09013_, _09012_, _09009_);
  and (_09014_, _09013_, _03137_);
  and (_09015_, _08951_, _03135_);
  and (_09016_, _09015_, _09010_);
  or (_09017_, _09016_, _02965_);
  or (_09019_, _09017_, _09014_);
  not (_09020_, _04645_);
  nor (_09021_, _05765_, _09020_);
  or (_09022_, _08936_, _05783_);
  or (_09023_, _09022_, _09021_);
  and (_09024_, _09023_, _05788_);
  and (_09025_, _09024_, _09019_);
  nor (_09026_, _05773_, _09020_);
  or (_09027_, _09026_, _08936_);
  and (_09028_, _09027_, _03123_);
  or (_09030_, _09028_, _03163_);
  or (_09031_, _09030_, _09025_);
  or (_09032_, _08948_, _03906_);
  and (_09033_, _09032_, _02498_);
  and (_09034_, _09033_, _09031_);
  and (_09035_, _08945_, _02497_);
  or (_09036_, _09035_, _02888_);
  or (_09037_, _09036_, _09034_);
  and (_09038_, _05235_, _04645_);
  or (_09039_, _08936_, _02890_);
  or (_09040_, _09039_, _09038_);
  and (_09041_, _09040_, _42668_);
  and (_09042_, _09041_, _09037_);
  or (_40495_, _09042_, _08935_);
  not (_09043_, _02937_);
  nor (_09044_, _08183_, _08176_);
  and (_09045_, _05254_, _02230_);
  and (_09046_, _09045_, \oc8051_golden_model_1.PC [7]);
  and (_09047_, _09046_, _06175_);
  and (_09048_, _09047_, \oc8051_golden_model_1.PC [11]);
  and (_09049_, _09048_, \oc8051_golden_model_1.PC [12]);
  and (_09050_, _09049_, \oc8051_golden_model_1.PC [13]);
  and (_09051_, _09050_, \oc8051_golden_model_1.PC [14]);
  nor (_09052_, _09051_, \oc8051_golden_model_1.PC [15]);
  and (_09053_, _09046_, \oc8051_golden_model_1.PC [8]);
  and (_09054_, _09053_, \oc8051_golden_model_1.PC [9]);
  and (_09055_, _09054_, \oc8051_golden_model_1.PC [10]);
  and (_09056_, _09055_, \oc8051_golden_model_1.PC [11]);
  and (_09057_, _09056_, \oc8051_golden_model_1.PC [12]);
  and (_09058_, _09057_, \oc8051_golden_model_1.PC [13]);
  and (_09059_, _09058_, \oc8051_golden_model_1.PC [14]);
  and (_09060_, _09059_, \oc8051_golden_model_1.PC [15]);
  nor (_09061_, _09060_, _09052_);
  nor (_09062_, _09061_, _09044_);
  and (_09063_, _07238_, _08024_);
  nor (_09064_, _09063_, _09061_);
  nor (_09065_, _07962_, _03133_);
  and (_09066_, _07322_, _07241_);
  nor (_09067_, _09066_, _09061_);
  and (_09068_, _02496_, _02964_);
  not (_09069_, _02535_);
  nor (_09070_, _03123_, _09069_);
  nor (_09071_, _09070_, _06205_);
  or (_09072_, _09071_, _09068_);
  nor (_09073_, _07935_, _07930_);
  and (_09074_, _09073_, _07926_);
  nor (_09075_, _09074_, _09061_);
  and (_09076_, _02496_, _02969_);
  nor (_09077_, _03135_, _03880_);
  nor (_09078_, _09077_, _06205_);
  or (_09079_, _09078_, _09076_);
  nor (_09080_, _07394_, _03138_);
  nor (_09081_, _07908_, _07911_);
  nor (_09082_, _09081_, _09061_);
  and (_09083_, _02496_, _02513_);
  and (_09084_, _08165_, _06205_);
  nor (_09085_, _06194_, \oc8051_golden_model_1.PC [14]);
  nor (_09086_, _09085_, _06195_);
  and (_09087_, _09086_, _02763_);
  nor (_09088_, _09086_, _02763_);
  nor (_09089_, _09088_, _09087_);
  not (_09090_, \oc8051_golden_model_1.PC [13]);
  and (_09091_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09092_, _09091_, _06174_);
  and (_09093_, _09092_, _05366_);
  and (_09094_, _09093_, \oc8051_golden_model_1.PC [12]);
  nor (_09095_, _09094_, _09090_);
  and (_09096_, _09094_, _09090_);
  or (_09097_, _09096_, _09095_);
  and (_09098_, _09097_, _02763_);
  nor (_09099_, _09097_, _02763_);
  nor (_09100_, _06192_, \oc8051_golden_model_1.PC [12]);
  nor (_09101_, _09100_, _06193_);
  and (_09102_, _09101_, _02763_);
  nor (_09103_, _06199_, \oc8051_golden_model_1.PC [11]);
  nor (_09104_, _09103_, _06200_);
  and (_09105_, _09104_, _02763_);
  nor (_09106_, _09104_, _02763_);
  nor (_09107_, _09106_, _09105_);
  nor (_09108_, _06198_, \oc8051_golden_model_1.PC [10]);
  nor (_09109_, _09108_, _06191_);
  and (_09110_, _09109_, _02763_);
  nor (_09111_, _09109_, _02763_);
  nor (_09112_, _09111_, _09110_);
  and (_09113_, _09112_, _09107_);
  nor (_09114_, _06197_, \oc8051_golden_model_1.PC [9]);
  nor (_09115_, _09114_, _06198_);
  and (_09116_, _09115_, _02763_);
  nor (_09117_, _09115_, _02763_);
  nor (_09118_, _09117_, _09116_);
  and (_09119_, _05368_, _02763_);
  nor (_09120_, _05368_, _02763_);
  and (_09121_, _05253_, _02626_);
  nor (_09122_, _09121_, \oc8051_golden_model_1.PC [6]);
  nor (_09123_, _09122_, _05365_);
  not (_09124_, _09123_);
  nor (_09125_, _09124_, _02927_);
  and (_09126_, _09124_, _02927_);
  nor (_09127_, _09126_, _09125_);
  and (_09128_, _02626_, \oc8051_golden_model_1.PC [4]);
  nor (_09129_, _09128_, \oc8051_golden_model_1.PC [5]);
  nor (_09130_, _09129_, _09121_);
  not (_09131_, _09130_);
  nor (_09132_, _09131_, _03211_);
  and (_09133_, _09131_, _03211_);
  nor (_09134_, _02626_, \oc8051_golden_model_1.PC [4]);
  nor (_09135_, _09134_, _09128_);
  not (_09136_, _09135_);
  nor (_09137_, _09136_, _03629_);
  nor (_09138_, _02794_, _02641_);
  and (_09139_, _02794_, _02641_);
  not (_09140_, _02648_);
  nor (_09141_, _03256_, _09140_);
  nor (_09142_, _03665_, \oc8051_golden_model_1.PC [1]);
  and (_09143_, _02835_, \oc8051_golden_model_1.PC [0]);
  and (_09144_, _03665_, \oc8051_golden_model_1.PC [1]);
  nor (_09145_, _09144_, _09142_);
  and (_09146_, _09145_, _09143_);
  nor (_09147_, _09146_, _09142_);
  and (_09148_, _03256_, _09140_);
  nor (_09149_, _09148_, _09141_);
  not (_09150_, _09149_);
  nor (_09151_, _09150_, _09147_);
  nor (_09152_, _09151_, _09141_);
  nor (_09153_, _09152_, _09139_);
  nor (_09154_, _09153_, _09138_);
  and (_09155_, _09136_, _03629_);
  nor (_09156_, _09155_, _09137_);
  not (_09157_, _09156_);
  nor (_09158_, _09157_, _09154_);
  nor (_09159_, _09158_, _09137_);
  nor (_09160_, _09159_, _09133_);
  nor (_09161_, _09160_, _09132_);
  not (_09162_, _09161_);
  and (_09163_, _09162_, _09127_);
  nor (_09164_, _09163_, _09125_);
  nor (_09165_, _09164_, _09120_);
  or (_09166_, _09165_, _09119_);
  nor (_09167_, _05366_, \oc8051_golden_model_1.PC [8]);
  nor (_09168_, _09167_, _06197_);
  and (_09169_, _09168_, _02763_);
  nor (_09170_, _09168_, _02763_);
  nor (_09171_, _09170_, _09169_);
  and (_09172_, _09171_, _09166_);
  and (_09173_, _09172_, _09118_);
  and (_09174_, _09173_, _09113_);
  nor (_09175_, _09169_, _09116_);
  not (_09176_, _09175_);
  and (_09177_, _09176_, _09113_);
  or (_09178_, _09177_, _09110_);
  or (_09179_, _09178_, _09174_);
  nor (_09180_, _09179_, _09105_);
  not (_09181_, _09180_);
  nor (_09182_, _09101_, _02763_);
  nor (_09183_, _09182_, _09102_);
  and (_09184_, _09183_, _09181_);
  nor (_09185_, _09184_, _09102_);
  nor (_09186_, _09185_, _09099_);
  nor (_09187_, _09186_, _09098_);
  not (_09188_, _09187_);
  and (_09189_, _09188_, _09089_);
  nor (_09190_, _09189_, _09087_);
  nor (_09191_, _06205_, _02763_);
  and (_09192_, _06205_, _02763_);
  nor (_09193_, _09192_, _09191_);
  and (_09194_, _09193_, _09190_);
  nor (_09195_, _09193_, _09190_);
  nor (_09196_, _09195_, _09194_);
  nor (_09197_, _09196_, _08165_);
  or (_09198_, _09197_, _09084_);
  and (_09199_, _09198_, _09083_);
  nor (_09200_, _06784_, _02546_);
  nor (_09201_, _09200_, _09061_);
  and (_09202_, _06189_, _02579_);
  not (_09203_, _09200_);
  nor (_09204_, _06205_, _02857_);
  or (_09205_, _09204_, _02579_);
  nor (_09206_, _06179_, \oc8051_golden_model_1.PC [14]);
  nor (_09207_, _09206_, _06180_);
  and (_09208_, _09207_, _05661_);
  nor (_09209_, _09207_, _05661_);
  nor (_09210_, _09209_, _09208_);
  nor (_09211_, _06185_, \oc8051_golden_model_1.PC [13]);
  nor (_09212_, _09211_, _06186_);
  not (_09213_, _09212_);
  nor (_09214_, _09213_, _05311_);
  and (_09215_, _09213_, _05311_);
  nor (_09216_, _06177_, \oc8051_golden_model_1.PC [12]);
  nor (_09217_, _09216_, _06178_);
  and (_09218_, _09217_, _05661_);
  not (_09219_, \oc8051_golden_model_1.PC [11]);
  nor (_09220_, _06176_, _09219_);
  and (_09221_, _06176_, _09219_);
  or (_09222_, _09221_, _09220_);
  not (_09223_, _09222_);
  nor (_09224_, _09223_, _05311_);
  and (_09225_, _09223_, _05311_);
  nor (_09226_, _09225_, _09224_);
  nor (_09227_, _06182_, \oc8051_golden_model_1.PC [10]);
  nor (_09228_, _09227_, _06183_);
  not (_09229_, _09228_);
  nor (_09230_, _09229_, _05311_);
  and (_09231_, _09229_, _05311_);
  nor (_09232_, _09231_, _09230_);
  and (_09233_, _09232_, _09226_);
  and (_09234_, _05257_, \oc8051_golden_model_1.PC [8]);
  nor (_09235_, _09234_, \oc8051_golden_model_1.PC [9]);
  nor (_09236_, _09235_, _06182_);
  not (_09237_, _09236_);
  nor (_09238_, _09237_, _05311_);
  and (_09239_, _09237_, _05311_);
  nor (_09240_, _09239_, _09238_);
  nor (_09241_, _05311_, _05260_);
  and (_09242_, _05311_, _05260_);
  and (_09243_, _05255_, _05253_);
  nor (_09244_, _09243_, \oc8051_golden_model_1.PC [6]);
  nor (_09245_, _09244_, _05256_);
  not (_09246_, _09245_);
  nor (_09247_, _09246_, _05649_);
  and (_09248_, _09246_, _05649_);
  nor (_09249_, _09248_, _09247_);
  and (_09250_, _05255_, \oc8051_golden_model_1.PC [4]);
  nor (_09251_, _09250_, \oc8051_golden_model_1.PC [5]);
  nor (_09252_, _09251_, _09243_);
  not (_09253_, _09252_);
  nor (_09254_, _09253_, _05613_);
  and (_09255_, _09253_, _05613_);
  nor (_09256_, _05255_, \oc8051_golden_model_1.PC [4]);
  nor (_09257_, _09256_, _09250_);
  not (_09258_, _09257_);
  nor (_09259_, _09258_, _05582_);
  and (_09260_, _02248_, \oc8051_golden_model_1.PC [2]);
  nor (_09261_, _09260_, \oc8051_golden_model_1.PC [3]);
  nor (_09262_, _09261_, _05255_);
  not (_09263_, _09262_);
  nor (_09264_, _09263_, _03057_);
  and (_09265_, _09263_, _03057_);
  nor (_09266_, _02248_, \oc8051_golden_model_1.PC [2]);
  nor (_09267_, _09266_, _09260_);
  not (_09268_, _09267_);
  nor (_09269_, _09268_, _03297_);
  not (_09270_, _02552_);
  nor (_09271_, _03698_, _09270_);
  nor (_09272_, _03486_, \oc8051_golden_model_1.PC [0]);
  and (_09273_, _03698_, _09270_);
  nor (_09274_, _09273_, _09271_);
  and (_09275_, _09274_, _09272_);
  nor (_09276_, _09275_, _09271_);
  and (_09277_, _09268_, _03297_);
  nor (_09278_, _09277_, _09269_);
  not (_09279_, _09278_);
  nor (_09280_, _09279_, _09276_);
  nor (_09281_, _09280_, _09269_);
  nor (_09282_, _09281_, _09265_);
  nor (_09283_, _09282_, _09264_);
  and (_09284_, _09258_, _05582_);
  nor (_09285_, _09284_, _09259_);
  not (_09286_, _09285_);
  nor (_09287_, _09286_, _09283_);
  nor (_09288_, _09287_, _09259_);
  nor (_09289_, _09288_, _09255_);
  nor (_09290_, _09289_, _09254_);
  not (_09291_, _09290_);
  and (_09292_, _09291_, _09249_);
  nor (_09293_, _09292_, _09247_);
  nor (_09294_, _09293_, _09242_);
  or (_09295_, _09294_, _09241_);
  nor (_09296_, _05257_, \oc8051_golden_model_1.PC [8]);
  nor (_09297_, _09296_, _09234_);
  not (_09298_, _09297_);
  nor (_09299_, _09298_, _05311_);
  and (_09300_, _09298_, _05311_);
  nor (_09301_, _09300_, _09299_);
  and (_09302_, _09301_, _09295_);
  and (_09303_, _09302_, _09240_);
  and (_09304_, _09303_, _09233_);
  nor (_09305_, _09299_, _09238_);
  not (_09306_, _09305_);
  and (_09307_, _09306_, _09233_);
  or (_09308_, _09307_, _09230_);
  or (_09309_, _09308_, _09304_);
  nor (_09310_, _09309_, _09224_);
  not (_09311_, _09310_);
  nor (_09312_, _09217_, _05661_);
  nor (_09313_, _09312_, _09218_);
  and (_09314_, _09313_, _09311_);
  nor (_09315_, _09314_, _09218_);
  nor (_09316_, _09315_, _09215_);
  nor (_09317_, _09316_, _09214_);
  not (_09318_, _09317_);
  and (_09319_, _09318_, _09210_);
  nor (_09320_, _09319_, _09208_);
  not (_09321_, _06189_);
  and (_09322_, _09321_, _05311_);
  nor (_09323_, _09321_, _05311_);
  nor (_09324_, _09323_, _09322_);
  and (_09325_, _09324_, _09320_);
  nor (_09326_, _09324_, _09320_);
  nor (_09327_, _09326_, _09325_);
  nor (_09328_, _05462_, _04551_);
  nor (_09329_, _09328_, _05513_);
  and (_09330_, _05849_, _02927_);
  nor (_09331_, _05849_, _02927_);
  nor (_09332_, _09331_, _09330_);
  and (_09333_, _09332_, _09329_);
  and (_09334_, _06078_, _04638_);
  and (_09335_, _06158_, _03211_);
  nor (_09336_, _09335_, _09334_);
  and (_09337_, _06123_, _04631_);
  and (_09338_, _06159_, _03629_);
  nor (_09339_, _09338_, _09337_);
  and (_09340_, _09339_, _09336_);
  and (_09341_, _09340_, _09333_);
  and (_09342_, _05986_, _02929_);
  and (_09343_, _06154_, _02794_);
  nor (_09344_, _09343_, _09342_);
  and (_09345_, _06031_, _04361_);
  and (_09346_, _06155_, _03256_);
  nor (_09347_, _09346_, _09345_);
  and (_09348_, _09347_, _09344_);
  and (_09349_, _06151_, _03665_);
  and (_09350_, _05895_, _03936_);
  nor (_09351_, _09350_, _09349_);
  and (_09352_, _06152_, _02837_);
  and (_09353_, _05940_, _02835_);
  nor (_09354_, _09353_, _09352_);
  and (_09355_, _09354_, _09351_);
  and (_09356_, _09355_, _09348_);
  and (_09357_, _09356_, _09341_);
  or (_09358_, _09357_, _09327_);
  nand (_09359_, _09357_, _06189_);
  and (_09360_, _09359_, _02978_);
  and (_09361_, _09360_, _09358_);
  nor (_09362_, _04604_, _04551_);
  not (_09363_, _09362_);
  and (_09364_, _09363_, _04605_);
  and (_09365_, _04770_, _02927_);
  nor (_09366_, _04770_, _02927_);
  nor (_09367_, _09366_, _09365_);
  and (_09368_, _09367_, _09364_);
  and (_09369_, _04877_, _03211_);
  nor (_09370_, _04877_, _03211_);
  nor (_09371_, _09370_, _09369_);
  nor (_09372_, _04982_, _03629_);
  and (_09373_, _04982_, _03629_);
  nor (_09374_, _09373_, _09372_);
  and (_09375_, _09374_, _09371_);
  and (_09376_, _09375_, _09368_);
  nor (_09377_, _04241_, _02794_);
  and (_09378_, _04241_, _02794_);
  nor (_09379_, _09378_, _09377_);
  nor (_09380_, _04435_, _03256_);
  and (_09381_, _04435_, _03256_);
  nor (_09382_, _09381_, _09380_);
  and (_09383_, _09382_, _09379_);
  and (_09384_, _04000_, _03665_);
  nor (_09385_, _04000_, _03665_);
  nor (_09386_, _09385_, _09384_);
  and (_09387_, _03808_, _02837_);
  nor (_09388_, _03808_, _02837_);
  nor (_09389_, _09388_, _09387_);
  and (_09390_, _09389_, _09386_);
  and (_09391_, _09390_, _09383_);
  and (_09392_, _09391_, _09376_);
  and (_09393_, _09392_, _09321_);
  and (_09394_, _02848_, _02868_);
  nor (_09395_, _09394_, _02954_);
  and (_09396_, _09395_, _02949_);
  not (_09397_, _09327_);
  nor (_09398_, _09392_, _09397_);
  or (_09399_, _09398_, _09396_);
  nor (_09400_, _09399_, _09393_);
  and (_09401_, _06205_, _03075_);
  and (_09402_, _03076_, _02609_);
  nor (_09403_, _09402_, _06205_);
  and (_09404_, _02879_, _02545_);
  nor (_09405_, _09404_, _07649_);
  not (_09406_, _09405_);
  and (_09407_, _04818_, _04714_);
  and (_09408_, _09407_, _05466_);
  not (_09409_, _05226_);
  and (_09410_, _09409_, _05178_);
  and (_09411_, _05468_, _09410_);
  and (_09412_, _09411_, _09408_);
  and (_09413_, _09412_, _09321_);
  nor (_09414_, _09397_, _09412_);
  or (_09415_, _09414_, _03810_);
  or (_09416_, _09415_, _09413_);
  and (_09417_, _05272_, _05270_);
  and (_09418_, _03808_, _04055_);
  and (_09419_, _09418_, _05244_);
  and (_09420_, _09419_, _09417_);
  nor (_09421_, _09420_, _09196_);
  and (_09422_, _09420_, _06205_);
  or (_09423_, _09422_, _05362_);
  nor (_09424_, _09423_, _09421_);
  not (_09425_, _02616_);
  not (_09426_, _07646_);
  nor (_09427_, _07633_, _03363_);
  nor (_09428_, _02852_, _02429_);
  nor (_09429_, _09428_, _02610_);
  nor (_09430_, _09429_, _07636_);
  and (_09431_, _09430_, _09427_);
  and (_09432_, _09431_, _09426_);
  or (_09433_, _09432_, _09061_);
  nor (_09434_, _03813_, _03818_);
  nand (_09435_, _09434_, _09427_);
  or (_09436_, _03072_, \oc8051_golden_model_1.PC [15]);
  or (_09437_, _07646_, _07636_);
  or (_09438_, _09437_, _09436_);
  or (_09439_, _09438_, _09429_);
  or (_09440_, _09439_, _09435_);
  and (_09441_, _09440_, _09433_);
  or (_09442_, _09441_, _09425_);
  not (_09443_, _06205_);
  and (_09444_, _09434_, _03387_);
  nand (_09445_, _09444_, _02616_);
  nand (_09446_, _09445_, _09443_);
  and (_09447_, _09446_, _09442_);
  nor (_09448_, _09447_, _05363_);
  nor (_09449_, _02886_, _02974_);
  not (_09450_, _09449_);
  or (_09451_, _09450_, _09448_);
  or (_09452_, _09451_, _09424_);
  and (_09453_, _09452_, _09416_);
  or (_09454_, _09453_, _09406_);
  not (_09455_, _09061_);
  and (_09456_, _09405_, _04265_);
  or (_09457_, _09456_, _09455_);
  and (_09458_, _09457_, _09402_);
  and (_09459_, _09458_, _09454_);
  nor (_09460_, _09459_, _09403_);
  nor (_09461_, _09428_, _02620_);
  nor (_09462_, _09461_, _09460_);
  not (_09463_, _09461_);
  nor (_09464_, _09463_, _09061_);
  nor (_09465_, _09464_, _03075_);
  not (_09466_, _09465_);
  nor (_09467_, _09466_, _09462_);
  nor (_09468_, _09467_, _09401_);
  and (_09469_, _02874_, _02545_);
  nor (_09470_, _09469_, _07692_);
  not (_09471_, _09470_);
  nor (_09472_, _09471_, _09468_);
  and (_09473_, _09471_, _09061_);
  not (_09474_, _02621_);
  nor (_09475_, _02875_, _09474_);
  and (_09476_, _09475_, _02877_);
  not (_09477_, _09476_);
  nor (_09478_, _09477_, _09473_);
  not (_09479_, _09478_);
  nor (_09480_, _09479_, _09472_);
  not (_09481_, _09396_);
  nor (_09482_, _09476_, _06205_);
  nor (_09483_, _09482_, _09481_);
  not (_09484_, _09483_);
  nor (_09485_, _09484_, _09480_);
  or (_09486_, _09485_, _02978_);
  nor (_09487_, _09486_, _09400_);
  or (_09488_, _09487_, _09361_);
  and (_09489_, _02868_, _02545_);
  not (_09490_, _09489_);
  and (_09491_, _09490_, _02953_);
  not (_09492_, _09491_);
  nor (_09493_, _09492_, _09488_);
  and (_09494_, _09489_, _09061_);
  not (_09495_, _09494_);
  nor (_09496_, _03059_, _04095_);
  and (_09497_, _09496_, _03064_);
  and (_09498_, _09497_, _03860_);
  and (_09499_, _09498_, _09495_);
  not (_09500_, _02950_);
  nor (_09501_, _07442_, \oc8051_golden_model_1.ACC [3]);
  and (_09502_, _07442_, \oc8051_golden_model_1.ACC [3]);
  nor (_09503_, _09502_, _09501_);
  and (_09504_, _09503_, _08087_);
  nor (_09505_, _07481_, \oc8051_golden_model_1.ACC [0]);
  and (_09506_, _07481_, \oc8051_golden_model_1.ACC [0]);
  nor (_09507_, _09506_, _09505_);
  and (_09508_, _09507_, _07576_);
  and (_09509_, _09508_, _09504_);
  and (_09510_, _08078_, _08082_);
  not (_09511_, _08070_);
  and (_09512_, _08074_, _09511_);
  and (_09513_, _09512_, _09510_);
  and (_09514_, _09513_, _09509_);
  nor (_09515_, _09514_, _09327_);
  and (_09516_, _09514_, _06189_);
  nor (_09517_, _09516_, _09515_);
  nor (_09518_, _09517_, _09500_);
  or (_09519_, _08125_, _08124_);
  and (_09520_, _09519_, _08128_);
  and (_09521_, _02837_, _02667_);
  nor (_09522_, _09521_, _08132_);
  nor (_09523_, _09522_, _08131_);
  and (_09524_, _09523_, _09520_);
  nor (_09525_, _08119_, _08123_);
  nor (_09526_, _08116_, _07896_);
  and (_09527_, _09526_, _09525_);
  and (_09528_, _09527_, _09524_);
  not (_09529_, _09528_);
  and (_09530_, _09529_, _09327_);
  not (_09531_, _02952_);
  and (_09532_, _09528_, _09321_);
  nor (_09533_, _09532_, _09531_);
  not (_09534_, _09533_);
  nor (_09535_, _09534_, _09530_);
  nor (_09536_, _09535_, _09518_);
  and (_09537_, _09536_, _09499_);
  not (_09538_, _09537_);
  nor (_09539_, _09538_, _09493_);
  and (_09540_, _03099_, _02578_);
  not (_09541_, _09540_);
  nor (_09542_, _08224_, _06247_);
  and (_09543_, _09542_, _09541_);
  not (_09544_, _09543_);
  nor (_09545_, _09498_, _06205_);
  nor (_09546_, _09545_, _09544_);
  not (_09547_, _09546_);
  nor (_09548_, _09547_, _09539_);
  nor (_09549_, _09543_, _09455_);
  not (_09550_, _03101_);
  not (_09551_, _02619_);
  nor (_09552_, _03100_, _09551_);
  and (_09553_, _09552_, _09550_);
  not (_09554_, _09553_);
  or (_09555_, _09554_, _09549_);
  or (_09556_, _09555_, _09548_);
  and (_09557_, _07718_, _07626_);
  or (_09558_, _09553_, _06205_);
  and (_09559_, _09558_, _09557_);
  and (_09560_, _09559_, _09556_);
  nor (_09561_, _07404_, _03106_);
  not (_09562_, _09561_);
  nor (_09563_, _09557_, _09455_);
  nor (_09564_, _09563_, _09562_);
  not (_09565_, _09564_);
  nor (_09566_, _09565_, _09560_);
  nor (_09567_, _09561_, _06205_);
  nor (_09568_, _09567_, _02583_);
  not (_09569_, _09568_);
  nor (_09570_, _09569_, _09566_);
  and (_09571_, _09061_, _02583_);
  nor (_09572_, _02863_, _02581_);
  not (_09573_, _09572_);
  nor (_09574_, _09573_, _09571_);
  not (_09575_, _09574_);
  nor (_09576_, _09575_, _09570_);
  nor (_09577_, _09572_, _06205_);
  nor (_09578_, _09577_, _02981_);
  not (_09580_, _09578_);
  nor (_09581_, _09580_, _09576_);
  not (_09582_, _02857_);
  and (_09583_, _06189_, _02981_);
  nor (_09584_, _09583_, _09582_);
  not (_09585_, _09584_);
  nor (_09586_, _09585_, _09581_);
  nor (_09587_, _09586_, _09205_);
  or (_09588_, _09587_, _09203_);
  nor (_09589_, _09588_, _09202_);
  nor (_09590_, _09589_, _09201_);
  nor (_09591_, _02933_, _02518_);
  not (_09592_, _09591_);
  nor (_09593_, _09592_, _09590_);
  and (_09594_, _02496_, _02517_);
  nor (_09595_, _09591_, _06205_);
  nor (_09596_, _09595_, _09594_);
  not (_09597_, _09596_);
  nor (_09598_, _09597_, _09593_);
  not (_09599_, _09594_);
  nor (_09601_, _09599_, _09196_);
  nor (_09602_, _09601_, _05754_);
  not (_09603_, _09602_);
  or (_09604_, _09603_, _09598_);
  nor (_09605_, _06205_, _05753_);
  nor (_09606_, _09605_, _02802_);
  nand (_09607_, _09606_, _09604_);
  and (_09608_, _06189_, _02802_);
  nor (_09609_, _09608_, _07859_);
  nand (_09610_, _09609_, _09607_);
  and (_09611_, _02545_, _02513_);
  nor (_09612_, _07860_, _06205_);
  nor (_09613_, _09612_, _09611_);
  nand (_09614_, _09613_, _09610_);
  and (_09615_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_09616_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_09617_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09618_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09619_, _09618_, _09617_);
  and (_09620_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09621_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09622_, _09621_, _09620_);
  not (_09623_, _09622_);
  and (_09624_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09625_, _02600_, _02596_);
  nor (_09626_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09627_, _09626_, _09624_);
  not (_09628_, _09627_);
  nor (_09629_, _09628_, _09625_);
  nor (_09630_, _09629_, _09624_);
  nor (_09631_, _09630_, _09623_);
  nor (_09632_, _09631_, _09620_);
  not (_09633_, _09632_);
  and (_09634_, _09633_, _09619_);
  nor (_09635_, _09634_, _09617_);
  nor (_09636_, _09635_, _09616_);
  or (_09637_, _09636_, _09615_);
  and (_09638_, _09637_, \oc8051_golden_model_1.DPH [0]);
  and (_09639_, _09638_, \oc8051_golden_model_1.DPH [1]);
  and (_09640_, _09639_, \oc8051_golden_model_1.DPH [2]);
  and (_09641_, _09640_, \oc8051_golden_model_1.DPH [3]);
  and (_09642_, _09641_, \oc8051_golden_model_1.DPH [4]);
  and (_09643_, _09642_, \oc8051_golden_model_1.DPH [5]);
  and (_09644_, _09643_, \oc8051_golden_model_1.DPH [6]);
  or (_09645_, _09644_, \oc8051_golden_model_1.DPH [7]);
  nand (_09646_, _09644_, \oc8051_golden_model_1.DPH [7]);
  and (_09647_, _09646_, _09645_);
  and (_09648_, _09647_, _09611_);
  nor (_09649_, _02932_, _02514_);
  not (_09650_, _09649_);
  nor (_09651_, _09650_, _09648_);
  nand (_09652_, _09651_, _09614_);
  nor (_09653_, _09649_, _06205_);
  nor (_09654_, _09653_, _09083_);
  and (_09655_, _09654_, _09652_);
  or (_09656_, _09655_, _09199_);
  and (_09657_, _07875_, _07880_);
  nand (_09658_, _09657_, _09656_);
  nor (_09659_, _09657_, _09455_);
  nor (_09660_, _07399_, _03129_);
  not (_09661_, _09660_);
  nor (_09662_, _09661_, _09659_);
  nand (_09663_, _09662_, _09658_);
  nor (_09664_, _09660_, _06205_);
  nor (_09665_, _09664_, _02980_);
  nand (_09666_, _09665_, _09663_);
  and (_09667_, _06189_, _02980_);
  nor (_09668_, _03127_, _02509_);
  not (_09669_, _09668_);
  nor (_09670_, _09669_, _09667_);
  nand (_09671_, _09670_, _09666_);
  and (_09672_, _02496_, _02508_);
  nor (_09673_, _09668_, _06205_);
  nor (_09674_, _09673_, _09672_);
  nand (_09675_, _09674_, _09671_);
  not (_09676_, _08165_);
  and (_09677_, _09676_, _06205_);
  nor (_09678_, _09196_, _09676_);
  or (_09679_, _09678_, _09677_);
  and (_09680_, _09679_, _09672_);
  not (_09681_, _09081_);
  nor (_09682_, _09681_, _09680_);
  and (_09683_, _09682_, _09675_);
  or (_09684_, _09683_, _09082_);
  nand (_09685_, _09684_, _09080_);
  nor (_09686_, _09080_, _06205_);
  nor (_09687_, _09686_, _02970_);
  nand (_09688_, _09687_, _09685_);
  not (_09689_, _09077_);
  and (_09690_, _06189_, _02970_);
  nor (_09691_, _09690_, _09689_);
  and (_09692_, _09691_, _09688_);
  or (_09693_, _09692_, _09079_);
  not (_09694_, _09074_);
  and (_09695_, _06205_, \oc8051_golden_model_1.PSW [7]);
  nor (_09696_, _09196_, \oc8051_golden_model_1.PSW [7]);
  or (_09697_, _09696_, _09695_);
  and (_09698_, _09697_, _09076_);
  nor (_09699_, _09698_, _09694_);
  and (_09700_, _09699_, _09693_);
  or (_09701_, _09700_, _09075_);
  nand (_09702_, _09701_, _07943_);
  nor (_09703_, _07943_, _06205_);
  nor (_09704_, _09703_, _02965_);
  nand (_09705_, _09704_, _09702_);
  not (_09706_, _09070_);
  and (_09707_, _06189_, _02965_);
  nor (_09708_, _09707_, _09706_);
  and (_09709_, _09708_, _09705_);
  or (_09710_, _09709_, _09072_);
  not (_09711_, _09066_);
  and (_09712_, _06205_, _07293_);
  nor (_09713_, _09196_, _07293_);
  or (_09714_, _09713_, _09712_);
  and (_09715_, _09714_, _09068_);
  nor (_09716_, _09715_, _09711_);
  and (_09717_, _09716_, _09710_);
  or (_09718_, _09717_, _09067_);
  nand (_09719_, _09718_, _09065_);
  nor (_09720_, _09065_, _06205_);
  nor (_09721_, _09720_, _07991_);
  and (_09722_, _09721_, _09719_);
  and (_09723_, _09061_, _07991_);
  or (_09724_, _09723_, _03145_);
  nor (_09725_, _09724_, _09722_);
  not (_09726_, _03145_);
  nor (_09727_, _04604_, _09726_);
  or (_09728_, _09727_, _09725_);
  nand (_09729_, _09728_, _02529_);
  nor (_09730_, _06205_, _02529_);
  nor (_09731_, _09730_, _02968_);
  nand (_09732_, _09731_, _09729_);
  not (_09733_, _04611_);
  and (_09734_, _05338_, \oc8051_golden_model_1.SCON [2]);
  and (_09735_, _05340_, \oc8051_golden_model_1.IE [2]);
  nor (_09736_, _09735_, _09734_);
  and (_09737_, _05320_, \oc8051_golden_model_1.TCON [2]);
  and (_09738_, _05349_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_09739_, _09738_, _09737_);
  and (_09740_, _09739_, _09736_);
  and (_09741_, _05331_, \oc8051_golden_model_1.PSW [2]);
  and (_09742_, _05333_, \oc8051_golden_model_1.B [2]);
  nor (_09743_, _09742_, _09741_);
  and (_09744_, _05328_, \oc8051_golden_model_1.IP [2]);
  and (_09745_, _05325_, \oc8051_golden_model_1.ACC [2]);
  nor (_09746_, _09745_, _09744_);
  and (_09747_, _09746_, _09743_);
  and (_09748_, _05344_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09749_, _05347_, \oc8051_golden_model_1.P2INREG [2]);
  and (_09750_, _04609_, \oc8051_golden_model_1.P0INREG [2]);
  or (_09751_, _09750_, _09749_);
  nor (_09752_, _09751_, _09748_);
  and (_09753_, _09752_, _09747_);
  and (_09754_, _09753_, _09740_);
  and (_09755_, _09754_, _05080_);
  nor (_09756_, _09755_, _09733_);
  not (_09757_, _04616_);
  and (_09758_, _05320_, \oc8051_golden_model_1.TCON [1]);
  and (_09759_, _05333_, \oc8051_golden_model_1.B [1]);
  nor (_09760_, _09759_, _09758_);
  and (_09761_, _05328_, \oc8051_golden_model_1.IP [1]);
  not (_09762_, _09761_);
  and (_09763_, _05331_, \oc8051_golden_model_1.PSW [1]);
  and (_09764_, _05325_, \oc8051_golden_model_1.ACC [1]);
  nor (_09765_, _09764_, _09763_);
  and (_09766_, _09765_, _09762_);
  and (_09767_, _09766_, _09760_);
  and (_09768_, _05338_, \oc8051_golden_model_1.SCON [1]);
  and (_09769_, _05340_, \oc8051_golden_model_1.IE [1]);
  nor (_09770_, _09769_, _09768_);
  and (_09771_, _04609_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09772_, _05347_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09773_, _09772_, _09771_);
  and (_09774_, _05344_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09775_, _05349_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09776_, _09775_, _09774_);
  and (_09777_, _09776_, _09773_);
  and (_09778_, _09777_, _09770_);
  and (_09779_, _09778_, _09767_);
  and (_09780_, _09779_, _05131_);
  nor (_09781_, _09780_, _09757_);
  nor (_09782_, _09781_, _09756_);
  and (_09783_, _04619_, _04361_);
  not (_09784_, _09783_);
  and (_09785_, _05320_, \oc8051_golden_model_1.TCON [4]);
  and (_09786_, _05325_, \oc8051_golden_model_1.ACC [4]);
  nor (_09787_, _09786_, _09785_);
  and (_09788_, _05328_, \oc8051_golden_model_1.IP [4]);
  not (_09789_, _09788_);
  and (_09790_, _05331_, \oc8051_golden_model_1.PSW [4]);
  and (_09791_, _05333_, \oc8051_golden_model_1.B [4]);
  nor (_09792_, _09791_, _09790_);
  and (_09793_, _09792_, _09789_);
  and (_09794_, _09793_, _09787_);
  and (_09795_, _05338_, \oc8051_golden_model_1.SCON [4]);
  and (_09796_, _05340_, \oc8051_golden_model_1.IE [4]);
  nor (_09797_, _09796_, _09795_);
  and (_09798_, _04609_, \oc8051_golden_model_1.P0INREG [4]);
  and (_09799_, _05347_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_09800_, _09799_, _09798_);
  and (_09801_, _05344_, \oc8051_golden_model_1.P1INREG [4]);
  and (_09802_, _05349_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09803_, _09802_, _09801_);
  and (_09804_, _09803_, _09800_);
  and (_09805_, _09804_, _09797_);
  and (_09806_, _09805_, _09794_);
  and (_09807_, _09806_, _04983_);
  nor (_09808_, _09807_, _09784_);
  nor (_09809_, _05527_, _05359_);
  nor (_09810_, _09809_, _09808_);
  and (_09811_, _09810_, _09782_);
  not (_09812_, _04620_);
  and (_09813_, _05320_, \oc8051_golden_model_1.TCON [0]);
  and (_09814_, _05325_, \oc8051_golden_model_1.ACC [0]);
  nor (_09815_, _09814_, _09813_);
  and (_09816_, _05331_, \oc8051_golden_model_1.PSW [0]);
  not (_09817_, _09816_);
  and (_09818_, _05328_, \oc8051_golden_model_1.IP [0]);
  and (_09819_, _05333_, \oc8051_golden_model_1.B [0]);
  nor (_09820_, _09819_, _09818_);
  and (_09821_, _09820_, _09817_);
  and (_09822_, _09821_, _09815_);
  and (_09823_, _05338_, \oc8051_golden_model_1.SCON [0]);
  and (_09824_, _05340_, \oc8051_golden_model_1.IE [0]);
  nor (_09825_, _09824_, _09823_);
  and (_09826_, _04609_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09827_, _05347_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09828_, _09827_, _09826_);
  and (_09829_, _05344_, \oc8051_golden_model_1.P1INREG [0]);
  and (_09830_, _05349_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09831_, _09830_, _09829_);
  and (_09832_, _09831_, _09828_);
  and (_09833_, _09832_, _09825_);
  and (_09834_, _09833_, _09822_);
  and (_09835_, _09834_, _05179_);
  nor (_09836_, _09835_, _09812_);
  and (_09837_, _04610_, _04361_);
  not (_09838_, _09837_);
  and (_09839_, _05338_, \oc8051_golden_model_1.SCON [6]);
  and (_09840_, _05340_, \oc8051_golden_model_1.IE [6]);
  nor (_09841_, _09840_, _09839_);
  and (_09842_, _05320_, \oc8051_golden_model_1.TCON [6]);
  and (_09843_, _05349_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09844_, _09843_, _09842_);
  and (_09845_, _09844_, _09841_);
  and (_09846_, _05331_, \oc8051_golden_model_1.PSW [6]);
  and (_09847_, _05333_, \oc8051_golden_model_1.B [6]);
  nor (_09848_, _09847_, _09846_);
  and (_09849_, _05328_, \oc8051_golden_model_1.IP [6]);
  and (_09850_, _05325_, \oc8051_golden_model_1.ACC [6]);
  nor (_09851_, _09850_, _09849_);
  and (_09852_, _09851_, _09848_);
  and (_09853_, _05344_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09854_, _05347_, \oc8051_golden_model_1.P2INREG [6]);
  and (_09855_, _04609_, \oc8051_golden_model_1.P0INREG [6]);
  or (_09856_, _09855_, _09854_);
  nor (_09857_, _09856_, _09853_);
  and (_09858_, _09857_, _09852_);
  and (_09859_, _09858_, _09845_);
  and (_09860_, _09859_, _04771_);
  nor (_09861_, _09860_, _09838_);
  nor (_09862_, _09861_, _09836_);
  not (_09863_, _04670_);
  and (_09864_, _05338_, \oc8051_golden_model_1.SCON [3]);
  and (_09865_, _05340_, \oc8051_golden_model_1.IE [3]);
  nor (_09866_, _09865_, _09864_);
  and (_09867_, _05320_, \oc8051_golden_model_1.TCON [3]);
  and (_09868_, _05349_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_09869_, _09868_, _09867_);
  and (_09870_, _09869_, _09866_);
  and (_09871_, _05331_, \oc8051_golden_model_1.PSW [3]);
  and (_09872_, _05325_, \oc8051_golden_model_1.ACC [3]);
  nor (_09873_, _09872_, _09871_);
  and (_09874_, _05328_, \oc8051_golden_model_1.IP [3]);
  and (_09875_, _05333_, \oc8051_golden_model_1.B [3]);
  nor (_09876_, _09875_, _09874_);
  and (_09877_, _09876_, _09873_);
  and (_09878_, _05344_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09879_, _05347_, \oc8051_golden_model_1.P2INREG [3]);
  and (_09880_, _04609_, \oc8051_golden_model_1.P0INREG [3]);
  or (_09881_, _09880_, _09879_);
  nor (_09882_, _09881_, _09878_);
  and (_09883_, _09882_, _09877_);
  and (_09884_, _09883_, _09870_);
  and (_09885_, _09884_, _05032_);
  nor (_09886_, _09885_, _09863_);
  and (_09887_, _04615_, _04361_);
  not (_09888_, _09887_);
  and (_09889_, _05320_, \oc8051_golden_model_1.TCON [5]);
  and (_09890_, _05325_, \oc8051_golden_model_1.ACC [5]);
  nor (_09891_, _09890_, _09889_);
  and (_09892_, _05331_, \oc8051_golden_model_1.PSW [5]);
  not (_09893_, _09892_);
  and (_09894_, _05328_, \oc8051_golden_model_1.IP [5]);
  and (_09895_, _05333_, \oc8051_golden_model_1.B [5]);
  nor (_09896_, _09895_, _09894_);
  and (_09897_, _09896_, _09893_);
  and (_09898_, _09897_, _09891_);
  and (_09899_, _05338_, \oc8051_golden_model_1.SCON [5]);
  and (_09900_, _05340_, \oc8051_golden_model_1.IE [5]);
  nor (_09901_, _09900_, _09899_);
  and (_09902_, _04609_, \oc8051_golden_model_1.P0INREG [5]);
  and (_09903_, _05347_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_09904_, _09903_, _09902_);
  and (_09905_, _05344_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09906_, _05349_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09907_, _09906_, _09905_);
  and (_09908_, _09907_, _09904_);
  and (_09909_, _09908_, _09901_);
  and (_09910_, _09909_, _09898_);
  and (_09911_, _09910_, _04878_);
  nor (_09912_, _09911_, _09888_);
  nor (_09913_, _09912_, _09886_);
  and (_09914_, _09913_, _09862_);
  and (_09915_, _09914_, _09811_);
  nor (_09916_, _09915_, _06189_);
  and (_09917_, _09915_, _09327_);
  or (_09918_, _09917_, _03561_);
  or (_09919_, _09918_, _09916_);
  and (_09920_, _09919_, _09063_);
  and (_09921_, _09920_, _09732_);
  or (_09922_, _09921_, _09064_);
  nand (_09923_, _09922_, _08066_);
  nor (_09924_, _08066_, _06205_);
  nor (_09925_, _09924_, _08111_);
  and (_09926_, _09925_, _09923_);
  and (_09927_, _09061_, _08111_);
  or (_09928_, _09927_, _02892_);
  nor (_09929_, _09928_, _09926_);
  nor (_09930_, _04604_, _02893_);
  or (_09931_, _09930_, _09929_);
  nand (_09932_, _09931_, _02537_);
  nor (_09933_, _06205_, _02537_);
  nor (_09934_, _09933_, _02940_);
  nand (_09935_, _09934_, _09932_);
  nor (_09936_, _09915_, _09397_);
  and (_09937_, _09915_, _09321_);
  nor (_09938_, _09937_, _09936_);
  and (_09939_, _09938_, _02940_);
  and (_09940_, _05268_, _05262_);
  and (_09941_, _09940_, _03909_);
  not (_09942_, _09941_);
  nor (_09943_, _09942_, _09939_);
  nand (_09944_, _09943_, _09935_);
  nor (_09945_, _09941_, _09061_);
  nor (_09946_, _09945_, _03163_);
  nand (_09947_, _09946_, _09944_);
  nor (_09948_, _08159_, _08154_);
  not (_09949_, _09948_);
  and (_09950_, _06205_, _03163_);
  nor (_09951_, _09950_, _09949_);
  nand (_09952_, _09951_, _09947_);
  nor (_09953_, _09061_, _09948_);
  nor (_09954_, _09953_, _02939_);
  and (_09955_, _09954_, _09952_);
  and (_09956_, _02939_, _02763_);
  or (_09957_, _09956_, _02525_);
  or (_09958_, _09957_, _09955_);
  nor (_09959_, _06205_, _02526_);
  nor (_09960_, _09959_, _02497_);
  nand (_09961_, _09960_, _09958_);
  and (_09962_, _09938_, _02497_);
  not (_09963_, _09428_);
  and (_09964_, _09963_, _02522_);
  nor (_09965_, _09964_, _09962_);
  nand (_09966_, _09965_, _09961_);
  and (_09967_, _09964_, _09455_);
  nor (_09968_, _09967_, _02888_);
  nand (_09969_, _09968_, _09966_);
  not (_09970_, _09044_);
  and (_09971_, _06205_, _02888_);
  nor (_09972_, _09971_, _09970_);
  and (_09973_, _09972_, _09969_);
  or (_09974_, _09973_, _09062_);
  nand (_09975_, _09974_, _09043_);
  nor (_09976_, _09043_, _02763_);
  nor (_09977_, _09976_, _02523_);
  nand (_09978_, _09977_, _09975_);
  and (_09979_, _02496_, _02522_);
  and (_09980_, _06205_, _02523_);
  nor (_09981_, _09980_, _09979_);
  and (_09982_, _09981_, _09978_);
  not (_09983_, _09979_);
  nor (_09984_, _09061_, _09983_);
  nor (_09985_, _09984_, _09982_);
  or (_09986_, _09985_, _42672_);
  or (_09987_, _42668_, \oc8051_golden_model_1.PC [15]);
  and (_09988_, _09987_, _43998_);
  and (_40497_, _09988_, _09986_);
  and (_09989_, _07323_, _05245_);
  nor (_09990_, _07327_, _05771_);
  or (_09991_, _09990_, _07389_);
  or (_09992_, _09991_, _09989_);
  nor (_09993_, _09992_, _07322_);
  nor (_09994_, _04690_, _07293_);
  and (_09995_, _05774_, _04690_);
  nor (_09996_, _09995_, _09994_);
  nor (_09997_, _09996_, _03128_);
  not (_09998_, _04690_);
  nor (_09999_, _05744_, _09998_);
  nor (_10000_, _09999_, _09994_);
  nor (_10001_, _10000_, _02838_);
  and (_10002_, _04690_, _04604_);
  nor (_10003_, _10002_, _09994_);
  and (_10004_, _10003_, _06770_);
  not (_10005_, _05497_);
  and (_10006_, _07520_, _10005_);
  and (_10007_, _07530_, _07526_);
  nor (_10008_, _10007_, _07524_);
  and (_10009_, _07964_, _07526_);
  not (_10010_, _10009_);
  nor (_10011_, _10010_, _07591_);
  not (_10012_, _10011_);
  and (_10013_, _10012_, _10008_);
  or (_10014_, _10013_, _10006_);
  and (_10015_, _10014_, _03106_);
  not (_10016_, _03100_);
  and (_10017_, _04609_, \oc8051_golden_model_1.P0 [2]);
  and (_10018_, _05344_, \oc8051_golden_model_1.P1 [2]);
  nor (_10019_, _10018_, _10017_);
  and (_10020_, _05349_, \oc8051_golden_model_1.P3 [2]);
  and (_10021_, _05347_, \oc8051_golden_model_1.P2 [2]);
  or (_10022_, _10021_, _10020_);
  nor (_10023_, _10022_, _09737_);
  and (_10024_, _10023_, _09747_);
  and (_10025_, _10024_, _09736_);
  and (_10026_, _10025_, _10019_);
  and (_10027_, _10026_, _05080_);
  nor (_10028_, _10027_, _09733_);
  and (_10029_, _05347_, \oc8051_golden_model_1.P2 [1]);
  and (_10030_, _05349_, \oc8051_golden_model_1.P3 [1]);
  nor (_10031_, _10030_, _10029_);
  and (_10032_, _04609_, \oc8051_golden_model_1.P0 [1]);
  and (_10033_, _05344_, \oc8051_golden_model_1.P1 [1]);
  nor (_10034_, _10033_, _10032_);
  and (_10035_, _10034_, _10031_);
  and (_10036_, _10035_, _09770_);
  and (_10037_, _10036_, _09767_);
  and (_10038_, _10037_, _05131_);
  nor (_10039_, _10038_, _09757_);
  nor (_10040_, _10039_, _10028_);
  and (_10041_, _05347_, \oc8051_golden_model_1.P2 [4]);
  and (_10042_, _05349_, \oc8051_golden_model_1.P3 [4]);
  nor (_10043_, _10042_, _10041_);
  and (_10044_, _04609_, \oc8051_golden_model_1.P0 [4]);
  and (_10045_, _05344_, \oc8051_golden_model_1.P1 [4]);
  nor (_10046_, _10045_, _10044_);
  and (_10047_, _10046_, _10043_);
  and (_10048_, _10047_, _09797_);
  and (_10049_, _10048_, _09794_);
  and (_10050_, _10049_, _04983_);
  nor (_10051_, _09784_, _10050_);
  nor (_10052_, _10051_, _05501_);
  and (_10053_, _10052_, _10040_);
  and (_10054_, _05347_, \oc8051_golden_model_1.P2 [0]);
  and (_10055_, _05349_, \oc8051_golden_model_1.P3 [0]);
  nor (_10056_, _10055_, _10054_);
  and (_10057_, _04609_, \oc8051_golden_model_1.P0 [0]);
  and (_10058_, _05344_, \oc8051_golden_model_1.P1 [0]);
  nor (_10059_, _10058_, _10057_);
  and (_10060_, _10059_, _10056_);
  and (_10061_, _10060_, _09825_);
  and (_10062_, _10061_, _09822_);
  and (_10063_, _10062_, _05179_);
  nor (_10064_, _10063_, _09812_);
  and (_10065_, _04609_, \oc8051_golden_model_1.P0 [6]);
  and (_10066_, _05344_, \oc8051_golden_model_1.P1 [6]);
  nor (_10067_, _10066_, _10065_);
  and (_10068_, _05349_, \oc8051_golden_model_1.P3 [6]);
  and (_10069_, _05347_, \oc8051_golden_model_1.P2 [6]);
  or (_10070_, _10069_, _10068_);
  nor (_10071_, _10070_, _09842_);
  and (_10072_, _10071_, _09852_);
  and (_10073_, _10072_, _09841_);
  and (_10074_, _10073_, _10067_);
  and (_10075_, _10074_, _04771_);
  nor (_10076_, _09838_, _10075_);
  nor (_10077_, _10076_, _10064_);
  and (_10078_, _04609_, \oc8051_golden_model_1.P0 [3]);
  and (_10079_, _05344_, \oc8051_golden_model_1.P1 [3]);
  nor (_10080_, _10079_, _10078_);
  and (_10081_, _05349_, \oc8051_golden_model_1.P3 [3]);
  and (_10082_, _05347_, \oc8051_golden_model_1.P2 [3]);
  or (_10083_, _10082_, _10081_);
  nor (_10084_, _10083_, _09867_);
  and (_10085_, _10084_, _09877_);
  and (_10086_, _10085_, _09866_);
  and (_10087_, _10086_, _10080_);
  and (_10088_, _10087_, _05032_);
  nor (_10089_, _10088_, _09863_);
  and (_10090_, _05347_, \oc8051_golden_model_1.P2 [5]);
  and (_10091_, _05349_, \oc8051_golden_model_1.P3 [5]);
  nor (_10092_, _10091_, _10090_);
  and (_10093_, _04609_, \oc8051_golden_model_1.P0 [5]);
  and (_10094_, _05344_, \oc8051_golden_model_1.P1 [5]);
  nor (_10095_, _10094_, _10093_);
  and (_10096_, _10095_, _10092_);
  and (_10097_, _10096_, _09901_);
  and (_10098_, _10097_, _09898_);
  and (_10099_, _10098_, _04878_);
  nor (_10100_, _09888_, _10099_);
  nor (_10101_, _10100_, _10089_);
  and (_10102_, _10101_, _10077_);
  and (_10103_, _10102_, _10053_);
  nor (_10104_, _10103_, \oc8051_golden_model_1.PSW [7]);
  nor (_10105_, _10104_, _10016_);
  not (_10106_, _07718_);
  nor (_10107_, _09915_, _09550_);
  and (_10108_, _05474_, _04690_);
  nor (_10109_, _10108_, _09994_);
  and (_10110_, _10109_, _02974_);
  and (_10111_, _04690_, \oc8051_golden_model_1.ACC [7]);
  nor (_10112_, _10111_, _09994_);
  nor (_10113_, _10112_, _03814_);
  nor (_10114_, _03813_, _07293_);
  or (_10115_, _10114_, _02974_);
  nor (_10116_, _10115_, _10113_);
  nor (_10117_, _10116_, _07649_);
  not (_10118_, _10117_);
  nor (_10119_, _10118_, _10110_);
  nor (_10120_, _07659_, \oc8051_golden_model_1.PSW [7]);
  not (_10121_, _10120_);
  nor (_10122_, _10121_, _07669_);
  not (_10123_, _10122_);
  and (_10124_, _10123_, _07649_);
  not (_10125_, _09404_);
  nand (_10126_, _10125_, _03076_);
  or (_10127_, _10126_, _10124_);
  or (_10128_, _10127_, _10119_);
  nor (_10129_, _05331_, _07293_);
  and (_10130_, _05360_, _05331_);
  nor (_10131_, _10130_, _10129_);
  and (_10132_, _10131_, _02880_);
  and (_10133_, _10003_, _03069_);
  nor (_10134_, _10133_, _10132_);
  and (_10135_, _10134_, _10128_);
  nor (_10136_, _10135_, _03075_);
  and (_10137_, _10112_, _03075_);
  or (_10138_, _09469_, _02876_);
  or (_10139_, _10138_, _10137_);
  nor (_10140_, _10139_, _10136_);
  and (_10141_, _05356_, _05331_);
  nor (_10142_, _10141_, _10129_);
  nor (_10143_, _10142_, _02877_);
  nor (_10144_, _10143_, _10140_);
  nor (_10145_, _10144_, _09481_);
  nand (_10146_, _09366_, _04605_);
  not (_10147_, _09376_);
  nor (_10148_, _09387_, _09384_);
  nor (_10149_, _09385_, _10148_);
  not (_10150_, _10149_);
  and (_10151_, _10150_, _09383_);
  and (_10152_, _09379_, _09380_);
  nor (_10153_, _10152_, _09377_);
  not (_10154_, _10153_);
  nor (_10155_, _10154_, _10151_);
  nor (_10156_, _10155_, _10147_);
  and (_10157_, _09371_, _09372_);
  or (_10158_, _10157_, _09370_);
  and (_10159_, _10158_, _09368_);
  or (_10160_, _10159_, _09362_);
  nor (_10161_, _10160_, _10156_);
  and (_10162_, _10161_, _10146_);
  or (_10163_, _09392_, _09396_);
  nor (_10164_, _10163_, _10162_);
  nor (_10165_, _10164_, _10145_);
  nor (_10166_, _10165_, _02978_);
  not (_10167_, _05513_);
  nor (_10168_, _09337_, _09334_);
  not (_10169_, _10168_);
  nor (_10170_, _09352_, _09349_);
  nor (_10171_, _09350_, _10170_);
  not (_10172_, _10171_);
  and (_10173_, _10172_, _09348_);
  and (_10174_, _09344_, _09345_);
  nor (_10175_, _10174_, _09342_);
  not (_10176_, _10175_);
  nor (_10177_, _10176_, _10173_);
  nor (_10178_, _10177_, _09338_);
  or (_10179_, _10178_, _10169_);
  nor (_10180_, _09335_, _09330_);
  and (_10181_, _10180_, _10179_);
  or (_10182_, _10181_, _09331_);
  and (_10183_, _10182_, _10167_);
  nor (_10184_, _10183_, _09328_);
  nor (_10185_, _09357_, _02979_);
  not (_10186_, _10185_);
  nor (_10187_, _10186_, _10184_);
  nor (_10188_, _10187_, _10166_);
  nor (_10189_, _10188_, _09492_);
  nand (_10190_, _09489_, \oc8051_golden_model_1.PSW [7]);
  nor (_10191_, _05497_, \oc8051_golden_model_1.ACC [7]);
  nor (_10192_, _08081_, _08076_);
  not (_10193_, _07576_);
  nor (_10194_, _09506_, _10193_);
  or (_10195_, _10194_, _07574_);
  and (_10196_, _10195_, _09504_);
  and (_10197_, _09503_, _08086_);
  nor (_10198_, _10197_, _09501_);
  not (_10199_, _10198_);
  nor (_10200_, _10199_, _10196_);
  or (_10201_, _10200_, _08080_);
  nand (_10202_, _10201_, _10192_);
  nor (_10203_, _08077_, _08072_);
  and (_10204_, _10203_, _10202_);
  or (_10205_, _10204_, _08073_);
  and (_10206_, _10205_, _09511_);
  nor (_10207_, _10206_, _10191_);
  nor (_10208_, _09514_, _09500_);
  not (_10209_, _10208_);
  nor (_10210_, _10209_, _10207_);
  nor (_10211_, _02927_, \oc8051_golden_model_1.ACC [6]);
  not (_10212_, _10211_);
  nor (_10213_, _10212_, _07896_);
  and (_10214_, _02763_, _05771_);
  and (_10215_, _03211_, \oc8051_golden_model_1.ACC [5]);
  nor (_10216_, _03211_, \oc8051_golden_model_1.ACC [5]);
  nor (_10217_, _03629_, \oc8051_golden_model_1.ACC [4]);
  nor (_10218_, _10217_, _10216_);
  nor (_10219_, _10218_, _10215_);
  and (_10220_, _10219_, _09526_);
  or (_10221_, _10220_, _10214_);
  nor (_10222_, _10221_, _10213_);
  and (_10223_, _02794_, \oc8051_golden_model_1.ACC [3]);
  nor (_10224_, _02794_, \oc8051_golden_model_1.ACC [3]);
  nor (_10225_, _03256_, \oc8051_golden_model_1.ACC [2]);
  nor (_10226_, _10225_, _10224_);
  nor (_10227_, _10226_, _10223_);
  nor (_10228_, _03665_, \oc8051_golden_model_1.ACC [1]);
  and (_10229_, _03665_, \oc8051_golden_model_1.ACC [1]);
  and (_10230_, _02837_, \oc8051_golden_model_1.ACC [0]);
  nor (_10231_, _10230_, _10229_);
  nor (_10232_, _10231_, _10228_);
  not (_10233_, _10232_);
  and (_10234_, _10233_, _09520_);
  or (_10235_, _10234_, _10227_);
  nand (_10236_, _10235_, _09527_);
  and (_10237_, _10236_, _10222_);
  or (_10238_, _09528_, _09531_);
  nor (_10239_, _10238_, _10237_);
  or (_10240_, _10239_, _09489_);
  or (_10241_, _10240_, _10210_);
  and (_10242_, _10241_, _10190_);
  nor (_10243_, _10242_, _10189_);
  nor (_10244_, _10243_, _03063_);
  nor (_10245_, _10129_, _05502_);
  or (_10246_, _10131_, _02870_);
  nor (_10247_, _10246_, _10245_);
  and (_10248_, _03062_, \oc8051_golden_model_1.PSW [7]);
  and (_10249_, _10248_, _10103_);
  nor (_10250_, _10249_, _10247_);
  not (_10251_, _10250_);
  nor (_10252_, _10251_, _10244_);
  nor (_10253_, _10252_, _06247_);
  and (_10254_, _10253_, _09550_);
  nor (_10255_, _10254_, _10107_);
  nor (_10256_, _10255_, _03100_);
  or (_10257_, _10256_, _10106_);
  nor (_10258_, _10257_, _10105_);
  and (_10259_, _07334_, _07330_);
  nor (_10260_, _10259_, _07328_);
  not (_10261_, _10260_);
  and (_10262_, _07336_, _07330_);
  not (_10263_, _10262_);
  nor (_10264_, _10263_, _07742_);
  nor (_10265_, _10264_, _10261_);
  nor (_10266_, _10265_, _09989_);
  and (_10267_, _10266_, _10106_);
  nor (_10268_, _10267_, _10258_);
  nor (_10269_, _10268_, _03434_);
  and (_10270_, _07253_, _07248_);
  nor (_10271_, _10270_, _07246_);
  and (_10272_, _07255_, _07248_);
  not (_10273_, _10272_);
  nor (_10274_, _10273_, _07619_);
  not (_10275_, _10274_);
  and (_10276_, _10275_, _10271_);
  and (_10277_, _07257_, _06158_);
  and (_10278_, _10277_, _05849_);
  and (_10279_, _10278_, _05462_);
  nor (_10280_, _10279_, _07626_);
  not (_10281_, _10280_);
  nor (_10282_, _10281_, _10276_);
  nor (_10283_, _10282_, _10269_);
  and (_10284_, _10283_, _03111_);
  or (_10285_, _10284_, _10015_);
  and (_10286_, _10285_, _07405_);
  and (_10287_, _07755_, _04695_);
  and (_10288_, _07769_, _07763_);
  and (_10289_, _10288_, _07818_);
  and (_10290_, _10288_, _07820_);
  not (_10291_, _10290_);
  and (_10292_, _07767_, _07763_);
  nor (_10293_, _10292_, _07761_);
  and (_10294_, _10293_, _10291_);
  not (_10295_, _10294_);
  nor (_10296_, _10295_, _10289_);
  nor (_10297_, _10296_, _10287_);
  nor (_10298_, _10297_, _07405_);
  nor (_10299_, _10298_, _06770_);
  not (_10300_, _10299_);
  nor (_10301_, _10300_, _10286_);
  nor (_10302_, _10301_, _10004_);
  nor (_10303_, _10302_, _02853_);
  and (_10304_, _04690_, _05462_);
  nor (_10305_, _09994_, _05540_);
  not (_10306_, _10305_);
  nor (_10307_, _10306_, _10304_);
  nor (_10308_, _10307_, _02579_);
  not (_10309_, _10308_);
  nor (_10310_, _10309_, _10303_);
  nor (_10311_, _10310_, _10001_);
  nor (_10312_, _10311_, _06784_);
  and (_10313_, _10312_, _03490_);
  nor (_10314_, _10103_, _07293_);
  and (_10315_, _10314_, _02933_);
  or (_10316_, _10315_, _02802_);
  or (_10317_, _10316_, _10313_);
  and (_10318_, _05661_, _04690_);
  nor (_10319_, _10318_, _09994_);
  nand (_10320_, _10319_, _02802_);
  and (_10321_, _10320_, _10317_);
  nor (_10322_, _10321_, _02932_);
  and (_10323_, _10103_, _07293_);
  and (_10324_, _10323_, _02932_);
  nor (_10325_, _10324_, _10322_);
  and (_10326_, _10325_, _03887_);
  and (_10327_, _05766_, _04690_);
  nor (_10328_, _10327_, _09994_);
  nor (_10329_, _10328_, _03887_);
  or (_10330_, _10329_, _10326_);
  and (_10331_, _10330_, _03128_);
  nor (_10332_, _10331_, _09997_);
  nor (_10333_, _10332_, _02970_);
  nor (_10334_, _09994_, _04715_);
  not (_10335_, _10334_);
  nor (_10336_, _10319_, _03883_);
  and (_10337_, _10336_, _10335_);
  nor (_10338_, _10337_, _10333_);
  nor (_10339_, _10338_, _03135_);
  nor (_10340_, _10112_, _03137_);
  and (_10341_, _10340_, _10335_);
  or (_10342_, _10341_, _10339_);
  and (_10343_, _10342_, _05783_);
  nor (_10344_, _05765_, _09998_);
  nor (_10345_, _10344_, _09994_);
  nor (_10346_, _10345_, _05783_);
  or (_10347_, _10346_, _10343_);
  and (_10348_, _10347_, _05788_);
  not (_10349_, _07322_);
  nor (_10350_, _05773_, _09998_);
  nor (_10351_, _10350_, _09994_);
  nor (_10352_, _10351_, _05788_);
  nor (_10353_, _10352_, _10349_);
  not (_10354_, _10353_);
  nor (_10355_, _10354_, _10348_);
  nor (_10356_, _10355_, _09993_);
  nor (_10357_, _10356_, _07240_);
  nor (_10358_, _07245_, _05771_);
  or (_10359_, _10358_, _07310_);
  or (_10360_, _10279_, _07241_);
  or (_10361_, _10360_, _10359_);
  and (_10362_, _10361_, _03134_);
  not (_10363_, _10362_);
  nor (_10364_, _10363_, _10357_);
  not (_10365_, _09065_);
  nor (_10366_, _07523_, _05771_);
  or (_10367_, _07962_, _10006_);
  or (_10368_, _10367_, _10366_);
  or (_10369_, _10368_, _07985_);
  and (_10370_, _10369_, _10365_);
  nor (_10371_, _10370_, _10364_);
  nor (_10372_, _07760_, _05771_);
  nor (_10373_, _10372_, _08013_);
  nor (_10374_, _10287_, _07993_);
  and (_10375_, _10374_, _10373_);
  or (_10376_, _10375_, _07991_);
  nor (_10377_, _10376_, _10371_);
  not (_10378_, _07238_);
  and (_10379_, _07991_, \oc8051_golden_model_1.ACC [7]);
  nor (_10380_, _10379_, _10378_);
  not (_10381_, _10380_);
  nor (_10382_, _10381_, _10377_);
  nor (_10383_, _07192_, _07190_);
  nor (_10384_, _10383_, _07189_);
  and (_10385_, _07224_, _07191_);
  or (_10386_, _10385_, _07238_);
  nor (_10387_, _10386_, _10384_);
  nor (_10388_, _10387_, _10382_);
  nor (_10389_, _10388_, _07188_);
  nor (_10390_, _08025_, _07885_);
  nor (_10391_, _10390_, _07884_);
  and (_10392_, _08057_, _07886_);
  or (_10393_, _10392_, _08024_);
  nor (_10394_, _10393_, _10391_);
  or (_10395_, _10394_, _02894_);
  nor (_10396_, _10395_, _10389_);
  not (_10397_, _08069_);
  and (_10398_, _08104_, _10397_);
  nor (_10399_, _10398_, _08068_);
  and (_10400_, _10399_, _02894_);
  or (_10401_, _10400_, _10396_);
  and (_10402_, _10401_, _08113_);
  not (_10403_, _07894_);
  nor (_10404_, _08114_, _07895_);
  not (_10405_, _10404_);
  or (_10406_, _10405_, _08143_);
  and (_10407_, _10406_, _10403_);
  and (_10408_, _10407_, _08065_);
  or (_10409_, _10408_, _10402_);
  nor (_10410_, _10409_, _03163_);
  and (_10411_, _10109_, _03163_);
  nor (_10412_, _10411_, _08159_);
  not (_10413_, _10412_);
  nor (_10414_, _10413_, _10410_);
  and (_10415_, _08159_, \oc8051_golden_model_1.ACC [0]);
  or (_10416_, _10415_, _10414_);
  and (_10417_, _10416_, _02498_);
  nor (_10418_, _10142_, _02498_);
  or (_10419_, _10418_, _10417_);
  nor (_10420_, _10419_, _02888_);
  and (_10421_, _05235_, _04690_);
  nor (_10422_, _10421_, _09994_);
  and (_10423_, _10422_, _02888_);
  nor (_10424_, _10423_, _10420_);
  or (_10425_, _10424_, _42672_);
  or (_10426_, _42668_, \oc8051_golden_model_1.PSW [7]);
  and (_10427_, _10426_, _43998_);
  and (_40498_, _10427_, _10425_);
  not (_10428_, \oc8051_golden_model_1.PCON [7]);
  nor (_10429_, _04685_, _10428_);
  and (_10430_, _05774_, _04685_);
  nor (_10431_, _10430_, _10429_);
  nor (_10432_, _10431_, _03128_);
  and (_10433_, _04685_, _04604_);
  nor (_10434_, _10433_, _10429_);
  and (_10435_, _10434_, _06770_);
  and (_10436_, _04685_, \oc8051_golden_model_1.ACC [7]);
  nor (_10437_, _10436_, _10429_);
  nor (_10438_, _10437_, _03814_);
  nor (_10439_, _03813_, _10428_);
  or (_10440_, _10439_, _10438_);
  and (_10441_, _10440_, _03810_);
  and (_10442_, _05474_, _04685_);
  nor (_10443_, _10442_, _10429_);
  nor (_10444_, _10443_, _03810_);
  or (_10445_, _10444_, _10441_);
  and (_10446_, _10445_, _03336_);
  nor (_10447_, _10434_, _03336_);
  nor (_10448_, _10447_, _10446_);
  nor (_10449_, _10448_, _03075_);
  nor (_10450_, _10437_, _03084_);
  nor (_10451_, _10450_, _06770_);
  not (_10452_, _10451_);
  nor (_10453_, _10452_, _10449_);
  nor (_10454_, _10453_, _10435_);
  nor (_10455_, _10454_, _02853_);
  and (_10456_, _04685_, _05462_);
  nor (_10457_, _10429_, _05540_);
  not (_10458_, _10457_);
  nor (_10459_, _10458_, _10456_);
  or (_10460_, _10459_, _02579_);
  nor (_10461_, _10460_, _10455_);
  not (_10462_, _04685_);
  nor (_10463_, _05744_, _10462_);
  nor (_10464_, _10463_, _10429_);
  nor (_10465_, _10464_, _02838_);
  or (_10466_, _10465_, _02802_);
  or (_10467_, _10466_, _10461_);
  and (_10468_, _05661_, _04685_);
  nor (_10469_, _10468_, _10429_);
  nand (_10470_, _10469_, _02802_);
  and (_10471_, _10470_, _10467_);
  and (_10472_, _10471_, _03887_);
  and (_10473_, _05766_, _04685_);
  nor (_10474_, _10473_, _10429_);
  nor (_10475_, _10474_, _03887_);
  or (_10476_, _10475_, _10472_);
  and (_10477_, _10476_, _03128_);
  nor (_10478_, _10477_, _10432_);
  nor (_10479_, _10478_, _02970_);
  nor (_10480_, _10429_, _04715_);
  not (_10481_, _10480_);
  nor (_10482_, _10469_, _03883_);
  and (_10483_, _10482_, _10481_);
  nor (_10484_, _10483_, _10479_);
  nor (_10485_, _10484_, _03135_);
  nor (_10486_, _10437_, _03137_);
  and (_10487_, _10486_, _10481_);
  or (_10488_, _10487_, _10485_);
  and (_10489_, _10488_, _05783_);
  nor (_10490_, _05765_, _10462_);
  nor (_10491_, _10490_, _10429_);
  nor (_10492_, _10491_, _05783_);
  or (_10493_, _10492_, _10489_);
  and (_10494_, _10493_, _05788_);
  nor (_10495_, _05773_, _10462_);
  nor (_10496_, _10495_, _10429_);
  nor (_10497_, _10496_, _05788_);
  or (_10498_, _10497_, _03163_);
  nor (_10499_, _10498_, _10494_);
  and (_10500_, _10443_, _03163_);
  or (_10501_, _10500_, _02888_);
  nor (_10502_, _10501_, _10499_);
  and (_10503_, _05235_, _04685_);
  nor (_10504_, _10503_, _10429_);
  nor (_10505_, _10504_, _02890_);
  or (_10506_, _10505_, _10502_);
  or (_10507_, _10506_, _42672_);
  or (_10508_, _42668_, \oc8051_golden_model_1.PCON [7]);
  and (_10509_, _10508_, _43998_);
  and (_40499_, _10509_, _10507_);
  not (_10510_, \oc8051_golden_model_1.SBUF [7]);
  nor (_10511_, _04700_, _10510_);
  and (_10512_, _05774_, _04700_);
  nor (_10513_, _10512_, _10511_);
  nor (_10514_, _10513_, _03128_);
  and (_10515_, _04700_, \oc8051_golden_model_1.ACC [7]);
  nor (_10516_, _10515_, _10511_);
  nor (_10517_, _10516_, _03084_);
  nor (_10518_, _10516_, _03814_);
  nor (_10519_, _03813_, _10510_);
  or (_10520_, _10519_, _10518_);
  and (_10521_, _10520_, _03810_);
  and (_10522_, _05474_, _04700_);
  nor (_10523_, _10522_, _10511_);
  nor (_10524_, _10523_, _03810_);
  or (_10525_, _10524_, _10521_);
  and (_10526_, _10525_, _03336_);
  and (_10527_, _04700_, _04604_);
  nor (_10528_, _10527_, _10511_);
  nor (_10529_, _10528_, _03336_);
  nor (_10530_, _10529_, _10526_);
  nor (_10531_, _10530_, _03075_);
  or (_10532_, _10531_, _06770_);
  nor (_10533_, _10532_, _10517_);
  and (_10534_, _10528_, _06770_);
  nor (_10535_, _10534_, _10533_);
  nor (_10536_, _10535_, _02853_);
  and (_10537_, _04700_, _05462_);
  nor (_10538_, _10511_, _05540_);
  not (_10539_, _10538_);
  nor (_10540_, _10539_, _10537_);
  or (_10541_, _10540_, _02579_);
  nor (_10542_, _10541_, _10536_);
  not (_10543_, _04700_);
  nor (_10544_, _05744_, _10543_);
  nor (_10545_, _10544_, _10511_);
  nor (_10546_, _10545_, _02838_);
  or (_10547_, _10546_, _02802_);
  or (_10548_, _10547_, _10542_);
  and (_10549_, _05661_, _04700_);
  nor (_10550_, _10549_, _10511_);
  nand (_10551_, _10550_, _02802_);
  and (_10552_, _10551_, _10548_);
  and (_10553_, _10552_, _03887_);
  and (_10554_, _05766_, _04700_);
  nor (_10555_, _10554_, _10511_);
  nor (_10556_, _10555_, _03887_);
  or (_10557_, _10556_, _10553_);
  and (_10558_, _10557_, _03128_);
  nor (_10559_, _10558_, _10514_);
  nor (_10560_, _10559_, _02970_);
  nor (_10561_, _10511_, _04715_);
  not (_10562_, _10561_);
  nor (_10563_, _10550_, _03883_);
  and (_10564_, _10563_, _10562_);
  nor (_10565_, _10564_, _10560_);
  nor (_10566_, _10565_, _03135_);
  nor (_10567_, _10516_, _03137_);
  and (_10568_, _10567_, _10562_);
  nor (_10569_, _10568_, _02965_);
  not (_10570_, _10569_);
  nor (_10571_, _10570_, _10566_);
  nor (_10572_, _05765_, _10543_);
  or (_10573_, _10511_, _05783_);
  nor (_10574_, _10573_, _10572_);
  or (_10575_, _10574_, _03123_);
  nor (_10576_, _10575_, _10571_);
  nor (_10577_, _05773_, _10543_);
  nor (_10578_, _10577_, _10511_);
  nor (_10579_, _10578_, _05788_);
  or (_10580_, _10579_, _03163_);
  nor (_10581_, _10580_, _10576_);
  and (_10582_, _10523_, _03163_);
  or (_10583_, _10582_, _02888_);
  nor (_10584_, _10583_, _10581_);
  and (_10585_, _05235_, _04700_);
  nor (_10586_, _10585_, _10511_);
  nor (_10587_, _10586_, _02890_);
  or (_10588_, _10587_, _10584_);
  or (_10589_, _10588_, _42672_);
  or (_10590_, _42668_, \oc8051_golden_model_1.SBUF [7]);
  and (_10591_, _10590_, _43998_);
  and (_40500_, _10591_, _10589_);
  not (_10592_, \oc8051_golden_model_1.SCON [7]);
  nor (_10593_, _04666_, _10592_);
  and (_10594_, _05774_, _04666_);
  nor (_10595_, _10594_, _10593_);
  nor (_10596_, _10595_, _03128_);
  and (_10597_, _04666_, _04604_);
  nor (_10598_, _10597_, _10593_);
  and (_10599_, _10598_, _06770_);
  nor (_10600_, _05338_, _10592_);
  and (_10601_, _05356_, _05338_);
  nor (_10602_, _10601_, _10600_);
  nor (_10603_, _10602_, _02877_);
  and (_10604_, _04666_, \oc8051_golden_model_1.ACC [7]);
  nor (_10605_, _10604_, _10593_);
  nor (_10606_, _10605_, _03814_);
  nor (_10607_, _03813_, _10592_);
  or (_10608_, _10607_, _10606_);
  and (_10609_, _10608_, _03810_);
  and (_10610_, _05474_, _04666_);
  nor (_10611_, _10610_, _10593_);
  nor (_10612_, _10611_, _03810_);
  or (_10613_, _10612_, _10609_);
  and (_10614_, _10613_, _02881_);
  and (_10615_, _05360_, _05338_);
  nor (_10616_, _10615_, _10600_);
  nor (_10617_, _10616_, _02881_);
  or (_10618_, _10617_, _03069_);
  or (_10619_, _10618_, _10614_);
  nand (_10620_, _10598_, _03069_);
  and (_10621_, _10620_, _10619_);
  and (_10622_, _10621_, _03084_);
  nor (_10623_, _10605_, _03084_);
  or (_10624_, _10623_, _10622_);
  and (_10625_, _10624_, _02877_);
  nor (_10626_, _10625_, _10603_);
  nor (_10627_, _10626_, _02869_);
  and (_10628_, _05503_, _05338_);
  nor (_10629_, _10628_, _10600_);
  nor (_10630_, _10629_, _02870_);
  nor (_10631_, _10630_, _10627_);
  nor (_10632_, _10631_, _02863_);
  not (_10633_, _05338_);
  nor (_10634_, _05530_, _10633_);
  nor (_10635_, _10634_, _10600_);
  nor (_10636_, _10635_, _02864_);
  nor (_10637_, _10636_, _06770_);
  not (_10638_, _10637_);
  nor (_10639_, _10638_, _10632_);
  nor (_10640_, _10639_, _10599_);
  nor (_10641_, _10640_, _02853_);
  and (_10642_, _04666_, _05462_);
  nor (_10643_, _10593_, _05540_);
  not (_10644_, _10643_);
  nor (_10645_, _10644_, _10642_);
  nor (_10646_, _10645_, _02579_);
  not (_10647_, _10646_);
  nor (_10648_, _10647_, _10641_);
  not (_10649_, _04666_);
  nor (_10650_, _05744_, _10649_);
  nor (_10651_, _10650_, _10593_);
  nor (_10652_, _10651_, _02838_);
  or (_10653_, _10652_, _02802_);
  or (_10654_, _10653_, _10648_);
  and (_10655_, _05661_, _04666_);
  nor (_10656_, _10655_, _10593_);
  nand (_10657_, _10656_, _02802_);
  and (_10658_, _10657_, _10654_);
  and (_10659_, _10658_, _03887_);
  and (_10660_, _05766_, _04666_);
  nor (_10661_, _10660_, _10593_);
  nor (_10662_, _10661_, _03887_);
  or (_10663_, _10662_, _10659_);
  and (_10664_, _10663_, _03128_);
  nor (_10665_, _10664_, _10596_);
  nor (_10666_, _10665_, _02970_);
  nor (_10667_, _10593_, _04715_);
  not (_10668_, _10667_);
  nor (_10669_, _10656_, _03883_);
  and (_10670_, _10669_, _10668_);
  nor (_10671_, _10670_, _10666_);
  nor (_10672_, _10671_, _03135_);
  nor (_10673_, _10605_, _03137_);
  and (_10674_, _10673_, _10668_);
  nor (_10675_, _10674_, _02965_);
  not (_10676_, _10675_);
  nor (_10677_, _10676_, _10672_);
  nor (_10678_, _05765_, _10649_);
  or (_10679_, _10593_, _05783_);
  nor (_10680_, _10679_, _10678_);
  or (_10681_, _10680_, _03123_);
  nor (_10682_, _10681_, _10677_);
  nor (_10683_, _05773_, _10649_);
  nor (_10684_, _10683_, _10593_);
  nor (_10685_, _10684_, _05788_);
  or (_10686_, _10685_, _10682_);
  and (_10687_, _10686_, _03906_);
  nor (_10688_, _10611_, _03906_);
  or (_10689_, _10688_, _10687_);
  and (_10690_, _10689_, _02498_);
  nor (_10691_, _10602_, _02498_);
  or (_10692_, _10691_, _10690_);
  and (_10693_, _10692_, _02890_);
  and (_10694_, _05235_, _04666_);
  nor (_10695_, _10694_, _10593_);
  nor (_10696_, _10695_, _02890_);
  or (_10697_, _10696_, _10693_);
  or (_10698_, _10697_, _42672_);
  or (_10699_, _42668_, \oc8051_golden_model_1.SCON [7]);
  and (_10700_, _10699_, _43998_);
  and (_40501_, _10700_, _10698_);
  and (_10701_, _04247_, \oc8051_golden_model_1.SP [4]);
  and (_10702_, _10701_, \oc8051_golden_model_1.SP [5]);
  and (_10703_, _10702_, \oc8051_golden_model_1.SP [6]);
  nor (_10704_, _10703_, \oc8051_golden_model_1.SP [7]);
  and (_10705_, _10703_, \oc8051_golden_model_1.SP [7]);
  nor (_10706_, _10705_, _10704_);
  nor (_10707_, _10706_, _03915_);
  not (_10708_, \oc8051_golden_model_1.SP [7]);
  nor (_10709_, _04617_, _10708_);
  and (_10710_, _05774_, _04617_);
  nor (_10711_, _10710_, _10709_);
  nor (_10712_, _10711_, _03128_);
  and (_10713_, _05474_, _04617_);
  nor (_10714_, _10713_, _10709_);
  and (_10715_, _10714_, _02974_);
  and (_10716_, _04617_, \oc8051_golden_model_1.ACC [7]);
  nor (_10717_, _10716_, _10709_);
  or (_10718_, _10717_, _03814_);
  nand (_10719_, _09434_, \oc8051_golden_model_1.SP [7]);
  not (_10720_, _10706_);
  nor (_10721_, _10720_, _02611_);
  nor (_10722_, _10721_, _02974_);
  and (_10723_, _10722_, _10719_);
  and (_10724_, _10723_, _10718_);
  nor (_10725_, _10724_, _04252_);
  not (_10727_, _10725_);
  nor (_10728_, _10727_, _10715_);
  nor (_10729_, _10720_, _02609_);
  or (_10730_, _10729_, _03069_);
  nor (_10731_, _10730_, _10728_);
  not (_10732_, \oc8051_golden_model_1.SP [6]);
  not (_10733_, \oc8051_golden_model_1.SP [5]);
  not (_10734_, \oc8051_golden_model_1.SP [4]);
  and (_10735_, _05380_, _10734_);
  and (_10736_, _10735_, _10733_);
  and (_10738_, _10736_, _10732_);
  and (_10739_, _10738_, _02866_);
  nor (_10740_, _10739_, _10708_);
  and (_10741_, _10739_, _10708_);
  nor (_10742_, _10741_, _10740_);
  and (_10743_, _10742_, _03069_);
  nor (_10744_, _10743_, _10731_);
  and (_10745_, _10744_, _03084_);
  nor (_10746_, _10717_, _03084_);
  or (_10747_, _10746_, _10745_);
  and (_10749_, _10747_, _03941_);
  and (_10750_, _03320_, _02501_);
  and (_10751_, _10703_, \oc8051_golden_model_1.SP [0]);
  nor (_10752_, _10751_, _10708_);
  and (_10753_, _10751_, _10708_);
  nor (_10754_, _10753_, _10752_);
  nor (_10755_, _10754_, _03941_);
  or (_10756_, _10755_, _10750_);
  nor (_10757_, _10756_, _10749_);
  nand (_10758_, _10720_, _10750_);
  and (_10760_, _10758_, _05535_);
  not (_10761_, _10760_);
  nor (_10762_, _10761_, _10757_);
  and (_10763_, _04617_, _04604_);
  nor (_10764_, _10763_, _10709_);
  nor (_10765_, _10764_, _05535_);
  nor (_10766_, _10765_, _02853_);
  not (_10767_, _10766_);
  nor (_10768_, _10767_, _10762_);
  and (_10769_, _04617_, _05462_);
  nor (_10771_, _10709_, _05540_);
  not (_10772_, _10771_);
  nor (_10773_, _10772_, _10769_);
  nor (_10774_, _10773_, _02579_);
  not (_10775_, _10774_);
  nor (_10776_, _10775_, _10768_);
  not (_10777_, _04617_);
  nor (_10778_, _05744_, _10777_);
  nor (_10779_, _10778_, _10709_);
  nor (_10780_, _10779_, _02838_);
  or (_10782_, _10780_, _02802_);
  or (_10783_, _10782_, _10776_);
  and (_10784_, _05661_, _04617_);
  nor (_10785_, _10784_, _10709_);
  nand (_10786_, _10785_, _02802_);
  and (_10787_, _10786_, _10783_);
  nor (_10788_, _10787_, _02514_);
  and (_10789_, _10720_, _02514_);
  nor (_10790_, _10789_, _10788_);
  and (_10791_, _10790_, _03887_);
  and (_10793_, _05766_, _04617_);
  nor (_10794_, _10793_, _10709_);
  nor (_10795_, _10794_, _03887_);
  or (_10796_, _10795_, _10791_);
  and (_10797_, _10796_, _03128_);
  nor (_10798_, _10797_, _10712_);
  nor (_10799_, _10798_, _02970_);
  nor (_10800_, _10709_, _04715_);
  not (_10801_, _10800_);
  nor (_10802_, _10785_, _03883_);
  and (_10803_, _10802_, _10801_);
  nor (_10804_, _10803_, _10799_);
  nor (_10805_, _10804_, _09689_);
  nor (_10806_, _10720_, _02532_);
  or (_10807_, _10800_, _03137_);
  nor (_10808_, _10807_, _10717_);
  nor (_10809_, _10808_, _10806_);
  and (_10810_, _10809_, _05783_);
  not (_10811_, _10810_);
  nor (_10812_, _10811_, _10805_);
  nor (_10813_, _05765_, _10777_);
  or (_10814_, _10709_, _05783_);
  nor (_10815_, _10814_, _10813_);
  nor (_10816_, _10815_, _10812_);
  and (_10817_, _10816_, _05788_);
  nor (_10818_, _05773_, _10777_);
  nor (_10819_, _10818_, _10709_);
  nor (_10820_, _10819_, _05788_);
  or (_10821_, _10820_, _10817_);
  and (_10822_, _10821_, _09726_);
  nor (_10823_, _10738_, \oc8051_golden_model_1.SP [7]);
  and (_10824_, _10738_, \oc8051_golden_model_1.SP [7]);
  nor (_10825_, _10824_, _10823_);
  and (_10826_, _10825_, _03145_);
  or (_10827_, _10826_, _03898_);
  nor (_10828_, _10827_, _10822_);
  nor (_10829_, _10706_, _02529_);
  nor (_10830_, _10829_, _10828_);
  and (_10831_, _10830_, _02893_);
  and (_10832_, _10825_, _02892_);
  or (_10833_, _10832_, _10831_);
  and (_10834_, _10833_, _03906_);
  nor (_10835_, _10714_, _03906_);
  nor (_10836_, _10835_, _04337_);
  not (_10837_, _10836_);
  nor (_10838_, _10837_, _10834_);
  nor (_10839_, _10838_, _10707_);
  and (_10840_, _10839_, _02890_);
  and (_10841_, _05235_, _04617_);
  nor (_10842_, _10841_, _10709_);
  nor (_10843_, _10842_, _02890_);
  or (_10844_, _10843_, _10840_);
  or (_10845_, _10844_, _42672_);
  or (_10846_, _42668_, \oc8051_golden_model_1.SP [7]);
  and (_10847_, _10846_, _43998_);
  and (_40503_, _10847_, _10845_);
  not (_10848_, \oc8051_golden_model_1.TCON [7]);
  nor (_10849_, _04622_, _10848_);
  and (_10850_, _05774_, _04622_);
  nor (_10851_, _10850_, _10849_);
  nor (_10852_, _10851_, _03128_);
  and (_10853_, _04622_, _04604_);
  nor (_10854_, _10853_, _10849_);
  and (_10855_, _10854_, _06770_);
  nor (_10856_, _05320_, _10848_);
  and (_10857_, _05356_, _05320_);
  nor (_10858_, _10857_, _10856_);
  nor (_10859_, _10858_, _02877_);
  and (_10860_, _04622_, \oc8051_golden_model_1.ACC [7]);
  nor (_10861_, _10860_, _10849_);
  nor (_10862_, _10861_, _03814_);
  nor (_10863_, _03813_, _10848_);
  or (_10864_, _10863_, _10862_);
  and (_10865_, _10864_, _03810_);
  and (_10866_, _05474_, _04622_);
  nor (_10867_, _10866_, _10849_);
  nor (_10868_, _10867_, _03810_);
  or (_10869_, _10868_, _10865_);
  and (_10870_, _10869_, _02881_);
  and (_10871_, _05360_, _05320_);
  nor (_10872_, _10871_, _10856_);
  nor (_10873_, _10872_, _02881_);
  or (_10874_, _10873_, _03069_);
  or (_10875_, _10874_, _10870_);
  nand (_10876_, _10854_, _03069_);
  and (_10877_, _10876_, _10875_);
  and (_10878_, _10877_, _03084_);
  nor (_10879_, _10861_, _03084_);
  or (_10880_, _10879_, _10878_);
  and (_10881_, _10880_, _02877_);
  nor (_10882_, _10881_, _10859_);
  nor (_10883_, _10882_, _02869_);
  nor (_10884_, _10856_, _05502_);
  or (_10885_, _10872_, _02870_);
  nor (_10886_, _10885_, _10884_);
  nor (_10887_, _10886_, _10883_);
  nor (_10888_, _10887_, _02863_);
  not (_10889_, _05320_);
  nor (_10890_, _05530_, _10889_);
  nor (_10891_, _10890_, _10856_);
  nor (_10892_, _10891_, _02864_);
  nor (_10893_, _10892_, _06770_);
  not (_10894_, _10893_);
  nor (_10895_, _10894_, _10888_);
  nor (_10896_, _10895_, _10855_);
  nor (_10897_, _10896_, _02853_);
  and (_10898_, _04622_, _05462_);
  nor (_10899_, _10849_, _05540_);
  not (_10900_, _10899_);
  nor (_10901_, _10900_, _10898_);
  nor (_10902_, _10901_, _02579_);
  not (_10903_, _10902_);
  nor (_10904_, _10903_, _10897_);
  not (_10905_, _04622_);
  nor (_10906_, _05744_, _10905_);
  nor (_10907_, _10906_, _10849_);
  nor (_10908_, _10907_, _02838_);
  or (_10909_, _10908_, _02802_);
  or (_10910_, _10909_, _10904_);
  and (_10911_, _05661_, _04622_);
  nor (_10912_, _10911_, _10849_);
  nand (_10913_, _10912_, _02802_);
  and (_10914_, _10913_, _10910_);
  and (_10915_, _10914_, _03887_);
  and (_10916_, _05766_, _04622_);
  nor (_10917_, _10916_, _10849_);
  nor (_10918_, _10917_, _03887_);
  or (_10919_, _10918_, _10915_);
  and (_10920_, _10919_, _03128_);
  nor (_10921_, _10920_, _10852_);
  nor (_10922_, _10921_, _02970_);
  nor (_10923_, _10849_, _04715_);
  not (_10924_, _10923_);
  nor (_10925_, _10912_, _03883_);
  and (_10926_, _10925_, _10924_);
  nor (_10927_, _10926_, _10922_);
  nor (_10928_, _10927_, _03135_);
  nor (_10929_, _10861_, _03137_);
  and (_10930_, _10929_, _10924_);
  or (_10931_, _10930_, _10928_);
  and (_10932_, _10931_, _05783_);
  nor (_10933_, _05765_, _10905_);
  nor (_10934_, _10933_, _10849_);
  nor (_10935_, _10934_, _05783_);
  or (_10936_, _10935_, _10932_);
  and (_10937_, _10936_, _05788_);
  nor (_10938_, _05773_, _10905_);
  nor (_10939_, _10938_, _10849_);
  nor (_10940_, _10939_, _05788_);
  or (_10941_, _10940_, _10937_);
  and (_10942_, _10941_, _03906_);
  nor (_10943_, _10867_, _03906_);
  or (_10944_, _10943_, _10942_);
  and (_10945_, _10944_, _02498_);
  nor (_10946_, _10858_, _02498_);
  or (_10947_, _10946_, _10945_);
  and (_10948_, _10947_, _02890_);
  and (_10949_, _05235_, _04622_);
  nor (_10950_, _10949_, _10849_);
  nor (_10951_, _10950_, _02890_);
  or (_10952_, _10951_, _10948_);
  or (_10953_, _10952_, _42672_);
  or (_10954_, _42668_, \oc8051_golden_model_1.TCON [7]);
  and (_10955_, _10954_, _43998_);
  and (_40504_, _10955_, _10953_);
  not (_10956_, \oc8051_golden_model_1.TH0 [7]);
  nor (_10957_, _04679_, _10956_);
  and (_10958_, _05774_, _04679_);
  nor (_10959_, _10958_, _10957_);
  nor (_10960_, _10959_, _03128_);
  and (_10961_, _04679_, \oc8051_golden_model_1.ACC [7]);
  nor (_10962_, _10961_, _10957_);
  nor (_10963_, _10962_, _03084_);
  nor (_10964_, _10962_, _03814_);
  nor (_10965_, _03813_, _10956_);
  or (_10966_, _10965_, _10964_);
  and (_10967_, _10966_, _03810_);
  and (_10968_, _05474_, _04679_);
  nor (_10969_, _10968_, _10957_);
  nor (_10970_, _10969_, _03810_);
  or (_10971_, _10970_, _10967_);
  and (_10972_, _10971_, _03336_);
  and (_10973_, _04679_, _04604_);
  nor (_10974_, _10973_, _10957_);
  nor (_10975_, _10974_, _03336_);
  nor (_10976_, _10975_, _10972_);
  nor (_10977_, _10976_, _03075_);
  or (_10978_, _10977_, _06770_);
  nor (_10979_, _10978_, _10963_);
  and (_10980_, _10974_, _06770_);
  nor (_10981_, _10980_, _10979_);
  nor (_10982_, _10981_, _02853_);
  and (_10983_, _04679_, _05462_);
  nor (_10984_, _10957_, _05540_);
  not (_10985_, _10984_);
  nor (_10986_, _10985_, _10983_);
  or (_10987_, _10986_, _02579_);
  nor (_10988_, _10987_, _10982_);
  not (_10989_, _04679_);
  nor (_10990_, _05744_, _10989_);
  nor (_10991_, _10990_, _10957_);
  nor (_10992_, _10991_, _02838_);
  or (_10993_, _10992_, _02802_);
  or (_10994_, _10993_, _10988_);
  and (_10995_, _05661_, _04679_);
  nor (_10996_, _10995_, _10957_);
  nand (_10997_, _10996_, _02802_);
  and (_10998_, _10997_, _10994_);
  and (_10999_, _10998_, _03887_);
  and (_11000_, _05766_, _04679_);
  nor (_11001_, _11000_, _10957_);
  nor (_11002_, _11001_, _03887_);
  or (_11003_, _11002_, _10999_);
  and (_11004_, _11003_, _03128_);
  nor (_11005_, _11004_, _10960_);
  nor (_11006_, _11005_, _02970_);
  nor (_11007_, _10957_, _04715_);
  not (_11008_, _11007_);
  nor (_11009_, _10996_, _03883_);
  and (_11010_, _11009_, _11008_);
  nor (_11011_, _11010_, _11006_);
  nor (_11012_, _11011_, _03135_);
  nor (_11013_, _10962_, _03137_);
  and (_11014_, _11013_, _11008_);
  nor (_11015_, _11014_, _02965_);
  not (_11016_, _11015_);
  nor (_11017_, _11016_, _11012_);
  nor (_11018_, _05765_, _10989_);
  or (_11019_, _10957_, _05783_);
  nor (_11020_, _11019_, _11018_);
  or (_11021_, _11020_, _03123_);
  nor (_11022_, _11021_, _11017_);
  nor (_11023_, _05773_, _10989_);
  nor (_11024_, _11023_, _10957_);
  nor (_11025_, _11024_, _05788_);
  or (_11026_, _11025_, _03163_);
  nor (_11027_, _11026_, _11022_);
  and (_11028_, _10969_, _03163_);
  or (_11029_, _11028_, _02888_);
  nor (_11030_, _11029_, _11027_);
  and (_11031_, _05235_, _04679_);
  nor (_11032_, _11031_, _10957_);
  nor (_11033_, _11032_, _02890_);
  or (_11034_, _11033_, _11030_);
  or (_11035_, _11034_, _42672_);
  or (_11036_, _42668_, \oc8051_golden_model_1.TH0 [7]);
  and (_11037_, _11036_, _43998_);
  and (_40505_, _11037_, _11035_);
  not (_11038_, \oc8051_golden_model_1.TH1 [7]);
  nor (_11039_, _04660_, _11038_);
  and (_11040_, _05774_, _04660_);
  nor (_11041_, _11040_, _11039_);
  nor (_11042_, _11041_, _03128_);
  and (_11043_, _04660_, _04604_);
  nor (_11044_, _11043_, _11039_);
  and (_11045_, _11044_, _06770_);
  and (_11046_, _04660_, \oc8051_golden_model_1.ACC [7]);
  nor (_11047_, _11046_, _11039_);
  nor (_11048_, _11047_, _03084_);
  nor (_11049_, _11047_, _03814_);
  nor (_11050_, _03813_, _11038_);
  or (_11051_, _11050_, _11049_);
  and (_11052_, _11051_, _03810_);
  and (_11053_, _05474_, _04660_);
  nor (_11054_, _11053_, _11039_);
  nor (_11055_, _11054_, _03810_);
  or (_11056_, _11055_, _11052_);
  and (_11057_, _11056_, _03336_);
  nor (_11058_, _11044_, _03336_);
  nor (_11059_, _11058_, _11057_);
  nor (_11060_, _11059_, _03075_);
  or (_11061_, _11060_, _06770_);
  nor (_11062_, _11061_, _11048_);
  nor (_11063_, _11062_, _11045_);
  nor (_11064_, _11063_, _02853_);
  and (_11065_, _04660_, _05462_);
  nor (_11066_, _11039_, _05540_);
  not (_11067_, _11066_);
  nor (_11068_, _11067_, _11065_);
  or (_11069_, _11068_, _02579_);
  nor (_11070_, _11069_, _11064_);
  not (_11071_, _04660_);
  nor (_11072_, _05744_, _11071_);
  nor (_11073_, _11072_, _11039_);
  nor (_11074_, _11073_, _02838_);
  or (_11075_, _11074_, _02802_);
  or (_11076_, _11075_, _11070_);
  and (_11077_, _05661_, _04660_);
  nor (_11078_, _11077_, _11039_);
  nand (_11079_, _11078_, _02802_);
  and (_11080_, _11079_, _11076_);
  and (_11081_, _11080_, _03887_);
  and (_11082_, _05766_, _04660_);
  nor (_11083_, _11082_, _11039_);
  nor (_11084_, _11083_, _03887_);
  or (_11085_, _11084_, _11081_);
  and (_11086_, _11085_, _03128_);
  nor (_11087_, _11086_, _11042_);
  nor (_11088_, _11087_, _02970_);
  nor (_11089_, _11039_, _04715_);
  not (_11090_, _11089_);
  nor (_11091_, _11078_, _03883_);
  and (_11092_, _11091_, _11090_);
  nor (_11093_, _11092_, _11088_);
  nor (_11094_, _11093_, _03135_);
  nor (_11095_, _11047_, _03137_);
  and (_11096_, _11095_, _11090_);
  or (_11097_, _11096_, _11094_);
  and (_11098_, _11097_, _05783_);
  nor (_11099_, _05765_, _11071_);
  nor (_11100_, _11099_, _11039_);
  nor (_11101_, _11100_, _05783_);
  or (_11102_, _11101_, _11098_);
  and (_11103_, _11102_, _05788_);
  nor (_11104_, _05773_, _11071_);
  nor (_11105_, _11104_, _11039_);
  nor (_11106_, _11105_, _05788_);
  or (_11107_, _11106_, _03163_);
  nor (_11108_, _11107_, _11103_);
  and (_11109_, _11054_, _03163_);
  or (_11110_, _11109_, _02888_);
  nor (_11111_, _11110_, _11108_);
  and (_11112_, _05235_, _04660_);
  nor (_11113_, _11112_, _11039_);
  nor (_11114_, _11113_, _02890_);
  or (_11115_, _11114_, _11111_);
  or (_11116_, _11115_, _42672_);
  or (_11117_, _42668_, \oc8051_golden_model_1.TH1 [7]);
  and (_11118_, _11117_, _43998_);
  and (_40506_, _11118_, _11116_);
  not (_11119_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11120_, _04676_, _11119_);
  and (_11121_, _05774_, _04676_);
  nor (_11122_, _11121_, _11120_);
  nor (_11123_, _11122_, _03128_);
  and (_11124_, _04676_, \oc8051_golden_model_1.ACC [7]);
  nor (_11125_, _11124_, _11120_);
  nor (_11126_, _11125_, _03084_);
  nor (_11127_, _11125_, _03814_);
  nor (_11128_, _03813_, _11119_);
  or (_11129_, _11128_, _11127_);
  and (_11130_, _11129_, _03810_);
  and (_11131_, _05474_, _04676_);
  nor (_11132_, _11131_, _11120_);
  nor (_11133_, _11132_, _03810_);
  or (_11134_, _11133_, _11130_);
  and (_11135_, _11134_, _03336_);
  and (_11136_, _04676_, _04604_);
  nor (_11137_, _11136_, _11120_);
  nor (_11138_, _11137_, _03336_);
  nor (_11139_, _11138_, _11135_);
  nor (_11140_, _11139_, _03075_);
  or (_11141_, _11140_, _06770_);
  nor (_11142_, _11141_, _11126_);
  and (_11143_, _11137_, _06770_);
  nor (_11144_, _11143_, _11142_);
  nor (_11145_, _11144_, _02853_);
  and (_11146_, _04676_, _05462_);
  nor (_11147_, _11120_, _05540_);
  not (_11148_, _11147_);
  nor (_11149_, _11148_, _11146_);
  or (_11150_, _11149_, _02579_);
  nor (_11151_, _11150_, _11145_);
  not (_11152_, _04676_);
  nor (_11153_, _05744_, _11152_);
  nor (_11154_, _11153_, _11120_);
  nor (_11155_, _11154_, _02838_);
  or (_11156_, _11155_, _02802_);
  or (_11157_, _11156_, _11151_);
  and (_11158_, _05661_, _04676_);
  nor (_11159_, _11158_, _11120_);
  nand (_11160_, _11159_, _02802_);
  and (_11161_, _11160_, _11157_);
  and (_11162_, _11161_, _03887_);
  and (_11163_, _05766_, _04676_);
  nor (_11164_, _11163_, _11120_);
  nor (_11165_, _11164_, _03887_);
  or (_11166_, _11165_, _11162_);
  and (_11167_, _11166_, _03128_);
  nor (_11168_, _11167_, _11123_);
  nor (_11169_, _11168_, _02970_);
  nor (_11170_, _11120_, _04715_);
  not (_11171_, _11170_);
  nor (_11172_, _11159_, _03883_);
  and (_11173_, _11172_, _11171_);
  nor (_11174_, _11173_, _11169_);
  nor (_11175_, _11174_, _03135_);
  nor (_11176_, _11125_, _03137_);
  and (_11177_, _11176_, _11171_);
  or (_11178_, _11177_, _11175_);
  and (_11179_, _11178_, _05783_);
  nor (_11180_, _05765_, _11152_);
  nor (_11181_, _11180_, _11120_);
  nor (_11182_, _11181_, _05783_);
  or (_11183_, _11182_, _11179_);
  and (_11184_, _11183_, _05788_);
  nor (_11185_, _05773_, _11152_);
  nor (_11186_, _11185_, _11120_);
  nor (_11187_, _11186_, _05788_);
  or (_11188_, _11187_, _03163_);
  nor (_11189_, _11188_, _11184_);
  and (_11190_, _11132_, _03163_);
  or (_11191_, _11190_, _02888_);
  nor (_11192_, _11191_, _11189_);
  and (_11193_, _05235_, _04676_);
  nor (_11194_, _11193_, _11120_);
  nor (_11195_, _11194_, _02890_);
  or (_11196_, _11195_, _11192_);
  or (_11197_, _11196_, _42672_);
  or (_11198_, _42668_, \oc8051_golden_model_1.TL0 [7]);
  and (_11199_, _11198_, _43998_);
  and (_40507_, _11199_, _11197_);
  not (_11200_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11201_, _04656_, _11200_);
  and (_11202_, _05774_, _04656_);
  nor (_11203_, _11202_, _11201_);
  nor (_11204_, _11203_, _03128_);
  and (_11205_, _04656_, \oc8051_golden_model_1.ACC [7]);
  nor (_11206_, _11205_, _11201_);
  nor (_11207_, _11206_, _03084_);
  nor (_11208_, _11206_, _03814_);
  nor (_11209_, _03813_, _11200_);
  or (_11210_, _11209_, _11208_);
  and (_11211_, _11210_, _03810_);
  and (_11212_, _05474_, _04656_);
  nor (_11213_, _11212_, _11201_);
  nor (_11214_, _11213_, _03810_);
  or (_11215_, _11214_, _11211_);
  and (_11216_, _11215_, _03336_);
  and (_11217_, _04656_, _04604_);
  nor (_11218_, _11217_, _11201_);
  nor (_11219_, _11218_, _03336_);
  nor (_11220_, _11219_, _11216_);
  nor (_11221_, _11220_, _03075_);
  or (_11222_, _11221_, _06770_);
  nor (_11223_, _11222_, _11207_);
  and (_11224_, _11218_, _06770_);
  nor (_11225_, _11224_, _11223_);
  nor (_11226_, _11225_, _02853_);
  and (_11227_, _04656_, _05462_);
  nor (_11228_, _11201_, _05540_);
  not (_11229_, _11228_);
  nor (_11230_, _11229_, _11227_);
  or (_11231_, _11230_, _02579_);
  nor (_11232_, _11231_, _11226_);
  not (_11233_, _04656_);
  nor (_11234_, _05744_, _11233_);
  nor (_11235_, _11234_, _11201_);
  nor (_11236_, _11235_, _02838_);
  or (_11237_, _11236_, _02802_);
  or (_11238_, _11237_, _11232_);
  and (_11239_, _05661_, _04656_);
  nor (_11240_, _11239_, _11201_);
  nand (_11241_, _11240_, _02802_);
  and (_11242_, _11241_, _11238_);
  and (_11243_, _11242_, _03887_);
  and (_11244_, _05766_, _04656_);
  nor (_11245_, _11244_, _11201_);
  nor (_11246_, _11245_, _03887_);
  or (_11247_, _11246_, _11243_);
  and (_11248_, _11247_, _03128_);
  nor (_11249_, _11248_, _11204_);
  nor (_11250_, _11249_, _02970_);
  nor (_11251_, _11201_, _04715_);
  not (_11252_, _11251_);
  nor (_11253_, _11240_, _03883_);
  and (_11254_, _11253_, _11252_);
  nor (_11255_, _11254_, _11250_);
  nor (_11256_, _11255_, _03135_);
  nor (_11257_, _11206_, _03137_);
  and (_11258_, _11257_, _11252_);
  or (_11259_, _11258_, _11256_);
  and (_11260_, _11259_, _05783_);
  nor (_11261_, _05765_, _11233_);
  nor (_11262_, _11261_, _11201_);
  nor (_11263_, _11262_, _05783_);
  or (_11264_, _11263_, _11260_);
  and (_11265_, _11264_, _05788_);
  nor (_11266_, _05773_, _11233_);
  nor (_11267_, _11266_, _11201_);
  nor (_11268_, _11267_, _05788_);
  or (_11269_, _11268_, _03163_);
  nor (_11270_, _11269_, _11265_);
  and (_11271_, _11213_, _03163_);
  or (_11272_, _11271_, _02888_);
  nor (_11273_, _11272_, _11270_);
  and (_11274_, _05235_, _04656_);
  nor (_11275_, _11274_, _11201_);
  nor (_11276_, _11275_, _02890_);
  or (_11277_, _11276_, _11273_);
  or (_11278_, _11277_, _42672_);
  or (_11279_, _42668_, \oc8051_golden_model_1.TL1 [7]);
  and (_11280_, _11279_, _43998_);
  and (_40508_, _11280_, _11278_);
  not (_11281_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11282_, _04664_, _11281_);
  and (_11283_, _05774_, _04664_);
  nor (_11284_, _11283_, _11282_);
  nor (_11285_, _11284_, _03128_);
  and (_11286_, _04664_, _04604_);
  nor (_11287_, _11286_, _11282_);
  and (_11288_, _11287_, _06770_);
  and (_11289_, _04664_, \oc8051_golden_model_1.ACC [7]);
  nor (_11290_, _11289_, _11282_);
  nor (_11291_, _11290_, _03814_);
  nor (_11292_, _03813_, _11281_);
  or (_11293_, _11292_, _11291_);
  and (_11294_, _11293_, _03810_);
  and (_11295_, _05474_, _04664_);
  nor (_11296_, _11295_, _11282_);
  nor (_11297_, _11296_, _03810_);
  or (_11298_, _11297_, _11294_);
  and (_11299_, _11298_, _03336_);
  nor (_11300_, _11287_, _03336_);
  nor (_11301_, _11300_, _11299_);
  nor (_11302_, _11301_, _03075_);
  nor (_11303_, _11290_, _03084_);
  nor (_11304_, _11303_, _06770_);
  not (_11305_, _11304_);
  nor (_11306_, _11305_, _11302_);
  nor (_11307_, _11306_, _11288_);
  nor (_11308_, _11307_, _02853_);
  and (_11309_, _04664_, _05462_);
  nor (_11310_, _11282_, _05540_);
  not (_11311_, _11310_);
  nor (_11312_, _11311_, _11309_);
  or (_11313_, _11312_, _02579_);
  nor (_11314_, _11313_, _11308_);
  not (_11315_, _04664_);
  nor (_11316_, _05744_, _11315_);
  nor (_11317_, _11316_, _11282_);
  nor (_11318_, _11317_, _02838_);
  or (_11319_, _11318_, _02802_);
  or (_11320_, _11319_, _11314_);
  and (_11321_, _05661_, _04664_);
  nor (_11322_, _11321_, _11282_);
  nand (_11323_, _11322_, _02802_);
  and (_11324_, _11323_, _11320_);
  and (_11325_, _11324_, _03887_);
  and (_11326_, _05766_, _04664_);
  nor (_11327_, _11326_, _11282_);
  nor (_11328_, _11327_, _03887_);
  or (_11329_, _11328_, _11325_);
  and (_11330_, _11329_, _03128_);
  nor (_11331_, _11330_, _11285_);
  nor (_11332_, _11331_, _02970_);
  nor (_11333_, _11282_, _04715_);
  not (_11334_, _11333_);
  nor (_11335_, _11322_, _03883_);
  and (_11336_, _11335_, _11334_);
  nor (_11337_, _11336_, _11332_);
  nor (_11338_, _11337_, _03135_);
  nor (_11339_, _11290_, _03137_);
  and (_11340_, _11339_, _11334_);
  nor (_11341_, _11340_, _02965_);
  not (_11342_, _11341_);
  nor (_11343_, _11342_, _11338_);
  nor (_11344_, _05765_, _11315_);
  or (_11345_, _11282_, _05783_);
  nor (_11346_, _11345_, _11344_);
  or (_11347_, _11346_, _03123_);
  nor (_11348_, _11347_, _11343_);
  nor (_11349_, _05773_, _11315_);
  nor (_11350_, _11349_, _11282_);
  nor (_11351_, _11350_, _05788_);
  or (_11352_, _11351_, _03163_);
  nor (_11353_, _11352_, _11348_);
  and (_11354_, _11296_, _03163_);
  or (_11355_, _11354_, _02888_);
  nor (_11356_, _11355_, _11353_);
  and (_11357_, _05235_, _04664_);
  nor (_11358_, _11357_, _11282_);
  nor (_11359_, _11358_, _02890_);
  or (_11360_, _11359_, _11356_);
  or (_11361_, _11360_, _42672_);
  or (_11362_, _42668_, \oc8051_golden_model_1.TMOD [7]);
  and (_11363_, _11362_, _43998_);
  and (_40509_, _11363_, _11361_);
  and (_11364_, _42672_, \oc8051_golden_model_1.P0INREG [7]);
  or (_11365_, _11364_, _00685_);
  and (_40510_, _11365_, _43998_);
  and (_11366_, _42672_, \oc8051_golden_model_1.P1INREG [7]);
  or (_11367_, _11366_, _00573_);
  and (_40511_, _11367_, _43998_);
  and (_11368_, _42672_, \oc8051_golden_model_1.P2INREG [7]);
  or (_11369_, _11368_, _00755_);
  and (_40512_, _11369_, _43998_);
  and (_11370_, _42672_, \oc8051_golden_model_1.P3INREG [7]);
  or (_11371_, _11370_, _00480_);
  and (_40514_, _11371_, _43998_);
  not (_11372_, _00000_);
  nor (_11373_, _04181_, _11372_);
  not (_11374_, _11373_);
  nor (_11375_, _11374_, _03929_);
  nor (_11376_, _11374_, _04092_);
  nor (_11377_, _11376_, _11375_);
  nor (_11378_, _04351_, _11374_);
  nor (_11379_, _04531_, _11374_);
  nor (_11380_, _11379_, _11378_);
  and (_11381_, _11380_, _11373_);
  and (_11382_, _11381_, _11377_);
  or (_11383_, _11382_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_11384_, _04543_, _11372_);
  not (_11385_, _11384_);
  not (_11386_, _03933_);
  and (_11387_, _11384_, _04539_);
  and (_11388_, _11384_, _04542_);
  or (_11389_, _11388_, _11387_);
  or (_11390_, _11389_, _11386_);
  or (_11391_, _11390_, _11385_);
  and (_11392_, _11391_, _11383_);
  not (_11393_, _11382_);
  and (_11394_, _05226_, _03923_);
  not (_11395_, _05789_);
  and (_11396_, _05226_, _03486_);
  nor (_11397_, _11396_, _05790_);
  nor (_11398_, _05226_, _03486_);
  nor (_11399_, _11398_, _11396_);
  and (_11400_, _11399_, _03888_);
  not (_11401_, _05536_);
  or (_11402_, _03808_, _11401_);
  nand (_11403_, _07481_, _03059_);
  nand (_11404_, _07481_, _02875_);
  nor (_11405_, _10063_, _04620_);
  or (_11406_, _11405_, _05315_);
  and (_11407_, _05226_, _03811_);
  nand (_11408_, _05363_, _03808_);
  nor (_11409_, _02611_, _02244_);
  and (_11410_, _02611_, \oc8051_golden_model_1.ACC [0]);
  nor (_11411_, _11410_, _11409_);
  and (_11412_, _11411_, _05362_);
  nor (_11413_, _11412_, _03811_);
  and (_11414_, _11413_, _11408_);
  or (_11415_, _11414_, _11407_);
  and (_11416_, _11415_, _05358_);
  nand (_11417_, _10063_, _09812_);
  and (_11418_, _11417_, _02883_);
  or (_11419_, _11418_, _04252_);
  or (_11420_, _11419_, _11416_);
  nor (_11421_, _02609_, \oc8051_golden_model_1.PC [0]);
  nor (_11422_, _11421_, _03836_);
  and (_11423_, _11422_, _11420_);
  and (_11424_, _03808_, _03836_);
  or (_11425_, _11424_, _03844_);
  or (_11426_, _11425_, _11423_);
  and (_11427_, _11426_, _11406_);
  or (_11428_, _11427_, _02875_);
  and (_11429_, _11428_, _11404_);
  or (_11430_, _11429_, _02872_);
  not (_11431_, _10064_);
  and (_11432_, _11417_, _11431_);
  or (_11433_, _11432_, _02873_);
  and (_11434_, _11433_, _02614_);
  and (_11435_, _11434_, _11430_);
  nor (_11436_, _02614_, _02244_);
  or (_11437_, _03059_, _11436_);
  or (_11438_, _11437_, _11435_);
  and (_11439_, _11438_, _11403_);
  or (_11440_, _11439_, _03859_);
  and (_11441_, _06152_, _04551_);
  nand (_11442_, _07480_, _03859_);
  or (_11443_, _11442_, _11441_);
  and (_11444_, _11443_, _11440_);
  or (_11445_, _11444_, _03858_);
  nor (_11446_, _09835_, _04620_);
  and (_11447_, _04620_, \oc8051_golden_model_1.PSW [7]);
  nor (_11448_, _11447_, _11446_);
  nand (_11449_, _11448_, _03858_);
  and (_11450_, _11449_, _04251_);
  and (_11451_, _11450_, _11445_);
  and (_11452_, _02581_, \oc8051_golden_model_1.PC [0]);
  or (_11453_, _05536_, _11452_);
  or (_11454_, _11453_, _11451_);
  and (_11455_, _11454_, _11402_);
  or (_11456_, _11455_, _05541_);
  or (_11457_, _06152_, _05546_);
  and (_11458_, _11457_, _05545_);
  and (_11459_, _11458_, _11456_);
  and (_11460_, _05311_, _03808_);
  and (_11461_, _05655_, \oc8051_golden_model_1.B [0]);
  and (_11462_, _05652_, \oc8051_golden_model_1.ACC [0]);
  nor (_11463_, _11462_, _11461_);
  and (_11464_, _05664_, \oc8051_golden_model_1.IP [0]);
  and (_11465_, _05668_, \oc8051_golden_model_1.PSW [0]);
  nor (_11466_, _11465_, _11464_);
  and (_11467_, _11466_, _11463_);
  and (_11468_, _05717_, \oc8051_golden_model_1.P1INREG [0]);
  not (_11469_, _11468_);
  and (_11470_, _05710_, \oc8051_golden_model_1.P0INREG [0]);
  not (_11471_, _11470_);
  and (_11472_, _05720_, \oc8051_golden_model_1.P2INREG [0]);
  and (_11473_, _08669_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_11474_, _11473_, _11472_);
  and (_11475_, _11474_, _11471_);
  and (_11476_, _11475_, _11469_);
  and (_11477_, _11476_, _11467_);
  and (_11478_, _05726_, \oc8051_golden_model_1.IE [0]);
  and (_11479_, _05729_, \oc8051_golden_model_1.SBUF [0]);
  and (_11480_, _05731_, \oc8051_golden_model_1.SCON [0]);
  or (_11481_, _11480_, _11479_);
  nor (_11482_, _11481_, _11478_);
  and (_11483_, _05678_, \oc8051_golden_model_1.TH1 [0]);
  and (_11484_, _05737_, \oc8051_golden_model_1.DPH [0]);
  nor (_11485_, _11484_, _11483_);
  and (_11486_, _11485_, _11482_);
  and (_11487_, _11486_, _11477_);
  and (_11488_, _05692_, \oc8051_golden_model_1.TH0 [0]);
  and (_11489_, _05696_, \oc8051_golden_model_1.TL1 [0]);
  nor (_11490_, _11489_, _11488_);
  and (_11491_, _05699_, \oc8051_golden_model_1.TCON [0]);
  and (_11492_, _05703_, \oc8051_golden_model_1.PCON [0]);
  nor (_11493_, _11492_, _11491_);
  and (_11494_, _11493_, _11490_);
  and (_11495_, _05707_, \oc8051_golden_model_1.DPL [0]);
  and (_11496_, _05687_, \oc8051_golden_model_1.TL0 [0]);
  nor (_11497_, _11496_, _11495_);
  and (_11498_, _05682_, \oc8051_golden_model_1.SP [0]);
  and (_11499_, _05735_, \oc8051_golden_model_1.TMOD [0]);
  nor (_11500_, _11499_, _11498_);
  and (_11501_, _11500_, _11497_);
  and (_11502_, _11501_, _11494_);
  and (_11503_, _11502_, _11487_);
  not (_11504_, _11503_);
  nor (_11505_, _11504_, _11460_);
  nor (_11506_, _11505_, _05545_);
  or (_11507_, _11506_, _05754_);
  or (_11508_, _11507_, _11459_);
  and (_11509_, _05754_, _02837_);
  nor (_11510_, _11509_, _02804_);
  and (_11511_, _11510_, _11508_);
  and (_11512_, _05672_, _02804_);
  or (_11513_, _11512_, _02514_);
  or (_11514_, _11513_, _11511_);
  and (_11515_, _02514_, _02244_);
  nor (_11516_, _11515_, _03888_);
  and (_11517_, _11516_, _11514_);
  or (_11518_, _11517_, _11400_);
  and (_11519_, _11518_, _05770_);
  and (_11520_, _05226_, _02667_);
  nor (_11521_, _05226_, _02667_);
  nor (_11522_, _11521_, _11520_);
  and (_11523_, _11522_, _03886_);
  or (_11524_, _11523_, _11519_);
  and (_11525_, _11524_, _03885_);
  and (_11526_, _11398_, _03884_);
  or (_11527_, _11526_, _11525_);
  and (_11528_, _11527_, _03882_);
  and (_11529_, _11521_, _03881_);
  or (_11530_, _11529_, _03880_);
  or (_11531_, _11530_, _11528_);
  nor (_11532_, _02532_, \oc8051_golden_model_1.PC [0]);
  nor (_11533_, _11532_, _05784_);
  and (_11534_, _11533_, _11531_);
  or (_11535_, _11534_, _11397_);
  and (_11536_, _11535_, _11395_);
  nor (_11537_, _11520_, _11395_);
  or (_11538_, _11537_, _03898_);
  or (_11539_, _11538_, _11536_);
  or (_11540_, _02529_, \oc8051_golden_model_1.PC [0]);
  and (_11541_, _11540_, _09940_);
  and (_11542_, _11541_, _11539_);
  nor (_11543_, _09940_, _03808_);
  or (_11544_, _11543_, _11542_);
  and (_11545_, _11544_, _03909_);
  and (_11546_, _05940_, _03575_);
  or (_11547_, _11546_, _03908_);
  or (_11548_, _11547_, _11545_);
  or (_11549_, _05226_, _04333_);
  and (_11550_, _11549_, _03915_);
  and (_11551_, _11550_, _11548_);
  and (_11552_, _02525_, \oc8051_golden_model_1.PC [0]);
  and (_11553_, _02939_, _02244_);
  or (_11554_, _11553_, _11552_);
  or (_11555_, _11554_, _02797_);
  or (_11556_, _11555_, _11551_);
  or (_11557_, _11446_, _02798_);
  and (_11558_, _11557_, _05237_);
  and (_11559_, _11558_, _11556_);
  nor (_11560_, _05237_, _03808_);
  or (_11561_, _11560_, _03920_);
  or (_11562_, _11561_, _11559_);
  or (_11563_, _05940_, _03921_);
  and (_11564_, _11563_, _06150_);
  and (_11565_, _11564_, _11562_);
  or (_11566_, _11565_, _11394_);
  or (_11567_, _11566_, _11393_);
  and (_11568_, _11567_, _11392_);
  and (_11569_, _04544_, _04539_);
  nor (_11570_, _11569_, _04545_);
  and (_11571_, _04544_, _03933_);
  and (_11572_, _11571_, _11570_);
  nand (_11573_, _09298_, _02939_);
  or (_11574_, _09168_, _02939_);
  and (_11575_, _11574_, _11573_);
  and (_11576_, _11575_, _04544_);
  and (_11577_, _11576_, _11572_);
  or (_40542_, _11577_, _11568_);
  nor (_11578_, _04185_, _03929_);
  nor (_11579_, _11578_, _04186_);
  nor (_11580_, _04185_, _04351_);
  or (_11581_, _11580_, _04532_);
  nor (_11582_, _11581_, _04185_);
  nand (_11583_, _11582_, _11579_);
  nor (_11584_, _05271_, _05239_);
  nand (_11585_, _11584_, _04514_);
  and (_11586_, _04149_, _02367_);
  nor (_11587_, _05178_, _02551_);
  or (_11588_, _11587_, _03882_);
  or (_11589_, _11401_, _04000_);
  nand (_11590_, _07467_, _03059_);
  not (_11591_, _10039_);
  nand (_11592_, _10038_, _09757_);
  and (_11593_, _11592_, _02872_);
  and (_11594_, _11593_, _11591_);
  nor (_11595_, _10038_, _04616_);
  or (_11596_, _11595_, _05315_);
  nand (_11597_, _11584_, _05363_);
  nor (_11598_, _02611_, \oc8051_golden_model_1.PC [1]);
  and (_11599_, _02611_, \oc8051_golden_model_1.ACC [1]);
  or (_11600_, _11599_, _11598_);
  nor (_11601_, _11600_, _04143_);
  nand (_11602_, _11601_, _04011_);
  or (_11603_, _11602_, _03729_);
  and (_11604_, _11603_, _11597_);
  and (_11605_, _11604_, _03812_);
  nor (_11606_, _05227_, _05467_);
  nor (_11607_, _11606_, _03812_);
  or (_11608_, _11607_, _11605_);
  or (_11609_, _11608_, _02883_);
  or (_11610_, _11592_, _05358_);
  and (_11611_, _11610_, _11609_);
  or (_11612_, _11611_, _04252_);
  nor (_11613_, _02609_, _02215_);
  nor (_11614_, _11613_, _03836_);
  and (_11615_, _11614_, _11612_);
  and (_11616_, _03836_, _04000_);
  or (_11617_, _11616_, _03844_);
  or (_11618_, _11617_, _11615_);
  and (_11619_, _11618_, _11596_);
  or (_11620_, _11619_, _02875_);
  nand (_11621_, _07467_, _02875_);
  and (_11622_, _11621_, _02873_);
  and (_11623_, _11622_, _11620_);
  or (_11624_, _11623_, _11594_);
  and (_11625_, _11624_, _02614_);
  nor (_11626_, _02614_, \oc8051_golden_model_1.PC [1]);
  or (_11627_, _03059_, _11626_);
  or (_11628_, _11627_, _11625_);
  and (_11629_, _11628_, _11590_);
  or (_11630_, _11629_, _03859_);
  and (_11631_, _06151_, _04551_);
  nand (_11632_, _07466_, _03859_);
  or (_11633_, _11632_, _11631_);
  and (_11634_, _11633_, _11630_);
  or (_11635_, _11634_, _03858_);
  nor (_11636_, _09780_, _04616_);
  and (_11637_, _04616_, \oc8051_golden_model_1.PSW [7]);
  nor (_11638_, _11637_, _11636_);
  nand (_11639_, _11638_, _03858_);
  and (_11640_, _11639_, _04251_);
  and (_11641_, _11640_, _11635_);
  and (_11642_, _02581_, _02215_);
  or (_11643_, _05536_, _11642_);
  or (_11644_, _11643_, _11641_);
  and (_11645_, _11644_, _11589_);
  or (_11646_, _11645_, _05541_);
  or (_11647_, _06151_, _05546_);
  and (_11648_, _11647_, _05545_);
  and (_11649_, _11648_, _11646_);
  and (_11650_, _05311_, _04000_);
  and (_11651_, _05717_, \oc8051_golden_model_1.P1INREG [1]);
  not (_11652_, _11651_);
  and (_11653_, _05710_, \oc8051_golden_model_1.P0INREG [1]);
  not (_11654_, _11653_);
  and (_11655_, _05720_, \oc8051_golden_model_1.P2INREG [1]);
  and (_11656_, _08669_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_11657_, _11656_, _11655_);
  and (_11658_, _11657_, _11654_);
  and (_11659_, _11658_, _11652_);
  and (_11660_, _05682_, \oc8051_golden_model_1.SP [1]);
  and (_11661_, _05687_, \oc8051_golden_model_1.TL0 [1]);
  nor (_11662_, _11661_, _11660_);
  and (_11663_, _11662_, _11659_);
  and (_11664_, _05664_, \oc8051_golden_model_1.IP [1]);
  and (_11665_, _05655_, \oc8051_golden_model_1.B [1]);
  nor (_11666_, _11665_, _11664_);
  and (_11667_, _05668_, \oc8051_golden_model_1.PSW [1]);
  and (_11668_, _05652_, \oc8051_golden_model_1.ACC [1]);
  nor (_11669_, _11668_, _11667_);
  and (_11670_, _11669_, _11666_);
  and (_11671_, _05726_, \oc8051_golden_model_1.IE [1]);
  and (_11672_, _05729_, \oc8051_golden_model_1.SBUF [1]);
  and (_11673_, _05731_, \oc8051_golden_model_1.SCON [1]);
  or (_11674_, _11673_, _11672_);
  nor (_11675_, _11674_, _11671_);
  and (_11676_, _11675_, _11670_);
  and (_11677_, _11676_, _11663_);
  and (_11678_, _05692_, \oc8051_golden_model_1.TH0 [1]);
  and (_11679_, _05696_, \oc8051_golden_model_1.TL1 [1]);
  nor (_11680_, _11679_, _11678_);
  and (_11681_, _05699_, \oc8051_golden_model_1.TCON [1]);
  and (_11682_, _05703_, \oc8051_golden_model_1.PCON [1]);
  nor (_11683_, _11682_, _11681_);
  and (_11684_, _11683_, _11680_);
  and (_11685_, _05737_, \oc8051_golden_model_1.DPH [1]);
  and (_11686_, _05735_, \oc8051_golden_model_1.TMOD [1]);
  nor (_11687_, _11686_, _11685_);
  and (_11688_, _05707_, \oc8051_golden_model_1.DPL [1]);
  and (_11689_, _05678_, \oc8051_golden_model_1.TH1 [1]);
  nor (_11690_, _11689_, _11688_);
  and (_11691_, _11690_, _11687_);
  and (_11692_, _11691_, _11684_);
  and (_11693_, _11692_, _11677_);
  not (_11694_, _11693_);
  nor (_11695_, _11694_, _11650_);
  nor (_11696_, _11695_, _05545_);
  or (_11697_, _11696_, _05754_);
  or (_11698_, _11697_, _11649_);
  and (_11699_, _05754_, _03665_);
  nor (_11700_, _11699_, _02804_);
  and (_11701_, _11700_, _11698_);
  and (_11702_, _05684_, _02804_);
  or (_11703_, _11702_, _02514_);
  or (_11704_, _11703_, _11701_);
  and (_11705_, _02514_, \oc8051_golden_model_1.PC [1]);
  nor (_11706_, _11705_, _03888_);
  and (_11707_, _11706_, _11704_);
  and (_11708_, _05178_, _03698_);
  nor (_11709_, _05178_, _03698_);
  nor (_11710_, _11709_, _11708_);
  and (_11711_, _11710_, _03888_);
  or (_11712_, _11711_, _03886_);
  or (_11713_, _11712_, _11707_);
  and (_11714_, _05178_, _02551_);
  nor (_11715_, _11714_, _11587_);
  or (_11716_, _11715_, _05770_);
  and (_11717_, _11716_, _03885_);
  and (_11718_, _11717_, _11713_);
  and (_11719_, _11709_, _03884_);
  or (_11720_, _11719_, _03881_);
  or (_11721_, _11720_, _11718_);
  and (_11722_, _11721_, _11588_);
  or (_11723_, _11722_, _03880_);
  nor (_11724_, _02532_, _02215_);
  nor (_11725_, _11724_, _05784_);
  and (_11726_, _11725_, _11723_);
  nor (_11727_, _11708_, _05790_);
  or (_11728_, _11727_, _05789_);
  or (_11729_, _11728_, _11726_);
  nand (_11730_, _11714_, _05789_);
  and (_11731_, _11730_, _02529_);
  and (_11732_, _11731_, _11729_);
  nor (_11733_, _02529_, \oc8051_golden_model_1.PC [1]);
  or (_11734_, _03317_, _11733_);
  or (_11735_, _11734_, _11732_);
  and (_11736_, _11584_, _03317_);
  nor (_11737_, _11736_, _03303_);
  and (_11738_, _11737_, _11735_);
  or (_11739_, _11738_, _11586_);
  and (_11740_, _11739_, _11585_);
  and (_11741_, _03368_, _02367_);
  nor (_11742_, _11741_, _03303_);
  nor (_11743_, _11742_, _11584_);
  or (_11744_, _11743_, _03575_);
  or (_11745_, _11744_, _11740_);
  or (_11746_, _05941_, _06153_);
  or (_11747_, _11746_, _03909_);
  and (_11748_, _11747_, _04333_);
  and (_11749_, _11748_, _11745_);
  nor (_11750_, _11606_, _04333_);
  or (_11751_, _11750_, _02939_);
  or (_11752_, _11751_, _11749_);
  nand (_11753_, _02939_, _09270_);
  and (_11754_, _11753_, _02526_);
  and (_11755_, _11754_, _11752_);
  and (_11756_, _02525_, _02215_);
  or (_11757_, _02797_, _11756_);
  or (_11758_, _11757_, _11755_);
  or (_11759_, _11636_, _02798_);
  and (_11760_, _11759_, _05237_);
  and (_11761_, _11760_, _11758_);
  and (_11762_, _03920_, _02543_);
  not (_11763_, _05237_);
  and (_11764_, _11584_, _11763_);
  or (_11765_, _11764_, _11762_);
  or (_11766_, _11765_, _11761_);
  not (_11767_, _03585_);
  and (_11768_, _05747_, _02522_);
  not (_11769_, _11768_);
  nor (_11770_, _05941_, _06153_);
  or (_11771_, _11770_, _11769_);
  and (_11772_, _11771_, _11767_);
  and (_11773_, _11772_, _11766_);
  and (_11774_, _11770_, _03585_);
  or (_11775_, _11774_, _03923_);
  or (_11776_, _11775_, _11773_);
  or (_11777_, _11606_, _06150_);
  and (_11778_, _11777_, _04184_);
  and (_11779_, _11778_, _11776_);
  or (_11780_, _11779_, _11583_);
  and (_11781_, _11583_, _03943_);
  nor (_11782_, _11781_, _11572_);
  and (_11783_, _11782_, _11780_);
  nand (_11784_, _09237_, _02939_);
  or (_11785_, _09115_, _02939_);
  and (_11786_, _11785_, _11784_);
  and (_11787_, _11786_, _04544_);
  and (_11788_, _11787_, _11572_);
  or (_40543_, _11788_, _11783_);
  or (_11789_, _11382_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_11790_, _11789_, _11391_);
  nor (_11791_, _05239_, _04435_);
  nor (_11792_, _11791_, _07352_);
  or (_11793_, _11792_, _04119_);
  and (_11794_, _11793_, _11763_);
  nor (_11795_, _09140_, _02529_);
  or (_11796_, _04435_, _11401_);
  nor (_11797_, _10027_, _04611_);
  or (_11798_, _11797_, _05315_);
  and (_11799_, _05467_, _05129_);
  nor (_11800_, _05467_, _05129_);
  nor (_11801_, _11800_, _11799_);
  nand (_11802_, _11801_, _03811_);
  and (_11803_, _05271_, _04494_);
  nor (_11804_, _05271_, _04494_);
  or (_11805_, _11804_, _11803_);
  and (_11806_, _11805_, _05363_);
  nor (_11807_, _09140_, _02611_);
  and (_11808_, _02611_, \oc8051_golden_model_1.ACC [2]);
  or (_11809_, _11808_, _11807_);
  and (_11810_, _11809_, _05362_);
  or (_11811_, _11810_, _03811_);
  or (_11812_, _11811_, _11806_);
  and (_11813_, _11812_, _05358_);
  and (_11814_, _11813_, _11802_);
  nand (_11815_, _10027_, _09733_);
  and (_11816_, _11815_, _02883_);
  or (_11817_, _11816_, _04252_);
  or (_11818_, _11817_, _11814_);
  nor (_11819_, _02648_, _02609_);
  nor (_11820_, _11819_, _03836_);
  and (_11821_, _11820_, _11818_);
  and (_11822_, _04435_, _03836_);
  or (_11823_, _11822_, _03844_);
  or (_11824_, _11823_, _11821_);
  and (_11825_, _11824_, _11798_);
  or (_11826_, _11825_, _02875_);
  nand (_11827_, _07453_, _02875_);
  and (_11828_, _11827_, _02873_);
  and (_11829_, _11828_, _11826_);
  not (_11830_, _10028_);
  and (_11831_, _11815_, _11830_);
  and (_11832_, _11831_, _02872_);
  or (_11833_, _11832_, _11829_);
  and (_11834_, _11833_, _02614_);
  nor (_11835_, _09140_, _02614_);
  or (_11836_, _03059_, _11835_);
  or (_11837_, _11836_, _11834_);
  nand (_11838_, _07453_, _03059_);
  and (_11839_, _11838_, _11837_);
  or (_11840_, _11839_, _03859_);
  and (_11841_, _06155_, _04551_);
  nand (_11842_, _07452_, _03859_);
  or (_11843_, _11842_, _11841_);
  and (_11844_, _11843_, _11840_);
  or (_11845_, _11844_, _03858_);
  nor (_11846_, _09755_, _04611_);
  and (_11847_, _04611_, \oc8051_golden_model_1.PSW [7]);
  nor (_11848_, _11847_, _11846_);
  nand (_11849_, _11848_, _03858_);
  and (_11850_, _11849_, _04251_);
  and (_11851_, _11850_, _11845_);
  and (_11852_, _02648_, _02581_);
  or (_11853_, _05536_, _11852_);
  or (_11854_, _11853_, _11851_);
  and (_11855_, _11854_, _11796_);
  or (_11856_, _11855_, _05541_);
  or (_11857_, _06155_, _05546_);
  and (_11858_, _11857_, _05545_);
  and (_11859_, _11858_, _11856_);
  and (_11860_, _05311_, _04435_);
  not (_11861_, _11860_);
  and (_11862_, _05731_, \oc8051_golden_model_1.SCON [2]);
  and (_11863_, _05726_, \oc8051_golden_model_1.IE [2]);
  nor (_11864_, _11863_, _11862_);
  and (_11865_, _05699_, \oc8051_golden_model_1.TCON [2]);
  and (_11866_, _05729_, \oc8051_golden_model_1.SBUF [2]);
  nor (_11867_, _11866_, _11865_);
  and (_11868_, _11867_, _11864_);
  and (_11869_, _05703_, \oc8051_golden_model_1.PCON [2]);
  and (_11870_, _05692_, \oc8051_golden_model_1.TH0 [2]);
  nor (_11871_, _11870_, _11869_);
  and (_11872_, _05707_, \oc8051_golden_model_1.DPL [2]);
  and (_11873_, _05696_, \oc8051_golden_model_1.TL1 [2]);
  nor (_11874_, _11873_, _11872_);
  and (_11875_, _11874_, _11871_);
  and (_11876_, _11875_, _11868_);
  and (_11877_, _05682_, \oc8051_golden_model_1.SP [2]);
  not (_11878_, _11877_);
  and (_11879_, _05717_, \oc8051_golden_model_1.P1INREG [2]);
  not (_11880_, _11879_);
  and (_11881_, _05710_, \oc8051_golden_model_1.P0INREG [2]);
  not (_11882_, _11881_);
  and (_11883_, _05720_, \oc8051_golden_model_1.P2INREG [2]);
  and (_11884_, _08669_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_11885_, _11884_, _11883_);
  and (_11886_, _11885_, _11882_);
  and (_11887_, _11886_, _11880_);
  and (_11888_, _11887_, _11878_);
  and (_11889_, _05655_, \oc8051_golden_model_1.B [2]);
  and (_11890_, _05652_, \oc8051_golden_model_1.ACC [2]);
  nor (_11891_, _11890_, _11889_);
  and (_11892_, _05664_, \oc8051_golden_model_1.IP [2]);
  and (_11893_, _05668_, \oc8051_golden_model_1.PSW [2]);
  nor (_11894_, _11893_, _11892_);
  and (_11895_, _11894_, _11891_);
  and (_11896_, _05735_, \oc8051_golden_model_1.TMOD [2]);
  and (_11897_, _05737_, \oc8051_golden_model_1.DPH [2]);
  nor (_11898_, _11897_, _11896_);
  and (_11899_, _05687_, \oc8051_golden_model_1.TL0 [2]);
  and (_11900_, _05678_, \oc8051_golden_model_1.TH1 [2]);
  nor (_11901_, _11900_, _11899_);
  and (_11902_, _11901_, _11898_);
  and (_11903_, _11902_, _11895_);
  and (_11904_, _11903_, _11888_);
  and (_11905_, _11904_, _11876_);
  and (_11906_, _11905_, _11861_);
  nor (_11907_, _11906_, _05545_);
  or (_11908_, _11907_, _05754_);
  or (_11909_, _11908_, _11859_);
  and (_11910_, _05754_, _03256_);
  nor (_11911_, _11910_, _02804_);
  and (_11912_, _11911_, _11909_);
  and (_11913_, _05701_, _02804_);
  or (_11914_, _11913_, _02514_);
  or (_11915_, _11914_, _11912_);
  and (_11916_, _09140_, _02514_);
  nor (_11917_, _11916_, _03888_);
  and (_11918_, _11917_, _11915_);
  and (_11919_, _05129_, _03297_);
  nor (_11920_, _05129_, _03297_);
  nor (_11921_, _11920_, _11919_);
  and (_11922_, _11921_, _03888_);
  or (_11923_, _11922_, _11918_);
  and (_11924_, _11923_, _05770_);
  nor (_11925_, _05129_, _06964_);
  and (_11926_, _05129_, _06964_);
  nor (_11927_, _11926_, _11925_);
  and (_11928_, _11927_, _03886_);
  or (_11929_, _11928_, _03884_);
  or (_11930_, _11929_, _11924_);
  or (_11931_, _11920_, _03885_);
  and (_11932_, _11931_, _03882_);
  and (_11933_, _11932_, _11930_);
  and (_11934_, _11925_, _03881_);
  or (_11935_, _11934_, _03880_);
  or (_11936_, _11935_, _11933_);
  nor (_11937_, _02648_, _02532_);
  nor (_11938_, _11937_, _05784_);
  and (_11939_, _11938_, _11936_);
  nor (_11940_, _11919_, _05790_);
  or (_11941_, _11940_, _05789_);
  or (_11942_, _11941_, _11939_);
  nand (_11943_, _11926_, _05789_);
  and (_11944_, _11943_, _02529_);
  and (_11945_, _11944_, _11942_);
  or (_11946_, _11945_, _11795_);
  and (_11947_, _11946_, _05265_);
  not (_11948_, _11741_);
  nor (_11949_, _11586_, _05266_);
  and (_11950_, _11949_, _11948_);
  nand (_11951_, _11805_, _05264_);
  nand (_11952_, _11951_, _11950_);
  or (_11953_, _11952_, _11947_);
  or (_11954_, _11805_, _11950_);
  and (_11955_, _11954_, _03909_);
  and (_11956_, _11955_, _11953_);
  and (_11957_, _05941_, _06031_);
  nor (_11958_, _05941_, _06031_);
  or (_11959_, _11958_, _11957_);
  and (_11960_, _11959_, _03575_);
  or (_11961_, _11960_, _11956_);
  and (_11962_, _11961_, _04333_);
  nor (_11963_, _11801_, _04333_);
  or (_11964_, _11963_, _02939_);
  or (_11965_, _11964_, _11962_);
  nand (_11966_, _09268_, _02939_);
  and (_11967_, _11966_, _02526_);
  and (_11968_, _11967_, _11965_);
  and (_11969_, _02648_, _02525_);
  or (_11970_, _02797_, _11969_);
  or (_11971_, _11970_, _11968_);
  or (_11972_, _11846_, _02798_);
  and (_11973_, _11972_, _06141_);
  and (_11974_, _11973_, _11971_);
  or (_11975_, _11974_, _11794_);
  or (_11976_, _11792_, _05238_);
  and (_11977_, _11976_, _03921_);
  and (_11978_, _11977_, _11975_);
  or (_11979_, _06155_, _06153_);
  nor (_11980_, _07272_, _03921_);
  and (_11981_, _11980_, _11979_);
  or (_11982_, _11981_, _03923_);
  or (_11983_, _11982_, _11978_);
  nor (_11984_, _05227_, _05130_);
  nor (_11985_, _11984_, _05228_);
  or (_11986_, _11985_, _06150_);
  and (_11987_, _11986_, _11373_);
  and (_11988_, _11987_, _11983_);
  or (_11989_, _11988_, _11393_);
  and (_11990_, _11989_, _11790_);
  nand (_11991_, _09229_, _02939_);
  or (_11992_, _09109_, _02939_);
  and (_11993_, _11992_, _11991_);
  and (_11994_, _11993_, _04544_);
  and (_11995_, _11994_, _11572_);
  or (_40545_, _11995_, _11990_);
  or (_11996_, _11382_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_11997_, _11996_, _11391_);
  or (_11998_, _07352_, _04241_);
  nor (_11999_, _05241_, _05237_);
  and (_12000_, _11999_, _11998_);
  nor (_12001_, _11957_, _05986_);
  or (_12002_, _12001_, _06033_);
  and (_12003_, _12002_, _03575_);
  nor (_12004_, _02641_, _02529_);
  nor (_12005_, _10088_, _04670_);
  or (_12006_, _12005_, _05315_);
  nor (_12007_, _11803_, _04311_);
  or (_12008_, _12007_, _05273_);
  or (_12009_, _12008_, _05362_);
  nor (_12010_, _02611_, _02641_);
  nand (_12011_, _02611_, \oc8051_golden_model_1.ACC [3]);
  nand (_12012_, _12011_, _05362_);
  or (_12013_, _12012_, _12010_);
  and (_12014_, _12013_, _12009_);
  and (_12015_, _12014_, _03812_);
  nor (_12016_, _11799_, _05078_);
  nor (_12017_, _12016_, _05469_);
  nor (_12018_, _12017_, _03812_);
  or (_12019_, _12018_, _12015_);
  or (_12020_, _12019_, _02883_);
  nand (_12021_, _10088_, _09863_);
  or (_12022_, _12021_, _05358_);
  and (_12023_, _12022_, _12020_);
  or (_12024_, _12023_, _04252_);
  nor (_12025_, _02609_, _02629_);
  nor (_12026_, _12025_, _03836_);
  and (_12027_, _12026_, _12024_);
  and (_12028_, _04241_, _03836_);
  or (_12029_, _12028_, _03844_);
  or (_12030_, _12029_, _12027_);
  and (_12031_, _12030_, _12006_);
  or (_12032_, _12031_, _02875_);
  nand (_12033_, _07442_, _02875_);
  and (_12034_, _12033_, _02873_);
  and (_12035_, _12034_, _12032_);
  not (_12036_, _10089_);
  and (_12037_, _12021_, _12036_);
  and (_12038_, _12037_, _02872_);
  or (_12039_, _12038_, _12035_);
  and (_12040_, _12039_, _02614_);
  nor (_12041_, _02614_, _02641_);
  or (_12042_, _03059_, _12041_);
  or (_12043_, _12042_, _12040_);
  nand (_12044_, _07442_, _03059_);
  and (_12045_, _12044_, _12043_);
  or (_12046_, _12045_, _03859_);
  or (_12047_, _05986_, _02763_);
  nand (_12048_, _12047_, _07441_);
  or (_12049_, _12048_, _03860_);
  and (_12050_, _12049_, _04298_);
  and (_12051_, _12050_, _12046_);
  and (_12052_, _04670_, \oc8051_golden_model_1.PSW [7]);
  nor (_12053_, _09885_, _04670_);
  nor (_12054_, _12053_, _12052_);
  nor (_12055_, _12054_, _04298_);
  or (_12056_, _12055_, _02581_);
  or (_12057_, _12056_, _12051_);
  and (_12058_, _02581_, _02641_);
  nor (_12059_, _12058_, _05536_);
  and (_12060_, _12059_, _12057_);
  and (_12061_, _04241_, _05536_);
  or (_12062_, _12061_, _05541_);
  or (_12063_, _12062_, _12060_);
  or (_12064_, _06154_, _05546_);
  and (_12065_, _12064_, _05545_);
  and (_12066_, _12065_, _12063_);
  and (_12067_, _05311_, _04241_);
  not (_12068_, _12067_);
  and (_12069_, _05717_, \oc8051_golden_model_1.P1INREG [3]);
  not (_12070_, _12069_);
  and (_12071_, _05710_, \oc8051_golden_model_1.P0INREG [3]);
  not (_12072_, _12071_);
  and (_12073_, _05720_, \oc8051_golden_model_1.P2INREG [3]);
  and (_12074_, _08669_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_12075_, _12074_, _12073_);
  and (_12076_, _12075_, _12072_);
  and (_12077_, _12076_, _12070_);
  and (_12078_, _05682_, \oc8051_golden_model_1.SP [3]);
  and (_12079_, _05687_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12080_, _12079_, _12078_);
  and (_12081_, _12080_, _12077_);
  and (_12082_, _05664_, \oc8051_golden_model_1.IP [3]);
  and (_12083_, _05655_, \oc8051_golden_model_1.B [3]);
  nor (_12084_, _12083_, _12082_);
  and (_12085_, _05668_, \oc8051_golden_model_1.PSW [3]);
  and (_12086_, _05652_, \oc8051_golden_model_1.ACC [3]);
  nor (_12087_, _12086_, _12085_);
  and (_12088_, _12087_, _12084_);
  and (_12089_, _05726_, \oc8051_golden_model_1.IE [3]);
  and (_12090_, _05729_, \oc8051_golden_model_1.SBUF [3]);
  and (_12091_, _05731_, \oc8051_golden_model_1.SCON [3]);
  or (_12092_, _12091_, _12090_);
  nor (_12093_, _12092_, _12089_);
  and (_12094_, _12093_, _12088_);
  and (_12095_, _12094_, _12081_);
  and (_12096_, _05692_, \oc8051_golden_model_1.TH0 [3]);
  and (_12097_, _05696_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12098_, _12097_, _12096_);
  and (_12099_, _05699_, \oc8051_golden_model_1.TCON [3]);
  and (_12100_, _05703_, \oc8051_golden_model_1.PCON [3]);
  nor (_12101_, _12100_, _12099_);
  and (_12102_, _12101_, _12098_);
  and (_12103_, _05737_, \oc8051_golden_model_1.DPH [3]);
  and (_12104_, _05735_, \oc8051_golden_model_1.TMOD [3]);
  nor (_12105_, _12104_, _12103_);
  and (_12106_, _05707_, \oc8051_golden_model_1.DPL [3]);
  and (_12107_, _05678_, \oc8051_golden_model_1.TH1 [3]);
  nor (_12108_, _12107_, _12106_);
  and (_12109_, _12108_, _12105_);
  and (_12110_, _12109_, _12102_);
  and (_12111_, _12110_, _12095_);
  and (_12112_, _12111_, _12068_);
  nor (_12113_, _12112_, _05545_);
  or (_12114_, _12113_, _05754_);
  or (_12115_, _12114_, _12066_);
  and (_12116_, _05754_, _02794_);
  nor (_12117_, _12116_, _02804_);
  and (_12118_, _12117_, _12115_);
  and (_12119_, _05658_, _02804_);
  or (_12120_, _12119_, _02514_);
  or (_12121_, _12120_, _12118_);
  and (_12122_, _02641_, _02514_);
  nor (_12123_, _12122_, _03888_);
  and (_12124_, _12123_, _12121_);
  and (_12125_, _05078_, _03057_);
  nor (_12126_, _05078_, _03057_);
  nor (_12127_, _12126_, _12125_);
  and (_12128_, _12127_, _03888_);
  or (_12129_, _12128_, _12124_);
  and (_12130_, _12129_, _05770_);
  nor (_12131_, _05078_, _02564_);
  and (_12132_, _05078_, _02564_);
  nor (_12133_, _12132_, _12131_);
  and (_12134_, _12133_, _03886_);
  or (_12135_, _12134_, _03884_);
  or (_12136_, _12135_, _12130_);
  or (_12137_, _12126_, _03885_);
  and (_12138_, _12137_, _03882_);
  and (_12139_, _12138_, _12136_);
  and (_12140_, _12131_, _03881_);
  or (_12141_, _12140_, _03880_);
  or (_12142_, _12141_, _12139_);
  nor (_12143_, _02629_, _02532_);
  nor (_12144_, _12143_, _05784_);
  and (_12145_, _12144_, _12142_);
  nor (_12146_, _12125_, _05790_);
  or (_12147_, _12146_, _05789_);
  or (_12148_, _12147_, _12145_);
  nand (_12149_, _12132_, _05789_);
  and (_12150_, _12149_, _02529_);
  and (_12151_, _12150_, _12148_);
  or (_12152_, _12151_, _12004_);
  and (_12153_, _12152_, _05268_);
  not (_12154_, _05268_);
  and (_12155_, _12008_, _12154_);
  or (_12156_, _12155_, _04153_);
  or (_12157_, _12156_, _12153_);
  or (_12158_, _12008_, _05262_);
  and (_12159_, _12158_, _03909_);
  and (_12160_, _12159_, _12157_);
  or (_12161_, _12160_, _12003_);
  and (_12162_, _12161_, _04333_);
  nor (_12163_, _12017_, _04333_);
  or (_12164_, _12163_, _02939_);
  or (_12165_, _12164_, _12162_);
  nand (_12166_, _09263_, _02939_);
  and (_12167_, _12166_, _02526_);
  and (_12168_, _12167_, _12165_);
  and (_12169_, _02629_, _02525_);
  or (_12170_, _02797_, _12169_);
  or (_12171_, _12170_, _12168_);
  or (_12172_, _12053_, _02798_);
  and (_12173_, _12172_, _05237_);
  and (_12174_, _12173_, _12171_);
  or (_12175_, _12174_, _12000_);
  and (_12176_, _12175_, _03921_);
  or (_12177_, _07272_, _06154_);
  nor (_12178_, _06157_, _03921_);
  and (_12179_, _12178_, _12177_);
  or (_12180_, _12179_, _03923_);
  or (_12181_, _12180_, _12176_);
  nor (_12182_, _05228_, _05079_);
  nor (_12183_, _12182_, _05229_);
  or (_12184_, _12183_, _06150_);
  and (_12185_, _12184_, _04184_);
  and (_12186_, _12185_, _12181_);
  or (_12187_, _12186_, _11583_);
  and (_12188_, _12187_, _11997_);
  nand (_12189_, _09223_, _02939_);
  or (_12190_, _09104_, _02939_);
  and (_12191_, _12190_, _12189_);
  and (_12192_, _12191_, _04544_);
  and (_12193_, _12192_, _11572_);
  or (_40546_, _12193_, _12188_);
  or (_12194_, _11382_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_12195_, _12194_, _11391_);
  and (_12196_, _06033_, _06123_);
  nor (_12197_, _06033_, _06123_);
  or (_12198_, _12197_, _12196_);
  and (_12199_, _12198_, _03575_);
  not (_12200_, _04982_);
  nor (_12201_, _05273_, _12200_);
  and (_12202_, _05273_, _12200_);
  or (_12203_, _12202_, _12201_);
  or (_12204_, _12203_, _05268_);
  nor (_12205_, _05030_, _06867_);
  and (_12206_, _05030_, _06867_);
  nor (_12207_, _12206_, _12205_);
  and (_12208_, _12207_, _03886_);
  and (_12209_, _05030_, _05582_);
  nor (_12210_, _05030_, _05582_);
  nor (_12211_, _12210_, _12209_);
  and (_12212_, _12211_, _03888_);
  nor (_12213_, _09783_, _10050_);
  or (_12214_, _12213_, _05315_);
  and (_12215_, _05469_, _05030_);
  nor (_12216_, _05469_, _05030_);
  nor (_12217_, _12216_, _12215_);
  nor (_12218_, _12217_, _03812_);
  or (_12219_, _06159_, _04265_);
  and (_12220_, _12203_, _05363_);
  or (_12221_, _09135_, _02611_);
  nand (_12222_, _02611_, _06867_);
  and (_12223_, _12222_, _12221_);
  and (_12224_, _12223_, _05362_);
  or (_12225_, _12224_, _02886_);
  or (_12226_, _12225_, _12220_);
  and (_12227_, _12226_, _03812_);
  and (_12228_, _12227_, _12219_);
  or (_12229_, _12228_, _12218_);
  and (_12230_, _12229_, _05358_);
  nand (_12231_, _09784_, _10050_);
  and (_12232_, _12231_, _02883_);
  or (_12233_, _12232_, _04252_);
  or (_12234_, _12233_, _12230_);
  nor (_12235_, _09135_, _02609_);
  nor (_12236_, _12235_, _03836_);
  and (_12237_, _12236_, _12234_);
  and (_12238_, _04982_, _03836_);
  or (_12239_, _12238_, _03844_);
  or (_12240_, _12239_, _12237_);
  and (_12241_, _12240_, _12214_);
  or (_12242_, _12241_, _02875_);
  nand (_12243_, _07517_, _02875_);
  and (_12244_, _12243_, _02873_);
  and (_12245_, _12244_, _12242_);
  not (_12246_, _10051_);
  and (_12247_, _12231_, _12246_);
  and (_12248_, _12247_, _02872_);
  or (_12249_, _12248_, _12245_);
  and (_12250_, _12249_, _02614_);
  nor (_12251_, _09136_, _02614_);
  or (_12252_, _12251_, _03059_);
  or (_12253_, _12252_, _12250_);
  nand (_12254_, _07517_, _03059_);
  and (_12255_, _12254_, _12253_);
  or (_12256_, _12255_, _03859_);
  and (_12257_, _06159_, _04551_);
  nand (_12258_, _07516_, _03859_);
  or (_12259_, _12258_, _12257_);
  and (_12260_, _12259_, _04298_);
  and (_12261_, _12260_, _12256_);
  nor (_12262_, _09807_, _09783_);
  and (_12263_, _09783_, \oc8051_golden_model_1.PSW [7]);
  nor (_12264_, _12263_, _12262_);
  nor (_12265_, _12264_, _04298_);
  or (_12266_, _12265_, _02581_);
  or (_12267_, _12266_, _12261_);
  and (_12268_, _09136_, _02581_);
  nor (_12269_, _12268_, _05536_);
  and (_12270_, _12269_, _12267_);
  and (_12271_, _04982_, _05536_);
  or (_12272_, _12271_, _05541_);
  or (_12273_, _12272_, _12270_);
  or (_12274_, _06159_, _05546_);
  and (_12275_, _12274_, _05545_);
  and (_12276_, _12275_, _12273_);
  and (_12277_, _05311_, _04982_);
  not (_12278_, _12277_);
  and (_12279_, _05682_, \oc8051_golden_model_1.SP [4]);
  and (_12280_, _05735_, \oc8051_golden_model_1.TMOD [4]);
  nor (_12281_, _12280_, _12279_);
  and (_12282_, _05707_, \oc8051_golden_model_1.DPL [4]);
  and (_12283_, _05687_, \oc8051_golden_model_1.TL0 [4]);
  nor (_12284_, _12283_, _12282_);
  and (_12285_, _12284_, _12281_);
  and (_12286_, _05726_, \oc8051_golden_model_1.IE [4]);
  and (_12287_, _05729_, \oc8051_golden_model_1.SBUF [4]);
  and (_12288_, _05731_, \oc8051_golden_model_1.SCON [4]);
  or (_12289_, _12288_, _12287_);
  nor (_12290_, _12289_, _12286_);
  and (_12291_, _05710_, \oc8051_golden_model_1.P0INREG [4]);
  not (_12292_, _12291_);
  nand (_12293_, _05714_, \oc8051_golden_model_1.P3INREG [4]);
  and (_12294_, _05717_, \oc8051_golden_model_1.P1INREG [4]);
  and (_12295_, _05720_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_12296_, _12295_, _12294_);
  and (_12297_, _12296_, _12293_);
  and (_12298_, _12297_, _12292_);
  and (_12299_, _12298_, _12290_);
  and (_12300_, _12299_, _12285_);
  and (_12301_, _05692_, \oc8051_golden_model_1.TH0 [4]);
  and (_12302_, _05696_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12303_, _12302_, _12301_);
  and (_12304_, _05699_, \oc8051_golden_model_1.TCON [4]);
  and (_12305_, _05703_, \oc8051_golden_model_1.PCON [4]);
  nor (_12306_, _12305_, _12304_);
  and (_12307_, _12306_, _12303_);
  and (_12308_, _05664_, \oc8051_golden_model_1.IP [4]);
  and (_12309_, _05655_, \oc8051_golden_model_1.B [4]);
  nor (_12310_, _12309_, _12308_);
  and (_12311_, _05668_, \oc8051_golden_model_1.PSW [4]);
  and (_12312_, _05652_, \oc8051_golden_model_1.ACC [4]);
  nor (_12313_, _12312_, _12311_);
  and (_12314_, _12313_, _12310_);
  and (_12315_, _05678_, \oc8051_golden_model_1.TH1 [4]);
  and (_12316_, _05737_, \oc8051_golden_model_1.DPH [4]);
  nor (_12317_, _12316_, _12315_);
  and (_12318_, _12317_, _12314_);
  and (_12319_, _12318_, _12307_);
  and (_12320_, _12319_, _12300_);
  and (_12321_, _12320_, _12278_);
  nor (_12322_, _12321_, _05545_);
  or (_12323_, _12322_, _05754_);
  or (_12324_, _12323_, _12276_);
  and (_12325_, _05754_, _03629_);
  nor (_12326_, _12325_, _02804_);
  and (_12327_, _12326_, _12324_);
  and (_12328_, _05666_, _02804_);
  or (_12329_, _12328_, _02514_);
  or (_12330_, _12329_, _12327_);
  and (_12331_, _09136_, _02514_);
  nor (_12332_, _12331_, _03888_);
  and (_12333_, _12332_, _12330_);
  or (_12334_, _12333_, _12212_);
  and (_12335_, _12334_, _05770_);
  or (_12336_, _12335_, _12208_);
  and (_12337_, _12336_, _03885_);
  and (_12338_, _12210_, _03884_);
  or (_12339_, _12338_, _12337_);
  and (_12340_, _12339_, _03882_);
  and (_12341_, _12205_, _03881_);
  or (_12342_, _12341_, _03880_);
  or (_12343_, _12342_, _12340_);
  nor (_12344_, _09135_, _02532_);
  nor (_12345_, _12344_, _05784_);
  and (_12346_, _12345_, _12343_);
  nor (_12347_, _12209_, _05790_);
  or (_12348_, _12347_, _05789_);
  or (_12349_, _12348_, _12346_);
  nand (_12350_, _12206_, _05789_);
  and (_12351_, _12350_, _02529_);
  and (_12352_, _12351_, _12349_);
  or (_12353_, _09136_, _02529_);
  nand (_12354_, _12353_, _05268_);
  or (_12355_, _12354_, _12352_);
  and (_12356_, _12355_, _12204_);
  or (_12357_, _12356_, _04153_);
  or (_12358_, _12203_, _05262_);
  and (_12359_, _12358_, _03909_);
  and (_12360_, _12359_, _12357_);
  or (_12361_, _12360_, _12199_);
  and (_12362_, _12361_, _04333_);
  nor (_12363_, _12217_, _04333_);
  or (_12364_, _12363_, _02939_);
  or (_12365_, _12364_, _12362_);
  nand (_12366_, _09258_, _02939_);
  and (_12367_, _12366_, _02526_);
  and (_12368_, _12367_, _12365_);
  and (_12369_, _09135_, _02525_);
  or (_12370_, _12369_, _02797_);
  or (_12371_, _12370_, _12368_);
  or (_12372_, _12262_, _02798_);
  and (_12373_, _12372_, _05237_);
  and (_12374_, _12373_, _12371_);
  or (_12375_, _05241_, _04982_);
  nor (_12376_, _05242_, _05237_);
  and (_12377_, _12376_, _12375_);
  or (_12378_, _12377_, _11762_);
  or (_12379_, _12378_, _12374_);
  nor (_12380_, _06159_, _06157_);
  nor (_12381_, _12380_, _07256_);
  or (_12382_, _12381_, _11769_);
  and (_12383_, _12382_, _11767_);
  and (_12384_, _12383_, _12379_);
  and (_12385_, _12381_, _03585_);
  or (_12386_, _12385_, _03923_);
  or (_12387_, _12386_, _12384_);
  nor (_12388_, _05229_, _05031_);
  nor (_12389_, _12388_, _05230_);
  or (_12390_, _12389_, _06150_);
  and (_12391_, _12390_, _04184_);
  and (_12392_, _12391_, _12387_);
  or (_12393_, _12392_, _11583_);
  and (_12394_, _12393_, _12195_);
  not (_12395_, _09101_);
  nor (_12396_, _12395_, _02939_);
  and (_12397_, _09217_, _02939_);
  or (_12398_, _12397_, _12396_);
  and (_12399_, _12398_, _04544_);
  and (_12400_, _12399_, _11572_);
  or (_40547_, _12400_, _12394_);
  or (_12401_, _11382_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_12402_, _12401_, _11391_);
  nor (_12403_, _05242_, _04877_);
  nor (_12404_, _12403_, _05243_);
  and (_12405_, _12404_, _11763_);
  nor (_12406_, _12215_, _04923_);
  nor (_12407_, _12406_, _05470_);
  nand (_12408_, _12407_, _03908_);
  nor (_12409_, _04923_, _06861_);
  and (_12410_, _04923_, _06861_);
  nor (_12411_, _12410_, _12409_);
  and (_12412_, _12411_, _03886_);
  and (_12413_, _04923_, _05613_);
  nor (_12414_, _04923_, _05613_);
  nor (_12415_, _12414_, _12413_);
  and (_12416_, _12415_, _03888_);
  nor (_12417_, _09887_, _10099_);
  or (_12418_, _12417_, _05315_);
  nor (_12419_, _12407_, _03812_);
  or (_12420_, _06158_, _04265_);
  not (_12421_, _04877_);
  nor (_12422_, _12202_, _12421_);
  or (_12423_, _12422_, _05274_);
  and (_12424_, _12423_, _05363_);
  or (_12425_, _09130_, _02611_);
  nand (_12426_, _02611_, _06861_);
  and (_12427_, _12426_, _12425_);
  and (_12428_, _12427_, _05362_);
  or (_12429_, _12428_, _02886_);
  or (_12430_, _12429_, _12424_);
  and (_12431_, _12430_, _03812_);
  and (_12432_, _12431_, _12420_);
  or (_12433_, _12432_, _12419_);
  and (_12434_, _12433_, _05358_);
  nand (_12435_, _09888_, _10099_);
  and (_12436_, _12435_, _02883_);
  or (_12437_, _12436_, _04252_);
  or (_12438_, _12437_, _12434_);
  nor (_12439_, _09130_, _02609_);
  nor (_12440_, _12439_, _03836_);
  and (_12441_, _12440_, _12438_);
  and (_12442_, _04877_, _03836_);
  or (_12443_, _12442_, _03844_);
  or (_12444_, _12443_, _12441_);
  and (_12445_, _12444_, _12418_);
  or (_12446_, _12445_, _02875_);
  nand (_12447_, _07504_, _02875_);
  and (_12448_, _12447_, _02873_);
  and (_12449_, _12448_, _12446_);
  not (_12450_, _10100_);
  and (_12451_, _12435_, _12450_);
  and (_12452_, _12451_, _02872_);
  or (_12453_, _12452_, _12449_);
  and (_12454_, _12453_, _02614_);
  nor (_12455_, _09131_, _02614_);
  or (_12456_, _12455_, _03059_);
  or (_12457_, _12456_, _12454_);
  nand (_12458_, _07504_, _03059_);
  and (_12459_, _12458_, _12457_);
  or (_12460_, _12459_, _03859_);
  and (_12461_, _06158_, _04551_);
  nand (_12462_, _07503_, _03859_);
  or (_12463_, _12462_, _12461_);
  and (_12464_, _12463_, _04298_);
  and (_12465_, _12464_, _12460_);
  nor (_12466_, _09911_, _09887_);
  and (_12467_, _09887_, \oc8051_golden_model_1.PSW [7]);
  nor (_12468_, _12467_, _12466_);
  nor (_12469_, _12468_, _04298_);
  or (_12470_, _12469_, _02581_);
  or (_12471_, _12470_, _12465_);
  and (_12472_, _09131_, _02581_);
  nor (_12473_, _12472_, _05536_);
  and (_12474_, _12473_, _12471_);
  and (_12475_, _04877_, _05536_);
  or (_12476_, _12475_, _05541_);
  or (_12477_, _12476_, _12474_);
  or (_12478_, _06158_, _05546_);
  and (_12479_, _12478_, _05545_);
  and (_12480_, _12479_, _12477_);
  and (_12481_, _05311_, _04877_);
  not (_12482_, _12481_);
  and (_12483_, _05655_, \oc8051_golden_model_1.B [5]);
  and (_12484_, _05652_, \oc8051_golden_model_1.ACC [5]);
  nor (_12485_, _12484_, _12483_);
  and (_12486_, _05664_, \oc8051_golden_model_1.IP [5]);
  and (_12487_, _05668_, \oc8051_golden_model_1.PSW [5]);
  nor (_12488_, _12487_, _12486_);
  and (_12489_, _12488_, _12485_);
  and (_12490_, _05735_, \oc8051_golden_model_1.TMOD [5]);
  and (_12491_, _05737_, \oc8051_golden_model_1.DPH [5]);
  nor (_12492_, _12491_, _12490_);
  and (_12493_, _05687_, \oc8051_golden_model_1.TL0 [5]);
  and (_12494_, _05678_, \oc8051_golden_model_1.TH1 [5]);
  nor (_12495_, _12494_, _12493_);
  and (_12496_, _12495_, _12492_);
  and (_12497_, _12496_, _12489_);
  and (_12498_, _05714_, \oc8051_golden_model_1.P3INREG [5]);
  not (_12499_, _12498_);
  and (_12500_, _05717_, \oc8051_golden_model_1.P1INREG [5]);
  and (_12501_, _05720_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_12502_, _12501_, _12500_);
  and (_12503_, _12502_, _12499_);
  and (_12504_, _05726_, \oc8051_golden_model_1.IE [5]);
  not (_12505_, _12504_);
  and (_12506_, _05731_, \oc8051_golden_model_1.SCON [5]);
  and (_12507_, _05729_, \oc8051_golden_model_1.SBUF [5]);
  nor (_12508_, _12507_, _12506_);
  and (_12509_, _12508_, _12505_);
  and (_12510_, _12509_, _12503_);
  and (_12511_, _05692_, \oc8051_golden_model_1.TH0 [5]);
  and (_12512_, _05696_, \oc8051_golden_model_1.TL1 [5]);
  nor (_12513_, _12512_, _12511_);
  and (_12514_, _05699_, \oc8051_golden_model_1.TCON [5]);
  and (_12515_, _05703_, \oc8051_golden_model_1.PCON [5]);
  nor (_12516_, _12515_, _12514_);
  and (_12517_, _12516_, _12513_);
  and (_12518_, _05707_, \oc8051_golden_model_1.DPL [5]);
  not (_12519_, _12518_);
  and (_12520_, _05682_, \oc8051_golden_model_1.SP [5]);
  and (_12521_, _05710_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_12522_, _12521_, _12520_);
  and (_12523_, _12522_, _12519_);
  and (_12524_, _12523_, _12517_);
  and (_12525_, _12524_, _12510_);
  and (_12526_, _12525_, _12497_);
  and (_12527_, _12526_, _12482_);
  nor (_12528_, _12527_, _05545_);
  or (_12529_, _12528_, _05754_);
  or (_12530_, _12529_, _12480_);
  and (_12531_, _05754_, _03211_);
  nor (_12532_, _12531_, _02804_);
  and (_12533_, _12532_, _12530_);
  and (_12534_, _05614_, _02804_);
  or (_12535_, _12534_, _02514_);
  or (_12536_, _12535_, _12533_);
  and (_12537_, _09131_, _02514_);
  nor (_12538_, _12537_, _03888_);
  and (_12539_, _12538_, _12536_);
  or (_12540_, _12539_, _12416_);
  and (_12541_, _12540_, _05770_);
  or (_12542_, _12541_, _12412_);
  and (_12543_, _12542_, _03885_);
  and (_12544_, _12414_, _03884_);
  or (_12545_, _12544_, _12543_);
  and (_12546_, _12545_, _03882_);
  and (_12547_, _12409_, _03881_);
  or (_12548_, _12547_, _03880_);
  or (_12549_, _12548_, _12546_);
  nor (_12550_, _09130_, _02532_);
  nor (_12551_, _12550_, _05784_);
  and (_12552_, _12551_, _12549_);
  nor (_12553_, _12413_, _05790_);
  or (_12554_, _12553_, _05789_);
  or (_12555_, _12554_, _12552_);
  nand (_12556_, _12410_, _05789_);
  and (_12557_, _12556_, _02529_);
  and (_12558_, _12557_, _12555_);
  or (_12559_, _09131_, _02529_);
  nand (_12560_, _12559_, _09940_);
  or (_12561_, _12560_, _12558_);
  or (_12562_, _12423_, _09940_);
  and (_12563_, _12562_, _03909_);
  and (_12564_, _12563_, _12561_);
  nor (_12565_, _12196_, _06078_);
  or (_12566_, _12565_, _06125_);
  and (_12567_, _12566_, _03575_);
  or (_12568_, _12567_, _03908_);
  or (_12569_, _12568_, _12564_);
  and (_12570_, _12569_, _12408_);
  or (_12571_, _12570_, _02939_);
  nand (_12572_, _09253_, _02939_);
  and (_12573_, _12572_, _02526_);
  and (_12574_, _12573_, _12571_);
  and (_12575_, _09130_, _02525_);
  or (_12576_, _12575_, _02797_);
  or (_12577_, _12576_, _12574_);
  or (_12578_, _12466_, _02798_);
  and (_12579_, _12578_, _05237_);
  and (_12580_, _12579_, _12577_);
  or (_12581_, _12580_, _12405_);
  and (_12582_, _12581_, _03921_);
  or (_12583_, _07256_, _06158_);
  nor (_12584_, _06161_, _03921_);
  and (_12585_, _12584_, _12583_);
  or (_12586_, _12585_, _03923_);
  or (_12587_, _12586_, _12582_);
  nor (_12588_, _05230_, _04924_);
  nor (_12589_, _12588_, _05231_);
  or (_12590_, _12589_, _06150_);
  and (_12591_, _12590_, _11373_);
  and (_12592_, _12591_, _12587_);
  or (_12593_, _12592_, _11393_);
  and (_12594_, _12593_, _12402_);
  nand (_12595_, _09213_, _02939_);
  or (_12596_, _09097_, _02939_);
  and (_12597_, _12596_, _12595_);
  and (_12598_, _12597_, _04544_);
  and (_12599_, _12598_, _11572_);
  or (_40548_, _12599_, _12594_);
  or (_12600_, _11382_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_12601_, _12600_, _11391_);
  nor (_12602_, _05470_, _04818_);
  nor (_12603_, _12602_, _05471_);
  nor (_12604_, _12603_, _04333_);
  nor (_12605_, _06125_, _05850_);
  or (_12606_, _12605_, _06126_);
  and (_12607_, _12606_, _03575_);
  nor (_12608_, _05274_, _05269_);
  or (_12609_, _12608_, _05275_);
  or (_12610_, _12609_, _05268_);
  nor (_12611_, _04818_, _06806_);
  and (_12612_, _04818_, _06806_);
  nor (_12613_, _12612_, _12611_);
  and (_12614_, _12613_, _03886_);
  or (_12615_, _04770_, _11401_);
  nor (_12616_, _09837_, _10075_);
  or (_12617_, _12616_, _05315_);
  nand (_12618_, _09838_, _10075_);
  or (_12619_, _12618_, _05358_);
  or (_12620_, _12609_, _05362_);
  nor (_12621_, _09124_, _02611_);
  and (_12622_, _02611_, \oc8051_golden_model_1.ACC [6]);
  nor (_12623_, _12622_, _12621_);
  nand (_12624_, _12623_, _05362_);
  and (_12625_, _12624_, _12620_);
  or (_12626_, _12625_, _02886_);
  or (_12627_, _05849_, _04265_);
  and (_12628_, _12627_, _12626_);
  or (_12629_, _12628_, _03811_);
  nand (_12630_, _12603_, _03811_);
  and (_12631_, _12630_, _12629_);
  or (_12632_, _12631_, _02883_);
  and (_12633_, _12632_, _12619_);
  or (_12634_, _12633_, _04252_);
  nor (_12635_, _09123_, _02609_);
  nor (_12636_, _12635_, _03836_);
  and (_12637_, _12636_, _12634_);
  and (_12638_, _04770_, _03836_);
  or (_12639_, _12638_, _03844_);
  or (_12640_, _12639_, _12637_);
  and (_12641_, _12640_, _12617_);
  or (_12642_, _12641_, _02875_);
  nand (_12643_, _07424_, _02875_);
  and (_12644_, _12643_, _02873_);
  and (_12645_, _12644_, _12642_);
  not (_12646_, _10076_);
  and (_12647_, _12618_, _12646_);
  and (_12648_, _12647_, _02872_);
  or (_12649_, _12648_, _12645_);
  and (_12650_, _12649_, _02614_);
  nor (_12651_, _09124_, _02614_);
  or (_12652_, _12651_, _03059_);
  or (_12653_, _12652_, _12650_);
  nand (_12654_, _07424_, _03059_);
  and (_12655_, _12654_, _12653_);
  or (_12656_, _12655_, _03859_);
  and (_12657_, _05849_, _04551_);
  nand (_12658_, _07423_, _03859_);
  or (_12659_, _12658_, _12657_);
  and (_12660_, _12659_, _12656_);
  or (_12661_, _12660_, _03858_);
  nor (_12662_, _09860_, _09837_);
  and (_12663_, _09837_, \oc8051_golden_model_1.PSW [7]);
  nor (_12664_, _12663_, _12662_);
  nand (_12665_, _12664_, _03858_);
  and (_12666_, _12665_, _04251_);
  and (_12667_, _12666_, _12661_);
  and (_12668_, _09123_, _02581_);
  or (_12669_, _12668_, _05536_);
  or (_12670_, _12669_, _12667_);
  and (_12671_, _12670_, _12615_);
  or (_12672_, _12671_, _05541_);
  or (_12673_, _05849_, _05546_);
  and (_12674_, _12673_, _05545_);
  and (_12675_, _12674_, _12672_);
  and (_12676_, _05311_, _04770_);
  not (_12677_, _12676_);
  and (_12678_, _05664_, \oc8051_golden_model_1.IP [6]);
  and (_12679_, _05655_, \oc8051_golden_model_1.B [6]);
  nor (_12680_, _12679_, _12678_);
  and (_12681_, _05668_, \oc8051_golden_model_1.PSW [6]);
  and (_12682_, _05652_, \oc8051_golden_model_1.ACC [6]);
  nor (_12683_, _12682_, _12681_);
  and (_12684_, _12683_, _12680_);
  and (_12685_, _05678_, \oc8051_golden_model_1.TH1 [6]);
  not (_12686_, _12685_);
  and (_12687_, _05682_, \oc8051_golden_model_1.SP [6]);
  and (_12688_, _05687_, \oc8051_golden_model_1.TL0 [6]);
  nor (_12689_, _12688_, _12687_);
  and (_12690_, _12689_, _12686_);
  and (_12691_, _12690_, _12684_);
  and (_12692_, _05692_, \oc8051_golden_model_1.TH0 [6]);
  and (_12693_, _05696_, \oc8051_golden_model_1.TL1 [6]);
  nor (_12694_, _12693_, _12692_);
  and (_12695_, _05699_, \oc8051_golden_model_1.TCON [6]);
  and (_12696_, _05703_, \oc8051_golden_model_1.PCON [6]);
  nor (_12697_, _12696_, _12695_);
  and (_12698_, _12697_, _12694_);
  and (_12699_, _05707_, \oc8051_golden_model_1.DPL [6]);
  not (_12700_, _12699_);
  and (_12701_, _05710_, \oc8051_golden_model_1.P0INREG [6]);
  not (_12702_, _12701_);
  nand (_12703_, _05714_, \oc8051_golden_model_1.P3INREG [6]);
  and (_12704_, _05717_, \oc8051_golden_model_1.P1INREG [6]);
  and (_12705_, _05720_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_12706_, _12705_, _12704_);
  and (_12707_, _12706_, _12703_);
  and (_12708_, _12707_, _12702_);
  and (_12709_, _12708_, _12700_);
  and (_12710_, _05726_, \oc8051_golden_model_1.IE [6]);
  and (_12711_, _05729_, \oc8051_golden_model_1.SBUF [6]);
  and (_12712_, _05731_, \oc8051_golden_model_1.SCON [6]);
  or (_12713_, _12712_, _12711_);
  nor (_12714_, _12713_, _12710_);
  and (_12715_, _05735_, \oc8051_golden_model_1.TMOD [6]);
  and (_12716_, _05737_, \oc8051_golden_model_1.DPH [6]);
  nor (_12717_, _12716_, _12715_);
  and (_12718_, _12717_, _12714_);
  and (_12719_, _12718_, _12709_);
  and (_12720_, _12719_, _12698_);
  and (_12721_, _12720_, _12691_);
  and (_12722_, _12721_, _12677_);
  nor (_12723_, _12722_, _05545_);
  or (_12724_, _12723_, _05754_);
  or (_12725_, _12724_, _12675_);
  and (_12726_, _05754_, _02927_);
  nor (_12727_, _12726_, _02804_);
  and (_12728_, _12727_, _12725_);
  not (_12729_, _05649_);
  and (_12730_, _12729_, _02804_);
  or (_12731_, _12730_, _02514_);
  or (_12732_, _12731_, _12728_);
  and (_12733_, _09124_, _02514_);
  nor (_12734_, _12733_, _03888_);
  and (_12735_, _12734_, _12732_);
  and (_12737_, _04818_, _05649_);
  nor (_12738_, _04818_, _05649_);
  nor (_12739_, _12738_, _12737_);
  and (_12740_, _12739_, _03888_);
  or (_12741_, _12740_, _12735_);
  and (_12742_, _12741_, _05770_);
  or (_12743_, _12742_, _12614_);
  and (_12744_, _12743_, _03885_);
  and (_12745_, _12738_, _03884_);
  or (_12746_, _12745_, _12744_);
  and (_12747_, _12746_, _03882_);
  and (_12748_, _12611_, _03881_);
  or (_12749_, _12748_, _03880_);
  or (_12750_, _12749_, _12747_);
  nor (_12751_, _09123_, _02532_);
  nor (_12752_, _12751_, _05784_);
  and (_12753_, _12752_, _12750_);
  nor (_12754_, _12737_, _05790_);
  or (_12755_, _12754_, _05789_);
  or (_12756_, _12755_, _12753_);
  nand (_12758_, _12612_, _05789_);
  and (_12759_, _12758_, _02529_);
  and (_12760_, _12759_, _12756_);
  or (_12761_, _09124_, _02529_);
  nand (_12762_, _12761_, _05268_);
  or (_12763_, _12762_, _12760_);
  and (_12764_, _12763_, _12610_);
  or (_12765_, _12764_, _04153_);
  or (_12766_, _12609_, _05262_);
  and (_12767_, _12766_, _03909_);
  and (_12768_, _12767_, _12765_);
  or (_12769_, _12768_, _12607_);
  and (_12770_, _12769_, _04333_);
  or (_12771_, _12770_, _12604_);
  and (_12772_, _12771_, _06173_);
  and (_12773_, _09245_, _02939_);
  or (_12774_, _12773_, _02525_);
  or (_12775_, _12774_, _12772_);
  and (_12776_, _09124_, _02525_);
  nor (_12777_, _12776_, _02797_);
  and (_12778_, _12777_, _12775_);
  and (_12779_, _12662_, _02797_);
  or (_12780_, _12779_, _11763_);
  or (_12781_, _12780_, _12778_);
  nor (_12782_, _05269_, _05243_);
  and (_12783_, _05269_, _05243_);
  or (_12784_, _12783_, _12782_);
  or (_12785_, _12784_, _05237_);
  and (_12786_, _12785_, _03921_);
  and (_12787_, _12786_, _12781_);
  nor (_12788_, _06161_, _05849_);
  nor (_12789_, _12788_, _06162_);
  and (_12790_, _12789_, _03920_);
  or (_12791_, _12790_, _03923_);
  or (_12792_, _12791_, _12787_);
  nor (_12793_, _05231_, _04819_);
  nor (_12794_, _12793_, _05232_);
  or (_12795_, _12794_, _06150_);
  and (_12796_, _12795_, _11373_);
  and (_12797_, _12796_, _12792_);
  or (_12798_, _12797_, _11393_);
  and (_12799_, _12798_, _12601_);
  not (_12800_, _09086_);
  nor (_12801_, _12800_, _02939_);
  and (_12802_, _09207_, _02939_);
  or (_12803_, _12802_, _12801_);
  and (_12804_, _12803_, _04544_);
  and (_12805_, _12804_, _11572_);
  or (_40549_, _12805_, _12799_);
  or (_12806_, _11382_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_12807_, _12806_, _11391_);
  or (_12808_, _11583_, _06170_);
  and (_12809_, _12808_, _12807_);
  and (_12810_, _11572_, _06208_);
  or (_40550_, _12810_, _12809_);
  and (_12811_, _11375_, _04092_);
  and (_12812_, _12811_, _11380_);
  or (_12813_, _12812_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_12814_, _04243_);
  or (_12815_, _11389_, _12814_);
  or (_12816_, _12815_, _11385_);
  and (_12817_, _12816_, _12813_);
  and (_12818_, _11566_, _04184_);
  nand (_12819_, _11578_, _04092_);
  or (_12820_, _12819_, _11581_);
  or (_12821_, _12820_, _12818_);
  and (_12822_, _12821_, _12817_);
  and (_12823_, _04544_, _04243_);
  and (_12824_, _12823_, _11570_);
  and (_12825_, _12824_, _11576_);
  or (_40554_, _12825_, _12822_);
  or (_12826_, _12812_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_12827_, _12826_, _12816_);
  and (_12828_, _11777_, _11373_);
  and (_12829_, _12828_, _11776_);
  not (_12830_, _12812_);
  or (_12831_, _12830_, _12829_);
  and (_12832_, _12831_, _12827_);
  and (_12833_, _12824_, _11787_);
  or (_40555_, _12833_, _12832_);
  or (_12834_, _12812_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_12835_, _12834_, _12816_);
  or (_12836_, _12830_, _11988_);
  and (_12837_, _12836_, _12835_);
  and (_12838_, _12824_, _11994_);
  or (_40556_, _12838_, _12837_);
  or (_12839_, _12812_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_12840_, _12839_, _12816_);
  or (_12841_, _12820_, _12186_);
  and (_12842_, _12841_, _12840_);
  and (_12843_, _12824_, _12192_);
  or (_40557_, _12843_, _12842_);
  or (_12844_, _12812_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_12845_, _12844_, _12816_);
  or (_12846_, _12820_, _12392_);
  and (_12847_, _12846_, _12845_);
  and (_12848_, _12824_, _12399_);
  or (_40559_, _12848_, _12847_);
  or (_12849_, _12812_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_12850_, _12849_, _12816_);
  or (_12851_, _12830_, _12592_);
  and (_12852_, _12851_, _12850_);
  and (_12853_, _12824_, _12598_);
  or (_40560_, _12853_, _12852_);
  or (_12854_, _12812_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_12855_, _12854_, _12816_);
  or (_12856_, _12830_, _12797_);
  and (_12857_, _12856_, _12855_);
  and (_12858_, _12824_, _12804_);
  or (_40561_, _12858_, _12857_);
  or (_12859_, _12812_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_12860_, _12859_, _12816_);
  or (_12861_, _12820_, _06170_);
  and (_12862_, _12861_, _12860_);
  and (_12863_, _12824_, _06208_);
  or (_40562_, _12863_, _12862_);
  and (_12864_, _11376_, _03929_);
  and (_12865_, _12864_, _11380_);
  or (_12866_, _12865_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_12867_, _05376_);
  or (_12868_, _11389_, _12867_);
  or (_12869_, _12868_, _11385_);
  and (_12870_, _12869_, _12866_);
  and (_12871_, _04186_, _03929_);
  not (_12872_, _12871_);
  nor (_12873_, _12872_, _11581_);
  not (_12874_, _12873_);
  or (_12875_, _12874_, _12818_);
  and (_12876_, _12875_, _12870_);
  and (_12877_, _05376_, _04544_);
  and (_12878_, _12877_, _11570_);
  and (_12879_, _12878_, _11576_);
  or (_40566_, _12879_, _12876_);
  or (_12880_, _12865_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_12881_, _12880_, _12869_);
  or (_12882_, _12874_, _11779_);
  and (_12883_, _12882_, _12881_);
  and (_12884_, _12878_, _11787_);
  or (_40567_, _12884_, _12883_);
  and (_12885_, _11986_, _04184_);
  and (_12886_, _12885_, _11983_);
  or (_12887_, _12874_, _12886_);
  nor (_12888_, _12873_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_12889_, _12888_, _12878_);
  and (_12890_, _12889_, _12887_);
  and (_12891_, _12878_, _11994_);
  or (_40568_, _12891_, _12890_);
  or (_12892_, _12865_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_12893_, _12892_, _12869_);
  or (_12894_, _12874_, _12186_);
  and (_12895_, _12894_, _12893_);
  and (_12896_, _12878_, _12192_);
  or (_40569_, _12896_, _12895_);
  or (_12897_, _12865_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_12898_, _12897_, _12869_);
  or (_12899_, _12874_, _12392_);
  and (_12900_, _12899_, _12898_);
  and (_12901_, _12878_, _12399_);
  or (_40570_, _12901_, _12900_);
  or (_12902_, _12865_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_12903_, _12902_, _12869_);
  and (_12904_, _12590_, _04184_);
  and (_12905_, _12904_, _12587_);
  or (_12906_, _12874_, _12905_);
  and (_12907_, _12906_, _12903_);
  and (_12908_, _12878_, _12598_);
  or (_40571_, _12908_, _12907_);
  or (_12909_, _12865_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_12910_, _12909_, _12869_);
  and (_12911_, _12795_, _04184_);
  and (_12912_, _12911_, _12792_);
  or (_12913_, _12874_, _12912_);
  and (_12914_, _12913_, _12910_);
  and (_12915_, _12878_, _12804_);
  or (_40573_, _12915_, _12914_);
  or (_12916_, _12865_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_12917_, _12916_, _12869_);
  or (_12918_, _12874_, _06170_);
  and (_12919_, _12918_, _12917_);
  and (_12920_, _12878_, _06208_);
  or (_40574_, _12920_, _12919_);
  not (_12921_, _04092_);
  and (_12922_, _11375_, _12921_);
  and (_12923_, _11380_, _12922_);
  or (_12924_, _12923_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_12925_, _03932_);
  or (_12926_, _11389_, _12925_);
  or (_12927_, _12926_, _11385_);
  and (_12928_, _12927_, _12924_);
  not (_12929_, _04187_);
  nor (_12930_, _11581_, _12929_);
  not (_12931_, _12930_);
  or (_12932_, _12931_, _12818_);
  and (_12933_, _12932_, _12928_);
  and (_12934_, _04544_, _03932_);
  and (_12935_, _12934_, _11570_);
  and (_12936_, _12935_, _11576_);
  or (_40577_, _12936_, _12933_);
  or (_12937_, _12923_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_12938_, _12937_, _12927_);
  or (_12939_, _12931_, _11779_);
  and (_12940_, _12939_, _12938_);
  and (_12941_, _12935_, _11787_);
  or (_40578_, _12941_, _12940_);
  or (_12942_, _12931_, _12886_);
  nor (_12943_, _12930_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_12944_, _12943_, _12935_);
  and (_12945_, _12944_, _12942_);
  and (_12946_, _12935_, _11994_);
  or (_40579_, _12946_, _12945_);
  or (_12947_, _12923_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_12948_, _12947_, _12927_);
  or (_12949_, _12931_, _12186_);
  and (_12950_, _12949_, _12948_);
  and (_12951_, _12935_, _12192_);
  or (_40580_, _12951_, _12950_);
  or (_12952_, _12923_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_12953_, _12952_, _12927_);
  or (_12954_, _12931_, _12392_);
  and (_12955_, _12954_, _12953_);
  and (_12956_, _12935_, _12399_);
  or (_40582_, _12956_, _12955_);
  or (_12957_, _12923_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_12958_, _12957_, _12927_);
  or (_12959_, _12931_, _12905_);
  and (_12960_, _12959_, _12958_);
  and (_12961_, _12935_, _12598_);
  or (_40583_, _12961_, _12960_);
  or (_12962_, _12923_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_12963_, _12962_, _12927_);
  or (_12964_, _12931_, _12912_);
  and (_12965_, _12964_, _12963_);
  and (_12966_, _12935_, _12804_);
  or (_40584_, _12966_, _12965_);
  or (_12967_, _12923_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_12968_, _12967_, _12927_);
  or (_12969_, _12931_, _06170_);
  and (_12970_, _12969_, _12968_);
  and (_12971_, _12935_, _06208_);
  or (_40585_, _12971_, _12970_);
  and (_12972_, _04532_, _04351_);
  and (_12973_, _12972_, _11579_);
  not (_12974_, _12973_);
  or (_12975_, _12974_, _12818_);
  not (_12976_, _04542_);
  and (_12977_, _11569_, _12976_);
  and (_12978_, _12977_, _03933_);
  nor (_12979_, _12973_, \oc8051_golden_model_1.IRAM[4] [0]);
  nor (_12980_, _12979_, _12978_);
  and (_12981_, _12980_, _12975_);
  and (_12982_, _12978_, _11576_);
  or (_40588_, _12982_, _12981_);
  or (_12983_, _12974_, _11779_);
  nor (_12984_, _12973_, \oc8051_golden_model_1.IRAM[4] [1]);
  nor (_12985_, _12984_, _12978_);
  and (_12986_, _12985_, _12983_);
  and (_12987_, _12978_, _11787_);
  or (_40590_, _12987_, _12986_);
  or (_12988_, _12974_, _12886_);
  nor (_12989_, _12973_, \oc8051_golden_model_1.IRAM[4] [2]);
  nor (_12990_, _12989_, _12978_);
  and (_12991_, _12990_, _12988_);
  and (_12992_, _12978_, _11994_);
  or (_40591_, _12992_, _12991_);
  or (_12993_, _12974_, _12186_);
  nor (_12994_, _12973_, \oc8051_golden_model_1.IRAM[4] [3]);
  nor (_12995_, _12994_, _12978_);
  and (_12996_, _12995_, _12993_);
  and (_12997_, _12978_, _12192_);
  or (_40592_, _12997_, _12996_);
  or (_12998_, _12974_, _12392_);
  and (_12999_, _11387_, _12976_);
  nand (_13000_, _12999_, _03933_);
  or (_13001_, _12973_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13002_, _13001_, _13000_);
  and (_13003_, _13002_, _12998_);
  and (_13004_, _12978_, _12399_);
  or (_40593_, _13004_, _13003_);
  or (_13005_, _12973_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_13006_, _13005_, _13000_);
  or (_13007_, _12974_, _12592_);
  and (_13008_, _13007_, _13006_);
  and (_13009_, _12978_, _12598_);
  or (_40594_, _13009_, _13008_);
  or (_13010_, _12974_, _12797_);
  or (_13011_, _12973_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13012_, _13011_, _13000_);
  and (_13013_, _13012_, _13010_);
  and (_13014_, _12978_, _12804_);
  or (_40596_, _13014_, _13013_);
  or (_13015_, _12974_, _06170_);
  or (_13016_, _12973_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13017_, _13016_, _13000_);
  and (_13018_, _13017_, _13015_);
  and (_13019_, _12978_, _06208_);
  or (_40597_, _13019_, _13018_);
  not (_13020_, _12972_);
  nor (_13021_, _13020_, _12819_);
  not (_13022_, _13021_);
  or (_13023_, _13022_, _12818_);
  and (_13024_, _12999_, _04243_);
  not (_13025_, _13024_);
  or (_13026_, _13021_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_13027_, _13026_, _13025_);
  and (_13028_, _13027_, _13023_);
  and (_13029_, _13024_, _11576_);
  or (_40600_, _13029_, _13028_);
  or (_13030_, _13022_, _11779_);
  or (_13031_, _13021_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13032_, _13031_, _13025_);
  and (_13033_, _13032_, _13030_);
  and (_13034_, _13024_, _11787_);
  or (_40601_, _13034_, _13033_);
  or (_13035_, _13022_, _12886_);
  or (_13036_, _13021_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13037_, _13036_, _13025_);
  and (_13038_, _13037_, _13035_);
  and (_13039_, _13024_, _11994_);
  or (_40602_, _13039_, _13038_);
  or (_13040_, _13022_, _12186_);
  or (_13041_, _13021_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_13042_, _13041_, _13025_);
  and (_13043_, _13042_, _13040_);
  and (_13044_, _13024_, _12192_);
  or (_40603_, _13044_, _13043_);
  and (_13045_, _13024_, _12399_);
  or (_13046_, _13021_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13047_, _13046_, _13025_);
  or (_13048_, _13022_, _12392_);
  and (_13049_, _13048_, _13047_);
  or (_40604_, _13049_, _13045_);
  and (_13050_, _13024_, _12598_);
  or (_13051_, _13021_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_13052_, _13051_, _13025_);
  or (_13053_, _13022_, _12905_);
  and (_13054_, _13053_, _13052_);
  or (_40606_, _13054_, _13050_);
  and (_13055_, _13024_, _12804_);
  or (_13056_, _13021_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13057_, _13056_, _13025_);
  or (_13058_, _13022_, _12912_);
  and (_13059_, _13058_, _13057_);
  or (_40607_, _13059_, _13055_);
  and (_13060_, _13024_, _06208_);
  or (_13061_, _13021_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_13062_, _13061_, _13025_);
  or (_13063_, _13022_, _06170_);
  and (_13064_, _13063_, _13062_);
  or (_40608_, _13064_, _13060_);
  and (_13065_, _12972_, _12871_);
  not (_13066_, _13065_);
  or (_13067_, _13066_, _12818_);
  and (_13068_, _12977_, _05376_);
  nor (_13069_, _13065_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_13070_, _13069_, _13068_);
  and (_13071_, _13070_, _13067_);
  and (_13072_, _13068_, _11576_);
  or (_40611_, _13072_, _13071_);
  or (_13073_, _13066_, _11779_);
  nor (_13074_, _13065_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_13075_, _13074_, _13068_);
  and (_13076_, _13075_, _13073_);
  and (_13077_, _13068_, _11787_);
  or (_40612_, _13077_, _13076_);
  or (_13078_, _13066_, _12886_);
  nor (_13079_, _13065_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_13080_, _13079_, _13068_);
  and (_13081_, _13080_, _13078_);
  and (_13082_, _13068_, _11994_);
  or (_40613_, _13082_, _13081_);
  or (_13083_, _13066_, _12186_);
  nor (_13084_, _13065_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_13085_, _13084_, _13068_);
  and (_13086_, _13085_, _13083_);
  and (_13087_, _13068_, _12192_);
  or (_40614_, _13087_, _13086_);
  nand (_13088_, _12999_, _05376_);
  or (_13089_, _13065_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13090_, _13089_, _13088_);
  or (_13091_, _13066_, _12392_);
  and (_13092_, _13091_, _13090_);
  and (_13093_, _13068_, _12399_);
  or (_40615_, _13093_, _13092_);
  or (_13094_, _13065_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_13095_, _13094_, _13088_);
  or (_13096_, _13066_, _12905_);
  and (_13097_, _13096_, _13095_);
  and (_13098_, _13068_, _12598_);
  or (_40617_, _13098_, _13097_);
  or (_13099_, _13065_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13100_, _13099_, _13088_);
  or (_13101_, _13066_, _12912_);
  and (_13102_, _13101_, _13100_);
  and (_13103_, _13068_, _12804_);
  or (_40618_, _13103_, _13102_);
  or (_13104_, _13065_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13105_, _13104_, _13088_);
  or (_13106_, _13066_, _06170_);
  and (_13107_, _13106_, _13105_);
  and (_13108_, _13068_, _06208_);
  or (_40619_, _13108_, _13107_);
  and (_13109_, _12972_, _04187_);
  not (_13110_, _13109_);
  or (_13111_, _13110_, _12818_);
  and (_13112_, _12977_, _03932_);
  nor (_13113_, _13109_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_13114_, _13113_, _13112_);
  and (_13115_, _13114_, _13111_);
  and (_13116_, _13112_, _11576_);
  or (_40622_, _13116_, _13115_);
  or (_13117_, _13110_, _11779_);
  nor (_13118_, _13109_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_13119_, _13118_, _13112_);
  and (_13120_, _13119_, _13117_);
  and (_13121_, _13112_, _11787_);
  or (_40623_, _13121_, _13120_);
  or (_13122_, _13110_, _12886_);
  nor (_13123_, _13109_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_13124_, _13123_, _13112_);
  and (_13125_, _13124_, _13122_);
  and (_13126_, _13112_, _11994_);
  or (_40624_, _13126_, _13125_);
  or (_13127_, _13110_, _12186_);
  nor (_13128_, _13109_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_13129_, _13128_, _13112_);
  and (_13130_, _13129_, _13127_);
  and (_13131_, _13112_, _12192_);
  or (_40625_, _13131_, _13130_);
  nand (_13132_, _12999_, _03932_);
  or (_13133_, _13109_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13134_, _13133_, _13132_);
  or (_13135_, _13110_, _12392_);
  and (_13136_, _13135_, _13134_);
  and (_13137_, _13112_, _12399_);
  or (_40627_, _13137_, _13136_);
  or (_13138_, _13109_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_13139_, _13138_, _13132_);
  or (_13140_, _13110_, _12905_);
  and (_13141_, _13140_, _13139_);
  and (_13142_, _13112_, _12598_);
  or (_40628_, _13142_, _13141_);
  or (_13143_, _13109_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13144_, _13143_, _13132_);
  or (_13145_, _13110_, _12912_);
  and (_13146_, _13145_, _13144_);
  and (_13147_, _13112_, _12804_);
  or (_40629_, _13147_, _13146_);
  or (_13148_, _13109_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13149_, _13148_, _13132_);
  or (_13150_, _13110_, _06170_);
  and (_13151_, _13150_, _13149_);
  and (_13152_, _13112_, _06208_);
  or (_40630_, _13152_, _13151_);
  and (_13153_, _11378_, _04531_);
  and (_13154_, _13153_, _11377_);
  or (_13155_, _13154_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_13156_, _04539_);
  and (_13157_, _04545_, _13156_);
  and (_13158_, _13157_, _03933_);
  not (_13159_, _13158_);
  and (_13160_, _13159_, _13155_);
  and (_13161_, _11580_, _04531_);
  and (_13162_, _13161_, _11579_);
  not (_13163_, _13162_);
  or (_13164_, _13163_, _12818_);
  and (_13165_, _13164_, _13160_);
  and (_13166_, _13158_, _11576_);
  or (_40633_, _13166_, _13165_);
  or (_13167_, _13163_, _11779_);
  or (_13168_, _13162_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13169_, _13168_, _13159_);
  and (_13170_, _13169_, _13167_);
  and (_13171_, _13158_, _11787_);
  or (_40634_, _13171_, _13170_);
  or (_13172_, _13163_, _12886_);
  or (_13173_, _13162_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13174_, _13173_, _13159_);
  and (_13175_, _13174_, _13172_);
  and (_13176_, _13158_, _11994_);
  or (_40635_, _13176_, _13175_);
  or (_13177_, _13163_, _12186_);
  or (_13178_, _13162_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13179_, _13178_, _13159_);
  and (_13180_, _13179_, _13177_);
  and (_13181_, _13158_, _12192_);
  or (_40636_, _13181_, _13180_);
  or (_13182_, _13154_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13183_, _13182_, _13159_);
  or (_13184_, _13163_, _12392_);
  and (_13185_, _13184_, _13183_);
  and (_13186_, _13158_, _12399_);
  or (_40637_, _13186_, _13185_);
  or (_13187_, _13154_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13188_, _13187_, _13159_);
  not (_13189_, _13154_);
  or (_13190_, _13189_, _12592_);
  and (_13191_, _13190_, _13188_);
  and (_13192_, _13158_, _12598_);
  or (_40638_, _13192_, _13191_);
  or (_13193_, _13154_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13194_, _13193_, _13159_);
  or (_13195_, _13189_, _12797_);
  and (_13196_, _13195_, _13194_);
  and (_13197_, _13158_, _12804_);
  or (_40640_, _13197_, _13196_);
  or (_13198_, _13154_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_13199_, _13198_, _13159_);
  or (_13200_, _13163_, _06170_);
  and (_13201_, _13200_, _13199_);
  and (_13202_, _13158_, _06208_);
  or (_40641_, _13202_, _13201_);
  and (_13203_, _13153_, _12811_);
  or (_13204_, _13203_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_13205_, _11388_, _04244_);
  and (_13206_, _13205_, _13204_);
  not (_13207_, _13161_);
  or (_13208_, _13207_, _12819_);
  or (_13209_, _13208_, _12818_);
  and (_13210_, _13209_, _13206_);
  and (_13211_, _13157_, _04243_);
  and (_13212_, _13211_, _11576_);
  or (_40645_, _13212_, _13210_);
  or (_13213_, _13203_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13214_, _13213_, _13205_);
  not (_13215_, _13203_);
  or (_13216_, _13215_, _12829_);
  and (_13217_, _13216_, _13214_);
  and (_13218_, _13211_, _11787_);
  or (_40646_, _13218_, _13217_);
  or (_13219_, _13203_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13220_, _13219_, _13205_);
  or (_13221_, _13215_, _11988_);
  and (_13222_, _13221_, _13220_);
  and (_13223_, _13211_, _11994_);
  or (_40647_, _13223_, _13222_);
  nor (_13224_, _13208_, _12186_);
  nor (_13225_, _13203_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_13226_, _13225_, _13211_);
  nor (_13227_, _13226_, _13224_);
  and (_13228_, _13211_, _12192_);
  or (_40648_, _13228_, _13227_);
  or (_13229_, _13203_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13230_, _13229_, _13205_);
  or (_13231_, _13208_, _12392_);
  and (_13232_, _13231_, _13230_);
  and (_13233_, _13211_, _12399_);
  or (_40649_, _13233_, _13232_);
  or (_13234_, _13203_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_13235_, _13234_, _13205_);
  or (_13236_, _13215_, _12592_);
  and (_13237_, _13236_, _13235_);
  and (_13238_, _13211_, _12598_);
  or (_40651_, _13238_, _13237_);
  or (_13239_, _13203_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13240_, _13239_, _13205_);
  or (_13241_, _13215_, _12797_);
  and (_13242_, _13241_, _13240_);
  and (_13243_, _13211_, _12804_);
  or (_40652_, _13243_, _13242_);
  or (_13244_, _13203_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13245_, _13244_, _13205_);
  or (_13246_, _13208_, _06170_);
  and (_13247_, _13246_, _13245_);
  and (_13248_, _13211_, _06208_);
  or (_40653_, _13248_, _13247_);
  and (_13249_, _13161_, _12871_);
  or (_13250_, _13249_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13251_, _13157_, _05376_);
  not (_13252_, _13251_);
  and (_13253_, _13252_, _13250_);
  not (_13254_, _13249_);
  or (_13255_, _13254_, _12818_);
  and (_13256_, _13255_, _13253_);
  and (_13257_, _13251_, _11576_);
  or (_40656_, _13257_, _13256_);
  or (_13258_, _13254_, _11779_);
  or (_13259_, _13249_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13260_, _13259_, _13252_);
  and (_13261_, _13260_, _13258_);
  and (_13262_, _13251_, _11787_);
  or (_40657_, _13262_, _13261_);
  or (_13263_, _13254_, _12886_);
  or (_13264_, _13249_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13265_, _13264_, _13252_);
  and (_13266_, _13265_, _13263_);
  and (_13267_, _13251_, _11994_);
  or (_40658_, _13267_, _13266_);
  or (_13268_, _13254_, _12186_);
  or (_13269_, _13249_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13270_, _13269_, _13252_);
  and (_13271_, _13270_, _13268_);
  and (_13272_, _13251_, _12192_);
  or (_40659_, _13272_, _13271_);
  or (_13273_, _13249_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13274_, _13273_, _13252_);
  or (_13275_, _13254_, _12392_);
  and (_13276_, _13275_, _13274_);
  and (_13277_, _13251_, _12399_);
  or (_40660_, _13277_, _13276_);
  or (_13278_, _13249_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13279_, _13278_, _13252_);
  or (_13280_, _13254_, _12905_);
  and (_13281_, _13280_, _13279_);
  and (_13282_, _13251_, _12598_);
  or (_40662_, _13282_, _13281_);
  or (_13283_, _13249_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13284_, _13283_, _13252_);
  or (_13285_, _13254_, _12912_);
  and (_13286_, _13285_, _13284_);
  and (_13287_, _13251_, _12804_);
  or (_40663_, _13287_, _13286_);
  or (_13288_, _13249_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13289_, _13288_, _13252_);
  or (_13290_, _13254_, _06170_);
  and (_13291_, _13290_, _13289_);
  and (_13292_, _13251_, _06208_);
  or (_40664_, _13292_, _13291_);
  and (_13293_, _13161_, _04187_);
  not (_13294_, _13293_);
  or (_13295_, _13294_, _12818_);
  and (_13296_, _13157_, _03932_);
  not (_13297_, _13296_);
  or (_13298_, _13293_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13299_, _13298_, _13297_);
  and (_13300_, _13299_, _13295_);
  and (_13301_, _13296_, _11576_);
  or (_40667_, _13301_, _13300_);
  and (_13302_, _13153_, _12922_);
  or (_13303_, _13302_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13304_, _13303_, _13297_);
  not (_13305_, _13302_);
  or (_13306_, _13305_, _12829_);
  and (_13307_, _13306_, _13304_);
  and (_13308_, _13296_, _11787_);
  or (_40668_, _13308_, _13307_);
  or (_13309_, _13302_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13310_, _13309_, _13297_);
  or (_13311_, _13305_, _11988_);
  and (_13312_, _13311_, _13310_);
  and (_13313_, _13296_, _11994_);
  or (_40669_, _13313_, _13312_);
  or (_13314_, _13294_, _12186_);
  or (_13315_, _13302_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13316_, _13315_, _13297_);
  and (_13317_, _13316_, _13314_);
  and (_13318_, _13296_, _12192_);
  or (_40670_, _13318_, _13317_);
  or (_13319_, _13302_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13320_, _13319_, _13297_);
  or (_13321_, _13294_, _12392_);
  and (_13322_, _13321_, _13320_);
  and (_13323_, _13296_, _12399_);
  or (_40672_, _13323_, _13322_);
  or (_13324_, _13302_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_13325_, _13324_, _13297_);
  or (_13326_, _13305_, _12592_);
  and (_13327_, _13326_, _13325_);
  and (_13328_, _13296_, _12598_);
  or (_40673_, _13328_, _13327_);
  or (_13329_, _13302_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_13330_, _13329_, _13297_);
  or (_13331_, _13305_, _12797_);
  and (_13332_, _13331_, _13330_);
  and (_13333_, _13296_, _12804_);
  or (_40674_, _13333_, _13332_);
  or (_13334_, _13302_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_13335_, _13334_, _13297_);
  or (_13336_, _13294_, _06170_);
  and (_13337_, _13336_, _13335_);
  and (_13338_, _13296_, _06208_);
  or (_40675_, _13338_, _13337_);
  and (_13339_, _11579_, _04533_);
  not (_13340_, _13339_);
  or (_13341_, _13340_, _12818_);
  and (_13342_, _04546_, _03933_);
  not (_13343_, _13342_);
  or (_13344_, _13339_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_13345_, _13344_, _13343_);
  and (_13346_, _13345_, _13341_);
  and (_13347_, _13342_, _11576_);
  or (_40678_, _13347_, _13346_);
  or (_13348_, _13340_, _11779_);
  or (_13349_, _13339_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_13350_, _13349_, _13343_);
  and (_13351_, _13350_, _13348_);
  and (_13352_, _13342_, _11787_);
  or (_40679_, _13352_, _13351_);
  or (_13353_, _13340_, _12886_);
  or (_13354_, _13339_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_13355_, _13354_, _13343_);
  and (_13356_, _13355_, _13353_);
  and (_13357_, _13342_, _11994_);
  or (_40680_, _13357_, _13356_);
  or (_13358_, _13340_, _12186_);
  or (_13359_, _13339_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_13360_, _13359_, _13343_);
  and (_13361_, _13360_, _13358_);
  and (_13362_, _13342_, _12192_);
  or (_40681_, _13362_, _13361_);
  or (_13363_, _13339_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_13364_, _13363_, _13343_);
  or (_13365_, _13340_, _12392_);
  and (_13366_, _13365_, _13364_);
  and (_13367_, _13342_, _12399_);
  or (_40682_, _13367_, _13366_);
  or (_13368_, _13339_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_13369_, _13368_, _13343_);
  or (_13370_, _13340_, _12905_);
  and (_13371_, _13370_, _13369_);
  and (_13372_, _13342_, _12598_);
  or (_40683_, _13372_, _13371_);
  or (_13373_, _13339_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_13374_, _13373_, _13343_);
  or (_13375_, _13340_, _12912_);
  and (_13376_, _13375_, _13374_);
  and (_13377_, _13342_, _12804_);
  or (_40684_, _13377_, _13376_);
  or (_13378_, _13339_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_13379_, _13378_, _13343_);
  or (_13380_, _13340_, _06170_);
  and (_13381_, _13380_, _13379_);
  and (_13382_, _13342_, _06208_);
  or (_40685_, _13382_, _13381_);
  not (_13383_, _04533_);
  nor (_13384_, _12819_, _13383_);
  not (_13385_, _13384_);
  or (_13386_, _13385_, _12818_);
  and (_13387_, _04546_, _04243_);
  not (_13388_, _13387_);
  or (_13389_, _13384_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_13390_, _13389_, _13388_);
  and (_13391_, _13390_, _13386_);
  and (_13392_, _13387_, _11576_);
  or (_40688_, _13392_, _13391_);
  not (_13393_, _04531_);
  and (_13394_, _11378_, _13393_);
  nand (_13395_, _12811_, _13394_);
  nand (_13396_, _13395_, _03992_);
  and (_13397_, _13396_, _13388_);
  or (_13398_, _13395_, _12829_);
  and (_13399_, _13398_, _13397_);
  and (_13400_, _13387_, _11787_);
  or (_40689_, _13400_, _13399_);
  nand (_13401_, _13395_, _04427_);
  and (_13402_, _13401_, _13388_);
  or (_13403_, _13395_, _11988_);
  and (_13404_, _13403_, _13402_);
  and (_13405_, _13387_, _11994_);
  or (_40691_, _13405_, _13404_);
  or (_13406_, _13385_, _12186_);
  nand (_13407_, _13395_, _04233_);
  and (_13408_, _13407_, _13388_);
  and (_13409_, _13408_, _13406_);
  and (_13410_, _13387_, _12192_);
  or (_40692_, _13410_, _13409_);
  nand (_13411_, _13395_, _04974_);
  and (_13412_, _13411_, _13388_);
  or (_13413_, _13385_, _12392_);
  and (_13414_, _13413_, _13412_);
  and (_13415_, _13387_, _12399_);
  or (_40693_, _13415_, _13414_);
  nand (_13416_, _13395_, _04869_);
  and (_13417_, _13416_, _13388_);
  or (_13418_, _13395_, _12592_);
  and (_13419_, _13418_, _13417_);
  and (_13420_, _13387_, _12598_);
  or (_40694_, _13420_, _13419_);
  nand (_13421_, _13395_, _04762_);
  and (_13422_, _13421_, _13388_);
  or (_13423_, _13395_, _12797_);
  and (_13424_, _13423_, _13422_);
  and (_13425_, _13387_, _12804_);
  or (_40695_, _13425_, _13424_);
  or (_13426_, _13384_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_13427_, _13426_, _13388_);
  or (_13428_, _13385_, _06170_);
  and (_13429_, _13428_, _13427_);
  and (_13430_, _13387_, _06208_);
  or (_40697_, _13430_, _13429_);
  and (_13431_, _12871_, _04533_);
  not (_13432_, _13431_);
  or (_13433_, _13432_, _12818_);
  and (_13434_, _05376_, _04546_);
  not (_13435_, _13434_);
  or (_13436_, _13431_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_13437_, _13436_, _13435_);
  and (_13438_, _13437_, _13433_);
  and (_13439_, _13434_, _11576_);
  or (_40699_, _13439_, _13438_);
  or (_13440_, _13432_, _11779_);
  or (_13441_, _13431_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_13442_, _13441_, _13435_);
  and (_13443_, _13442_, _13440_);
  and (_13444_, _13434_, _11787_);
  or (_40700_, _13444_, _13443_);
  or (_13445_, _13432_, _12886_);
  or (_13446_, _13431_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_13447_, _13446_, _13435_);
  and (_13448_, _13447_, _13445_);
  and (_13449_, _13434_, _11994_);
  or (_40702_, _13449_, _13448_);
  or (_13450_, _13432_, _12186_);
  or (_13451_, _13431_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_13452_, _13451_, _13435_);
  and (_13453_, _13452_, _13450_);
  and (_13454_, _13434_, _12192_);
  or (_40703_, _13454_, _13453_);
  or (_13455_, _13431_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_13456_, _13455_, _13435_);
  or (_13457_, _13432_, _12392_);
  and (_13458_, _13457_, _13456_);
  and (_13459_, _13434_, _12399_);
  or (_40704_, _13459_, _13458_);
  or (_13460_, _13431_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_13461_, _13460_, _13435_);
  or (_13462_, _13432_, _12905_);
  and (_13463_, _13462_, _13461_);
  and (_13464_, _13434_, _12598_);
  or (_40705_, _13464_, _13463_);
  or (_13465_, _13431_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_13466_, _13465_, _13435_);
  or (_13467_, _13432_, _12912_);
  and (_13468_, _13467_, _13466_);
  and (_13469_, _13434_, _12804_);
  or (_40706_, _13469_, _13468_);
  or (_13470_, _13431_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_13471_, _13470_, _13435_);
  or (_13472_, _13432_, _06170_);
  and (_13473_, _13472_, _13471_);
  and (_13474_, _13434_, _06208_);
  or (_40707_, _13474_, _13473_);
  or (_13475_, _12818_, _04550_);
  or (_13476_, _04534_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_13477_, _13476_, _04548_);
  and (_13478_, _13477_, _13475_);
  and (_13479_, _11576_, _04547_);
  or (_40710_, _13479_, _13478_);
  or (_13480_, _11779_, _04550_);
  or (_13481_, _04534_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_13482_, _13481_, _04548_);
  and (_13483_, _13482_, _13480_);
  and (_13484_, _11787_, _04547_);
  or (_40711_, _13484_, _13483_);
  or (_13485_, _12886_, _04550_);
  or (_13486_, _04534_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_13487_, _13486_, _04548_);
  and (_13488_, _13487_, _13485_);
  and (_13489_, _11994_, _04547_);
  or (_40712_, _13489_, _13488_);
  or (_13490_, _12186_, _04550_);
  or (_13491_, _04534_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_13492_, _13491_, _04548_);
  and (_13493_, _13492_, _13490_);
  and (_13494_, _12192_, _04547_);
  or (_40713_, _13494_, _13493_);
  or (_13495_, _04534_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_13496_, _13495_, _04548_);
  or (_13497_, _12392_, _04550_);
  and (_13498_, _13497_, _13496_);
  and (_13499_, _12399_, _04547_);
  or (_40714_, _13499_, _13498_);
  or (_13500_, _12905_, _04550_);
  or (_13501_, _04534_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_13502_, _13501_, _04548_);
  and (_13503_, _13502_, _13500_);
  and (_13504_, _12598_, _04547_);
  or (_40715_, _13504_, _13503_);
  or (_13505_, _12912_, _04550_);
  or (_13506_, _04534_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_13507_, _13506_, _04548_);
  and (_13508_, _13507_, _13505_);
  and (_13509_, _12804_, _04547_);
  or (_40716_, _13509_, _13508_);
  nor (_13510_, _42668_, _06825_);
  nor (_13511_, _04696_, _06825_);
  and (_13512_, _11522_, _04696_);
  or (_13513_, _13512_, _13511_);
  and (_13514_, _13513_, _03127_);
  and (_13515_, _04696_, _05672_);
  or (_13516_, _13515_, _13511_);
  or (_13517_, _13516_, _02803_);
  and (_13518_, _04696_, _03808_);
  or (_13519_, _13518_, _13511_);
  or (_13520_, _13519_, _05535_);
  and (_13521_, _05226_, _04696_);
  or (_13522_, _13521_, _13511_);
  or (_13523_, _13522_, _03810_);
  and (_13524_, _04696_, \oc8051_golden_model_1.ACC [0]);
  or (_13525_, _13524_, _13511_);
  and (_13526_, _13525_, _03813_);
  nor (_13527_, _03813_, _06825_);
  or (_13528_, _13527_, _02974_);
  or (_13529_, _13528_, _13526_);
  and (_13530_, _13529_, _02881_);
  and (_13531_, _13530_, _13523_);
  and (_13532_, _11417_, _05333_);
  nor (_13533_, _05333_, _06825_);
  or (_13534_, _13533_, _13532_);
  and (_13535_, _13534_, _02880_);
  or (_13536_, _13535_, _13531_);
  and (_13537_, _13536_, _03336_);
  and (_13538_, _13519_, _03069_);
  or (_13539_, _13538_, _03075_);
  or (_13540_, _13539_, _13537_);
  or (_13541_, _13525_, _03084_);
  and (_13542_, _13541_, _02877_);
  and (_13543_, _13542_, _13540_);
  and (_13544_, _13511_, _02876_);
  or (_13545_, _13544_, _02869_);
  or (_13546_, _13545_, _13543_);
  or (_13547_, _13522_, _02870_);
  and (_13548_, _13547_, _13546_);
  or (_13549_, _13548_, _06247_);
  nor (_13550_, _06729_, _06727_);
  nor (_13551_, _13550_, _06730_);
  or (_13552_, _13551_, _06253_);
  and (_13553_, _13552_, _02864_);
  and (_13554_, _13553_, _13549_);
  nor (_13555_, _11448_, _06771_);
  or (_13556_, _13555_, _13533_);
  and (_13558_, _13556_, _02863_);
  or (_13559_, _13558_, _06770_);
  or (_13560_, _13559_, _13554_);
  and (_13561_, _13560_, _13520_);
  or (_13562_, _13561_, _02853_);
  and (_13563_, _04696_, _06152_);
  or (_13564_, _13511_, _05540_);
  or (_13565_, _13564_, _13563_);
  and (_13566_, _13565_, _13562_);
  or (_13567_, _13566_, _02579_);
  nor (_13569_, _11505_, _06785_);
  or (_13570_, _13511_, _02838_);
  or (_13571_, _13570_, _13569_);
  and (_13572_, _13571_, _06791_);
  and (_13573_, _13572_, _13567_);
  nor (_13574_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_13575_, _13574_, _06708_);
  or (_13576_, _07138_, _13575_);
  nand (_13577_, _07138_, _02667_);
  and (_13578_, _13577_, _06784_);
  and (_13580_, _13578_, _13576_);
  or (_13581_, _13580_, _02802_);
  or (_13582_, _13581_, _13573_);
  and (_13583_, _13582_, _13517_);
  or (_13584_, _13583_, _02980_);
  and (_13585_, _11399_, _04696_);
  or (_13586_, _13511_, _03887_);
  or (_13587_, _13586_, _13585_);
  and (_13588_, _13587_, _03128_);
  and (_13589_, _13588_, _13584_);
  or (_13591_, _13589_, _13514_);
  and (_13592_, _13591_, _03883_);
  nand (_13593_, _13516_, _02970_);
  nor (_13594_, _13593_, _13521_);
  or (_13595_, _13594_, _13592_);
  and (_13596_, _13595_, _03137_);
  or (_13597_, _13511_, _09409_);
  and (_13598_, _13525_, _03135_);
  and (_13599_, _13598_, _13597_);
  or (_13600_, _13599_, _02965_);
  or (_13602_, _13600_, _13596_);
  nor (_13603_, _11396_, _06785_);
  or (_13604_, _13511_, _05783_);
  or (_13605_, _13604_, _13603_);
  and (_13606_, _13605_, _05788_);
  and (_13607_, _13606_, _13602_);
  nor (_13608_, _11520_, _06785_);
  or (_13609_, _13608_, _13511_);
  and (_13610_, _13609_, _03123_);
  or (_13611_, _13610_, _03163_);
  or (_13613_, _13611_, _13607_);
  or (_13614_, _13522_, _03906_);
  and (_13615_, _13614_, _02498_);
  and (_13616_, _13615_, _13613_);
  and (_13617_, _13511_, _02497_);
  or (_13618_, _13617_, _02888_);
  or (_13619_, _13618_, _13616_);
  or (_13620_, _13522_, _02890_);
  and (_13621_, _13620_, _42668_);
  and (_13622_, _13621_, _13619_);
  or (_13624_, _13622_, _13510_);
  and (_43414_, _13624_, _43998_);
  nor (_13625_, _42668_, _06796_);
  or (_13626_, _04696_, \oc8051_golden_model_1.B [1]);
  nand (_13627_, _04696_, _03698_);
  and (_13628_, _13627_, _02802_);
  and (_13629_, _13628_, _13626_);
  nor (_13630_, _05333_, _06796_);
  and (_13631_, _11595_, _05333_);
  or (_13632_, _13631_, _13630_);
  and (_13634_, _13632_, _02876_);
  nor (_13635_, _04696_, _06796_);
  and (_13636_, _04696_, _04000_);
  or (_13637_, _13636_, _13635_);
  or (_13638_, _13637_, _03336_);
  and (_13639_, _11606_, _04696_);
  not (_13640_, _13639_);
  and (_13641_, _13640_, _13626_);
  or (_13642_, _13641_, _03810_);
  nand (_13643_, _04696_, _02551_);
  and (_13645_, _13643_, _13626_);
  and (_13646_, _13645_, _03813_);
  nor (_13647_, _03813_, _06796_);
  or (_13648_, _13647_, _02974_);
  or (_13649_, _13648_, _13646_);
  and (_13650_, _13649_, _02881_);
  and (_13651_, _13650_, _13642_);
  and (_13652_, _11592_, _05333_);
  or (_13653_, _13652_, _13630_);
  and (_13654_, _13653_, _02880_);
  or (_13656_, _13654_, _03069_);
  or (_13657_, _13656_, _13651_);
  and (_13658_, _13657_, _13638_);
  or (_13659_, _13658_, _03075_);
  or (_13660_, _13645_, _03084_);
  and (_13661_, _13660_, _02877_);
  and (_13662_, _13661_, _13659_);
  or (_13663_, _13662_, _13634_);
  and (_13664_, _13663_, _02870_);
  and (_13665_, _13652_, _11591_);
  or (_13667_, _13665_, _13630_);
  and (_13668_, _13667_, _02869_);
  or (_13669_, _13668_, _06247_);
  or (_13670_, _13669_, _13664_);
  nor (_13671_, _06733_, _06675_);
  nor (_13672_, _13671_, _06734_);
  or (_13673_, _13672_, _06253_);
  and (_13674_, _13673_, _02864_);
  and (_13675_, _13674_, _13670_);
  nor (_13676_, _11638_, _06771_);
  or (_13678_, _13676_, _13630_);
  and (_13679_, _13678_, _02863_);
  or (_13680_, _13679_, _06770_);
  or (_13681_, _13680_, _13675_);
  or (_13682_, _13637_, _05535_);
  and (_13683_, _13682_, _13681_);
  or (_13684_, _13683_, _02853_);
  and (_13685_, _04696_, _06151_);
  or (_13686_, _13635_, _05540_);
  or (_13687_, _13686_, _13685_);
  and (_13689_, _13687_, _02838_);
  and (_13690_, _13689_, _13684_);
  nand (_13691_, _11695_, _04696_);
  and (_13692_, _13626_, _02579_);
  and (_13693_, _13692_, _13691_);
  or (_13694_, _13693_, _06784_);
  or (_13695_, _13694_, _13690_);
  nor (_13696_, _07133_, _07132_);
  or (_13697_, _13696_, _07134_);
  nor (_13698_, _13697_, _07138_);
  and (_13700_, _07138_, _07104_);
  or (_13701_, _13700_, _13698_);
  or (_13702_, _13701_, _06791_);
  and (_13703_, _13702_, _02803_);
  and (_13704_, _13703_, _13695_);
  or (_13705_, _13704_, _13629_);
  and (_13706_, _13705_, _03887_);
  or (_13707_, _11710_, _06785_);
  and (_13708_, _13626_, _02980_);
  and (_13709_, _13708_, _13707_);
  or (_13710_, _13709_, _13706_);
  and (_13711_, _13710_, _03128_);
  or (_13712_, _11715_, _06785_);
  and (_13713_, _13626_, _03127_);
  and (_13714_, _13713_, _13712_);
  or (_13715_, _13714_, _13711_);
  and (_13716_, _13715_, _03883_);
  or (_13717_, _11709_, _06785_);
  and (_13718_, _13626_, _02970_);
  and (_13719_, _13718_, _13717_);
  or (_13720_, _13719_, _13716_);
  and (_13721_, _13720_, _03137_);
  not (_13722_, _05178_);
  or (_13723_, _13635_, _13722_);
  and (_13724_, _13645_, _03135_);
  and (_13725_, _13724_, _13723_);
  or (_13726_, _13725_, _13721_);
  and (_13727_, _13726_, _03124_);
  or (_13728_, _13643_, _13722_);
  and (_13729_, _13626_, _03123_);
  and (_13730_, _13729_, _13728_);
  or (_13731_, _13627_, _13722_);
  and (_13732_, _13626_, _02965_);
  and (_13733_, _13732_, _13731_);
  or (_13734_, _13733_, _03163_);
  or (_13735_, _13734_, _13730_);
  or (_13736_, _13735_, _13727_);
  or (_13737_, _13641_, _03906_);
  and (_13738_, _13737_, _02498_);
  and (_13739_, _13738_, _13736_);
  and (_13740_, _13632_, _02497_);
  or (_13741_, _13740_, _02888_);
  or (_13742_, _13741_, _13739_);
  or (_13743_, _13635_, _02890_);
  or (_13744_, _13743_, _13639_);
  and (_13745_, _13744_, _42668_);
  and (_13746_, _13745_, _13742_);
  or (_13747_, _13746_, _13625_);
  and (_43415_, _13747_, _43998_);
  nor (_13748_, _42668_, _06850_);
  nor (_13749_, _04696_, _06850_);
  and (_13750_, _11927_, _04696_);
  or (_13751_, _13750_, _13749_);
  and (_13752_, _13751_, _03127_);
  and (_13753_, _04696_, _05701_);
  or (_13754_, _13753_, _13749_);
  or (_13755_, _13754_, _02803_);
  and (_13756_, _04696_, _04435_);
  or (_13757_, _13756_, _13749_);
  or (_13758_, _13757_, _05535_);
  and (_13759_, _11815_, _05333_);
  and (_13760_, _13759_, _11830_);
  nor (_13761_, _05333_, _06850_);
  or (_13762_, _13761_, _02870_);
  or (_13763_, _13762_, _13760_);
  or (_13764_, _13757_, _03336_);
  nor (_13765_, _11801_, _06785_);
  or (_13766_, _13765_, _13749_);
  or (_13767_, _13766_, _03810_);
  and (_13768_, _04696_, \oc8051_golden_model_1.ACC [2]);
  or (_13769_, _13768_, _13749_);
  and (_13770_, _13769_, _03813_);
  nor (_13771_, _03813_, _06850_);
  or (_13772_, _13771_, _02974_);
  or (_13773_, _13772_, _13770_);
  and (_13774_, _13773_, _02881_);
  and (_13775_, _13774_, _13767_);
  or (_13776_, _13761_, _13759_);
  and (_13777_, _13776_, _02880_);
  or (_13778_, _13777_, _03069_);
  or (_13779_, _13778_, _13775_);
  and (_13780_, _13779_, _13764_);
  or (_13781_, _13780_, _03075_);
  or (_13782_, _13769_, _03084_);
  and (_13783_, _13782_, _02877_);
  and (_13784_, _13783_, _13781_);
  and (_13785_, _11797_, _05333_);
  or (_13786_, _13785_, _13761_);
  and (_13787_, _13786_, _02876_);
  or (_13788_, _13787_, _02869_);
  or (_13789_, _13788_, _13784_);
  and (_13790_, _13789_, _13763_);
  or (_13791_, _13790_, _06247_);
  nor (_13792_, _06736_, _06630_);
  nor (_13793_, _13792_, _06737_);
  or (_13794_, _13793_, _06253_);
  and (_13795_, _13794_, _02864_);
  and (_13796_, _13795_, _13791_);
  nor (_13797_, _11848_, _06771_);
  or (_13798_, _13797_, _13761_);
  and (_13799_, _13798_, _02863_);
  or (_13800_, _13799_, _06770_);
  or (_13801_, _13800_, _13796_);
  and (_13802_, _13801_, _13758_);
  or (_13803_, _13802_, _02853_);
  and (_13804_, _04696_, _06155_);
  or (_13805_, _13749_, _05540_);
  or (_13806_, _13805_, _13804_);
  and (_13807_, _13806_, _13803_);
  or (_13808_, _13807_, _02579_);
  nor (_13809_, _11906_, _06785_);
  or (_13810_, _13749_, _02838_);
  or (_13811_, _13810_, _13809_);
  and (_13812_, _13811_, _06791_);
  and (_13813_, _13812_, _13808_);
  nor (_13814_, _07134_, _07105_);
  not (_13815_, _13814_);
  and (_13816_, _13815_, _07097_);
  nor (_13817_, _13815_, _07097_);
  nor (_13818_, _13817_, _13816_);
  or (_13819_, _13818_, _07138_);
  not (_13820_, _07138_);
  or (_13821_, _13820_, _07094_);
  and (_13822_, _13821_, _06784_);
  and (_13823_, _13822_, _13819_);
  or (_13824_, _13823_, _02802_);
  or (_13825_, _13824_, _13813_);
  and (_13826_, _13825_, _13755_);
  or (_13827_, _13826_, _02980_);
  and (_13828_, _11921_, _04696_);
  or (_13829_, _13749_, _03887_);
  or (_13830_, _13829_, _13828_);
  and (_13831_, _13830_, _03128_);
  and (_13832_, _13831_, _13827_);
  or (_13833_, _13832_, _13752_);
  and (_13834_, _13833_, _03883_);
  or (_13835_, _13749_, _05130_);
  and (_13836_, _13754_, _02970_);
  and (_13837_, _13836_, _13835_);
  or (_13838_, _13837_, _13834_);
  and (_13839_, _13838_, _03137_);
  and (_13840_, _13769_, _03135_);
  and (_13841_, _13840_, _13835_);
  or (_13842_, _13841_, _02965_);
  or (_13843_, _13842_, _13839_);
  nor (_13844_, _11919_, _06785_);
  or (_13845_, _13749_, _05783_);
  or (_13846_, _13845_, _13844_);
  and (_13847_, _13846_, _05788_);
  and (_13848_, _13847_, _13843_);
  nor (_13849_, _11926_, _06785_);
  or (_13850_, _13849_, _13749_);
  and (_13851_, _13850_, _03123_);
  or (_13852_, _13851_, _03163_);
  or (_13853_, _13852_, _13848_);
  or (_13854_, _13766_, _03906_);
  and (_13855_, _13854_, _02498_);
  and (_13856_, _13855_, _13853_);
  and (_13857_, _13786_, _02497_);
  or (_13858_, _13857_, _02888_);
  or (_13859_, _13858_, _13856_);
  and (_13860_, _11985_, _04696_);
  or (_13861_, _13749_, _02890_);
  or (_13862_, _13861_, _13860_);
  and (_13863_, _13862_, _42668_);
  and (_13864_, _13863_, _13859_);
  or (_13865_, _13864_, _13748_);
  and (_43416_, _13865_, _43998_);
  nor (_13866_, _42668_, _06836_);
  nor (_13867_, _04696_, _06836_);
  and (_13868_, _12133_, _04696_);
  or (_13869_, _13868_, _13867_);
  and (_13870_, _13869_, _03127_);
  and (_13871_, _04696_, _05658_);
  or (_13872_, _13871_, _13867_);
  or (_13873_, _13872_, _02803_);
  nor (_13874_, _12112_, _06785_);
  or (_13875_, _13874_, _13867_);
  and (_13876_, _13875_, _02579_);
  nor (_13877_, _05333_, _06836_);
  and (_13878_, _12021_, _05333_);
  or (_13879_, _13878_, _13877_);
  or (_13880_, _13877_, _12036_);
  and (_13881_, _13880_, _13879_);
  or (_13882_, _13881_, _02870_);
  nor (_13883_, _12017_, _06785_);
  or (_13884_, _13883_, _13867_);
  or (_13885_, _13884_, _03810_);
  and (_13886_, _04696_, \oc8051_golden_model_1.ACC [3]);
  or (_13887_, _13886_, _13867_);
  and (_13888_, _13887_, _03813_);
  nor (_13889_, _03813_, _06836_);
  or (_13890_, _13889_, _02974_);
  or (_13891_, _13890_, _13888_);
  and (_13892_, _13891_, _02881_);
  and (_13893_, _13892_, _13885_);
  and (_13894_, _13879_, _02880_);
  or (_13895_, _13894_, _03069_);
  or (_13896_, _13895_, _13893_);
  and (_13897_, _04696_, _04241_);
  or (_13898_, _13897_, _13867_);
  or (_13899_, _13898_, _03336_);
  and (_13900_, _13899_, _13896_);
  or (_13901_, _13900_, _03075_);
  or (_13902_, _13887_, _03084_);
  and (_13903_, _13902_, _02877_);
  and (_13904_, _13903_, _13901_);
  and (_13905_, _12005_, _05333_);
  or (_13906_, _13905_, _13877_);
  and (_13907_, _13906_, _02876_);
  or (_13908_, _13907_, _02869_);
  or (_13909_, _13908_, _13904_);
  and (_13910_, _13909_, _13882_);
  or (_13911_, _13910_, _06247_);
  nor (_13912_, _06739_, _06572_);
  nor (_13913_, _13912_, _06740_);
  or (_13914_, _13913_, _06253_);
  and (_13915_, _13914_, _02864_);
  and (_13916_, _13915_, _13911_);
  nor (_13917_, _12054_, _06771_);
  or (_13918_, _13917_, _13877_);
  and (_13919_, _13918_, _02863_);
  or (_13920_, _13919_, _06770_);
  or (_13921_, _13920_, _13916_);
  or (_13922_, _13898_, _05535_);
  and (_13923_, _13922_, _13921_);
  or (_13924_, _13923_, _02853_);
  and (_13925_, _04696_, _06154_);
  or (_13926_, _13867_, _05540_);
  or (_13927_, _13926_, _13925_);
  and (_13928_, _13927_, _02838_);
  and (_13929_, _13928_, _13924_);
  or (_13930_, _13929_, _13876_);
  and (_13931_, _13930_, _06791_);
  nor (_13932_, _13816_, _07096_);
  nor (_13933_, _13932_, _07089_);
  and (_13934_, _13932_, _07089_);
  or (_13935_, _13934_, _13933_);
  or (_13936_, _13935_, _07138_);
  or (_13937_, _13820_, _07086_);
  and (_13938_, _13937_, _06784_);
  and (_13939_, _13938_, _13936_);
  or (_13940_, _13939_, _02802_);
  or (_13941_, _13940_, _13931_);
  and (_13942_, _13941_, _13873_);
  or (_13943_, _13942_, _02980_);
  and (_13944_, _12127_, _04696_);
  or (_13945_, _13867_, _03887_);
  or (_13946_, _13945_, _13944_);
  and (_13947_, _13946_, _03128_);
  and (_13948_, _13947_, _13943_);
  or (_13949_, _13948_, _13870_);
  and (_13950_, _13949_, _03883_);
  or (_13951_, _13867_, _05079_);
  and (_13952_, _13872_, _02970_);
  and (_13953_, _13952_, _13951_);
  or (_13954_, _13953_, _13950_);
  and (_13955_, _13954_, _03137_);
  and (_13956_, _13887_, _03135_);
  and (_13957_, _13956_, _13951_);
  or (_13958_, _13957_, _02965_);
  or (_13959_, _13958_, _13955_);
  nor (_13960_, _12125_, _06785_);
  or (_13961_, _13867_, _05783_);
  or (_13962_, _13961_, _13960_);
  and (_13963_, _13962_, _05788_);
  and (_13964_, _13963_, _13959_);
  nor (_13965_, _12132_, _06785_);
  or (_13966_, _13965_, _13867_);
  and (_13967_, _13966_, _03123_);
  or (_13968_, _13967_, _03163_);
  or (_13969_, _13968_, _13964_);
  or (_13970_, _13884_, _03906_);
  and (_13971_, _13970_, _02498_);
  and (_13972_, _13971_, _13969_);
  and (_13973_, _13906_, _02497_);
  or (_13974_, _13973_, _02888_);
  or (_13975_, _13974_, _13972_);
  and (_13976_, _12183_, _04696_);
  or (_13977_, _13867_, _02890_);
  or (_13978_, _13977_, _13976_);
  and (_13979_, _13978_, _42668_);
  and (_13980_, _13979_, _13975_);
  or (_13981_, _13980_, _13866_);
  and (_43417_, _13981_, _43998_);
  nor (_13982_, _42668_, _06931_);
  nor (_13983_, _04696_, _06931_);
  and (_13984_, _12207_, _04696_);
  or (_13985_, _13984_, _13983_);
  and (_13986_, _13985_, _03127_);
  and (_13987_, _05666_, _04696_);
  or (_13988_, _13987_, _13983_);
  or (_13989_, _13988_, _02803_);
  nor (_13990_, _12321_, _06785_);
  or (_13991_, _13990_, _13983_);
  and (_13992_, _13991_, _02579_);
  and (_13993_, _04696_, _04982_);
  or (_13994_, _13993_, _13983_);
  or (_13995_, _13994_, _05535_);
  nor (_13996_, _05333_, _06931_);
  and (_13997_, _12213_, _05333_);
  or (_13998_, _13997_, _13996_);
  and (_13999_, _13998_, _02876_);
  nor (_14000_, _12217_, _06785_);
  or (_14001_, _14000_, _13983_);
  or (_14002_, _14001_, _03810_);
  and (_14003_, _04696_, \oc8051_golden_model_1.ACC [4]);
  or (_14004_, _14003_, _13983_);
  and (_14005_, _14004_, _03813_);
  nor (_14006_, _03813_, _06931_);
  or (_14007_, _14006_, _02974_);
  or (_14008_, _14007_, _14005_);
  and (_14009_, _14008_, _02881_);
  and (_14010_, _14009_, _14002_);
  and (_14011_, _12231_, _05333_);
  or (_14012_, _14011_, _13996_);
  and (_14013_, _14012_, _02880_);
  or (_14014_, _14013_, _03069_);
  or (_14015_, _14014_, _14010_);
  or (_14016_, _13994_, _03336_);
  and (_14017_, _14016_, _14015_);
  or (_14018_, _14017_, _03075_);
  or (_14019_, _14004_, _03084_);
  and (_14020_, _14019_, _02877_);
  and (_14021_, _14020_, _14018_);
  or (_14022_, _14021_, _13999_);
  and (_14023_, _14022_, _02870_);
  or (_14024_, _13996_, _12246_);
  and (_14025_, _14024_, _02869_);
  and (_14026_, _14025_, _14012_);
  or (_14027_, _14026_, _06247_);
  or (_14028_, _14027_, _14023_);
  nor (_14029_, _06744_, _06742_);
  nor (_14030_, _14029_, _06745_);
  or (_14031_, _14030_, _06253_);
  and (_14032_, _14031_, _02864_);
  and (_14033_, _14032_, _14028_);
  nor (_14034_, _12264_, _06771_);
  or (_14035_, _14034_, _13996_);
  and (_14036_, _14035_, _02863_);
  or (_14037_, _14036_, _06770_);
  or (_14038_, _14037_, _14033_);
  and (_14039_, _14038_, _13995_);
  or (_14040_, _14039_, _02853_);
  and (_14041_, _04696_, _06159_);
  or (_14042_, _13983_, _05540_);
  or (_14043_, _14042_, _14041_);
  and (_14044_, _14043_, _02838_);
  and (_14045_, _14044_, _14040_);
  or (_14046_, _14045_, _13992_);
  and (_14047_, _14046_, _06791_);
  or (_14048_, _13820_, _07078_);
  nor (_14049_, _13932_, _07087_);
  or (_14050_, _14049_, _07088_);
  nand (_14051_, _14050_, _07127_);
  or (_14052_, _14050_, _07127_);
  and (_14053_, _14052_, _14051_);
  or (_14054_, _14053_, _07138_);
  and (_14055_, _14054_, _06784_);
  and (_14056_, _14055_, _14048_);
  or (_14057_, _14056_, _02802_);
  or (_14058_, _14057_, _14047_);
  and (_14059_, _14058_, _13989_);
  or (_14060_, _14059_, _02980_);
  and (_14061_, _12211_, _04696_);
  or (_14062_, _13983_, _03887_);
  or (_14063_, _14062_, _14061_);
  and (_14064_, _14063_, _03128_);
  and (_14065_, _14064_, _14060_);
  or (_14066_, _14065_, _13986_);
  and (_14067_, _14066_, _03883_);
  or (_14068_, _13983_, _05031_);
  and (_14069_, _13988_, _02970_);
  and (_14070_, _14069_, _14068_);
  or (_14071_, _14070_, _14067_);
  and (_14072_, _14071_, _03137_);
  and (_14073_, _14004_, _03135_);
  and (_14074_, _14073_, _14068_);
  or (_14075_, _14074_, _02965_);
  or (_14076_, _14075_, _14072_);
  nor (_14077_, _12209_, _06785_);
  or (_14078_, _13983_, _05783_);
  or (_14079_, _14078_, _14077_);
  and (_14080_, _14079_, _05788_);
  and (_14081_, _14080_, _14076_);
  nor (_14082_, _12206_, _06785_);
  or (_14083_, _14082_, _13983_);
  and (_14084_, _14083_, _03123_);
  or (_14085_, _14084_, _03163_);
  or (_14086_, _14085_, _14081_);
  or (_14087_, _14001_, _03906_);
  and (_14088_, _14087_, _02498_);
  and (_14089_, _14088_, _14086_);
  and (_14090_, _13998_, _02497_);
  or (_14091_, _14090_, _02888_);
  or (_14092_, _14091_, _14089_);
  and (_14093_, _12389_, _04696_);
  or (_14094_, _13983_, _02890_);
  or (_14095_, _14094_, _14093_);
  and (_14096_, _14095_, _42668_);
  and (_14097_, _14096_, _14092_);
  or (_14098_, _14097_, _13982_);
  and (_43418_, _14098_, _43998_);
  nor (_14099_, _42668_, _06922_);
  nor (_14100_, _04696_, _06922_);
  and (_14101_, _12411_, _04696_);
  or (_14102_, _14101_, _14100_);
  and (_14103_, _14102_, _03127_);
  and (_14104_, _05614_, _04696_);
  or (_14105_, _14104_, _14100_);
  or (_14106_, _14105_, _02803_);
  nor (_14107_, _12527_, _06785_);
  or (_14108_, _14107_, _14100_);
  and (_14109_, _14108_, _02579_);
  and (_14110_, _04696_, _04877_);
  or (_14111_, _14110_, _14100_);
  or (_14112_, _14111_, _05535_);
  nor (_14113_, _05333_, _06922_);
  and (_14114_, _12417_, _05333_);
  or (_14115_, _14114_, _14113_);
  and (_14116_, _14115_, _02876_);
  nor (_14117_, _12407_, _06785_);
  or (_14118_, _14117_, _14100_);
  or (_14119_, _14118_, _03810_);
  and (_14120_, _04696_, \oc8051_golden_model_1.ACC [5]);
  or (_14121_, _14120_, _14100_);
  and (_14122_, _14121_, _03813_);
  nor (_14123_, _03813_, _06922_);
  or (_14124_, _14123_, _02974_);
  or (_14125_, _14124_, _14122_);
  and (_14126_, _14125_, _02881_);
  and (_14127_, _14126_, _14119_);
  and (_14128_, _12435_, _05333_);
  or (_14129_, _14128_, _14113_);
  and (_14130_, _14129_, _02880_);
  or (_14131_, _14130_, _03069_);
  or (_14132_, _14131_, _14127_);
  or (_14133_, _14111_, _03336_);
  and (_14134_, _14133_, _14132_);
  or (_14135_, _14134_, _03075_);
  or (_14136_, _14121_, _03084_);
  and (_14137_, _14136_, _02877_);
  and (_14138_, _14137_, _14135_);
  or (_14139_, _14138_, _14116_);
  and (_14140_, _14139_, _02870_);
  or (_14141_, _14113_, _12450_);
  and (_14142_, _14129_, _02869_);
  and (_14143_, _14142_, _14141_);
  or (_14144_, _14143_, _06247_);
  or (_14145_, _14144_, _14140_);
  or (_14146_, _06444_, _06445_);
  not (_14147_, _14146_);
  nor (_14148_, _14147_, _06746_);
  and (_14149_, _14147_, _06746_);
  or (_14150_, _14149_, _14148_);
  or (_14151_, _14150_, _06253_);
  and (_14152_, _14151_, _02864_);
  and (_14153_, _14152_, _14145_);
  nor (_14154_, _12468_, _06771_);
  or (_14155_, _14154_, _14113_);
  and (_14156_, _14155_, _02863_);
  or (_14157_, _14156_, _06770_);
  or (_14158_, _14157_, _14153_);
  and (_14159_, _14158_, _14112_);
  or (_14160_, _14159_, _02853_);
  and (_14161_, _04696_, _06158_);
  or (_14162_, _14100_, _05540_);
  or (_14163_, _14162_, _14161_);
  and (_14164_, _14163_, _02838_);
  and (_14165_, _14164_, _14160_);
  or (_14166_, _14165_, _14109_);
  and (_14167_, _14166_, _06791_);
  or (_14168_, _13820_, _07070_);
  not (_14169_, _07116_);
  and (_14170_, _14051_, _14169_);
  nor (_14171_, _14170_, _07128_);
  and (_14172_, _14170_, _07128_);
  or (_14173_, _14172_, _14171_);
  or (_14174_, _14173_, _07138_);
  and (_14175_, _14174_, _06784_);
  and (_14176_, _14175_, _14168_);
  or (_14177_, _14176_, _02802_);
  or (_14178_, _14177_, _14167_);
  and (_14179_, _14178_, _14106_);
  or (_14180_, _14179_, _02980_);
  and (_14181_, _12415_, _04696_);
  or (_14182_, _14100_, _03887_);
  or (_14183_, _14182_, _14181_);
  and (_14184_, _14183_, _03128_);
  and (_14185_, _14184_, _14180_);
  or (_14186_, _14185_, _14103_);
  and (_14187_, _14186_, _03883_);
  or (_14188_, _14100_, _04924_);
  and (_14189_, _14105_, _02970_);
  and (_14190_, _14189_, _14188_);
  or (_14191_, _14190_, _14187_);
  and (_14192_, _14191_, _03137_);
  and (_14193_, _14121_, _03135_);
  and (_14194_, _14193_, _14188_);
  or (_14195_, _14194_, _02965_);
  or (_14196_, _14195_, _14192_);
  nor (_14197_, _12413_, _06785_);
  or (_14198_, _14100_, _05783_);
  or (_14199_, _14198_, _14197_);
  and (_14200_, _14199_, _05788_);
  and (_14201_, _14200_, _14196_);
  nor (_14202_, _12410_, _06785_);
  or (_14203_, _14202_, _14100_);
  and (_14204_, _14203_, _03123_);
  or (_14205_, _14204_, _03163_);
  or (_14206_, _14205_, _14201_);
  or (_14207_, _14118_, _03906_);
  and (_14208_, _14207_, _02498_);
  and (_14209_, _14208_, _14206_);
  and (_14210_, _14115_, _02497_);
  or (_14211_, _14210_, _02888_);
  or (_14212_, _14211_, _14209_);
  and (_14213_, _12589_, _04696_);
  or (_14214_, _14100_, _02890_);
  or (_14215_, _14214_, _14213_);
  and (_14216_, _14215_, _42668_);
  and (_14217_, _14216_, _14212_);
  or (_14218_, _14217_, _14099_);
  and (_43419_, _14218_, _43998_);
  nor (_14219_, _42668_, _07055_);
  nor (_14220_, _04696_, _07055_);
  and (_14221_, _12613_, _04696_);
  or (_14222_, _14221_, _14220_);
  and (_14223_, _14222_, _03127_);
  and (_14224_, _12729_, _04696_);
  or (_14225_, _14224_, _14220_);
  or (_14226_, _14225_, _02803_);
  nor (_14227_, _12722_, _06785_);
  or (_14228_, _14227_, _14220_);
  and (_14229_, _14228_, _02579_);
  and (_14230_, _04696_, _04770_);
  or (_14231_, _14230_, _14220_);
  or (_14232_, _14231_, _05535_);
  nor (_14233_, _05333_, _07055_);
  and (_14234_, _12616_, _05333_);
  or (_14235_, _14234_, _14233_);
  and (_14236_, _14235_, _02876_);
  nor (_14237_, _12603_, _06785_);
  or (_14238_, _14237_, _14220_);
  or (_14239_, _14238_, _03810_);
  and (_14240_, _04696_, \oc8051_golden_model_1.ACC [6]);
  or (_14241_, _14240_, _14220_);
  and (_14242_, _14241_, _03813_);
  nor (_14243_, _03813_, _07055_);
  or (_14244_, _14243_, _02974_);
  or (_14245_, _14244_, _14242_);
  and (_14246_, _14245_, _02881_);
  and (_14247_, _14246_, _14239_);
  and (_14248_, _12618_, _05333_);
  or (_14249_, _14248_, _14233_);
  and (_14250_, _14249_, _02880_);
  or (_14251_, _14250_, _03069_);
  or (_14252_, _14251_, _14247_);
  or (_14253_, _14231_, _03336_);
  and (_14254_, _14253_, _14252_);
  or (_14255_, _14254_, _03075_);
  or (_14256_, _14241_, _03084_);
  and (_14257_, _14256_, _02877_);
  and (_14258_, _14257_, _14255_);
  or (_14259_, _14258_, _14236_);
  and (_14260_, _14259_, _02870_);
  or (_14261_, _14233_, _12646_);
  and (_14262_, _14249_, _02869_);
  and (_14263_, _14262_, _14261_);
  or (_14264_, _14263_, _06247_);
  or (_14265_, _14264_, _14260_);
  nor (_14266_, _06762_, _06749_);
  nor (_14267_, _14266_, _06763_);
  or (_14268_, _14267_, _06253_);
  and (_14269_, _14268_, _02864_);
  and (_14270_, _14269_, _14265_);
  nor (_14271_, _12664_, _06771_);
  or (_14272_, _14271_, _14233_);
  and (_14273_, _14272_, _02863_);
  or (_14274_, _14273_, _06770_);
  or (_14275_, _14274_, _14270_);
  and (_14276_, _14275_, _14232_);
  or (_14277_, _14276_, _02853_);
  and (_14278_, _04696_, _05849_);
  or (_14279_, _14220_, _05540_);
  or (_14280_, _14279_, _14278_);
  and (_14281_, _14280_, _02838_);
  and (_14282_, _14281_, _14277_);
  or (_14283_, _14282_, _14229_);
  and (_14284_, _14283_, _06791_);
  or (_14285_, _13820_, _07061_);
  nor (_14286_, _14170_, _07071_);
  or (_14287_, _14286_, _07072_);
  or (_14288_, _14287_, _07125_);
  nand (_14289_, _14287_, _07125_);
  and (_14290_, _14289_, _14288_);
  or (_14291_, _14290_, _07138_);
  and (_14292_, _14291_, _06784_);
  and (_14293_, _14292_, _14285_);
  or (_14294_, _14293_, _02802_);
  or (_14295_, _14294_, _14284_);
  and (_14296_, _14295_, _14226_);
  or (_14297_, _14296_, _02980_);
  and (_14298_, _12739_, _04696_);
  or (_14299_, _14220_, _03887_);
  or (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _03128_);
  and (_14302_, _14301_, _14297_);
  or (_14303_, _14302_, _14223_);
  and (_14304_, _14303_, _03883_);
  or (_14305_, _14220_, _04819_);
  and (_14306_, _14225_, _02970_);
  and (_14307_, _14306_, _14305_);
  or (_14308_, _14307_, _14304_);
  and (_14309_, _14308_, _03137_);
  and (_14310_, _14241_, _03135_);
  and (_14311_, _14310_, _14305_);
  or (_14312_, _14311_, _02965_);
  or (_14313_, _14312_, _14309_);
  nor (_14314_, _12737_, _06785_);
  or (_14315_, _14220_, _05783_);
  or (_14316_, _14315_, _14314_);
  and (_14317_, _14316_, _05788_);
  and (_14318_, _14317_, _14313_);
  nor (_14319_, _12612_, _06785_);
  or (_14320_, _14319_, _14220_);
  and (_14321_, _14320_, _03123_);
  or (_14322_, _14321_, _03163_);
  or (_14323_, _14322_, _14318_);
  or (_14324_, _14238_, _03906_);
  and (_14325_, _14324_, _02498_);
  and (_14326_, _14325_, _14323_);
  and (_14327_, _14235_, _02497_);
  or (_14328_, _14327_, _02888_);
  or (_14329_, _14328_, _14326_);
  and (_14330_, _12794_, _04696_);
  or (_14331_, _14220_, _02890_);
  or (_14332_, _14331_, _14330_);
  and (_14333_, _14332_, _42668_);
  and (_14334_, _14333_, _14329_);
  or (_14335_, _14334_, _14219_);
  and (_43421_, _14335_, _43998_);
  nor (_14336_, _42668_, _02667_);
  nand (_14337_, _08111_, _05771_);
  nor (_14338_, _03808_, \oc8051_golden_model_1.ACC [0]);
  nor (_14339_, _14338_, _07213_);
  and (_14340_, _14339_, _10378_);
  nand (_14341_, _07614_, _07240_);
  nand (_14342_, _07942_, _09521_);
  not (_14343_, _03732_);
  nor (_14344_, _14338_, _14343_);
  or (_14345_, _08046_, _07912_);
  nor (_14346_, _04706_, _02667_);
  and (_14347_, _04706_, _03808_);
  nor (_14348_, _14347_, _14346_);
  nand (_14349_, _14348_, _06770_);
  nand (_14350_, _07804_, _07404_);
  nand (_14351_, _07737_, _03433_);
  or (_14352_, _07628_, _03808_);
  nor (_14353_, _03363_, _02886_);
  or (_14354_, _14353_, _06152_);
  or (_14355_, _07635_, _03808_);
  not (_14356_, _09427_);
  or (_14357_, _07636_, \oc8051_golden_model_1.ACC [0]);
  nand (_14358_, _07636_, \oc8051_golden_model_1.ACC [0]);
  and (_14359_, _14358_, _14357_);
  or (_14360_, _14359_, _14356_);
  and (_14361_, _14360_, _14355_);
  or (_14362_, _14361_, _03072_);
  nand (_14363_, _07481_, _03072_);
  and (_14364_, _14363_, _09426_);
  and (_14365_, _14364_, _14362_);
  or (_14366_, _14365_, _02886_);
  and (_14367_, _14366_, _03810_);
  and (_14368_, _14367_, _14354_);
  and (_14369_, _05226_, _04706_);
  nor (_14370_, _14369_, _14346_);
  nor (_14371_, _14370_, _03810_);
  or (_14372_, _14371_, _02880_);
  or (_14373_, _14372_, _14368_);
  nor (_14374_, _05325_, _02667_);
  and (_14375_, _11417_, _05325_);
  nor (_14376_, _14375_, _14374_);
  nand (_14377_, _14376_, _02880_);
  and (_14378_, _14377_, _03336_);
  and (_14379_, _14378_, _14373_);
  nor (_14380_, _14348_, _03336_);
  or (_14381_, _14380_, _07682_);
  or (_14382_, _14381_, _14379_);
  and (_14383_, _14382_, _14352_);
  or (_14384_, _14383_, _03399_);
  or (_14385_, _06152_, _03840_);
  and (_14386_, _14385_, _03084_);
  and (_14387_, _14386_, _14384_);
  nor (_14388_, _07481_, _03084_);
  or (_14389_, _14388_, _07692_);
  or (_14390_, _14389_, _14387_);
  nand (_14391_, _07692_, _06867_);
  and (_14392_, _14391_, _14390_);
  or (_14393_, _14392_, _02876_);
  or (_14394_, _14346_, _02877_);
  and (_14395_, _14394_, _02870_);
  and (_14396_, _14395_, _14393_);
  nor (_14397_, _14370_, _02870_);
  or (_14398_, _14397_, _06247_);
  or (_14399_, _14398_, _14396_);
  not (_14400_, _06708_);
  nand (_14401_, _14400_, _06247_);
  and (_14402_, _14401_, _07717_);
  and (_14403_, _14402_, _14399_);
  nor (_14404_, _07737_, _07717_);
  or (_14405_, _14404_, _03433_);
  or (_14406_, _14405_, _14403_);
  and (_14407_, _14406_, _14351_);
  or (_14408_, _14407_, _03434_);
  nand (_14409_, _07614_, _03434_);
  and (_14410_, _14409_, _03111_);
  and (_14411_, _14410_, _14408_);
  nand (_14412_, _07573_, _07405_);
  and (_14413_, _14412_, _09562_);
  or (_14414_, _14413_, _14411_);
  and (_14415_, _14414_, _14350_);
  or (_14416_, _14415_, _02583_);
  or (_14417_, _02835_, _02605_);
  and (_14418_, _14417_, _02864_);
  and (_14419_, _14418_, _14416_);
  nor (_14420_, _11448_, _07833_);
  nor (_14421_, _14420_, _14374_);
  nor (_14422_, _14421_, _02864_);
  or (_14423_, _14422_, _06770_);
  or (_14424_, _14423_, _14419_);
  and (_14425_, _14424_, _14349_);
  or (_14426_, _14425_, _02853_);
  and (_14427_, _04706_, _06152_);
  nor (_14428_, _14427_, _14346_);
  nand (_14429_, _14428_, _02853_);
  and (_14430_, _14429_, _02838_);
  and (_14431_, _14430_, _14426_);
  nor (_14432_, _11505_, _07846_);
  nor (_14433_, _14432_, _14346_);
  nor (_14434_, _14433_, _02838_);
  or (_14435_, _14434_, _06784_);
  or (_14436_, _14435_, _14431_);
  nand (_14437_, _07138_, _06784_);
  and (_14438_, _14437_, _14436_);
  and (_14439_, _14438_, _02635_);
  and (_14440_, _02835_, _02546_);
  or (_14441_, _14440_, _02802_);
  or (_14442_, _14441_, _14439_);
  and (_14443_, _04706_, _05672_);
  nor (_14444_, _14443_, _14346_);
  nand (_14445_, _14444_, _02802_);
  and (_14446_, _14445_, _07860_);
  and (_14447_, _14446_, _14442_);
  and (_14448_, _07859_, _02835_);
  or (_14449_, _14448_, _07876_);
  or (_14450_, _14449_, _14447_);
  and (_14451_, _14339_, _07880_);
  or (_14452_, _14451_, _09657_);
  and (_14453_, _14452_, _14450_);
  and (_14454_, _05940_, _02667_);
  nor (_14455_, _08046_, _14454_);
  and (_14456_, _14455_, _07879_);
  or (_14457_, _14456_, _03129_);
  or (_14458_, _14457_, _14453_);
  or (_14459_, _11522_, _07890_);
  and (_14460_, _14459_, _07897_);
  and (_14461_, _14460_, _14458_);
  and (_14462_, _07399_, _09522_);
  or (_14463_, _14462_, _02980_);
  or (_14464_, _14463_, _14461_);
  and (_14465_, _11399_, _04706_);
  nor (_14466_, _14465_, _14346_);
  nand (_14467_, _14466_, _02980_);
  and (_14468_, _14467_, _03128_);
  and (_14469_, _14468_, _14464_);
  and (_14470_, _02848_, _02969_);
  and (_14471_, _14346_, _03127_);
  or (_14472_, _14471_, _14470_);
  or (_14473_, _14472_, _14469_);
  and (_14474_, _02854_, _02969_);
  nor (_14475_, _03521_, _14474_);
  and (_14476_, _02947_, _02969_);
  nor (_14477_, _14476_, _03515_);
  and (_14478_, _14477_, _14475_);
  and (_14479_, _14478_, _07213_);
  or (_14480_, _14479_, _07907_);
  and (_14481_, _14480_, _14473_);
  not (_14482_, _07213_);
  nor (_14483_, _14478_, _14482_);
  or (_14484_, _14483_, _07911_);
  or (_14485_, _14484_, _14481_);
  and (_14486_, _14485_, _14345_);
  or (_14487_, _14486_, _03138_);
  or (_14488_, _11521_, _07396_);
  and (_14489_, _14488_, _07395_);
  and (_14490_, _14489_, _14487_);
  and (_14491_, _08132_, _07394_);
  or (_14492_, _14491_, _14490_);
  and (_14493_, _14492_, _03883_);
  nor (_14494_, _14444_, _14369_);
  and (_14495_, _14494_, _02970_);
  or (_14496_, _14495_, _07925_);
  or (_14497_, _14496_, _14493_);
  nor (_14498_, _14338_, _03732_);
  or (_14499_, _14498_, _07926_);
  and (_14500_, _14499_, _14497_);
  or (_14501_, _14500_, _14344_);
  and (_14502_, _14501_, _07931_);
  nor (_14503_, _14338_, _07931_);
  or (_14504_, _14503_, _07935_);
  or (_14505_, _14504_, _14502_);
  nand (_14506_, _14454_, _07935_);
  and (_14507_, _14506_, _03122_);
  and (_14508_, _14507_, _14505_);
  nand (_14509_, _11520_, _07945_);
  and (_14510_, _14509_, _07944_);
  or (_14511_, _14510_, _14508_);
  and (_14512_, _14511_, _14342_);
  or (_14513_, _14512_, _02965_);
  nor (_14514_, _11396_, _07846_);
  nor (_14515_, _14514_, _14346_);
  nand (_14516_, _14515_, _02965_);
  and (_14517_, _14516_, _07322_);
  and (_14518_, _14517_, _14513_);
  nor (_14519_, _07737_, _07322_);
  or (_14520_, _14519_, _07240_);
  or (_14521_, _14520_, _14518_);
  and (_14522_, _14521_, _14341_);
  or (_14523_, _14522_, _03133_);
  nand (_14524_, _07573_, _03133_);
  and (_14525_, _14524_, _07993_);
  and (_14526_, _14525_, _14523_);
  nor (_14527_, _07993_, _07804_);
  or (_14528_, _14527_, _07991_);
  or (_14529_, _14528_, _14526_);
  nand (_14530_, _07991_, _07293_);
  and (_14531_, _14530_, _07238_);
  and (_14532_, _14531_, _14529_);
  or (_14533_, _14532_, _14340_);
  and (_14534_, _14533_, _08024_);
  and (_14535_, _14455_, _07188_);
  or (_14536_, _14535_, _02894_);
  or (_14537_, _14536_, _14534_);
  nand (_14538_, _09507_, _02894_);
  and (_14539_, _14538_, _08113_);
  and (_14540_, _14539_, _14537_);
  and (_14541_, _08065_, _09522_);
  or (_14542_, _14541_, _08111_);
  or (_14543_, _14542_, _14540_);
  and (_14544_, _14543_, _14337_);
  or (_14545_, _14544_, _03163_);
  nand (_14546_, _14370_, _03163_);
  and (_14547_, _14546_, _08155_);
  and (_14548_, _14547_, _14545_);
  nor (_14549_, _08159_, _02667_);
  nor (_14550_, _14549_, _09948_);
  or (_14551_, _14550_, _14548_);
  nand (_14552_, _08159_, _02551_);
  and (_14553_, _14552_, _02498_);
  and (_14554_, _14553_, _14551_);
  and (_14555_, _14346_, _02497_);
  or (_14556_, _14555_, _02888_);
  or (_14557_, _14556_, _14554_);
  nand (_14558_, _14370_, _02888_);
  and (_14559_, _14558_, _08177_);
  and (_14560_, _14559_, _14557_);
  and (_14561_, _08176_, _02667_);
  or (_14562_, _14561_, _08183_);
  or (_14563_, _14562_, _14560_);
  nand (_14564_, _08183_, _02551_);
  and (_14565_, _14564_, _42668_);
  and (_14566_, _14565_, _14563_);
  or (_14567_, _14566_, _14336_);
  and (_43422_, _14567_, _43998_);
  nor (_14568_, _42668_, _02551_);
  nand (_14569_, _08111_, _02667_);
  nor (_14570_, _08046_, _08045_);
  nor (_14571_, _14570_, _08047_);
  or (_14572_, _14571_, _08024_);
  nand (_14573_, _07942_, _08130_);
  nand (_14574_, _07925_, _07211_);
  nor (_14575_, _04706_, _02551_);
  and (_14576_, _04706_, _04000_);
  nor (_14577_, _14576_, _14575_);
  nand (_14578_, _14577_, _06770_);
  not (_14579_, _07578_);
  and (_14580_, _14579_, _02835_);
  nor (_14581_, _14580_, _07577_);
  and (_14582_, _14581_, _08131_);
  nor (_14583_, _14581_, _08131_);
  nor (_14584_, _14583_, _14582_);
  nand (_14585_, _14584_, _07404_);
  or (_14586_, _07635_, _04000_);
  nor (_14587_, _07636_, \oc8051_golden_model_1.ACC [1]);
  and (_14588_, _07636_, \oc8051_golden_model_1.ACC [1]);
  or (_14589_, _14588_, _14587_);
  nand (_14590_, _14589_, _09427_);
  and (_14591_, _14590_, _14586_);
  or (_14592_, _14591_, _03072_);
  nand (_14593_, _07467_, _03072_);
  and (_14594_, _14593_, _09426_);
  and (_14595_, _14594_, _14592_);
  or (_14596_, _14595_, _02886_);
  or (_14597_, _14353_, _06151_);
  and (_14598_, _14597_, _14596_);
  and (_14599_, _14598_, _03810_);
  nor (_14600_, _04706_, \oc8051_golden_model_1.ACC [1]);
  and (_14601_, _11606_, _04706_);
  nor (_14602_, _14601_, _14600_);
  and (_14603_, _14602_, _02974_);
  or (_14604_, _14603_, _07649_);
  or (_14605_, _14604_, _14599_);
  nor (_14606_, _07656_, \oc8051_golden_model_1.PSW [6]);
  nor (_14607_, _14606_, \oc8051_golden_model_1.ACC [1]);
  and (_14608_, _14606_, \oc8051_golden_model_1.ACC [1]);
  nor (_14609_, _14608_, _14607_);
  nand (_14610_, _14609_, _07649_);
  and (_14611_, _14610_, _03076_);
  and (_14612_, _14611_, _14605_);
  nor (_14613_, _05325_, _02551_);
  and (_14614_, _11592_, _05325_);
  nor (_14615_, _14614_, _14613_);
  nor (_14616_, _14615_, _02881_);
  nor (_14617_, _14577_, _03336_);
  or (_14618_, _14617_, _07682_);
  or (_14619_, _14618_, _14616_);
  or (_14620_, _14619_, _14612_);
  or (_14621_, _07628_, _04000_);
  and (_14622_, _14621_, _14620_);
  or (_14623_, _14622_, _03399_);
  or (_14624_, _06151_, _03840_);
  and (_14625_, _14624_, _03084_);
  and (_14626_, _14625_, _14623_);
  nor (_14627_, _07467_, _03084_);
  or (_14628_, _14627_, _07692_);
  or (_14629_, _14628_, _14626_);
  nand (_14630_, _07692_, _06861_);
  and (_14631_, _14630_, _14629_);
  or (_14632_, _14631_, _02876_);
  and (_14633_, _11595_, _05325_);
  nor (_14634_, _14633_, _14613_);
  nand (_14635_, _14634_, _02876_);
  and (_14636_, _14635_, _02870_);
  and (_14637_, _14636_, _14632_);
  and (_14638_, _14614_, _11591_);
  nor (_14639_, _14638_, _14613_);
  nor (_14640_, _14639_, _02870_);
  or (_14641_, _14640_, _06247_);
  or (_14642_, _14641_, _14637_);
  and (_14643_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_14644_, _14643_, _07100_);
  nor (_14645_, _14644_, _06709_);
  or (_14646_, _14645_, _06253_);
  and (_14647_, _14646_, _07718_);
  and (_14648_, _14647_, _14642_);
  not (_14649_, _09557_);
  and (_14650_, _14579_, _03808_);
  nor (_14651_, _14650_, _07577_);
  and (_14652_, _14651_, _07212_);
  nor (_14653_, _14651_, _07212_);
  or (_14654_, _14653_, _14652_);
  or (_14655_, _14654_, _03434_);
  and (_14656_, _14655_, _14649_);
  or (_14657_, _14656_, _14648_);
  and (_14658_, _14579_, _06152_);
  nor (_14659_, _14658_, _07577_);
  and (_14660_, _14659_, _08045_);
  nor (_14661_, _14659_, _08045_);
  or (_14662_, _14661_, _14660_);
  or (_14663_, _14662_, _07626_);
  and (_14664_, _14663_, _03111_);
  and (_14665_, _14664_, _14657_);
  nand (_14666_, _07583_, _07405_);
  and (_14667_, _14666_, _09562_);
  or (_14668_, _14667_, _14665_);
  and (_14669_, _14668_, _14585_);
  or (_14670_, _14669_, _02583_);
  nand (_14671_, _03665_, _02583_);
  and (_14672_, _14671_, _02864_);
  and (_14674_, _14672_, _14670_);
  nor (_14675_, _11638_, _07833_);
  nor (_14676_, _14675_, _14613_);
  nor (_14677_, _14676_, _02864_);
  or (_14678_, _14677_, _06770_);
  or (_14679_, _14678_, _14674_);
  and (_14680_, _14679_, _14578_);
  or (_14681_, _14680_, _02853_);
  and (_14682_, _04706_, _06151_);
  nor (_14683_, _14682_, _14575_);
  nand (_14685_, _14683_, _02853_);
  and (_14686_, _14685_, _02838_);
  and (_14687_, _14686_, _14681_);
  nor (_14688_, _11695_, _07846_);
  nor (_14689_, _14688_, _14575_);
  nor (_14690_, _14689_, _02838_);
  or (_14691_, _14690_, _06784_);
  or (_14692_, _14691_, _14687_);
  nand (_14693_, _07048_, _06784_);
  and (_14694_, _14693_, _14692_);
  and (_14696_, _14694_, _02635_);
  nor (_14697_, _03665_, _02635_);
  or (_14698_, _14697_, _02802_);
  or (_14699_, _14698_, _14696_);
  and (_14700_, _04706_, _03698_);
  nor (_14701_, _14700_, _14600_);
  or (_14702_, _14701_, _02803_);
  and (_14703_, _14702_, _07860_);
  and (_14704_, _14703_, _14699_);
  nor (_14705_, _07860_, _03665_);
  or (_14707_, _14705_, _07869_);
  or (_14708_, _14707_, _14704_);
  or (_14709_, _07870_, _07212_);
  nor (_14710_, _03735_, _03503_);
  and (_14711_, _14710_, _14709_);
  and (_14712_, _14711_, _14708_);
  and (_14713_, _02854_, _02508_);
  not (_14714_, _14710_);
  and (_14715_, _14714_, _07212_);
  or (_14716_, _14715_, _14713_);
  or (_14718_, _14716_, _14712_);
  not (_14719_, _14713_);
  or (_14720_, _14719_, _07212_);
  and (_14721_, _14720_, _07880_);
  and (_14722_, _14721_, _14718_);
  and (_14723_, _08045_, _07879_);
  or (_14724_, _14723_, _03129_);
  or (_14725_, _14724_, _14722_);
  or (_14726_, _11715_, _07890_);
  and (_14727_, _14726_, _14725_);
  or (_14729_, _14727_, _07399_);
  or (_14730_, _07897_, _08131_);
  and (_14731_, _14730_, _14729_);
  or (_14732_, _14731_, _02980_);
  and (_14733_, _11710_, _04706_);
  nor (_14734_, _14733_, _14575_);
  nand (_14735_, _14734_, _02980_);
  and (_14736_, _14735_, _03128_);
  and (_14737_, _14736_, _14732_);
  and (_14738_, _14575_, _03127_);
  or (_14740_, _14738_, _09681_);
  or (_14741_, _14740_, _14737_);
  or (_14742_, _08043_, _07912_);
  or (_14743_, _07907_, _07210_);
  and (_14744_, _14743_, _14742_);
  and (_14745_, _14744_, _14741_);
  or (_14746_, _14745_, _03138_);
  or (_14747_, _11587_, _07396_);
  and (_14748_, _14747_, _07395_);
  and (_14749_, _14748_, _14746_);
  and (_14751_, _08129_, _07394_);
  or (_14752_, _14751_, _14749_);
  and (_14753_, _14752_, _03883_);
  and (_14754_, _11709_, _04706_);
  nor (_14755_, _14754_, _14575_);
  nor (_14756_, _14755_, _03883_);
  or (_14757_, _14756_, _07925_);
  or (_14758_, _14757_, _14753_);
  and (_14759_, _14758_, _14574_);
  and (_14760_, _04009_, _02964_);
  nor (_14762_, _14760_, _03732_);
  not (_14763_, _14762_);
  or (_14764_, _14763_, _14759_);
  nand (_14765_, _14763_, _07211_);
  and (_14766_, _14765_, _03529_);
  and (_14767_, _14766_, _14764_);
  nor (_14768_, _07211_, _03529_);
  or (_14769_, _14768_, _07935_);
  or (_14770_, _14769_, _14767_);
  nand (_14771_, _08044_, _07935_);
  and (_14773_, _14771_, _03122_);
  and (_14774_, _14773_, _14770_);
  nand (_14775_, _11714_, _07945_);
  and (_14776_, _14775_, _07944_);
  or (_14777_, _14776_, _14774_);
  and (_14778_, _14777_, _14573_);
  or (_14779_, _14778_, _02965_);
  nor (_14780_, _11708_, _07846_);
  or (_14781_, _14780_, _14575_);
  or (_14782_, _14781_, _05783_);
  and (_14784_, _14782_, _07322_);
  and (_14785_, _14784_, _14779_);
  and (_14786_, _07376_, _07372_);
  nor (_14787_, _14786_, _07377_);
  and (_14788_, _14787_, _10349_);
  or (_14789_, _14788_, _07240_);
  or (_14790_, _14789_, _14785_);
  and (_14791_, _07297_, _07292_);
  nor (_14792_, _14791_, _07298_);
  or (_14793_, _14792_, _07241_);
  and (_14795_, _14793_, _03134_);
  and (_14796_, _14795_, _14790_);
  and (_14797_, _07972_, _07970_);
  nor (_14798_, _14797_, _07973_);
  and (_14799_, _14798_, _03133_);
  or (_14800_, _14799_, _07962_);
  or (_14801_, _14800_, _14796_);
  and (_14802_, _08000_, _07798_);
  nor (_14803_, _14802_, _08001_);
  or (_14804_, _14803_, _07993_);
  and (_14806_, _14804_, _14801_);
  or (_14807_, _14806_, _07991_);
  nand (_14808_, _07991_, _02667_);
  and (_14809_, _14808_, _07238_);
  and (_14810_, _14809_, _14807_);
  nor (_14811_, _07213_, _07212_);
  nor (_14812_, _14811_, _07214_);
  and (_14813_, _14812_, _10378_);
  or (_14814_, _14813_, _07188_);
  or (_14815_, _14814_, _14810_);
  and (_14817_, _14815_, _14572_);
  or (_14818_, _14817_, _02894_);
  and (_14819_, _08090_, _07576_);
  nor (_14820_, _14819_, _08091_);
  or (_14821_, _14820_, _02896_);
  and (_14822_, _14821_, _08113_);
  and (_14823_, _14822_, _14818_);
  nor (_14824_, _08132_, _08131_);
  nor (_14825_, _14824_, _08133_);
  and (_14826_, _14825_, _08065_);
  or (_14828_, _14826_, _08111_);
  or (_14829_, _14828_, _14823_);
  and (_14830_, _14829_, _14569_);
  or (_14831_, _14830_, _03163_);
  or (_14832_, _14602_, _03906_);
  and (_14833_, _14832_, _08155_);
  and (_14834_, _14833_, _14831_);
  nor (_14835_, _08184_, _08160_);
  not (_14836_, _14835_);
  nor (_14837_, _14836_, _08159_);
  nor (_14839_, _14837_, _09948_);
  or (_14840_, _14839_, _14834_);
  nand (_14841_, _08159_, _06964_);
  and (_14842_, _14841_, _02498_);
  and (_14843_, _14842_, _14840_);
  nor (_14844_, _14634_, _02498_);
  or (_14845_, _14844_, _02888_);
  or (_14846_, _14845_, _14843_);
  nor (_14847_, _14601_, _14575_);
  nand (_14848_, _14847_, _02888_);
  and (_14849_, _14848_, _08177_);
  and (_14850_, _14849_, _14846_);
  and (_14851_, _14835_, _08176_);
  or (_14852_, _14851_, _08183_);
  or (_14853_, _14852_, _14850_);
  nand (_14854_, _08183_, _06964_);
  and (_14855_, _14854_, _42668_);
  and (_14856_, _14855_, _14853_);
  or (_14857_, _14856_, _14568_);
  and (_43423_, _14857_, _43998_);
  nor (_14859_, _42668_, _06964_);
  nand (_14860_, _08111_, _02551_);
  nand (_14861_, _07942_, _08127_);
  not (_14862_, _07206_);
  or (_14863_, _03309_, _02531_);
  not (_14864_, _14863_);
  nor (_14865_, _14864_, _03738_);
  nor (_14866_, _14865_, _14862_);
  nor (_14867_, _04706_, _06964_);
  and (_14868_, _14867_, _03127_);
  and (_14870_, _04706_, _04435_);
  nor (_14871_, _14870_, _14867_);
  nand (_14872_, _14871_, _06770_);
  or (_14873_, _07628_, _04435_);
  and (_14874_, _07636_, _06964_);
  or (_14875_, _07636_, _06964_);
  nand (_14876_, _14875_, _09427_);
  or (_14877_, _14876_, _14874_);
  or (_14878_, _07635_, _04435_);
  and (_14879_, _14878_, _14877_);
  or (_14881_, _14879_, _03072_);
  nand (_14882_, _07453_, _03072_);
  and (_14883_, _14882_, _09426_);
  and (_14884_, _14883_, _14881_);
  or (_14885_, _14884_, _02886_);
  or (_14886_, _14353_, _06155_);
  and (_14887_, _14886_, _14885_);
  and (_14888_, _14887_, _03810_);
  nor (_14889_, _11801_, _07846_);
  nor (_14890_, _14889_, _14867_);
  nor (_14892_, _14890_, _03810_);
  or (_14893_, _14892_, _07649_);
  or (_14894_, _14893_, _14888_);
  nand (_14895_, _14606_, \oc8051_golden_model_1.ACC [2]);
  and (_14896_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_14897_, _14896_, _07655_);
  or (_14898_, _14897_, _14606_);
  and (_14899_, _14898_, _14895_);
  nand (_14900_, _14899_, _07649_);
  and (_14901_, _14900_, _03076_);
  and (_14903_, _14901_, _14894_);
  nor (_14904_, _05325_, _06964_);
  and (_14905_, _11815_, _05325_);
  nor (_14906_, _14905_, _14904_);
  nor (_14907_, _14906_, _02881_);
  nor (_14908_, _14871_, _03336_);
  or (_14909_, _14908_, _07682_);
  or (_14910_, _14909_, _14907_);
  or (_14911_, _14910_, _14903_);
  and (_14912_, _14911_, _14873_);
  or (_14914_, _14912_, _03399_);
  or (_14915_, _06155_, _03840_);
  and (_14916_, _14915_, _03084_);
  and (_14917_, _14916_, _14914_);
  nor (_14918_, _07453_, _03084_);
  or (_14919_, _14918_, _07692_);
  or (_14920_, _14919_, _14917_);
  nand (_14921_, _07692_, _06806_);
  and (_14922_, _14921_, _14920_);
  or (_14923_, _14922_, _02876_);
  and (_14925_, _11797_, _05325_);
  nor (_14926_, _14925_, _14904_);
  nand (_14927_, _14926_, _02876_);
  and (_14928_, _14927_, _02870_);
  and (_14929_, _14928_, _14923_);
  and (_14930_, _14905_, _11830_);
  nor (_14931_, _14930_, _14904_);
  nor (_14932_, _14931_, _02870_);
  or (_14933_, _14932_, _06247_);
  or (_14934_, _14933_, _14929_);
  nor (_14935_, _06711_, _06709_);
  nor (_14936_, _14935_, _06712_);
  or (_14937_, _14936_, _06253_);
  and (_14938_, _14937_, _14934_);
  or (_14939_, _14938_, _10106_);
  nor (_14940_, _04000_, _02551_);
  and (_14941_, _03808_, _02667_);
  nor (_14942_, _14941_, _07212_);
  nor (_14943_, _14942_, _14940_);
  nor (_14944_, _14943_, _07208_);
  and (_14947_, _14943_, _07208_);
  nor (_14948_, _14947_, _14944_);
  nor (_14949_, _14339_, _07212_);
  not (_14950_, _14949_);
  or (_14951_, _14950_, _14948_);
  and (_14952_, _14951_, \oc8051_golden_model_1.PSW [7]);
  nor (_14953_, _14948_, \oc8051_golden_model_1.PSW [7]);
  or (_14954_, _14953_, _14952_);
  nand (_14955_, _14950_, _14948_);
  and (_14956_, _14955_, _14954_);
  nor (_14958_, _14956_, _03434_);
  or (_14959_, _14958_, _09557_);
  and (_14960_, _14959_, _14939_);
  and (_14961_, _05895_, \oc8051_golden_model_1.ACC [1]);
  and (_14962_, _06152_, _02667_);
  nor (_14963_, _14962_, _08045_);
  nor (_14964_, _14963_, _14961_);
  nor (_14965_, _08041_, _14964_);
  and (_14966_, _08041_, _14964_);
  nor (_14967_, _14966_, _14965_);
  nor (_14969_, _14455_, _08045_);
  and (_14970_, _14969_, \oc8051_golden_model_1.PSW [7]);
  not (_14971_, _14970_);
  nor (_14972_, _14971_, _14967_);
  and (_14973_, _14971_, _14967_);
  nor (_14974_, _14973_, _14972_);
  nor (_14975_, _14974_, _07626_);
  or (_14976_, _14975_, _03106_);
  or (_14977_, _14976_, _14960_);
  nor (_14978_, _09505_, _07574_);
  or (_14980_, _14978_, _07575_);
  and (_14981_, _08087_, _14980_);
  nor (_14982_, _08087_, _14980_);
  nor (_14983_, _14982_, _14981_);
  and (_14984_, _09508_, \oc8051_golden_model_1.PSW [7]);
  not (_14985_, _14984_);
  nor (_14986_, _14985_, _14983_);
  and (_14987_, _14985_, _14983_);
  nor (_14988_, _14987_, _14986_);
  nand (_14989_, _14988_, _03106_);
  and (_14991_, _14989_, _07405_);
  and (_14992_, _14991_, _14977_);
  and (_14993_, _02835_, _02667_);
  nor (_14994_, _14993_, _08131_);
  nor (_14995_, _14994_, _10229_);
  not (_14996_, _08128_);
  nor (_14997_, _14996_, _14995_);
  and (_14998_, _14996_, _14995_);
  nor (_14999_, _14998_, _14997_);
  and (_15000_, _09523_, \oc8051_golden_model_1.PSW [7]);
  and (_15002_, _15000_, _14999_);
  nor (_15003_, _15000_, _14999_);
  or (_15004_, _15003_, _15002_);
  nor (_15005_, _15004_, _07405_);
  or (_15006_, _15005_, _02583_);
  or (_15007_, _15006_, _14992_);
  nand (_15008_, _03256_, _02583_);
  and (_15009_, _15008_, _02864_);
  and (_15010_, _15009_, _15007_);
  nor (_15011_, _11848_, _07833_);
  nor (_15013_, _15011_, _14904_);
  nor (_15014_, _15013_, _02864_);
  or (_15015_, _15014_, _06770_);
  or (_15016_, _15015_, _15010_);
  and (_15017_, _15016_, _14872_);
  or (_15018_, _15017_, _02853_);
  and (_15019_, _04706_, _06155_);
  nor (_15020_, _15019_, _14867_);
  nand (_15021_, _15020_, _02853_);
  and (_15022_, _15021_, _02838_);
  and (_15024_, _15022_, _15018_);
  nor (_15025_, _11906_, _07846_);
  nor (_15026_, _15025_, _14867_);
  nor (_15027_, _15026_, _02838_);
  or (_15028_, _15027_, _06784_);
  or (_15029_, _15028_, _15024_);
  or (_15030_, _06984_, _06791_);
  and (_15031_, _15030_, _15029_);
  and (_15032_, _15031_, _02635_);
  nor (_15033_, _03256_, _02635_);
  or (_15035_, _15033_, _02802_);
  or (_15036_, _15035_, _15032_);
  and (_15037_, _04706_, _05701_);
  nor (_15038_, _15037_, _14867_);
  nand (_15039_, _15038_, _02802_);
  and (_15040_, _15039_, _07860_);
  and (_15041_, _15040_, _15036_);
  nor (_15042_, _07860_, _03256_);
  or (_15043_, _15042_, _07869_);
  or (_15044_, _15043_, _15041_);
  or (_15046_, _07870_, _07208_);
  and (_15047_, _15046_, _14710_);
  and (_15048_, _15047_, _15044_);
  and (_15049_, _14714_, _07208_);
  or (_15050_, _15049_, _14713_);
  or (_15051_, _15050_, _15048_);
  or (_15052_, _14719_, _07208_);
  and (_15053_, _15052_, _07880_);
  and (_15054_, _15053_, _15051_);
  and (_15055_, _08041_, _07879_);
  or (_15057_, _15055_, _03129_);
  or (_15058_, _15057_, _15054_);
  or (_15059_, _11927_, _07890_);
  and (_15060_, _15059_, _07897_);
  and (_15061_, _15060_, _15058_);
  nor (_15062_, _07897_, _08128_);
  or (_15063_, _15062_, _02980_);
  or (_15064_, _15063_, _15061_);
  and (_15065_, _11921_, _04706_);
  nor (_15066_, _15065_, _14867_);
  nand (_15068_, _15066_, _02980_);
  and (_15069_, _15068_, _03128_);
  and (_15070_, _15069_, _15064_);
  or (_15071_, _15070_, _14868_);
  and (_15072_, _15071_, _14865_);
  nor (_15073_, _15072_, _14866_);
  nor (_15074_, _15073_, _14474_);
  and (_15075_, _07206_, _14474_);
  or (_15076_, _15075_, _15074_);
  and (_15077_, _15076_, _07912_);
  and (_15079_, _08039_, _07911_);
  or (_15080_, _15079_, _03138_);
  or (_15081_, _15080_, _15077_);
  or (_15082_, _11925_, _07396_);
  and (_15083_, _15082_, _07395_);
  and (_15084_, _15083_, _15081_);
  and (_15085_, _08126_, _07394_);
  or (_15086_, _15085_, _15084_);
  and (_15087_, _15086_, _03883_);
  or (_15088_, _15038_, _11926_);
  nor (_15090_, _15088_, _03883_);
  or (_15091_, _15090_, _07925_);
  or (_15092_, _15091_, _15087_);
  nand (_15093_, _07925_, _07207_);
  and (_15094_, _15093_, _14343_);
  and (_15095_, _15094_, _15092_);
  nor (_15096_, _07207_, _14343_);
  or (_15097_, _15096_, _15095_);
  and (_15098_, _15097_, _07931_);
  nor (_15099_, _07207_, _07931_);
  or (_15101_, _15099_, _07935_);
  or (_15102_, _15101_, _15098_);
  nand (_15103_, _08040_, _07935_);
  and (_15104_, _15103_, _03122_);
  and (_15105_, _15104_, _15102_);
  nand (_15106_, _11926_, _07945_);
  and (_15107_, _15106_, _07944_);
  or (_15108_, _15107_, _15105_);
  and (_15109_, _15108_, _14861_);
  or (_15110_, _15109_, _02965_);
  nor (_15112_, _11919_, _07846_);
  nor (_15113_, _15112_, _14867_);
  nand (_15114_, _15113_, _02965_);
  and (_15115_, _15114_, _07322_);
  and (_15116_, _15115_, _15110_);
  and (_15117_, _07378_, _07365_);
  nor (_15118_, _15117_, _07379_);
  and (_15119_, _15118_, _10349_);
  or (_15120_, _15119_, _07240_);
  or (_15121_, _15120_, _15116_);
  and (_15123_, _07299_, _07285_);
  nor (_15124_, _15123_, _07300_);
  or (_15125_, _15124_, _07241_);
  and (_15126_, _15125_, _03134_);
  and (_15127_, _15126_, _15121_);
  and (_15128_, _07974_, _07556_);
  nor (_15129_, _15128_, _07975_);
  or (_15130_, _15129_, _07962_);
  and (_15131_, _15130_, _10365_);
  or (_15132_, _15131_, _15127_);
  and (_15134_, _08002_, _07791_);
  nor (_15135_, _15134_, _08003_);
  or (_15136_, _15135_, _07993_);
  and (_15137_, _15136_, _15132_);
  or (_15138_, _15137_, _07991_);
  nand (_15139_, _07991_, _02551_);
  and (_15140_, _15139_, _07238_);
  and (_15141_, _15140_, _15138_);
  and (_15142_, _07215_, _07209_);
  nor (_15143_, _15142_, _07216_);
  and (_15145_, _15143_, _10378_);
  or (_15146_, _15145_, _07188_);
  or (_15147_, _15146_, _15141_);
  and (_15148_, _08048_, _08042_);
  nor (_15149_, _15148_, _08049_);
  or (_15150_, _15149_, _08024_);
  and (_15151_, _15150_, _15147_);
  or (_15152_, _15151_, _02894_);
  and (_15153_, _08092_, _08087_);
  nor (_15154_, _15153_, _08093_);
  or (_15156_, _15154_, _02896_);
  and (_15157_, _15156_, _08113_);
  and (_15158_, _15157_, _15152_);
  and (_15159_, _08134_, _08128_);
  nor (_15160_, _15159_, _08135_);
  and (_15161_, _15160_, _08065_);
  or (_15162_, _15161_, _08111_);
  or (_15163_, _15162_, _15158_);
  and (_15164_, _15163_, _14860_);
  or (_15165_, _15164_, _03163_);
  nand (_15167_, _14890_, _03163_);
  and (_15168_, _15167_, _08155_);
  and (_15169_, _15168_, _15165_);
  and (_15170_, _07655_, _02667_);
  nor (_15171_, _08160_, _06964_);
  or (_15172_, _15171_, _15170_);
  and (_15173_, _15172_, _08154_);
  or (_15174_, _15173_, _08159_);
  or (_15175_, _15174_, _15169_);
  nand (_15176_, _08159_, _02564_);
  and (_15178_, _15176_, _02498_);
  and (_15179_, _15178_, _15175_);
  nor (_15180_, _14926_, _02498_);
  or (_15181_, _15180_, _02888_);
  or (_15182_, _15181_, _15179_);
  and (_15183_, _11985_, _04706_);
  nor (_15184_, _15183_, _14867_);
  nand (_15185_, _15184_, _02888_);
  and (_15186_, _15185_, _08177_);
  and (_15187_, _15186_, _15182_);
  and (_15189_, _08184_, \oc8051_golden_model_1.ACC [2]);
  nor (_15190_, _08184_, \oc8051_golden_model_1.ACC [2]);
  nor (_15191_, _15190_, _15189_);
  nor (_15192_, _15191_, _08183_);
  nor (_15193_, _15192_, _09044_);
  or (_15194_, _15193_, _15187_);
  nand (_15195_, _08183_, _02564_);
  and (_15196_, _15195_, _42668_);
  and (_15197_, _15196_, _15194_);
  or (_15198_, _15197_, _14859_);
  and (_43424_, _15198_, _43998_);
  nor (_15200_, _42668_, _02564_);
  nor (_15201_, _07202_, _07204_);
  nor (_15202_, _15201_, _07217_);
  and (_15203_, _15201_, _07217_);
  nor (_15204_, _15203_, _15202_);
  nand (_15205_, _15204_, _10378_);
  or (_15206_, _14760_, _03535_);
  not (_15207_, _03323_);
  and (_15208_, _02947_, _02964_);
  nor (_15210_, _15208_, _03308_);
  and (_15211_, _15210_, _15207_);
  not (_15212_, _15211_);
  nand (_15213_, _15212_, _07202_);
  nor (_15214_, _04706_, _02564_);
  and (_15215_, _12127_, _04706_);
  nor (_15216_, _15215_, _15214_);
  nand (_15217_, _15216_, _02980_);
  and (_15218_, _04706_, _04241_);
  nor (_15219_, _15218_, _15214_);
  nand (_15221_, _15219_, _06770_);
  not (_15222_, _14969_);
  or (_15223_, _15222_, _14967_);
  and (_15224_, _15223_, \oc8051_golden_model_1.PSW [7]);
  and (_15225_, _06031_, \oc8051_golden_model_1.ACC [2]);
  nor (_15226_, _14965_, _15225_);
  nor (_15227_, _08037_, _08035_);
  nor (_15228_, _15227_, _15226_);
  and (_15229_, _15227_, _15226_);
  nor (_15230_, _15229_, _15228_);
  and (_15232_, _15230_, \oc8051_golden_model_1.PSW [7]);
  nor (_15233_, _15230_, \oc8051_golden_model_1.PSW [7]);
  nor (_15234_, _15233_, _15232_);
  and (_15235_, _15234_, _15224_);
  nor (_15236_, _15234_, _15224_);
  or (_15237_, _15236_, _15235_);
  nor (_15238_, _15237_, _07626_);
  nor (_15239_, _05325_, _02564_);
  and (_15240_, _12021_, _05325_);
  and (_15241_, _15240_, _12036_);
  nor (_15243_, _15241_, _15239_);
  nor (_15244_, _15243_, _02870_);
  or (_15245_, _07628_, _04241_);
  or (_15246_, _14353_, _06154_);
  nor (_15247_, _07442_, _03387_);
  or (_15248_, _07635_, _04241_);
  and (_15249_, _07636_, _02564_);
  or (_15250_, _07636_, _02564_);
  nand (_15251_, _15250_, _09427_);
  or (_15252_, _15251_, _15249_);
  and (_15254_, _15252_, _03387_);
  and (_15255_, _15254_, _15248_);
  or (_15256_, _15255_, _15247_);
  and (_15257_, _15256_, _09426_);
  or (_15258_, _15257_, _02886_);
  and (_15259_, _15258_, _03810_);
  and (_15260_, _15259_, _15246_);
  nor (_15261_, _12017_, _07846_);
  nor (_15262_, _15261_, _15214_);
  nor (_15263_, _15262_, _03810_);
  or (_15265_, _15263_, _07649_);
  or (_15266_, _15265_, _15260_);
  not (_15267_, \oc8051_golden_model_1.PSW [6]);
  nor (_15268_, _07655_, _15267_);
  nor (_15269_, _15268_, \oc8051_golden_model_1.ACC [3]);
  nor (_15270_, _15269_, _07656_);
  not (_15271_, _15270_);
  nand (_15272_, _15271_, _07649_);
  and (_15273_, _15272_, _15266_);
  or (_15274_, _15273_, _02880_);
  nor (_15276_, _15240_, _15239_);
  nand (_15277_, _15276_, _02880_);
  and (_15278_, _15277_, _03336_);
  and (_15279_, _15278_, _15274_);
  nor (_15280_, _15219_, _03336_);
  or (_15281_, _15280_, _07682_);
  or (_15282_, _15281_, _15279_);
  and (_15283_, _15282_, _15245_);
  or (_15284_, _15283_, _03399_);
  or (_15285_, _06154_, _03840_);
  and (_15287_, _15285_, _03084_);
  and (_15288_, _15287_, _15284_);
  nor (_15289_, _07442_, _03084_);
  or (_15290_, _15289_, _07692_);
  or (_15291_, _15290_, _15288_);
  nand (_15292_, _07692_, _05771_);
  and (_15293_, _15292_, _15291_);
  or (_15294_, _15293_, _02876_);
  and (_15295_, _12005_, _05325_);
  nor (_15296_, _15295_, _15239_);
  nand (_15298_, _15296_, _02876_);
  and (_15299_, _15298_, _02870_);
  and (_15300_, _15299_, _15294_);
  or (_15301_, _15300_, _15244_);
  and (_15302_, _15301_, _06253_);
  nor (_15303_, _06714_, _06712_);
  nor (_15304_, _15303_, _06715_);
  nand (_15305_, _15304_, _06247_);
  nand (_15306_, _15305_, _07718_);
  or (_15307_, _15306_, _15302_);
  nor (_15309_, _04435_, _06964_);
  nor (_15310_, _14944_, _15309_);
  and (_15311_, _15310_, _15201_);
  nor (_15312_, _15310_, _15201_);
  or (_15313_, _15312_, _15311_);
  nor (_15314_, _15313_, _07293_);
  and (_15315_, _15313_, _07293_);
  nor (_15316_, _15315_, _15314_);
  and (_15317_, _15316_, _14952_);
  nor (_15318_, _15316_, _14952_);
  nor (_15320_, _15318_, _15317_);
  or (_15321_, _15320_, _07718_);
  and (_15322_, _15321_, _07626_);
  and (_15323_, _15322_, _15307_);
  or (_15324_, _15323_, _15238_);
  and (_15325_, _15324_, _03111_);
  nor (_15326_, _14981_, _08085_);
  nor (_15327_, _09503_, _15326_);
  and (_15328_, _09503_, _15326_);
  or (_15329_, _15328_, _15327_);
  not (_15331_, _14986_);
  nor (_15332_, _15331_, _15329_);
  and (_15333_, _15331_, _15329_);
  nor (_15334_, _15333_, _15332_);
  nand (_15335_, _15334_, _07405_);
  and (_15336_, _15335_, _09562_);
  or (_15337_, _15336_, _15325_);
  and (_15338_, _03256_, \oc8051_golden_model_1.ACC [2]);
  nor (_15339_, _14997_, _15338_);
  not (_15340_, _09519_);
  and (_15342_, _15340_, _15339_);
  nor (_15343_, _15340_, _15339_);
  nor (_15344_, _15343_, _15342_);
  not (_15345_, _15000_);
  nor (_15346_, _15345_, _14999_);
  not (_15347_, _15346_);
  or (_15348_, _15347_, _15344_);
  nand (_15349_, _15347_, _15344_);
  and (_15350_, _15349_, _15348_);
  nand (_15351_, _15350_, _07404_);
  and (_15353_, _15351_, _15337_);
  or (_15354_, _15353_, _02583_);
  nand (_15355_, _02794_, _02583_);
  and (_15356_, _15355_, _02864_);
  and (_15357_, _15356_, _15354_);
  nor (_15358_, _12054_, _07833_);
  nor (_15359_, _15358_, _15239_);
  nor (_15360_, _15359_, _02864_);
  or (_15361_, _15360_, _06770_);
  or (_15362_, _15361_, _15357_);
  and (_15364_, _15362_, _15221_);
  or (_15365_, _15364_, _02853_);
  and (_15366_, _04706_, _06154_);
  nor (_15367_, _15366_, _15214_);
  nand (_15368_, _15367_, _02853_);
  and (_15369_, _15368_, _02838_);
  and (_15370_, _15369_, _15365_);
  nor (_15371_, _12112_, _07846_);
  nor (_15372_, _15371_, _15214_);
  nor (_15373_, _15372_, _02838_);
  or (_15375_, _15373_, _06784_);
  or (_15376_, _15375_, _15370_);
  or (_15377_, _06928_, _06791_);
  and (_15378_, _15377_, _15376_);
  and (_15379_, _15378_, _02635_);
  nor (_15380_, _02794_, _02635_);
  or (_15381_, _15380_, _02802_);
  or (_15382_, _15381_, _15379_);
  and (_15383_, _04706_, _05658_);
  nor (_15384_, _15383_, _15214_);
  nand (_15386_, _15384_, _02802_);
  and (_15387_, _15386_, _07860_);
  and (_15388_, _15387_, _15382_);
  nor (_15389_, _07860_, _02794_);
  or (_15390_, _15389_, _07876_);
  or (_15391_, _15390_, _15388_);
  or (_15392_, _07875_, _15201_);
  and (_15393_, _15392_, _07880_);
  and (_15394_, _15393_, _15391_);
  and (_15395_, _15227_, _07879_);
  or (_15397_, _15395_, _03129_);
  or (_15398_, _15397_, _15394_);
  or (_15399_, _12133_, _07890_);
  and (_15400_, _15399_, _07897_);
  and (_15401_, _15400_, _15398_);
  nor (_15402_, _07897_, _09519_);
  or (_15403_, _15402_, _02980_);
  or (_15404_, _15403_, _15401_);
  and (_15405_, _15404_, _15217_);
  or (_15406_, _15405_, _03127_);
  and (_15408_, _04149_, _02969_);
  nor (_15409_, _14864_, _15408_);
  or (_15410_, _15214_, _03128_);
  and (_15411_, _15410_, _15409_);
  and (_15412_, _15411_, _15406_);
  nor (_15413_, _15409_, _07205_);
  or (_15414_, _15413_, _15412_);
  or (_15415_, _15414_, _03518_);
  nand (_15416_, _07205_, _03518_);
  and (_15417_, _15416_, _15415_);
  or (_15419_, _15417_, _07911_);
  or (_15420_, _08037_, _07912_);
  and (_15421_, _15420_, _15419_);
  or (_15422_, _15421_, _03138_);
  or (_15423_, _12131_, _07396_);
  and (_15424_, _15423_, _07395_);
  and (_15425_, _15424_, _15422_);
  and (_15426_, _08124_, _07394_);
  or (_15427_, _15426_, _15425_);
  and (_15428_, _15427_, _03883_);
  or (_15430_, _15384_, _12132_);
  nor (_15431_, _15430_, _03883_);
  or (_15432_, _15431_, _15212_);
  or (_15433_, _15432_, _15428_);
  and (_15434_, _15433_, _15213_);
  or (_15435_, _15434_, _15206_);
  nand (_15436_, _15206_, _07202_);
  and (_15437_, _15436_, _03529_);
  and (_15438_, _15437_, _15435_);
  or (_15439_, _07935_, _03528_);
  not (_15441_, _07935_);
  nand (_15442_, _07202_, _15441_);
  and (_15443_, _15442_, _15439_);
  or (_15444_, _15443_, _15438_);
  nand (_15445_, _08035_, _07935_);
  and (_15446_, _15445_, _03122_);
  and (_15447_, _15446_, _15444_);
  nor (_15448_, _12132_, _03122_);
  or (_15449_, _15448_, _07942_);
  or (_15450_, _15449_, _15447_);
  nand (_15452_, _07942_, _08125_);
  and (_15453_, _15452_, _05783_);
  and (_15454_, _15453_, _15450_);
  nor (_15455_, _12125_, _07846_);
  nor (_15456_, _15455_, _15214_);
  nor (_15457_, _15456_, _05783_);
  or (_15458_, _15457_, _09711_);
  or (_15459_, _15458_, _15454_);
  and (_15460_, _07301_, _07279_);
  nor (_15461_, _15460_, _07302_);
  or (_15463_, _15461_, _07241_);
  and (_15464_, _07380_, _07359_);
  nor (_15465_, _15464_, _07381_);
  or (_15466_, _15465_, _07322_);
  and (_15467_, _15466_, _03134_);
  and (_15468_, _15467_, _15463_);
  and (_15469_, _15468_, _15459_);
  and (_15470_, _07976_, _07551_);
  nor (_15471_, _15470_, _07977_);
  or (_15472_, _15471_, _07962_);
  and (_15474_, _15472_, _10365_);
  or (_15475_, _15474_, _15469_);
  and (_15476_, _08004_, _07786_);
  nor (_15477_, _15476_, _08005_);
  or (_15478_, _15477_, _07993_);
  and (_15479_, _15478_, _07992_);
  and (_15480_, _15479_, _15475_);
  nand (_15481_, _07991_, \oc8051_golden_model_1.ACC [2]);
  nand (_15482_, _15481_, _07238_);
  or (_15483_, _15482_, _15480_);
  and (_15485_, _15483_, _15205_);
  or (_15486_, _15485_, _07188_);
  nor (_15487_, _08050_, _15227_);
  and (_15488_, _08050_, _15227_);
  nor (_15489_, _15488_, _15487_);
  nand (_15490_, _15489_, _07188_);
  and (_15491_, _15490_, _02896_);
  and (_15492_, _15491_, _15486_);
  nor (_15493_, _08094_, _09503_);
  and (_15494_, _08094_, _09503_);
  nor (_15496_, _15494_, _15493_);
  or (_15497_, _15496_, _08065_);
  and (_15498_, _15497_, _08067_);
  or (_15499_, _15498_, _15492_);
  nor (_15500_, _08136_, _09519_);
  and (_15501_, _08136_, _09519_);
  nor (_15502_, _15501_, _15500_);
  or (_15503_, _15502_, _08113_);
  and (_15504_, _15503_, _08112_);
  and (_15505_, _15504_, _15499_);
  and (_15507_, _08111_, \oc8051_golden_model_1.ACC [2]);
  or (_15508_, _15507_, _03163_);
  or (_15509_, _15508_, _15505_);
  nand (_15510_, _15262_, _03163_);
  and (_15511_, _15510_, _08155_);
  and (_15512_, _15511_, _15509_);
  nor (_15513_, _15170_, _02564_);
  or (_15514_, _15513_, _08161_);
  and (_15515_, _15514_, _08154_);
  or (_15516_, _15515_, _08159_);
  or (_15518_, _15516_, _15512_);
  nand (_15519_, _08159_, _06867_);
  and (_15520_, _15519_, _02498_);
  and (_15521_, _15520_, _15518_);
  nor (_15522_, _15296_, _02498_);
  or (_15523_, _15522_, _02888_);
  or (_15524_, _15523_, _15521_);
  and (_15525_, _12183_, _04706_);
  nor (_15526_, _15525_, _15214_);
  nand (_15527_, _15526_, _02888_);
  and (_15529_, _15527_, _08177_);
  and (_15530_, _15529_, _15524_);
  or (_15531_, _15189_, \oc8051_golden_model_1.ACC [3]);
  and (_15532_, _15531_, _08185_);
  and (_15533_, _15532_, _08176_);
  or (_15534_, _15533_, _08183_);
  or (_15535_, _15534_, _15530_);
  nand (_15536_, _08183_, _06867_);
  and (_15537_, _15536_, _42668_);
  and (_15538_, _15537_, _15535_);
  or (_15540_, _15538_, _15200_);
  and (_43425_, _15540_, _43998_);
  nor (_15541_, _42668_, _06867_);
  nand (_15542_, _08111_, _02564_);
  and (_15543_, _08006_, _07780_);
  nor (_15544_, _15543_, _08007_);
  or (_15545_, _15544_, _07993_);
  nor (_15546_, _04706_, _06867_);
  and (_15547_, _05666_, _04706_);
  nor (_15548_, _15547_, _15546_);
  or (_15550_, _15548_, _12206_);
  nor (_15551_, _15550_, _03883_);
  and (_15552_, _12211_, _04706_);
  nor (_15553_, _15552_, _15546_);
  nand (_15554_, _15553_, _02980_);
  not (_15555_, _03504_);
  or (_15556_, _08034_, _15555_);
  and (_15557_, _04706_, _04982_);
  nor (_15558_, _15557_, _15546_);
  nand (_15559_, _15558_, _06770_);
  or (_15561_, _07628_, _04982_);
  nor (_15562_, _07517_, _03387_);
  or (_15563_, _06159_, _07631_);
  and (_15564_, _07633_, _04982_);
  and (_15565_, _07636_, _06867_);
  nor (_15566_, _07636_, _06867_);
  or (_15567_, _15566_, _15565_);
  and (_15568_, _15567_, _07635_);
  or (_15569_, _15568_, _03363_);
  or (_15570_, _15569_, _15564_);
  and (_15572_, _15570_, _03387_);
  and (_15573_, _15572_, _15563_);
  or (_15574_, _15573_, _15562_);
  and (_15575_, _15574_, _07647_);
  nor (_15576_, _12217_, _07846_);
  nor (_15577_, _15576_, _15546_);
  nor (_15578_, _15577_, _03810_);
  or (_15579_, _15578_, _07649_);
  or (_15580_, _15579_, _15575_);
  nor (_15581_, _07656_, \oc8051_golden_model_1.ACC [4]);
  nor (_15583_, _15581_, _07662_);
  not (_15584_, _15583_);
  nand (_15585_, _15584_, _07649_);
  and (_15586_, _15585_, _03076_);
  and (_15587_, _15586_, _15580_);
  nor (_15588_, _05325_, _06867_);
  and (_15589_, _12231_, _05325_);
  nor (_15590_, _15589_, _15588_);
  nor (_15591_, _15590_, _02881_);
  nor (_15592_, _15558_, _03336_);
  or (_15594_, _15592_, _07682_);
  or (_15595_, _15594_, _15591_);
  or (_15596_, _15595_, _15587_);
  and (_15597_, _15596_, _15561_);
  or (_15598_, _15597_, _03399_);
  or (_15599_, _06159_, _03840_);
  and (_15600_, _15599_, _03084_);
  and (_15601_, _15600_, _15598_);
  nor (_15602_, _07517_, _03084_);
  or (_15603_, _15602_, _07692_);
  or (_15605_, _15603_, _15601_);
  nand (_15606_, _07692_, _02667_);
  and (_15607_, _15606_, _15605_);
  or (_15608_, _15607_, _02876_);
  and (_15609_, _12213_, _05325_);
  nor (_15610_, _15609_, _15588_);
  nand (_15611_, _15610_, _02876_);
  and (_15612_, _15611_, _02870_);
  and (_15613_, _15612_, _15608_);
  and (_15614_, _15589_, _12246_);
  nor (_15616_, _15614_, _15588_);
  nor (_15617_, _15616_, _02870_);
  or (_15618_, _15617_, _06247_);
  or (_15619_, _15618_, _15613_);
  nor (_15620_, _06717_, _06715_);
  nor (_15621_, _15620_, _06718_);
  or (_15622_, _15621_, _06253_);
  and (_15623_, _15622_, _15619_);
  or (_15624_, _15623_, _10106_);
  or (_15625_, _15317_, _15314_);
  and (_15627_, _04241_, _02564_);
  or (_15628_, _04241_, _02564_);
  and (_15629_, _15310_, _15628_);
  or (_15630_, _15629_, _15627_);
  nor (_15631_, _15630_, _07201_);
  and (_15632_, _15630_, _07201_);
  nor (_15633_, _15632_, _15631_);
  and (_15634_, _15633_, \oc8051_golden_model_1.PSW [7]);
  nor (_15635_, _15633_, \oc8051_golden_model_1.PSW [7]);
  nor (_15636_, _15635_, _15634_);
  and (_15638_, _15636_, _15625_);
  nor (_15639_, _15636_, _15625_);
  nor (_15640_, _15639_, _15638_);
  and (_15641_, _15640_, _07626_);
  or (_15642_, _15641_, _09557_);
  and (_15643_, _15642_, _15624_);
  or (_15644_, _15235_, _15232_);
  and (_15645_, _06154_, _02564_);
  or (_15646_, _06154_, _02564_);
  and (_15647_, _15646_, _15226_);
  or (_15649_, _15647_, _15645_);
  nor (_15650_, _08034_, _15649_);
  and (_15651_, _08034_, _15649_);
  nor (_15652_, _15651_, _15650_);
  and (_15653_, _15652_, \oc8051_golden_model_1.PSW [7]);
  nor (_15654_, _15652_, \oc8051_golden_model_1.PSW [7]);
  nor (_15655_, _15654_, _15653_);
  and (_15656_, _15655_, _15644_);
  nor (_15657_, _15655_, _15644_);
  nor (_15658_, _15657_, _15656_);
  and (_15660_, _15658_, _03434_);
  or (_15661_, _15660_, _03106_);
  or (_15662_, _15661_, _15643_);
  nor (_15663_, _15326_, _09501_);
  or (_15664_, _15663_, _09502_);
  and (_15665_, _08082_, _15664_);
  nor (_15666_, _08082_, _15664_);
  nor (_15667_, _15666_, _15665_);
  or (_15668_, _15332_, _15667_);
  nand (_15669_, _15332_, _15667_);
  and (_15671_, _15669_, _15668_);
  or (_15672_, _15671_, _03111_);
  and (_15673_, _15672_, _07405_);
  and (_15674_, _15673_, _15662_);
  nor (_15675_, _09524_, _07293_);
  nor (_15676_, _15339_, _10224_);
  nor (_15677_, _15676_, _10223_);
  nor (_15678_, _08123_, _15677_);
  and (_15679_, _08123_, _15677_);
  nor (_15680_, _15679_, _15678_);
  and (_15682_, _15680_, \oc8051_golden_model_1.PSW [7]);
  nor (_15683_, _15680_, \oc8051_golden_model_1.PSW [7]);
  nor (_15684_, _15683_, _15682_);
  and (_15685_, _15684_, _15675_);
  nor (_15686_, _15684_, _15675_);
  nor (_15687_, _15686_, _15685_);
  and (_15688_, _15687_, _07404_);
  or (_15689_, _15688_, _02583_);
  or (_15690_, _15689_, _15674_);
  nand (_15691_, _03629_, _02583_);
  and (_15693_, _15691_, _02864_);
  and (_15694_, _15693_, _15690_);
  nor (_15695_, _12264_, _07833_);
  nor (_15696_, _15695_, _15588_);
  nor (_15697_, _15696_, _02864_);
  or (_15698_, _15697_, _06770_);
  or (_15699_, _15698_, _15694_);
  and (_15700_, _15699_, _15559_);
  or (_15701_, _15700_, _02853_);
  and (_15702_, _04706_, _06159_);
  nor (_15704_, _15702_, _15546_);
  nand (_15705_, _15704_, _02853_);
  and (_15706_, _15705_, _02838_);
  and (_15707_, _15706_, _15701_);
  nor (_15708_, _12321_, _07846_);
  nor (_15709_, _15708_, _15546_);
  nor (_15710_, _15709_, _02838_);
  or (_15711_, _15710_, _06784_);
  or (_15712_, _15711_, _15707_);
  or (_15713_, _06874_, _06791_);
  and (_15715_, _15713_, _15712_);
  and (_15716_, _15715_, _02635_);
  nor (_15717_, _03629_, _02635_);
  or (_15718_, _15717_, _02802_);
  or (_15719_, _15718_, _15716_);
  nand (_15720_, _15548_, _02802_);
  and (_15721_, _15720_, _07860_);
  and (_15722_, _15721_, _15719_);
  nor (_15723_, _07860_, _03629_);
  or (_15724_, _15723_, _07869_);
  or (_15726_, _15724_, _15722_);
  or (_15727_, _07870_, _07201_);
  and (_15728_, _15727_, _14710_);
  and (_15729_, _15728_, _15726_);
  and (_15730_, _14714_, _07201_);
  or (_15731_, _15730_, _14713_);
  or (_15732_, _15731_, _15729_);
  and (_15733_, _05747_, _02508_);
  not (_15734_, _15733_);
  or (_15735_, _14719_, _07201_);
  and (_15737_, _15735_, _15734_);
  and (_15738_, _15737_, _15732_);
  or (_15739_, _08034_, _02462_);
  and (_15740_, _15739_, _07879_);
  or (_15741_, _15740_, _15738_);
  and (_15742_, _15741_, _15556_);
  or (_15743_, _15742_, _03129_);
  or (_15744_, _12207_, _07890_);
  and (_15745_, _15744_, _07897_);
  and (_15746_, _15745_, _15743_);
  and (_15748_, _07399_, _08123_);
  or (_15749_, _15748_, _02980_);
  or (_15750_, _15749_, _15746_);
  and (_15751_, _15750_, _15554_);
  or (_15752_, _15751_, _03127_);
  or (_15753_, _15546_, _03128_);
  and (_15754_, _15753_, _09081_);
  and (_15755_, _15754_, _15752_);
  and (_15756_, _08032_, _07911_);
  and (_15757_, _07908_, _07199_);
  or (_15759_, _15757_, _03138_);
  or (_15760_, _15759_, _15756_);
  or (_15761_, _15760_, _15755_);
  or (_15762_, _12205_, _07396_);
  and (_15763_, _15762_, _15761_);
  or (_15764_, _15763_, _07394_);
  or (_15765_, _08121_, _07395_);
  and (_15766_, _15765_, _03883_);
  and (_15767_, _15766_, _15764_);
  or (_15768_, _15767_, _15551_);
  and (_15770_, _15768_, _15211_);
  nor (_15771_, _15211_, _07200_);
  or (_15772_, _15771_, _15206_);
  or (_15773_, _15772_, _15770_);
  nand (_15774_, _15206_, _07200_);
  and (_15775_, _15774_, _03529_);
  and (_15776_, _15775_, _15773_);
  nand (_15777_, _07200_, _15441_);
  and (_15778_, _15777_, _15439_);
  or (_15779_, _15778_, _15776_);
  nand (_15781_, _08033_, _07935_);
  and (_15782_, _15781_, _03122_);
  and (_15783_, _15782_, _15779_);
  nor (_15784_, _12206_, _03122_);
  or (_15785_, _15784_, _07942_);
  or (_15786_, _15785_, _15783_);
  nand (_15787_, _07942_, _08122_);
  and (_15788_, _15787_, _15786_);
  or (_15789_, _15788_, _02965_);
  nor (_15790_, _12209_, _07846_);
  nor (_15792_, _15790_, _15546_);
  nand (_15793_, _15792_, _02965_);
  and (_15794_, _15793_, _07322_);
  and (_15795_, _15794_, _15789_);
  and (_15796_, _07382_, _07351_);
  nor (_15797_, _15796_, _07383_);
  and (_15798_, _15797_, _10349_);
  or (_15799_, _15798_, _07240_);
  or (_15800_, _15799_, _15795_);
  and (_15801_, _07303_, _07271_);
  nor (_15803_, _15801_, _07304_);
  or (_15804_, _15803_, _07241_);
  and (_15805_, _15804_, _03134_);
  and (_15806_, _15805_, _15800_);
  and (_15807_, _07978_, _07544_);
  nor (_15808_, _15807_, _07979_);
  or (_15809_, _15808_, _07962_);
  and (_15810_, _15809_, _10365_);
  or (_15811_, _15810_, _15806_);
  and (_15812_, _15811_, _15545_);
  or (_15814_, _15812_, _07991_);
  nand (_15815_, _07991_, _02564_);
  and (_15816_, _15815_, _07238_);
  and (_15817_, _15816_, _15814_);
  nor (_15818_, _07219_, _07201_);
  nor (_15819_, _15818_, _07220_);
  and (_15820_, _15819_, _10378_);
  or (_15821_, _15820_, _07188_);
  or (_15822_, _15821_, _15817_);
  nor (_15823_, _08052_, _08034_);
  nor (_15825_, _15823_, _08053_);
  or (_15826_, _15825_, _08024_);
  and (_15827_, _15826_, _15822_);
  or (_15828_, _15827_, _02894_);
  nor (_15829_, _08098_, _08083_);
  nor (_15830_, _15829_, _08099_);
  or (_15831_, _15830_, _02896_);
  and (_15832_, _15831_, _08113_);
  and (_15833_, _15832_, _15828_);
  nor (_15834_, _08138_, _08123_);
  nor (_15836_, _15834_, _08139_);
  and (_15837_, _15836_, _08065_);
  or (_15838_, _15837_, _08111_);
  or (_15839_, _15838_, _15833_);
  and (_15840_, _15839_, _15542_);
  or (_15841_, _15840_, _03163_);
  nand (_15842_, _15577_, _03163_);
  and (_15843_, _15842_, _08155_);
  and (_15844_, _15843_, _15841_);
  and (_15845_, _08161_, _06867_);
  nor (_15847_, _08161_, _06867_);
  nor (_15848_, _15847_, _15845_);
  not (_15849_, _15848_);
  and (_15850_, _15849_, _08154_);
  or (_15851_, _15850_, _08159_);
  or (_15852_, _15851_, _15844_);
  nand (_15853_, _08159_, _06861_);
  and (_15854_, _15853_, _02498_);
  and (_15855_, _15854_, _15852_);
  nor (_15856_, _15610_, _02498_);
  or (_15858_, _15856_, _02888_);
  or (_15859_, _15858_, _15855_);
  and (_15860_, _12389_, _04706_);
  nor (_15861_, _15860_, _15546_);
  nand (_15862_, _15861_, _02888_);
  and (_15863_, _15862_, _08177_);
  and (_15864_, _15863_, _15859_);
  and (_15865_, _08185_, _06867_);
  nor (_15866_, _15865_, _08186_);
  nor (_15867_, _15866_, _08183_);
  nor (_15869_, _15867_, _09044_);
  or (_15870_, _15869_, _15864_);
  nand (_15871_, _08183_, _06861_);
  and (_15872_, _15871_, _42668_);
  and (_15873_, _15872_, _15870_);
  or (_15874_, _15873_, _15541_);
  and (_43426_, _15874_, _43998_);
  nor (_15875_, _42668_, _06861_);
  and (_15876_, _07221_, _07198_);
  nor (_15877_, _15876_, _07222_);
  or (_15879_, _15877_, _07238_);
  or (_15880_, _08028_, _07912_);
  nor (_15881_, _04706_, _06861_);
  and (_15882_, _12415_, _04706_);
  nor (_15883_, _15882_, _15881_);
  nand (_15884_, _15883_, _02980_);
  or (_15885_, _08030_, _15555_);
  and (_15886_, _04706_, _04877_);
  nor (_15887_, _15886_, _15881_);
  nand (_15888_, _15887_, _06770_);
  and (_15890_, _03629_, \oc8051_golden_model_1.ACC [4]);
  nor (_15891_, _15678_, _15890_);
  nor (_15892_, _08119_, _15891_);
  and (_15893_, _08119_, _15891_);
  nor (_15894_, _15893_, _15892_);
  and (_15895_, _15894_, \oc8051_golden_model_1.PSW [7]);
  nor (_15896_, _15894_, \oc8051_golden_model_1.PSW [7]);
  nor (_15897_, _15896_, _15895_);
  nor (_15898_, _15685_, _15682_);
  not (_15899_, _15898_);
  and (_15901_, _15899_, _15897_);
  nor (_15902_, _15899_, _15897_);
  nor (_15903_, _15902_, _15901_);
  or (_15904_, _15903_, _07405_);
  and (_15905_, _06123_, \oc8051_golden_model_1.ACC [4]);
  nor (_15906_, _15650_, _15905_);
  and (_15907_, _08031_, _15906_);
  nor (_15908_, _08031_, _15906_);
  nor (_15909_, _15908_, _15907_);
  nor (_15910_, _15909_, _07293_);
  and (_15912_, _15909_, _07293_);
  nor (_15913_, _15912_, _15910_);
  nor (_15914_, _15656_, _15653_);
  not (_15915_, _15914_);
  and (_15916_, _15915_, _15913_);
  nor (_15917_, _15915_, _15913_);
  nor (_15918_, _15917_, _15916_);
  and (_15919_, _15918_, _03434_);
  nor (_15920_, _05325_, _06861_);
  and (_15921_, _12435_, _05325_);
  and (_15923_, _15921_, _12450_);
  nor (_15924_, _15923_, _15920_);
  nor (_15925_, _15924_, _02870_);
  or (_15926_, _07628_, _04877_);
  nor (_15927_, _07504_, _03387_);
  or (_15928_, _06158_, _07631_);
  and (_15929_, _07633_, _04877_);
  and (_15930_, _07636_, _06861_);
  nor (_15931_, _07636_, _06861_);
  or (_15932_, _15931_, _15930_);
  and (_15934_, _15932_, _07635_);
  or (_15935_, _15934_, _03363_);
  or (_15936_, _15935_, _15929_);
  and (_15937_, _15936_, _03387_);
  and (_15938_, _15937_, _15928_);
  or (_15939_, _15938_, _15927_);
  and (_15940_, _15939_, _07647_);
  nor (_15941_, _12407_, _07846_);
  nor (_15942_, _15941_, _15881_);
  nor (_15943_, _15942_, _03810_);
  or (_15945_, _15943_, _07649_);
  or (_15946_, _15945_, _15940_);
  and (_15947_, _10122_, _07664_);
  nor (_15948_, _10122_, _07664_);
  nor (_15949_, _15948_, _15947_);
  nand (_15950_, _15949_, _07649_);
  and (_15951_, _15950_, _03076_);
  and (_15952_, _15951_, _15946_);
  nor (_15953_, _15921_, _15920_);
  nor (_15954_, _15953_, _02881_);
  nor (_15956_, _15887_, _03336_);
  or (_15957_, _15956_, _07682_);
  or (_15958_, _15957_, _15954_);
  or (_15959_, _15958_, _15952_);
  and (_15960_, _15959_, _15926_);
  or (_15961_, _15960_, _03399_);
  or (_15962_, _06158_, _03840_);
  and (_15963_, _15962_, _03084_);
  and (_15964_, _15963_, _15961_);
  nor (_15965_, _07504_, _03084_);
  or (_15967_, _15965_, _07692_);
  or (_15968_, _15967_, _15964_);
  nand (_15969_, _07692_, _02551_);
  and (_15970_, _15969_, _15968_);
  or (_15971_, _15970_, _02876_);
  and (_15972_, _12417_, _05325_);
  nor (_15973_, _15972_, _15920_);
  nand (_15974_, _15973_, _02876_);
  and (_15975_, _15974_, _02870_);
  and (_15976_, _15975_, _15971_);
  or (_15978_, _15976_, _15925_);
  and (_15979_, _15978_, _06253_);
  nor (_15980_, _06720_, _06718_);
  nor (_15981_, _15980_, _06721_);
  and (_15982_, _15981_, _06247_);
  or (_15983_, _15982_, _10106_);
  or (_15984_, _15983_, _15979_);
  nor (_15985_, _04982_, _06867_);
  nor (_15986_, _15631_, _15985_);
  nor (_15987_, _15986_, _07197_);
  and (_15989_, _15986_, _07197_);
  nor (_15990_, _15989_, _15987_);
  and (_15991_, _15990_, \oc8051_golden_model_1.PSW [7]);
  nor (_15992_, _15990_, \oc8051_golden_model_1.PSW [7]);
  nor (_15993_, _15992_, _15991_);
  nor (_15994_, _15638_, _15634_);
  not (_15995_, _15994_);
  and (_15996_, _15995_, _15993_);
  nor (_15997_, _15995_, _15993_);
  nor (_15998_, _15997_, _15996_);
  or (_16000_, _15998_, _07718_);
  and (_16001_, _16000_, _07626_);
  and (_16002_, _16001_, _15984_);
  or (_16003_, _16002_, _15919_);
  and (_16004_, _16003_, _03111_);
  not (_16005_, _09509_);
  nor (_16006_, _16005_, _15667_);
  nor (_16007_, _16006_, _07293_);
  not (_16008_, _16007_);
  nor (_16009_, _15665_, _08080_);
  nor (_16011_, _08078_, _16009_);
  and (_16012_, _08078_, _16009_);
  or (_16013_, _16012_, _16011_);
  and (_16014_, _16013_, _07293_);
  nor (_16015_, _16013_, _07293_);
  nor (_16016_, _16015_, _16014_);
  and (_16017_, _16016_, _16008_);
  nor (_16018_, _16016_, _16008_);
  nor (_16019_, _16018_, _16017_);
  or (_16020_, _16019_, _07404_);
  and (_16022_, _16020_, _09562_);
  or (_16023_, _16022_, _16004_);
  and (_16024_, _16023_, _15904_);
  or (_16025_, _16024_, _02583_);
  nand (_16026_, _03211_, _02583_);
  and (_16027_, _16026_, _02864_);
  and (_16028_, _16027_, _16025_);
  nor (_16029_, _12468_, _07833_);
  nor (_16030_, _16029_, _15920_);
  nor (_16031_, _16030_, _02864_);
  or (_16033_, _16031_, _06770_);
  or (_16034_, _16033_, _16028_);
  and (_16035_, _16034_, _15888_);
  or (_16036_, _16035_, _02853_);
  and (_16037_, _04706_, _06158_);
  nor (_16038_, _16037_, _15881_);
  nand (_16039_, _16038_, _02853_);
  and (_16040_, _16039_, _02838_);
  and (_16041_, _16040_, _16036_);
  nor (_16042_, _12527_, _07846_);
  nor (_16044_, _16042_, _15881_);
  nor (_16045_, _16044_, _02838_);
  or (_16046_, _16045_, _06784_);
  or (_16047_, _16046_, _16041_);
  or (_16048_, _06844_, _06791_);
  and (_16049_, _16048_, _16047_);
  and (_16050_, _16049_, _02635_);
  nor (_16051_, _03211_, _02635_);
  or (_16052_, _16051_, _02802_);
  or (_16053_, _16052_, _16050_);
  and (_16055_, _05614_, _04706_);
  nor (_16056_, _16055_, _15881_);
  nand (_16057_, _16056_, _02802_);
  and (_16058_, _16057_, _07860_);
  and (_16059_, _16058_, _16053_);
  nor (_16060_, _07860_, _03211_);
  or (_16061_, _16060_, _07876_);
  or (_16062_, _16061_, _16059_);
  or (_16063_, _07875_, _07197_);
  and (_16064_, _16063_, _15734_);
  and (_16066_, _16064_, _16062_);
  or (_16067_, _08030_, _02462_);
  and (_16068_, _16067_, _07879_);
  or (_16069_, _16068_, _16066_);
  and (_16070_, _16069_, _15885_);
  or (_16071_, _16070_, _03129_);
  or (_16072_, _12411_, _07890_);
  and (_16073_, _16072_, _07897_);
  and (_16074_, _16073_, _16071_);
  and (_16075_, _07399_, _08119_);
  or (_16077_, _16075_, _02980_);
  or (_16078_, _16077_, _16074_);
  and (_16079_, _16078_, _15884_);
  or (_16080_, _16079_, _03127_);
  or (_16081_, _15881_, _03128_);
  and (_16082_, _16081_, _07907_);
  and (_16083_, _16082_, _16080_);
  and (_16084_, _07908_, _07195_);
  or (_16085_, _16084_, _07911_);
  or (_16086_, _16085_, _16083_);
  and (_16088_, _16086_, _15880_);
  or (_16089_, _16088_, _03138_);
  or (_16090_, _12409_, _07396_);
  and (_16091_, _16090_, _07395_);
  and (_16092_, _16091_, _16089_);
  and (_16093_, _08117_, _07394_);
  or (_16094_, _16093_, _16092_);
  and (_16095_, _16094_, _03883_);
  or (_16096_, _16056_, _12410_);
  nor (_16097_, _16096_, _03883_);
  or (_16099_, _16097_, _15212_);
  or (_16100_, _16099_, _16095_);
  nand (_16101_, _15212_, _07196_);
  nor (_16102_, _03535_, _07930_);
  and (_16103_, _16102_, _16101_);
  and (_16104_, _16103_, _16100_);
  nor (_16105_, _16102_, _07196_);
  or (_16106_, _16105_, _07935_);
  or (_16107_, _16106_, _16104_);
  nand (_16108_, _08029_, _07935_);
  and (_16110_, _16108_, _03122_);
  and (_16111_, _16110_, _16107_);
  nand (_16112_, _12410_, _07945_);
  and (_16113_, _16112_, _07944_);
  or (_16114_, _16113_, _16111_);
  nand (_16115_, _07942_, _08118_);
  and (_16116_, _16115_, _05783_);
  and (_16117_, _16116_, _16114_);
  nor (_16118_, _12413_, _07846_);
  nor (_16119_, _16118_, _15881_);
  or (_16121_, _16119_, _05783_);
  and (_16122_, _04009_, _02967_);
  not (_16123_, _16122_);
  and (_16124_, _07321_, _16123_);
  nand (_16125_, _16124_, _16121_);
  or (_16126_, _16125_, _16117_);
  not (_16127_, _03546_);
  and (_16128_, _07384_, _07343_);
  nor (_16129_, _16128_, _07385_);
  or (_16130_, _16129_, _16124_);
  and (_16132_, _16130_, _16127_);
  and (_16133_, _16132_, _16126_);
  and (_16134_, _16129_, _03546_);
  or (_16135_, _16134_, _07240_);
  or (_16136_, _16135_, _16133_);
  and (_16137_, _07305_, _07263_);
  nor (_16138_, _16137_, _07306_);
  or (_16139_, _16138_, _07241_);
  and (_16140_, _16139_, _03134_);
  and (_16141_, _16140_, _16136_);
  and (_16143_, _07980_, _07539_);
  nor (_16144_, _16143_, _07981_);
  or (_16145_, _16144_, _07962_);
  and (_16146_, _16145_, _10365_);
  or (_16147_, _16146_, _16141_);
  and (_16148_, _08008_, _07775_);
  nor (_16149_, _16148_, _08009_);
  or (_16150_, _16149_, _07993_);
  and (_16151_, _16150_, _07992_);
  and (_16152_, _16151_, _16147_);
  nand (_16154_, _07991_, \oc8051_golden_model_1.ACC [4]);
  nand (_16155_, _16154_, _07238_);
  or (_16156_, _16155_, _16152_);
  and (_16157_, _16156_, _15879_);
  or (_16158_, _16157_, _07188_);
  and (_16159_, _08054_, _08031_);
  nor (_16160_, _16159_, _08055_);
  or (_16161_, _16160_, _08024_);
  and (_16162_, _16161_, _02896_);
  and (_16163_, _16162_, _16158_);
  and (_16165_, _08100_, _08078_);
  nor (_16166_, _16165_, _08101_);
  or (_16167_, _16166_, _08065_);
  and (_16168_, _16167_, _08067_);
  or (_16169_, _16168_, _16163_);
  and (_16170_, _08140_, _08120_);
  nor (_16171_, _16170_, _08141_);
  or (_16172_, _16171_, _08113_);
  and (_16173_, _16172_, _08112_);
  and (_16174_, _16173_, _16169_);
  and (_16176_, _08111_, \oc8051_golden_model_1.ACC [4]);
  or (_16177_, _16176_, _03163_);
  or (_16178_, _16177_, _16174_);
  nand (_16179_, _15942_, _03163_);
  and (_16180_, _16179_, _08155_);
  and (_16181_, _16180_, _16178_);
  nor (_16182_, _15845_, _06861_);
  or (_16183_, _16182_, _08162_);
  nor (_16184_, _16183_, _08159_);
  nor (_16185_, _16184_, _09948_);
  or (_16187_, _16185_, _16181_);
  nand (_16188_, _08159_, _06806_);
  and (_16189_, _16188_, _02498_);
  and (_16190_, _16189_, _16187_);
  nor (_16191_, _15973_, _02498_);
  or (_16192_, _16191_, _02888_);
  or (_16193_, _16192_, _16190_);
  and (_16194_, _12589_, _04706_);
  nor (_16195_, _16194_, _15881_);
  nand (_16196_, _16195_, _02888_);
  and (_16198_, _16196_, _08177_);
  and (_16199_, _16198_, _16193_);
  nor (_16200_, _08186_, \oc8051_golden_model_1.ACC [5]);
  nor (_16201_, _16200_, _08187_);
  nor (_16202_, _16201_, _08183_);
  nor (_16203_, _16202_, _09044_);
  or (_16204_, _16203_, _16199_);
  nand (_16205_, _08183_, _06806_);
  and (_16206_, _16205_, _42668_);
  and (_16207_, _16206_, _16204_);
  or (_16209_, _16207_, _15875_);
  and (_43427_, _16209_, _43998_);
  nor (_16210_, _42668_, _06806_);
  nand (_16211_, _08111_, _06861_);
  and (_16212_, _08010_, _07769_);
  nor (_16213_, _16212_, _08011_);
  or (_16214_, _16213_, _07993_);
  nand (_16215_, _07925_, _07193_);
  nor (_16216_, _04706_, _06806_);
  and (_16217_, _12739_, _04706_);
  nor (_16219_, _16217_, _16216_);
  nand (_16220_, _16219_, _02980_);
  or (_16221_, _07871_, _07194_);
  and (_16222_, _04706_, _04770_);
  nor (_16223_, _16222_, _16216_);
  nand (_16224_, _16223_, _06770_);
  nor (_16225_, _16007_, _16013_);
  nor (_16226_, _16014_, _16225_);
  not (_16227_, _16226_);
  nor (_16228_, _16009_, _08076_);
  or (_16230_, _16228_, _08077_);
  and (_16231_, _16230_, _08074_);
  nor (_16232_, _16230_, _08074_);
  nor (_16233_, _16232_, _16231_);
  nor (_16234_, _16233_, \oc8051_golden_model_1.PSW [7]);
  and (_16235_, _16233_, \oc8051_golden_model_1.PSW [7]);
  or (_16236_, _16235_, _16234_);
  nor (_16237_, _16236_, _16227_);
  and (_16238_, _16236_, _16227_);
  nor (_16239_, _16238_, _16237_);
  or (_16241_, _16239_, _03111_);
  and (_16242_, _16241_, _07405_);
  or (_16243_, _06158_, _06861_);
  and (_16244_, _06158_, _06861_);
  or (_16245_, _15906_, _16244_);
  and (_16246_, _16245_, _16243_);
  nor (_16247_, _16246_, _08027_);
  and (_16248_, _16246_, _08027_);
  nor (_16249_, _16248_, _16247_);
  nor (_16250_, _15916_, _15910_);
  and (_16252_, _16250_, \oc8051_golden_model_1.PSW [7]);
  or (_16253_, _16252_, _16249_);
  nand (_16254_, _16252_, _16249_);
  and (_16255_, _16254_, _16253_);
  and (_16256_, _16255_, _03434_);
  or (_16257_, _07628_, _04770_);
  nor (_16258_, _07424_, _03387_);
  or (_16259_, _05849_, _07631_);
  or (_16260_, _07635_, _04770_);
  nor (_16261_, _07636_, \oc8051_golden_model_1.ACC [6]);
  and (_16263_, _07636_, \oc8051_golden_model_1.ACC [6]);
  or (_16264_, _16263_, _16261_);
  nand (_16265_, _16264_, _09427_);
  and (_16266_, _16265_, _16260_);
  and (_16267_, _16266_, _03387_);
  and (_16268_, _16267_, _16259_);
  or (_16269_, _16268_, _16258_);
  and (_16270_, _16269_, _07647_);
  nor (_16271_, _12603_, _07846_);
  nor (_16272_, _16271_, _16216_);
  nor (_16274_, _16272_, _03810_);
  or (_16275_, _16274_, _07649_);
  or (_16276_, _16275_, _16270_);
  not (_16277_, _07666_);
  nor (_16278_, _15948_, _16277_);
  and (_16279_, _10121_, _07667_);
  nor (_16280_, _16279_, _16278_);
  nand (_16281_, _16280_, _07649_);
  and (_16282_, _16281_, _03076_);
  and (_16283_, _16282_, _16276_);
  nor (_16285_, _05325_, _06806_);
  and (_16286_, _12618_, _05325_);
  nor (_16287_, _16286_, _16285_);
  nor (_16288_, _16287_, _02881_);
  nor (_16289_, _16223_, _03336_);
  or (_16290_, _16289_, _07682_);
  or (_16291_, _16290_, _16288_);
  or (_16292_, _16291_, _16283_);
  and (_16293_, _16292_, _16257_);
  or (_16294_, _16293_, _03399_);
  or (_16296_, _05849_, _03840_);
  and (_16297_, _16296_, _03084_);
  and (_16298_, _16297_, _16294_);
  nor (_16299_, _07424_, _03084_);
  or (_16300_, _16299_, _07692_);
  or (_16301_, _16300_, _16298_);
  nand (_16302_, _07692_, _06964_);
  and (_16303_, _16302_, _16301_);
  or (_16304_, _16303_, _02876_);
  and (_16305_, _12616_, _05325_);
  nor (_16307_, _16305_, _16285_);
  nand (_16308_, _16307_, _02876_);
  and (_16309_, _16308_, _02870_);
  and (_16310_, _16309_, _16304_);
  and (_16311_, _16286_, _12646_);
  nor (_16312_, _16311_, _16285_);
  nor (_16313_, _16312_, _02870_);
  or (_16314_, _16313_, _06247_);
  or (_16315_, _16314_, _16310_);
  nor (_16316_, _06723_, _06721_);
  nor (_16318_, _16316_, _06724_);
  or (_16319_, _16318_, _06253_);
  and (_16320_, _16319_, _16315_);
  or (_16321_, _16320_, _10106_);
  or (_16322_, _04877_, _06861_);
  and (_16323_, _04877_, _06861_);
  or (_16324_, _15986_, _16323_);
  and (_16325_, _16324_, _16322_);
  nor (_16326_, _16325_, _07194_);
  and (_16327_, _16325_, _07194_);
  nor (_16329_, _16327_, _16326_);
  nor (_16330_, _15996_, _15991_);
  and (_16331_, _16330_, \oc8051_golden_model_1.PSW [7]);
  nor (_16332_, _16331_, _16329_);
  and (_16333_, _16331_, _16329_);
  nor (_16334_, _16333_, _16332_);
  or (_16335_, _16334_, _07718_);
  and (_16336_, _16335_, _07626_);
  and (_16337_, _16336_, _16321_);
  or (_16338_, _16337_, _03106_);
  or (_16340_, _16338_, _16256_);
  and (_16341_, _16340_, _16242_);
  nor (_16342_, _15891_, _10216_);
  nor (_16343_, _16342_, _10215_);
  nor (_16344_, _16343_, _08116_);
  and (_16345_, _16343_, _08116_);
  nor (_16346_, _16345_, _16344_);
  nor (_16347_, _15901_, _15895_);
  and (_16348_, _16347_, \oc8051_golden_model_1.PSW [7]);
  or (_16349_, _16348_, _16346_);
  nand (_16351_, _16348_, _16346_);
  and (_16352_, _16351_, _16349_);
  and (_16353_, _16352_, _07404_);
  or (_16354_, _16353_, _02583_);
  or (_16355_, _16354_, _16341_);
  nand (_16356_, _02927_, _02583_);
  and (_16357_, _16356_, _02864_);
  and (_16358_, _16357_, _16355_);
  nor (_16359_, _12664_, _07833_);
  nor (_16360_, _16359_, _16285_);
  nor (_16362_, _16360_, _02864_);
  or (_16363_, _16362_, _06770_);
  or (_16364_, _16363_, _16358_);
  and (_16365_, _16364_, _16224_);
  or (_16366_, _16365_, _02853_);
  and (_16367_, _04706_, _05849_);
  nor (_16368_, _16367_, _16216_);
  nand (_16369_, _16368_, _02853_);
  and (_16370_, _16369_, _02838_);
  and (_16371_, _16370_, _16366_);
  nor (_16373_, _12722_, _07846_);
  nor (_16374_, _16373_, _16216_);
  nor (_16375_, _16374_, _02838_);
  or (_16376_, _16375_, _06784_);
  or (_16377_, _16376_, _16371_);
  not (_16378_, _06807_);
  and (_16379_, _06812_, _16378_);
  not (_16380_, _16379_);
  nand (_16381_, _16380_, _06784_);
  and (_16382_, _16381_, _16377_);
  and (_16384_, _16382_, _02635_);
  nor (_16385_, _02927_, _02635_);
  or (_16386_, _16385_, _02802_);
  or (_16387_, _16386_, _16384_);
  and (_16388_, _12729_, _04706_);
  nor (_16389_, _16388_, _16216_);
  nand (_16390_, _16389_, _02802_);
  and (_16391_, _16390_, _07860_);
  and (_16392_, _16391_, _16387_);
  nand (_16393_, _07871_, _03510_);
  nor (_16395_, _07860_, _02927_);
  or (_16396_, _16395_, _16393_);
  or (_16397_, _16396_, _16392_);
  and (_16398_, _16397_, _16221_);
  or (_16399_, _16398_, _14713_);
  and (_16400_, _07879_, _02543_);
  not (_16401_, _16400_);
  or (_16402_, _07874_, _07194_);
  and (_16403_, _16402_, _16401_);
  and (_16404_, _16403_, _16399_);
  and (_16406_, _15733_, _08027_);
  or (_16407_, _16406_, _16404_);
  and (_16408_, _16407_, _15555_);
  and (_16409_, _08027_, _03504_);
  or (_16410_, _16409_, _03129_);
  or (_16411_, _16410_, _16408_);
  or (_16412_, _12613_, _07890_);
  and (_16413_, _16412_, _07897_);
  and (_16414_, _16413_, _16411_);
  and (_16415_, _07399_, _08116_);
  or (_16417_, _16415_, _02980_);
  or (_16418_, _16417_, _16414_);
  and (_16419_, _16418_, _16220_);
  or (_16420_, _16419_, _03127_);
  or (_16421_, _16216_, _03128_);
  and (_16422_, _16421_, _07907_);
  and (_16423_, _16422_, _16420_);
  and (_16424_, _07908_, _07192_);
  or (_16425_, _16424_, _07911_);
  or (_16426_, _16425_, _16423_);
  or (_16428_, _08025_, _07912_);
  and (_16429_, _16428_, _16426_);
  or (_16430_, _16429_, _03138_);
  or (_16431_, _12611_, _07396_);
  and (_16432_, _16431_, _07395_);
  and (_16433_, _16432_, _16430_);
  and (_16434_, _08114_, _07394_);
  or (_16435_, _16434_, _16433_);
  and (_16436_, _16435_, _03883_);
  or (_16437_, _16389_, _12612_);
  nor (_16439_, _16437_, _03883_);
  or (_16440_, _16439_, _07925_);
  or (_16441_, _16440_, _16436_);
  and (_16442_, _16441_, _16215_);
  or (_16443_, _16442_, _14763_);
  nand (_16444_, _14763_, _07193_);
  and (_16445_, _16444_, _03529_);
  and (_16446_, _16445_, _16443_);
  nor (_16447_, _07193_, _03529_);
  or (_16448_, _16447_, _07935_);
  or (_16450_, _16448_, _16446_);
  nand (_16451_, _08026_, _07935_);
  and (_16452_, _16451_, _03122_);
  and (_16453_, _16452_, _16450_);
  nor (_16454_, _12612_, _03122_);
  or (_16455_, _16454_, _07942_);
  or (_16456_, _16455_, _16453_);
  nand (_16457_, _07942_, _08115_);
  and (_16458_, _16457_, _16456_);
  or (_16459_, _16458_, _02965_);
  nor (_16461_, _12737_, _07846_);
  nor (_16462_, _16461_, _16216_);
  nand (_16463_, _16462_, _02965_);
  and (_16464_, _16463_, _07322_);
  and (_16465_, _16464_, _16459_);
  and (_16466_, _07386_, _07336_);
  nor (_16467_, _16466_, _07387_);
  and (_16468_, _16467_, _10349_);
  or (_16469_, _16468_, _07240_);
  or (_16470_, _16469_, _16465_);
  and (_16472_, _07307_, _07255_);
  nor (_16473_, _16472_, _07308_);
  or (_16474_, _16473_, _07241_);
  and (_16475_, _16474_, _03134_);
  and (_16476_, _16475_, _16470_);
  and (_16477_, _07982_, _07964_);
  nor (_16478_, _16477_, _07983_);
  or (_16479_, _16478_, _07962_);
  and (_16480_, _16479_, _10365_);
  or (_16481_, _16480_, _16476_);
  and (_16483_, _16481_, _16214_);
  or (_16484_, _16483_, _07991_);
  nand (_16485_, _07991_, _06861_);
  and (_16486_, _16485_, _07238_);
  and (_16487_, _16486_, _16484_);
  nor (_16488_, _07223_, _07194_);
  nor (_16489_, _16488_, _07224_);
  and (_16490_, _16489_, _10378_);
  or (_16491_, _16490_, _16487_);
  and (_16492_, _16491_, _08024_);
  nor (_16494_, _08056_, _08027_);
  nor (_16495_, _16494_, _08057_);
  and (_16496_, _16495_, _07188_);
  or (_16497_, _16496_, _02894_);
  or (_16498_, _16497_, _16492_);
  and (_16499_, _08102_, _08074_);
  nor (_16500_, _16499_, _08103_);
  or (_16501_, _16500_, _02896_);
  and (_16502_, _16501_, _08113_);
  and (_16503_, _16502_, _16498_);
  nor (_16505_, _08142_, _08116_);
  nor (_16506_, _16505_, _08143_);
  and (_16507_, _16506_, _08065_);
  or (_16508_, _16507_, _08111_);
  or (_16509_, _16508_, _16503_);
  and (_16510_, _16509_, _16211_);
  or (_16511_, _16510_, _03163_);
  nand (_16512_, _16272_, _03163_);
  and (_16513_, _16512_, _08155_);
  and (_16514_, _16513_, _16511_);
  nor (_16516_, _08162_, _06806_);
  or (_16517_, _16516_, _08163_);
  nor (_16518_, _16517_, _08159_);
  nor (_16519_, _16518_, _09948_);
  or (_16520_, _16519_, _16514_);
  nand (_16521_, _08159_, _05771_);
  and (_16522_, _16521_, _02498_);
  and (_16523_, _16522_, _16520_);
  nor (_16524_, _16307_, _02498_);
  or (_16525_, _16524_, _02888_);
  or (_16527_, _16525_, _16523_);
  and (_16528_, _12794_, _04706_);
  nor (_16529_, _16528_, _16216_);
  nand (_16530_, _16529_, _02888_);
  and (_16531_, _16530_, _08177_);
  and (_16532_, _16531_, _16527_);
  nor (_16533_, _08187_, \oc8051_golden_model_1.ACC [6]);
  nor (_16534_, _16533_, _08188_);
  and (_16535_, _16534_, _08176_);
  or (_16536_, _16535_, _08183_);
  or (_16538_, _16536_, _16532_);
  nand (_16539_, _08183_, _05771_);
  and (_16540_, _16539_, _42668_);
  and (_16541_, _16540_, _16538_);
  or (_16542_, _16541_, _16210_);
  and (_43428_, _16542_, _43998_);
  not (_16543_, \oc8051_golden_model_1.DPL [0]);
  nor (_16544_, _42668_, _16543_);
  and (_16545_, _05226_, _04612_);
  nor (_16546_, _04612_, _16543_);
  and (_16548_, _04612_, _05672_);
  or (_16549_, _16548_, _16546_);
  nand (_16550_, _16549_, _02970_);
  nor (_16551_, _16550_, _16545_);
  and (_16552_, _11522_, _04612_);
  or (_16553_, _16552_, _16546_);
  and (_16554_, _16553_, _03127_);
  and (_16555_, _04612_, _06152_);
  or (_16556_, _16555_, _16546_);
  and (_16557_, _16556_, _02853_);
  and (_16559_, _08224_, _16543_);
  and (_16560_, _04612_, _03808_);
  or (_16561_, _16560_, _16546_);
  or (_16562_, _16561_, _03336_);
  or (_16563_, _16546_, _16545_);
  and (_16564_, _16563_, _02974_);
  nor (_16565_, _03813_, _16543_);
  and (_16566_, _04612_, \oc8051_golden_model_1.ACC [0]);
  or (_16567_, _16566_, _16546_);
  and (_16568_, _16567_, _03813_);
  or (_16570_, _16568_, _16565_);
  and (_16571_, _16570_, _03810_);
  or (_16572_, _16571_, _03069_);
  or (_16573_, _16572_, _16564_);
  and (_16574_, _16573_, _16562_);
  or (_16575_, _16574_, _03075_);
  or (_16576_, _16567_, _03084_);
  and (_16577_, _16576_, _08225_);
  and (_16578_, _16577_, _16575_);
  or (_16579_, _16578_, _16559_);
  and (_16581_, _16579_, _08209_);
  nor (_16582_, _03486_, _08209_);
  or (_16583_, _16582_, _06770_);
  or (_16584_, _16583_, _16581_);
  or (_16585_, _16561_, _05535_);
  and (_16586_, _16585_, _05540_);
  and (_16587_, _16586_, _16584_);
  or (_16588_, _16587_, _02579_);
  or (_16589_, _16588_, _16557_);
  nor (_16590_, _11505_, _08251_);
  or (_16592_, _16546_, _02838_);
  or (_16593_, _16592_, _16590_);
  and (_16594_, _16593_, _02803_);
  and (_16595_, _16594_, _16589_);
  and (_16596_, _16549_, _02802_);
  or (_16597_, _16596_, _02980_);
  or (_16598_, _16597_, _16595_);
  and (_16599_, _11399_, _04612_);
  or (_16600_, _16546_, _03887_);
  or (_16601_, _16600_, _16599_);
  and (_16603_, _16601_, _03128_);
  and (_16604_, _16603_, _16598_);
  or (_16605_, _16604_, _16554_);
  and (_16606_, _16605_, _03883_);
  or (_16607_, _16606_, _16551_);
  and (_16608_, _16607_, _03137_);
  or (_16609_, _16546_, _09409_);
  and (_16610_, _16567_, _03135_);
  and (_16611_, _16610_, _16609_);
  or (_16612_, _16611_, _02965_);
  or (_16614_, _16612_, _16608_);
  nor (_16615_, _11396_, _08251_);
  or (_16616_, _16546_, _05783_);
  or (_16617_, _16616_, _16615_);
  and (_16618_, _16617_, _05788_);
  and (_16619_, _16618_, _16614_);
  nor (_16620_, _11520_, _08251_);
  or (_16621_, _16620_, _16546_);
  and (_16622_, _16621_, _03123_);
  nor (_16623_, _03163_, _02888_);
  not (_16625_, _16623_);
  or (_16626_, _16625_, _16622_);
  or (_16627_, _16626_, _16619_);
  or (_16628_, _16623_, _16563_);
  and (_16629_, _16628_, _42668_);
  and (_16630_, _16629_, _16627_);
  or (_16631_, _16630_, _16544_);
  and (_43430_, _16631_, _43998_);
  not (_16632_, \oc8051_golden_model_1.DPL [1]);
  nor (_16633_, _42668_, _16632_);
  or (_16635_, _11715_, _08251_);
  or (_16636_, _04612_, \oc8051_golden_model_1.DPL [1]);
  and (_16637_, _16636_, _03127_);
  and (_16638_, _16637_, _16635_);
  nand (_16639_, _11695_, _04612_);
  and (_16640_, _16636_, _02579_);
  and (_16641_, _16640_, _16639_);
  nor (_16642_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_16643_, _16642_, _08229_);
  and (_16644_, _16643_, _08224_);
  and (_16646_, _11606_, _04612_);
  not (_16647_, _16646_);
  and (_16648_, _16647_, _16636_);
  or (_16649_, _16648_, _03810_);
  nand (_16650_, _04612_, _02551_);
  and (_16651_, _16650_, _16636_);
  and (_16652_, _16651_, _03813_);
  nor (_16653_, _03813_, _16632_);
  or (_16654_, _16653_, _02974_);
  or (_16655_, _16654_, _16652_);
  and (_16657_, _16655_, _03336_);
  and (_16658_, _16657_, _16649_);
  nor (_16659_, _04612_, _16632_);
  and (_16660_, _04612_, _04000_);
  or (_16661_, _16660_, _16659_);
  and (_16662_, _16661_, _03069_);
  or (_16663_, _16662_, _03075_);
  or (_16664_, _16663_, _16658_);
  or (_16665_, _16651_, _03084_);
  and (_16666_, _16665_, _08225_);
  and (_16668_, _16666_, _16664_);
  or (_16669_, _16668_, _16644_);
  and (_16670_, _16669_, _08209_);
  nor (_16671_, _03698_, _08209_);
  or (_16672_, _16671_, _06770_);
  or (_16673_, _16672_, _16670_);
  or (_16674_, _16661_, _05535_);
  and (_16675_, _16674_, _16673_);
  or (_16676_, _16675_, _02853_);
  and (_16677_, _04612_, _06151_);
  or (_16679_, _16659_, _05540_);
  or (_16680_, _16679_, _16677_);
  and (_16681_, _16680_, _02838_);
  and (_16682_, _16681_, _16676_);
  or (_16683_, _16682_, _16641_);
  and (_16684_, _16683_, _02803_);
  nand (_16685_, _04612_, _03698_);
  and (_16686_, _16636_, _02802_);
  and (_16687_, _16686_, _16685_);
  or (_16688_, _16687_, _16684_);
  and (_16691_, _16688_, _03887_);
  or (_16692_, _11710_, _08251_);
  and (_16693_, _16636_, _02980_);
  and (_16694_, _16693_, _16692_);
  or (_16695_, _16694_, _16691_);
  and (_16696_, _16695_, _03128_);
  or (_16697_, _16696_, _16638_);
  and (_16698_, _16697_, _03883_);
  or (_16699_, _11709_, _08251_);
  and (_16700_, _16636_, _02970_);
  and (_16702_, _16700_, _16699_);
  or (_16703_, _16702_, _16698_);
  and (_16704_, _16703_, _03137_);
  or (_16705_, _16659_, _13722_);
  and (_16706_, _16651_, _03135_);
  and (_16707_, _16706_, _16705_);
  or (_16708_, _16707_, _16704_);
  and (_16709_, _16708_, _03124_);
  or (_16710_, _16650_, _13722_);
  and (_16711_, _16636_, _03123_);
  and (_16713_, _16711_, _16710_);
  or (_16714_, _16713_, _03163_);
  or (_16715_, _16685_, _13722_);
  and (_16716_, _16636_, _02965_);
  and (_16717_, _16716_, _16715_);
  or (_16718_, _16717_, _16714_);
  or (_16719_, _16718_, _16709_);
  or (_16720_, _16648_, _03906_);
  and (_16721_, _16720_, _16719_);
  or (_16722_, _16721_, _02888_);
  or (_16724_, _16659_, _02890_);
  or (_16725_, _16724_, _16646_);
  and (_16726_, _16725_, _42668_);
  and (_16727_, _16726_, _16722_);
  or (_16728_, _16727_, _16633_);
  and (_43431_, _16728_, _43998_);
  or (_16729_, _42668_, \oc8051_golden_model_1.DPL [2]);
  and (_16730_, _16729_, _43998_);
  not (_16731_, \oc8051_golden_model_1.DPL [2]);
  nor (_16732_, _04612_, _16731_);
  and (_16734_, _11927_, _04612_);
  or (_16735_, _16734_, _16732_);
  and (_16736_, _16735_, _03127_);
  and (_16737_, _04612_, _04435_);
  or (_16738_, _16737_, _16732_);
  or (_16739_, _16738_, _05535_);
  or (_16740_, _16738_, _03336_);
  nor (_16741_, _11801_, _08251_);
  or (_16742_, _16741_, _16732_);
  and (_16743_, _16742_, _02974_);
  nor (_16745_, _03813_, _16731_);
  and (_16746_, _04612_, \oc8051_golden_model_1.ACC [2]);
  or (_16747_, _16746_, _16732_);
  and (_16748_, _16747_, _03813_);
  or (_16749_, _16748_, _16745_);
  and (_16750_, _16749_, _03810_);
  or (_16751_, _16750_, _03069_);
  or (_16752_, _16751_, _16743_);
  and (_16753_, _16752_, _16740_);
  or (_16754_, _16753_, _03075_);
  or (_16756_, _16747_, _03084_);
  and (_16757_, _16756_, _08225_);
  and (_16758_, _16757_, _16754_);
  nor (_16759_, _08229_, \oc8051_golden_model_1.DPL [2]);
  nor (_16760_, _16759_, _08230_);
  and (_16761_, _16760_, _08224_);
  or (_16762_, _16761_, _16758_);
  and (_16763_, _16762_, _08209_);
  nor (_16764_, _03297_, _08209_);
  or (_16765_, _16764_, _06770_);
  or (_16767_, _16765_, _16763_);
  and (_16768_, _16767_, _16739_);
  or (_16769_, _16768_, _02853_);
  and (_16770_, _04612_, _06155_);
  or (_16771_, _16732_, _05540_);
  or (_16772_, _16771_, _16770_);
  and (_16773_, _16772_, _02838_);
  and (_16774_, _16773_, _16769_);
  nor (_16775_, _11906_, _08251_);
  or (_16776_, _16775_, _16732_);
  and (_16778_, _16776_, _02579_);
  or (_16779_, _16778_, _02802_);
  or (_16780_, _16779_, _16774_);
  and (_16781_, _04612_, _05701_);
  or (_16782_, _16781_, _16732_);
  or (_16783_, _16782_, _02803_);
  and (_16784_, _16783_, _16780_);
  or (_16785_, _16784_, _02980_);
  and (_16786_, _11921_, _04612_);
  or (_16787_, _16732_, _03887_);
  or (_16789_, _16787_, _16786_);
  and (_16790_, _16789_, _03128_);
  and (_16791_, _16790_, _16785_);
  or (_16792_, _16791_, _16736_);
  and (_16793_, _16792_, _03883_);
  or (_16794_, _16732_, _05130_);
  and (_16795_, _16782_, _02970_);
  and (_16796_, _16795_, _16794_);
  or (_16797_, _16796_, _16793_);
  and (_16798_, _16797_, _03137_);
  and (_16800_, _16747_, _03135_);
  and (_16801_, _16800_, _16794_);
  or (_16802_, _16801_, _02965_);
  or (_16803_, _16802_, _16798_);
  nor (_16804_, _11919_, _08251_);
  or (_16805_, _16732_, _05783_);
  or (_16806_, _16805_, _16804_);
  and (_16807_, _16806_, _05788_);
  and (_16808_, _16807_, _16803_);
  nor (_16809_, _11926_, _08251_);
  or (_16811_, _16809_, _16732_);
  and (_16812_, _16811_, _03123_);
  or (_16813_, _16812_, _03163_);
  or (_16814_, _16813_, _16808_);
  or (_16815_, _16742_, _03906_);
  and (_16816_, _16815_, _02890_);
  and (_16817_, _16816_, _16814_);
  and (_16818_, _11985_, _04612_);
  or (_16819_, _16818_, _16732_);
  and (_16820_, _16819_, _02888_);
  or (_16822_, _16820_, _42672_);
  or (_16823_, _16822_, _16817_);
  and (_43432_, _16823_, _16730_);
  or (_16824_, _42668_, \oc8051_golden_model_1.DPL [3]);
  and (_16825_, _16824_, _43998_);
  and (_16826_, _08251_, \oc8051_golden_model_1.DPL [3]);
  and (_16827_, _12133_, _04612_);
  or (_16828_, _16827_, _16826_);
  and (_16829_, _16828_, _03127_);
  and (_16830_, _04612_, _04241_);
  or (_16832_, _16830_, _16826_);
  or (_16833_, _16832_, _05535_);
  nor (_16834_, _08230_, \oc8051_golden_model_1.DPL [3]);
  nor (_16835_, _16834_, _08231_);
  and (_16836_, _16835_, _08224_);
  nor (_16837_, _12017_, _08251_);
  or (_16838_, _16837_, _16826_);
  or (_16839_, _16838_, _03810_);
  and (_16840_, _04612_, \oc8051_golden_model_1.ACC [3]);
  or (_16841_, _16840_, _16826_);
  and (_16843_, _16841_, _03813_);
  and (_16844_, _03814_, \oc8051_golden_model_1.DPL [3]);
  or (_16845_, _16844_, _02974_);
  or (_16846_, _16845_, _16843_);
  and (_16847_, _16846_, _03336_);
  and (_16848_, _16847_, _16839_);
  and (_16849_, _16832_, _03069_);
  or (_16850_, _16849_, _03075_);
  or (_16851_, _16850_, _16848_);
  or (_16852_, _16841_, _03084_);
  and (_16854_, _16852_, _08225_);
  and (_16855_, _16854_, _16851_);
  or (_16856_, _16855_, _16836_);
  and (_16857_, _16856_, _08209_);
  nor (_16858_, _03057_, _08209_);
  or (_16859_, _16858_, _06770_);
  or (_16860_, _16859_, _16857_);
  and (_16861_, _16860_, _16833_);
  or (_16862_, _16861_, _02853_);
  and (_16863_, _04612_, _06154_);
  or (_16865_, _16826_, _05540_);
  or (_16866_, _16865_, _16863_);
  and (_16867_, _16866_, _02838_);
  and (_16868_, _16867_, _16862_);
  nor (_16869_, _12112_, _08251_);
  or (_16870_, _16869_, _16826_);
  and (_16871_, _16870_, _02579_);
  or (_16872_, _16871_, _02802_);
  or (_16873_, _16872_, _16868_);
  and (_16874_, _04612_, _05658_);
  or (_16876_, _16874_, _16826_);
  or (_16877_, _16876_, _02803_);
  and (_16878_, _16877_, _16873_);
  or (_16879_, _16878_, _02980_);
  and (_16880_, _12127_, _04612_);
  or (_16881_, _16826_, _03887_);
  or (_16882_, _16881_, _16880_);
  and (_16883_, _16882_, _03128_);
  and (_16884_, _16883_, _16879_);
  or (_16885_, _16884_, _16829_);
  and (_16887_, _16885_, _03883_);
  or (_16888_, _16826_, _05079_);
  and (_16889_, _16876_, _02970_);
  and (_16890_, _16889_, _16888_);
  or (_16891_, _16890_, _16887_);
  and (_16892_, _16891_, _03137_);
  and (_16893_, _16841_, _03135_);
  and (_16894_, _16893_, _16888_);
  or (_16895_, _16894_, _02965_);
  or (_16896_, _16895_, _16892_);
  nor (_16898_, _12125_, _08251_);
  or (_16899_, _16826_, _05783_);
  or (_16900_, _16899_, _16898_);
  and (_16901_, _16900_, _05788_);
  and (_16902_, _16901_, _16896_);
  nor (_16903_, _12132_, _08251_);
  or (_16904_, _16903_, _16826_);
  and (_16905_, _16904_, _03123_);
  or (_16906_, _16905_, _03163_);
  or (_16907_, _16906_, _16902_);
  or (_16909_, _16838_, _03906_);
  and (_16910_, _16909_, _02890_);
  and (_16911_, _16910_, _16907_);
  and (_16912_, _12183_, _04612_);
  or (_16913_, _16912_, _16826_);
  and (_16914_, _16913_, _02888_);
  or (_16915_, _16914_, _42672_);
  or (_16916_, _16915_, _16911_);
  and (_43433_, _16916_, _16825_);
  or (_16917_, _42668_, \oc8051_golden_model_1.DPL [4]);
  and (_16919_, _16917_, _43998_);
  and (_16920_, _08251_, \oc8051_golden_model_1.DPL [4]);
  and (_16921_, _12207_, _04612_);
  or (_16922_, _16921_, _16920_);
  and (_16923_, _16922_, _03127_);
  and (_16924_, _04612_, _04982_);
  or (_16925_, _16924_, _16920_);
  or (_16926_, _16925_, _05535_);
  nor (_16927_, _12217_, _08251_);
  or (_16928_, _16927_, _16920_);
  or (_16930_, _16928_, _03810_);
  and (_16931_, _04612_, \oc8051_golden_model_1.ACC [4]);
  or (_16932_, _16931_, _16920_);
  and (_16933_, _16932_, _03813_);
  and (_16934_, _03814_, \oc8051_golden_model_1.DPL [4]);
  or (_16935_, _16934_, _02974_);
  or (_16936_, _16935_, _16933_);
  and (_16937_, _16936_, _03336_);
  and (_16938_, _16937_, _16930_);
  and (_16939_, _16925_, _03069_);
  or (_16941_, _16939_, _03075_);
  or (_16942_, _16941_, _16938_);
  or (_16943_, _16932_, _03084_);
  and (_16944_, _16943_, _08225_);
  and (_16945_, _16944_, _16942_);
  nor (_16946_, _08231_, \oc8051_golden_model_1.DPL [4]);
  nor (_16947_, _16946_, _08232_);
  and (_16948_, _16947_, _08224_);
  or (_16949_, _16948_, _16945_);
  and (_16950_, _16949_, _08209_);
  nor (_16952_, _05582_, _08209_);
  or (_16953_, _16952_, _06770_);
  or (_16954_, _16953_, _16950_);
  and (_16955_, _16954_, _16926_);
  or (_16956_, _16955_, _02853_);
  and (_16957_, _04612_, _06159_);
  or (_16958_, _16920_, _05540_);
  or (_16959_, _16958_, _16957_);
  and (_16960_, _16959_, _02838_);
  and (_16961_, _16960_, _16956_);
  nor (_16963_, _12321_, _08251_);
  or (_16964_, _16963_, _16920_);
  and (_16965_, _16964_, _02579_);
  or (_16966_, _16965_, _02802_);
  or (_16967_, _16966_, _16961_);
  and (_16968_, _05666_, _04612_);
  or (_16969_, _16968_, _16920_);
  or (_16970_, _16969_, _02803_);
  and (_16971_, _16970_, _16967_);
  or (_16972_, _16971_, _02980_);
  and (_16974_, _12211_, _04612_);
  or (_16975_, _16920_, _03887_);
  or (_16976_, _16975_, _16974_);
  and (_16977_, _16976_, _03128_);
  and (_16978_, _16977_, _16972_);
  or (_16979_, _16978_, _16923_);
  and (_16980_, _16979_, _03883_);
  or (_16981_, _16920_, _05031_);
  and (_16982_, _16969_, _02970_);
  and (_16983_, _16982_, _16981_);
  or (_16985_, _16983_, _16980_);
  and (_16986_, _16985_, _03137_);
  and (_16987_, _16932_, _03135_);
  and (_16988_, _16987_, _16981_);
  or (_16989_, _16988_, _02965_);
  or (_16990_, _16989_, _16986_);
  nor (_16991_, _12209_, _08251_);
  or (_16992_, _16920_, _05783_);
  or (_16993_, _16992_, _16991_);
  and (_16994_, _16993_, _05788_);
  and (_16996_, _16994_, _16990_);
  nor (_16997_, _12206_, _08251_);
  or (_16998_, _16997_, _16920_);
  and (_16999_, _16998_, _03123_);
  or (_17000_, _16999_, _03163_);
  or (_17001_, _17000_, _16996_);
  or (_17002_, _16928_, _03906_);
  and (_17003_, _17002_, _02890_);
  and (_17004_, _17003_, _17001_);
  and (_17005_, _12389_, _04612_);
  or (_17007_, _17005_, _16920_);
  and (_17008_, _17007_, _02888_);
  or (_17009_, _17008_, _42672_);
  or (_17010_, _17009_, _17004_);
  and (_43434_, _17010_, _16919_);
  or (_17011_, _42668_, \oc8051_golden_model_1.DPL [5]);
  and (_17012_, _17011_, _43998_);
  and (_17013_, _08251_, \oc8051_golden_model_1.DPL [5]);
  and (_17014_, _12411_, _04612_);
  or (_17015_, _17014_, _17013_);
  and (_17017_, _17015_, _03127_);
  and (_17018_, _04612_, _04877_);
  or (_17019_, _17018_, _17013_);
  or (_17020_, _17019_, _05535_);
  nor (_17021_, _12407_, _08251_);
  or (_17022_, _17021_, _17013_);
  or (_17023_, _17022_, _03810_);
  and (_17024_, _04612_, \oc8051_golden_model_1.ACC [5]);
  or (_17025_, _17024_, _17013_);
  and (_17026_, _17025_, _03813_);
  and (_17028_, _03814_, \oc8051_golden_model_1.DPL [5]);
  or (_17029_, _17028_, _02974_);
  or (_17030_, _17029_, _17026_);
  and (_17031_, _17030_, _03336_);
  and (_17032_, _17031_, _17023_);
  and (_17033_, _17019_, _03069_);
  or (_17034_, _17033_, _03075_);
  or (_17035_, _17034_, _17032_);
  or (_17036_, _17025_, _03084_);
  and (_17037_, _17036_, _08225_);
  and (_17039_, _17037_, _17035_);
  nor (_17040_, _08232_, \oc8051_golden_model_1.DPL [5]);
  nor (_17041_, _17040_, _08233_);
  and (_17042_, _17041_, _08224_);
  or (_17043_, _17042_, _17039_);
  and (_17044_, _17043_, _08209_);
  nor (_17045_, _05613_, _08209_);
  or (_17046_, _17045_, _06770_);
  or (_17047_, _17046_, _17044_);
  and (_17048_, _17047_, _17020_);
  or (_17050_, _17048_, _02853_);
  and (_17051_, _04612_, _06158_);
  or (_17052_, _17013_, _05540_);
  or (_17053_, _17052_, _17051_);
  and (_17054_, _17053_, _02838_);
  and (_17055_, _17054_, _17050_);
  nor (_17056_, _12527_, _08251_);
  or (_17057_, _17056_, _17013_);
  and (_17058_, _17057_, _02579_);
  or (_17059_, _17058_, _02802_);
  or (_17061_, _17059_, _17055_);
  and (_17062_, _05614_, _04612_);
  or (_17063_, _17062_, _17013_);
  or (_17064_, _17063_, _02803_);
  and (_17065_, _17064_, _17061_);
  or (_17066_, _17065_, _02980_);
  and (_17067_, _12415_, _04612_);
  or (_17068_, _17013_, _03887_);
  or (_17069_, _17068_, _17067_);
  and (_17070_, _17069_, _03128_);
  and (_17072_, _17070_, _17066_);
  or (_17073_, _17072_, _17017_);
  and (_17074_, _17073_, _03883_);
  or (_17075_, _17013_, _04924_);
  and (_17076_, _17063_, _02970_);
  and (_17077_, _17076_, _17075_);
  or (_17078_, _17077_, _17074_);
  and (_17079_, _17078_, _03137_);
  and (_17080_, _17025_, _03135_);
  and (_17081_, _17080_, _17075_);
  or (_17083_, _17081_, _02965_);
  or (_17084_, _17083_, _17079_);
  nor (_17085_, _12413_, _08251_);
  or (_17086_, _17013_, _05783_);
  or (_17087_, _17086_, _17085_);
  and (_17088_, _17087_, _05788_);
  and (_17089_, _17088_, _17084_);
  nor (_17090_, _12410_, _08251_);
  or (_17091_, _17090_, _17013_);
  and (_17092_, _17091_, _03123_);
  or (_17094_, _17092_, _03163_);
  or (_17095_, _17094_, _17089_);
  or (_17096_, _17022_, _03906_);
  and (_17097_, _17096_, _02890_);
  and (_17098_, _17097_, _17095_);
  and (_17099_, _12589_, _04612_);
  or (_17100_, _17099_, _17013_);
  and (_17101_, _17100_, _02888_);
  or (_17102_, _17101_, _42672_);
  or (_17103_, _17102_, _17098_);
  and (_43435_, _17103_, _17012_);
  or (_17105_, _42668_, \oc8051_golden_model_1.DPL [6]);
  and (_17106_, _17105_, _43998_);
  not (_17107_, \oc8051_golden_model_1.DPL [6]);
  nor (_17108_, _04612_, _17107_);
  and (_17109_, _12613_, _04612_);
  or (_17110_, _17109_, _17108_);
  and (_17111_, _17110_, _03127_);
  and (_17112_, _04612_, _04770_);
  or (_17113_, _17112_, _17108_);
  or (_17115_, _17113_, _05535_);
  nor (_17116_, _12603_, _08251_);
  or (_17117_, _17116_, _17108_);
  or (_17118_, _17117_, _03810_);
  and (_17119_, _04612_, \oc8051_golden_model_1.ACC [6]);
  or (_17120_, _17119_, _17108_);
  and (_17121_, _17120_, _03813_);
  nor (_17122_, _03813_, _17107_);
  or (_17123_, _17122_, _02974_);
  or (_17124_, _17123_, _17121_);
  and (_17126_, _17124_, _03336_);
  and (_17127_, _17126_, _17118_);
  and (_17128_, _17113_, _03069_);
  or (_17129_, _17128_, _03075_);
  or (_17130_, _17129_, _17127_);
  or (_17131_, _17120_, _03084_);
  and (_17132_, _17131_, _08225_);
  and (_17133_, _17132_, _17130_);
  nor (_17134_, _08233_, \oc8051_golden_model_1.DPL [6]);
  nor (_17135_, _17134_, _08234_);
  and (_17137_, _17135_, _08224_);
  or (_17138_, _17137_, _17133_);
  and (_17139_, _17138_, _08209_);
  nor (_17140_, _05649_, _08209_);
  or (_17141_, _17140_, _06770_);
  or (_17142_, _17141_, _17139_);
  and (_17143_, _17142_, _17115_);
  or (_17144_, _17143_, _02853_);
  and (_17145_, _04612_, _05849_);
  or (_17146_, _17108_, _05540_);
  or (_17148_, _17146_, _17145_);
  and (_17149_, _17148_, _02838_);
  and (_17150_, _17149_, _17144_);
  nor (_17151_, _12722_, _08251_);
  or (_17152_, _17151_, _17108_);
  and (_17153_, _17152_, _02579_);
  or (_17154_, _17153_, _02802_);
  or (_17155_, _17154_, _17150_);
  and (_17156_, _12729_, _04612_);
  or (_17157_, _17156_, _17108_);
  or (_17159_, _17157_, _02803_);
  and (_17160_, _17159_, _17155_);
  or (_17161_, _17160_, _02980_);
  and (_17162_, _12739_, _04612_);
  or (_17163_, _17108_, _03887_);
  or (_17164_, _17163_, _17162_);
  and (_17165_, _17164_, _03128_);
  and (_17166_, _17165_, _17161_);
  or (_17167_, _17166_, _17111_);
  and (_17168_, _17167_, _03883_);
  or (_17170_, _17108_, _04819_);
  and (_17171_, _17157_, _02970_);
  and (_17172_, _17171_, _17170_);
  or (_17173_, _17172_, _17168_);
  and (_17174_, _17173_, _03137_);
  and (_17175_, _17120_, _03135_);
  and (_17176_, _17175_, _17170_);
  or (_17177_, _17176_, _02965_);
  or (_17178_, _17177_, _17174_);
  nor (_17179_, _12737_, _08251_);
  or (_17181_, _17108_, _05783_);
  or (_17182_, _17181_, _17179_);
  and (_17183_, _17182_, _05788_);
  and (_17184_, _17183_, _17178_);
  nor (_17185_, _12612_, _08251_);
  or (_17186_, _17185_, _17108_);
  and (_17187_, _17186_, _03123_);
  or (_17188_, _17187_, _03163_);
  or (_17189_, _17188_, _17184_);
  or (_17190_, _17117_, _03906_);
  and (_17192_, _17190_, _02890_);
  and (_17193_, _17192_, _17189_);
  and (_17194_, _12794_, _04612_);
  or (_17195_, _17194_, _17108_);
  and (_17196_, _17195_, _02888_);
  or (_17197_, _17196_, _42672_);
  or (_17198_, _17197_, _17193_);
  and (_43436_, _17198_, _17106_);
  not (_17199_, \oc8051_golden_model_1.DPH [0]);
  nor (_17200_, _42668_, _17199_);
  nor (_17202_, _04783_, _17199_);
  and (_17203_, _05226_, _04671_);
  or (_17204_, _17203_, _17202_);
  or (_17205_, _17204_, _03810_);
  and (_17206_, _04783_, \oc8051_golden_model_1.ACC [0]);
  or (_17207_, _17206_, _17202_);
  and (_17208_, _17207_, _03813_);
  nor (_17209_, _03813_, _17199_);
  or (_17210_, _17209_, _02974_);
  or (_17211_, _17210_, _17208_);
  and (_17213_, _17211_, _03336_);
  and (_17214_, _17213_, _17205_);
  and (_17215_, _04671_, _03808_);
  or (_17216_, _17215_, _17202_);
  and (_17217_, _17216_, _03069_);
  or (_17218_, _17217_, _03075_);
  or (_17219_, _17218_, _17214_);
  or (_17220_, _17207_, _03084_);
  and (_17221_, _17220_, _08225_);
  and (_17222_, _17221_, _17219_);
  nor (_17224_, _08236_, \oc8051_golden_model_1.DPH [0]);
  nor (_17225_, _17224_, _08323_);
  and (_17226_, _17225_, _08224_);
  or (_17227_, _17226_, _17222_);
  and (_17228_, _17227_, _08209_);
  and (_17229_, _02835_, _02981_);
  or (_17230_, _17229_, _06770_);
  or (_17231_, _17230_, _17228_);
  or (_17232_, _17216_, _05535_);
  and (_17233_, _17232_, _17231_);
  or (_17235_, _17233_, _02853_);
  and (_17236_, _04783_, _06152_);
  or (_17237_, _17202_, _05540_);
  or (_17238_, _17237_, _17236_);
  and (_17239_, _17238_, _17235_);
  or (_17240_, _17239_, _02579_);
  nor (_17241_, _11505_, _08373_);
  or (_17242_, _17202_, _02838_);
  or (_17243_, _17242_, _17241_);
  and (_17244_, _17243_, _02803_);
  and (_17246_, _17244_, _17240_);
  and (_17247_, _04783_, _05672_);
  or (_17248_, _17247_, _17202_);
  and (_17249_, _17248_, _02802_);
  or (_17250_, _17249_, _02980_);
  or (_17251_, _17250_, _17246_);
  and (_17252_, _11399_, _04783_);
  or (_17253_, _17252_, _17202_);
  or (_17254_, _17253_, _03887_);
  and (_17255_, _17254_, _17251_);
  or (_17257_, _17255_, _03127_);
  and (_17258_, _11522_, _04671_);
  or (_17259_, _17202_, _03128_);
  or (_17260_, _17259_, _17258_);
  and (_17261_, _17260_, _03883_);
  and (_17262_, _17261_, _17257_);
  nand (_17263_, _17248_, _02970_);
  nor (_17264_, _17263_, _17203_);
  or (_17265_, _17264_, _17262_);
  and (_17266_, _17265_, _03137_);
  or (_17268_, _17202_, _09409_);
  and (_17269_, _17207_, _03135_);
  and (_17270_, _17269_, _17268_);
  or (_17271_, _17270_, _02965_);
  or (_17272_, _17271_, _17266_);
  nor (_17273_, _11396_, _08346_);
  or (_17274_, _17273_, _17202_);
  or (_17275_, _17274_, _05783_);
  and (_17276_, _17275_, _05788_);
  and (_17277_, _17276_, _17272_);
  nor (_17279_, _11520_, _08373_);
  or (_17280_, _17279_, _17202_);
  and (_17281_, _17280_, _03123_);
  or (_17282_, _17281_, _16625_);
  or (_17283_, _17282_, _17277_);
  or (_17284_, _17204_, _16623_);
  and (_17285_, _17284_, _42668_);
  and (_17286_, _17285_, _17283_);
  or (_17287_, _17286_, _17200_);
  and (_43438_, _17287_, _43998_);
  not (_17289_, \oc8051_golden_model_1.DPH [1]);
  nor (_17290_, _42668_, _17289_);
  or (_17291_, _11715_, _08373_);
  or (_17292_, _04783_, \oc8051_golden_model_1.DPH [1]);
  and (_17293_, _17292_, _03127_);
  and (_17294_, _17293_, _17291_);
  and (_17295_, _17292_, _02802_);
  nand (_17296_, _04671_, _03698_);
  and (_17297_, _17296_, _17295_);
  nor (_17298_, _08323_, \oc8051_golden_model_1.DPH [1]);
  nor (_17300_, _17298_, _08324_);
  and (_17301_, _17300_, _08224_);
  nand (_17302_, _11606_, _04671_);
  and (_17303_, _17302_, _17292_);
  or (_17304_, _17303_, _03810_);
  nand (_17305_, _04671_, _02551_);
  and (_17306_, _17305_, _17292_);
  and (_17307_, _17306_, _03813_);
  nor (_17308_, _03813_, _17289_);
  or (_17309_, _17308_, _02974_);
  or (_17311_, _17309_, _17307_);
  and (_17312_, _17311_, _03336_);
  and (_17313_, _17312_, _17304_);
  nor (_17314_, _04783_, _17289_);
  and (_17315_, _04671_, _04000_);
  or (_17316_, _17315_, _17314_);
  and (_17317_, _17316_, _03069_);
  or (_17318_, _17317_, _03075_);
  or (_17319_, _17318_, _17313_);
  or (_17320_, _17306_, _03084_);
  and (_17322_, _17320_, _08225_);
  and (_17323_, _17322_, _17319_);
  or (_17324_, _17323_, _17301_);
  and (_17325_, _17324_, _08209_);
  nor (_17326_, _08209_, _03665_);
  or (_17327_, _17326_, _06770_);
  or (_17328_, _17327_, _17325_);
  or (_17329_, _17316_, _05535_);
  and (_17330_, _17329_, _17328_);
  or (_17331_, _17330_, _02853_);
  and (_17333_, _04783_, _06151_);
  or (_17334_, _17314_, _05540_);
  or (_17335_, _17334_, _17333_);
  and (_17336_, _17335_, _02838_);
  and (_17337_, _17336_, _17331_);
  and (_17338_, _17292_, _02579_);
  nand (_17339_, _11695_, _04671_);
  and (_17340_, _17339_, _17338_);
  or (_17341_, _17340_, _17337_);
  and (_17342_, _17341_, _02803_);
  or (_17344_, _17342_, _17297_);
  and (_17345_, _17344_, _03887_);
  or (_17346_, _11710_, _08373_);
  and (_17347_, _17292_, _02980_);
  and (_17348_, _17347_, _17346_);
  or (_17349_, _17348_, _17345_);
  and (_17350_, _17349_, _03128_);
  or (_17351_, _17350_, _17294_);
  and (_17352_, _17351_, _03883_);
  or (_17353_, _11709_, _08373_);
  and (_17355_, _17292_, _02970_);
  and (_17356_, _17355_, _17353_);
  or (_17357_, _17356_, _17352_);
  and (_17358_, _17357_, _03137_);
  or (_17359_, _17314_, _13722_);
  and (_17360_, _17306_, _03135_);
  and (_17361_, _17360_, _17359_);
  or (_17362_, _17361_, _17358_);
  and (_17363_, _17362_, _03124_);
  or (_17364_, _17305_, _13722_);
  and (_17366_, _17292_, _03123_);
  and (_17367_, _17366_, _17364_);
  or (_17368_, _17367_, _03163_);
  or (_17369_, _17296_, _13722_);
  and (_17370_, _17292_, _02965_);
  and (_17371_, _17370_, _17369_);
  or (_17372_, _17371_, _17368_);
  or (_17373_, _17372_, _17363_);
  or (_17374_, _17303_, _03906_);
  and (_17375_, _17374_, _17373_);
  or (_17377_, _17375_, _02888_);
  nor (_17378_, _17314_, _02890_);
  nand (_17379_, _17378_, _17302_);
  and (_17380_, _17379_, _42668_);
  and (_17381_, _17380_, _17377_);
  or (_17382_, _17381_, _17290_);
  and (_43439_, _17382_, _43998_);
  or (_17383_, _42668_, \oc8051_golden_model_1.DPH [2]);
  and (_17384_, _17383_, _43998_);
  not (_17385_, \oc8051_golden_model_1.DPH [2]);
  nor (_17387_, _04783_, _17385_);
  and (_17388_, _11927_, _04671_);
  or (_17389_, _17388_, _17387_);
  and (_17390_, _17389_, _03127_);
  and (_17391_, _04671_, _04435_);
  or (_17392_, _17391_, _17387_);
  or (_17393_, _17392_, _05535_);
  or (_17394_, _17392_, _03336_);
  nor (_17395_, _11801_, _08373_);
  or (_17396_, _17395_, _17387_);
  and (_17397_, _17396_, _02974_);
  nor (_17398_, _03813_, _17385_);
  and (_17399_, _04783_, \oc8051_golden_model_1.ACC [2]);
  or (_17400_, _17399_, _17387_);
  and (_17401_, _17400_, _03813_);
  or (_17402_, _17401_, _17398_);
  and (_17403_, _17402_, _03810_);
  or (_17404_, _17403_, _03069_);
  or (_17405_, _17404_, _17397_);
  and (_17406_, _17405_, _17394_);
  or (_17409_, _17406_, _03075_);
  or (_17410_, _17400_, _03084_);
  and (_17411_, _17410_, _08225_);
  and (_17412_, _17411_, _17409_);
  or (_17413_, _08324_, \oc8051_golden_model_1.DPH [2]);
  nor (_17414_, _08325_, _08225_);
  and (_17415_, _17414_, _17413_);
  or (_17416_, _17415_, _17412_);
  and (_17417_, _17416_, _08209_);
  nor (_17418_, _03256_, _08209_);
  or (_17419_, _17418_, _06770_);
  or (_17420_, _17419_, _17417_);
  and (_17421_, _17420_, _17393_);
  or (_17422_, _17421_, _02853_);
  or (_17423_, _17387_, _05540_);
  and (_17424_, _04783_, _06155_);
  or (_17425_, _17424_, _17423_);
  and (_17426_, _17425_, _02838_);
  and (_17427_, _17426_, _17422_);
  nor (_17428_, _11906_, _08346_);
  or (_17431_, _17428_, _17387_);
  and (_17432_, _17431_, _02579_);
  or (_17433_, _17432_, _02802_);
  or (_17434_, _17433_, _17427_);
  and (_17435_, _04783_, _05701_);
  or (_17436_, _17435_, _17387_);
  or (_17437_, _17436_, _02803_);
  and (_17438_, _17437_, _17434_);
  or (_17439_, _17438_, _02980_);
  and (_17440_, _11921_, _04671_);
  or (_17442_, _17387_, _03887_);
  or (_17443_, _17442_, _17440_);
  and (_17444_, _17443_, _03128_);
  and (_17445_, _17444_, _17439_);
  or (_17446_, _17445_, _17390_);
  and (_17447_, _17446_, _03883_);
  or (_17448_, _17387_, _05130_);
  and (_17449_, _17436_, _02970_);
  and (_17450_, _17449_, _17448_);
  or (_17451_, _17450_, _17447_);
  and (_17453_, _17451_, _03137_);
  and (_17454_, _17400_, _03135_);
  and (_17455_, _17454_, _17448_);
  or (_17456_, _17455_, _02965_);
  or (_17457_, _17456_, _17453_);
  nor (_17458_, _11919_, _08373_);
  or (_17459_, _17387_, _05783_);
  or (_17460_, _17459_, _17458_);
  and (_17461_, _17460_, _05788_);
  and (_17462_, _17461_, _17457_);
  nor (_17464_, _11926_, _08373_);
  or (_17465_, _17464_, _17387_);
  and (_17466_, _17465_, _03123_);
  or (_17467_, _17466_, _03163_);
  or (_17468_, _17467_, _17462_);
  or (_17469_, _17396_, _03906_);
  and (_17470_, _17469_, _02890_);
  and (_17471_, _17470_, _17468_);
  and (_17472_, _11985_, _04671_);
  or (_17473_, _17472_, _17387_);
  and (_17475_, _17473_, _02888_);
  or (_17476_, _17475_, _42672_);
  or (_17477_, _17476_, _17471_);
  and (_43440_, _17477_, _17384_);
  or (_17478_, _42668_, \oc8051_golden_model_1.DPH [3]);
  and (_17479_, _17478_, _43998_);
  and (_17480_, _08346_, \oc8051_golden_model_1.DPH [3]);
  and (_17481_, _12133_, _04671_);
  or (_17482_, _17481_, _17480_);
  and (_17483_, _17482_, _03127_);
  and (_17485_, _04671_, _04241_);
  or (_17486_, _17485_, _17480_);
  or (_17487_, _17486_, _05535_);
  or (_17488_, _08325_, \oc8051_golden_model_1.DPH [3]);
  nor (_17489_, _08326_, _08225_);
  and (_17490_, _17489_, _17488_);
  nor (_17491_, _12017_, _08373_);
  or (_17492_, _17491_, _17480_);
  or (_17493_, _17492_, _03810_);
  and (_17494_, _04783_, \oc8051_golden_model_1.ACC [3]);
  or (_17496_, _17494_, _17480_);
  and (_17497_, _17496_, _03813_);
  and (_17498_, _03814_, \oc8051_golden_model_1.DPH [3]);
  or (_17499_, _17498_, _02974_);
  or (_17500_, _17499_, _17497_);
  and (_17501_, _17500_, _03336_);
  and (_17502_, _17501_, _17493_);
  and (_17503_, _17486_, _03069_);
  or (_17504_, _17503_, _03075_);
  or (_17505_, _17504_, _17502_);
  or (_17507_, _17496_, _03084_);
  and (_17508_, _17507_, _08225_);
  and (_17509_, _17508_, _17505_);
  or (_17510_, _17509_, _17490_);
  and (_17511_, _17510_, _08209_);
  nor (_17512_, _08209_, _02794_);
  or (_17513_, _17512_, _06770_);
  or (_17514_, _17513_, _17511_);
  and (_17515_, _17514_, _17487_);
  or (_17516_, _17515_, _02853_);
  or (_17518_, _17480_, _05540_);
  and (_17519_, _04783_, _06154_);
  or (_17520_, _17519_, _17518_);
  and (_17521_, _17520_, _02838_);
  and (_17522_, _17521_, _17516_);
  nor (_17523_, _12112_, _08346_);
  or (_17524_, _17523_, _17480_);
  and (_17525_, _17524_, _02579_);
  or (_17526_, _17525_, _02802_);
  or (_17527_, _17526_, _17522_);
  and (_17529_, _04783_, _05658_);
  or (_17530_, _17529_, _17480_);
  or (_17531_, _17530_, _02803_);
  and (_17532_, _17531_, _17527_);
  or (_17533_, _17532_, _02980_);
  and (_17534_, _12127_, _04671_);
  or (_17535_, _17480_, _03887_);
  or (_17536_, _17535_, _17534_);
  and (_17537_, _17536_, _03128_);
  and (_17538_, _17537_, _17533_);
  or (_17540_, _17538_, _17483_);
  and (_17541_, _17540_, _03883_);
  or (_17542_, _17480_, _05079_);
  and (_17543_, _17530_, _02970_);
  and (_17544_, _17543_, _17542_);
  or (_17545_, _17544_, _17541_);
  and (_17546_, _17545_, _03137_);
  and (_17547_, _17496_, _03135_);
  and (_17548_, _17547_, _17542_);
  or (_17549_, _17548_, _02965_);
  or (_17551_, _17549_, _17546_);
  nor (_17552_, _12125_, _08373_);
  or (_17553_, _17480_, _05783_);
  or (_17554_, _17553_, _17552_);
  and (_17555_, _17554_, _05788_);
  and (_17556_, _17555_, _17551_);
  nor (_17557_, _12132_, _08373_);
  or (_17558_, _17557_, _17480_);
  and (_17559_, _17558_, _03123_);
  or (_17560_, _17559_, _03163_);
  or (_17562_, _17560_, _17556_);
  or (_17563_, _17492_, _03906_);
  and (_17564_, _17563_, _02890_);
  and (_17565_, _17564_, _17562_);
  and (_17566_, _12183_, _04671_);
  or (_17567_, _17566_, _17480_);
  and (_17568_, _17567_, _02888_);
  or (_17569_, _17568_, _42672_);
  or (_17570_, _17569_, _17565_);
  and (_43441_, _17570_, _17479_);
  or (_17572_, _42668_, \oc8051_golden_model_1.DPH [4]);
  and (_17573_, _17572_, _43998_);
  and (_17574_, _08346_, \oc8051_golden_model_1.DPH [4]);
  and (_17575_, _12207_, _04671_);
  or (_17576_, _17575_, _17574_);
  and (_17577_, _17576_, _03127_);
  and (_17578_, _04671_, _04982_);
  or (_17579_, _17578_, _17574_);
  or (_17580_, _17579_, _05535_);
  nor (_17581_, _12217_, _08373_);
  or (_17583_, _17581_, _17574_);
  or (_17584_, _17583_, _03810_);
  and (_17585_, _04783_, \oc8051_golden_model_1.ACC [4]);
  or (_17586_, _17585_, _17574_);
  and (_17587_, _17586_, _03813_);
  and (_17588_, _03814_, \oc8051_golden_model_1.DPH [4]);
  or (_17589_, _17588_, _02974_);
  or (_17590_, _17589_, _17587_);
  and (_17591_, _17590_, _03336_);
  and (_17592_, _17591_, _17584_);
  and (_17594_, _17579_, _03069_);
  or (_17595_, _17594_, _03075_);
  or (_17596_, _17595_, _17592_);
  or (_17597_, _17586_, _03084_);
  and (_17598_, _17597_, _08225_);
  and (_17599_, _17598_, _17596_);
  or (_17600_, _08326_, \oc8051_golden_model_1.DPH [4]);
  nor (_17601_, _08327_, _08225_);
  and (_17602_, _17601_, _17600_);
  or (_17603_, _17602_, _17599_);
  and (_17605_, _17603_, _08209_);
  nor (_17606_, _08209_, _03629_);
  or (_17607_, _17606_, _06770_);
  or (_17608_, _17607_, _17605_);
  and (_17609_, _17608_, _17580_);
  or (_17610_, _17609_, _02853_);
  or (_17611_, _17574_, _05540_);
  and (_17612_, _04783_, _06159_);
  or (_17613_, _17612_, _17611_);
  and (_17614_, _17613_, _02838_);
  and (_17616_, _17614_, _17610_);
  nor (_17617_, _12321_, _08346_);
  or (_17618_, _17617_, _17574_);
  and (_17619_, _17618_, _02579_);
  or (_17620_, _17619_, _02802_);
  or (_17621_, _17620_, _17616_);
  and (_17622_, _05666_, _04783_);
  or (_17623_, _17622_, _17574_);
  or (_17624_, _17623_, _02803_);
  and (_17625_, _17624_, _17621_);
  or (_17627_, _17625_, _02980_);
  and (_17628_, _12211_, _04671_);
  or (_17629_, _17574_, _03887_);
  or (_17630_, _17629_, _17628_);
  and (_17631_, _17630_, _03128_);
  and (_17632_, _17631_, _17627_);
  or (_17633_, _17632_, _17577_);
  and (_17634_, _17633_, _03883_);
  or (_17635_, _17574_, _05031_);
  and (_17636_, _17623_, _02970_);
  and (_17638_, _17636_, _17635_);
  or (_17639_, _17638_, _17634_);
  and (_17640_, _17639_, _03137_);
  and (_17641_, _17586_, _03135_);
  and (_17642_, _17641_, _17635_);
  or (_17643_, _17642_, _02965_);
  or (_17644_, _17643_, _17640_);
  nor (_17645_, _12209_, _08373_);
  or (_17646_, _17574_, _05783_);
  or (_17647_, _17646_, _17645_);
  and (_17649_, _17647_, _05788_);
  and (_17650_, _17649_, _17644_);
  nor (_17651_, _12206_, _08373_);
  or (_17652_, _17651_, _17574_);
  and (_17653_, _17652_, _03123_);
  or (_17654_, _17653_, _03163_);
  or (_17655_, _17654_, _17650_);
  or (_17656_, _17583_, _03906_);
  and (_17657_, _17656_, _02890_);
  and (_17658_, _17657_, _17655_);
  and (_17660_, _12389_, _04671_);
  or (_17661_, _17660_, _17574_);
  and (_17662_, _17661_, _02888_);
  or (_17663_, _17662_, _42672_);
  or (_17664_, _17663_, _17658_);
  and (_43443_, _17664_, _17573_);
  or (_17665_, _42668_, \oc8051_golden_model_1.DPH [5]);
  and (_17666_, _17665_, _43998_);
  not (_17667_, \oc8051_golden_model_1.DPH [5]);
  nor (_17668_, _04783_, _17667_);
  and (_17670_, _12411_, _04671_);
  or (_17671_, _17670_, _17668_);
  and (_17672_, _17671_, _03127_);
  and (_17673_, _04671_, _04877_);
  or (_17674_, _17673_, _17668_);
  or (_17675_, _17674_, _05535_);
  nor (_17676_, _12407_, _08373_);
  or (_17677_, _17676_, _17668_);
  or (_17678_, _17677_, _03810_);
  and (_17679_, _04783_, \oc8051_golden_model_1.ACC [5]);
  or (_17681_, _17679_, _17668_);
  and (_17682_, _17681_, _03813_);
  nor (_17683_, _03813_, _17667_);
  or (_17684_, _17683_, _02974_);
  or (_17685_, _17684_, _17682_);
  and (_17686_, _17685_, _03336_);
  and (_17687_, _17686_, _17678_);
  and (_17688_, _17674_, _03069_);
  or (_17689_, _17688_, _03075_);
  or (_17690_, _17689_, _17687_);
  or (_17692_, _17681_, _03084_);
  and (_17693_, _17692_, _08225_);
  and (_17694_, _17693_, _17690_);
  or (_17695_, _08327_, \oc8051_golden_model_1.DPH [5]);
  nor (_17696_, _08328_, _08225_);
  and (_17697_, _17696_, _17695_);
  or (_17698_, _17697_, _17694_);
  and (_17699_, _17698_, _08209_);
  nor (_17700_, _03211_, _08209_);
  or (_17701_, _17700_, _06770_);
  or (_17703_, _17701_, _17699_);
  and (_17704_, _17703_, _17675_);
  or (_17705_, _17704_, _02853_);
  or (_17706_, _17668_, _05540_);
  and (_17707_, _04783_, _06158_);
  or (_17708_, _17707_, _17706_);
  and (_17709_, _17708_, _02838_);
  and (_17710_, _17709_, _17705_);
  nor (_17711_, _12527_, _08346_);
  or (_17712_, _17711_, _17668_);
  and (_17714_, _17712_, _02579_);
  or (_17715_, _17714_, _02802_);
  or (_17716_, _17715_, _17710_);
  and (_17717_, _05614_, _04783_);
  or (_17718_, _17717_, _17668_);
  or (_17719_, _17718_, _02803_);
  and (_17720_, _17719_, _17716_);
  or (_17721_, _17720_, _02980_);
  and (_17722_, _12415_, _04671_);
  or (_17723_, _17668_, _03887_);
  or (_17725_, _17723_, _17722_);
  and (_17726_, _17725_, _03128_);
  and (_17727_, _17726_, _17721_);
  or (_17728_, _17727_, _17672_);
  and (_17729_, _17728_, _03883_);
  or (_17730_, _17668_, _04924_);
  and (_17731_, _17718_, _02970_);
  and (_17732_, _17731_, _17730_);
  or (_17733_, _17732_, _17729_);
  and (_17734_, _17733_, _03137_);
  and (_17736_, _17681_, _03135_);
  and (_17737_, _17736_, _17730_);
  or (_17738_, _17737_, _02965_);
  or (_17739_, _17738_, _17734_);
  nor (_17740_, _12413_, _08373_);
  or (_17741_, _17668_, _05783_);
  or (_17742_, _17741_, _17740_);
  and (_17743_, _17742_, _05788_);
  and (_17744_, _17743_, _17739_);
  nor (_17745_, _12410_, _08373_);
  or (_17747_, _17745_, _17668_);
  and (_17748_, _17747_, _03123_);
  or (_17749_, _17748_, _03163_);
  or (_17750_, _17749_, _17744_);
  or (_17751_, _17677_, _03906_);
  and (_17752_, _17751_, _02890_);
  and (_17753_, _17752_, _17750_);
  and (_17754_, _12589_, _04671_);
  or (_17755_, _17754_, _17668_);
  and (_17756_, _17755_, _02888_);
  or (_17758_, _17756_, _42672_);
  or (_17759_, _17758_, _17753_);
  and (_43444_, _17759_, _17666_);
  or (_17760_, _42668_, \oc8051_golden_model_1.DPH [6]);
  and (_17761_, _17760_, _43998_);
  not (_17762_, \oc8051_golden_model_1.DPH [6]);
  nor (_17763_, _04783_, _17762_);
  and (_17764_, _12613_, _04671_);
  or (_17765_, _17764_, _17763_);
  and (_17766_, _17765_, _03127_);
  and (_17768_, _04671_, _04770_);
  or (_17769_, _17768_, _17763_);
  or (_17770_, _17769_, _05535_);
  nor (_17771_, _12603_, _08373_);
  or (_17772_, _17771_, _17763_);
  or (_17773_, _17772_, _03810_);
  and (_17774_, _04783_, \oc8051_golden_model_1.ACC [6]);
  or (_17775_, _17774_, _17763_);
  and (_17776_, _17775_, _03813_);
  nor (_17777_, _03813_, _17762_);
  or (_17779_, _17777_, _02974_);
  or (_17780_, _17779_, _17776_);
  and (_17781_, _17780_, _03336_);
  and (_17782_, _17781_, _17773_);
  and (_17783_, _17769_, _03069_);
  or (_17784_, _17783_, _03075_);
  or (_17785_, _17784_, _17782_);
  or (_17786_, _17775_, _03084_);
  and (_17787_, _17786_, _08225_);
  and (_17788_, _17787_, _17785_);
  or (_17790_, _08328_, \oc8051_golden_model_1.DPH [6]);
  nor (_17791_, _08329_, _08225_);
  and (_17792_, _17791_, _17790_);
  or (_17793_, _17792_, _17788_);
  and (_17794_, _17793_, _08209_);
  nor (_17795_, _08209_, _02927_);
  or (_17796_, _17795_, _06770_);
  or (_17797_, _17796_, _17794_);
  and (_17798_, _17797_, _17770_);
  or (_17799_, _17798_, _02853_);
  or (_17801_, _17763_, _05540_);
  and (_17802_, _04783_, _05849_);
  or (_17803_, _17802_, _17801_);
  and (_17804_, _17803_, _02838_);
  and (_17805_, _17804_, _17799_);
  nor (_17806_, _12722_, _08346_);
  or (_17807_, _17806_, _17763_);
  and (_17808_, _17807_, _02579_);
  or (_17809_, _17808_, _02802_);
  or (_17810_, _17809_, _17805_);
  and (_17812_, _12729_, _04783_);
  or (_17813_, _17812_, _17763_);
  or (_17814_, _17813_, _02803_);
  and (_17815_, _17814_, _17810_);
  or (_17816_, _17815_, _02980_);
  and (_17817_, _12739_, _04671_);
  or (_17818_, _17763_, _03887_);
  or (_17819_, _17818_, _17817_);
  and (_17820_, _17819_, _03128_);
  and (_17821_, _17820_, _17816_);
  or (_17823_, _17821_, _17766_);
  and (_17824_, _17823_, _03883_);
  or (_17825_, _17763_, _04819_);
  and (_17826_, _17813_, _02970_);
  and (_17827_, _17826_, _17825_);
  or (_17828_, _17827_, _17824_);
  and (_17829_, _17828_, _03137_);
  and (_17830_, _17775_, _03135_);
  and (_17831_, _17830_, _17825_);
  or (_17832_, _17831_, _02965_);
  or (_17834_, _17832_, _17829_);
  nor (_17835_, _12737_, _08373_);
  or (_17836_, _17763_, _05783_);
  or (_17837_, _17836_, _17835_);
  and (_17838_, _17837_, _05788_);
  and (_17839_, _17838_, _17834_);
  nor (_17840_, _12612_, _08373_);
  or (_17841_, _17840_, _17763_);
  and (_17842_, _17841_, _03123_);
  or (_17843_, _17842_, _03163_);
  or (_17845_, _17843_, _17839_);
  or (_17846_, _17772_, _03906_);
  and (_17847_, _17846_, _02890_);
  and (_17848_, _17847_, _17845_);
  and (_17849_, _12794_, _04671_);
  or (_17850_, _17849_, _17763_);
  and (_17851_, _17850_, _02888_);
  or (_17852_, _17851_, _42672_);
  or (_17853_, _17852_, _17848_);
  and (_43445_, _17853_, _17761_);
  not (_17855_, \oc8051_golden_model_1.IE [0]);
  nor (_17856_, _04703_, _17855_);
  and (_17857_, _11522_, _04703_);
  nor (_17858_, _17857_, _17856_);
  nor (_17859_, _17858_, _03128_);
  and (_17860_, _04703_, _03808_);
  nor (_17861_, _17860_, _17856_);
  and (_17862_, _17861_, _06770_);
  and (_17863_, _04703_, \oc8051_golden_model_1.ACC [0]);
  nor (_17864_, _17863_, _17856_);
  nor (_17866_, _17864_, _03814_);
  nor (_17867_, _03813_, _17855_);
  or (_17868_, _17867_, _17866_);
  and (_17869_, _17868_, _03810_);
  and (_17870_, _05226_, _04703_);
  nor (_17871_, _17870_, _17856_);
  nor (_17872_, _17871_, _03810_);
  or (_17873_, _17872_, _17869_);
  and (_17874_, _17873_, _02881_);
  nor (_17875_, _05340_, _17855_);
  and (_17877_, _11417_, _05340_);
  nor (_17878_, _17877_, _17875_);
  nor (_17879_, _17878_, _02881_);
  nor (_17880_, _17879_, _17874_);
  nor (_17881_, _17880_, _03069_);
  nor (_17882_, _17861_, _03336_);
  or (_17883_, _17882_, _17881_);
  and (_17884_, _17883_, _03084_);
  nor (_17885_, _17864_, _03084_);
  or (_17886_, _17885_, _17884_);
  and (_17888_, _17886_, _02877_);
  and (_17889_, _17856_, _02876_);
  or (_17890_, _17889_, _17888_);
  and (_17891_, _17890_, _02870_);
  nor (_17892_, _17871_, _02870_);
  or (_17893_, _17892_, _17891_);
  and (_17894_, _17893_, _02864_);
  nor (_17895_, _11448_, _08433_);
  nor (_17896_, _17895_, _17875_);
  nor (_17897_, _17896_, _02864_);
  or (_17899_, _17897_, _06770_);
  nor (_17900_, _17899_, _17894_);
  nor (_17901_, _17900_, _17862_);
  nor (_17902_, _17901_, _02853_);
  and (_17903_, _04703_, _06152_);
  nor (_17904_, _17856_, _05540_);
  not (_17905_, _17904_);
  nor (_17906_, _17905_, _17903_);
  or (_17907_, _17906_, _02579_);
  nor (_17908_, _17907_, _17902_);
  nor (_17910_, _11505_, _08449_);
  nor (_17911_, _17910_, _17856_);
  nor (_17912_, _17911_, _02838_);
  or (_17913_, _17912_, _02802_);
  or (_17914_, _17913_, _17908_);
  and (_17915_, _04703_, _05672_);
  nor (_17916_, _17915_, _17856_);
  nand (_17917_, _17916_, _02802_);
  and (_17918_, _17917_, _17914_);
  and (_17919_, _17918_, _03887_);
  and (_17921_, _11399_, _04703_);
  nor (_17922_, _17921_, _17856_);
  nor (_17923_, _17922_, _03887_);
  or (_17924_, _17923_, _17919_);
  and (_17925_, _17924_, _03128_);
  nor (_17926_, _17925_, _17859_);
  nor (_17927_, _17926_, _02970_);
  or (_17928_, _17916_, _03883_);
  nor (_17929_, _17928_, _17870_);
  nor (_17930_, _17929_, _17927_);
  nor (_17932_, _17930_, _03135_);
  and (_17933_, _11521_, _04703_);
  or (_17934_, _17933_, _17856_);
  and (_17935_, _17934_, _03135_);
  or (_17936_, _17935_, _17932_);
  and (_17937_, _17936_, _05783_);
  nor (_17938_, _11396_, _08449_);
  nor (_17939_, _17938_, _17856_);
  nor (_17940_, _17939_, _05783_);
  or (_17941_, _17940_, _17937_);
  and (_17943_, _17941_, _05788_);
  nor (_17944_, _11520_, _08449_);
  nor (_17945_, _17944_, _17856_);
  nor (_17946_, _17945_, _05788_);
  or (_17947_, _17946_, _17943_);
  and (_17948_, _17947_, _03906_);
  nor (_17949_, _17871_, _03906_);
  or (_17950_, _17949_, _17948_);
  and (_17951_, _17950_, _02498_);
  and (_17952_, _17856_, _02497_);
  or (_17954_, _17952_, _17951_);
  and (_17955_, _17954_, _02890_);
  nor (_17956_, _17871_, _02890_);
  or (_17957_, _17956_, _17955_);
  or (_17958_, _17957_, _42672_);
  or (_17959_, _42668_, \oc8051_golden_model_1.IE [0]);
  and (_17960_, _17959_, _43998_);
  and (_43446_, _17960_, _17958_);
  not (_17961_, _03124_);
  not (_17962_, \oc8051_golden_model_1.IE [1]);
  nor (_17964_, _04703_, _17962_);
  nor (_17965_, _11695_, _08449_);
  or (_17966_, _17965_, _17964_);
  and (_17967_, _17966_, _02579_);
  and (_17968_, _04703_, _06151_);
  or (_17969_, _17968_, _17964_);
  and (_17970_, _17969_, _02853_);
  nor (_17971_, _04703_, \oc8051_golden_model_1.IE [1]);
  and (_17972_, _04703_, _02551_);
  nor (_17973_, _17972_, _17971_);
  and (_17975_, _17973_, _03813_);
  nor (_17976_, _03813_, _17962_);
  or (_17977_, _17976_, _17975_);
  and (_17978_, _17977_, _03810_);
  and (_17979_, _11606_, _04703_);
  nor (_17980_, _17979_, _17971_);
  and (_17981_, _17980_, _02974_);
  or (_17982_, _17981_, _17978_);
  and (_17983_, _17982_, _02881_);
  nor (_17984_, _05340_, _17962_);
  and (_17986_, _11592_, _05340_);
  nor (_17987_, _17986_, _17984_);
  nor (_17988_, _17987_, _02881_);
  or (_17989_, _17988_, _17983_);
  and (_17990_, _17989_, _03336_);
  and (_17991_, _04703_, _04000_);
  nor (_17992_, _17991_, _17964_);
  nor (_17993_, _17992_, _03336_);
  or (_17994_, _17993_, _17990_);
  and (_17995_, _17994_, _03084_);
  and (_17997_, _17973_, _03075_);
  or (_17998_, _17997_, _17995_);
  and (_17999_, _17998_, _02877_);
  and (_18000_, _11595_, _05340_);
  nor (_18001_, _18000_, _17984_);
  nor (_18002_, _18001_, _02877_);
  or (_18003_, _18002_, _17999_);
  and (_18004_, _18003_, _02870_);
  and (_18005_, _17986_, _11591_);
  or (_18006_, _18005_, _17984_);
  and (_18008_, _18006_, _02869_);
  or (_18009_, _18008_, _18004_);
  and (_18010_, _18009_, _02864_);
  nor (_18011_, _11638_, _08433_);
  nor (_18012_, _17984_, _18011_);
  nor (_18013_, _18012_, _02864_);
  or (_18014_, _18013_, _06770_);
  nor (_18015_, _18014_, _18010_);
  and (_18016_, _17992_, _06770_);
  or (_18017_, _18016_, _02853_);
  nor (_18019_, _18017_, _18015_);
  or (_18020_, _18019_, _17970_);
  and (_18021_, _18020_, _02838_);
  nor (_18022_, _18021_, _17967_);
  nor (_18023_, _18022_, _02802_);
  and (_18024_, _04703_, _03698_);
  not (_18025_, _18024_);
  nor (_18026_, _17971_, _02803_);
  and (_18027_, _18026_, _18025_);
  nor (_18028_, _18027_, _18023_);
  nor (_18030_, _18028_, _02980_);
  not (_18031_, _17971_);
  nor (_18032_, _11710_, _08449_);
  nor (_18033_, _18032_, _03887_);
  and (_18034_, _18033_, _18031_);
  nor (_18035_, _18034_, _18030_);
  nor (_18036_, _18035_, _03127_);
  nor (_18037_, _11715_, _08449_);
  nor (_18038_, _18037_, _03128_);
  and (_18039_, _18038_, _18031_);
  nor (_18041_, _18039_, _18036_);
  nor (_18042_, _18041_, _02970_);
  nor (_18043_, _11709_, _08449_);
  nor (_18044_, _18043_, _03883_);
  and (_18045_, _18044_, _18031_);
  nor (_18046_, _18045_, _18042_);
  nor (_18047_, _18046_, _03135_);
  nor (_18048_, _17964_, _13722_);
  nor (_18049_, _18048_, _03137_);
  and (_18050_, _18049_, _17973_);
  nor (_18052_, _18050_, _18047_);
  or (_18053_, _18052_, _17961_);
  and (_18054_, _11714_, _04703_);
  or (_18055_, _18054_, _05788_);
  or (_18056_, _18055_, _17971_);
  and (_18057_, _18056_, _03906_);
  and (_18058_, _18024_, _05178_);
  or (_18059_, _17971_, _05783_);
  or (_18060_, _18059_, _18058_);
  and (_18061_, _18060_, _18057_);
  and (_18063_, _18061_, _18053_);
  nor (_18064_, _17980_, _03906_);
  or (_18065_, _18064_, _02497_);
  nor (_18066_, _18065_, _18063_);
  nor (_18067_, _18001_, _02498_);
  or (_18068_, _18067_, _02888_);
  nor (_18069_, _18068_, _18066_);
  nor (_18070_, _17979_, _17964_);
  and (_18071_, _18070_, _02888_);
  nor (_18072_, _18071_, _18069_);
  or (_18074_, _18072_, _42672_);
  or (_18075_, _42668_, \oc8051_golden_model_1.IE [1]);
  and (_18076_, _18075_, _43998_);
  and (_43447_, _18076_, _18074_);
  not (_18077_, \oc8051_golden_model_1.IE [2]);
  nor (_18078_, _04703_, _18077_);
  and (_18079_, _11927_, _04703_);
  nor (_18080_, _18079_, _18078_);
  nor (_18081_, _18080_, _03128_);
  and (_18082_, _04703_, _04435_);
  nor (_18084_, _18082_, _18078_);
  and (_18085_, _18084_, _06770_);
  nor (_18086_, _18084_, _03336_);
  nor (_18087_, _05340_, _18077_);
  and (_18088_, _11815_, _05340_);
  nor (_18089_, _18088_, _18087_);
  and (_18090_, _18089_, _02880_);
  nor (_18091_, _11801_, _08449_);
  nor (_18092_, _18091_, _18078_);
  nor (_18093_, _18092_, _03810_);
  nor (_18095_, _03813_, _18077_);
  and (_18096_, _04703_, \oc8051_golden_model_1.ACC [2]);
  nor (_18097_, _18096_, _18078_);
  nor (_18098_, _18097_, _03814_);
  nor (_18099_, _18098_, _18095_);
  nor (_18100_, _18099_, _02974_);
  or (_18101_, _18100_, _02880_);
  nor (_18102_, _18101_, _18093_);
  nor (_18103_, _18102_, _18090_);
  and (_18104_, _18103_, _03336_);
  or (_18106_, _18104_, _18086_);
  and (_18107_, _18106_, _03084_);
  nor (_18108_, _18097_, _03084_);
  or (_18109_, _18108_, _18107_);
  and (_18110_, _18109_, _02877_);
  and (_18111_, _11797_, _05340_);
  nor (_18112_, _18111_, _18087_);
  nor (_18113_, _18112_, _02877_);
  or (_18114_, _18113_, _18110_);
  and (_18115_, _18114_, _02870_);
  nor (_18117_, _18087_, _11830_);
  nor (_18118_, _18117_, _18089_);
  and (_18119_, _18118_, _02869_);
  or (_18120_, _18119_, _18115_);
  and (_18121_, _18120_, _02864_);
  nor (_18122_, _11848_, _08433_);
  nor (_18123_, _18122_, _18087_);
  nor (_18124_, _18123_, _02864_);
  nor (_18125_, _18124_, _06770_);
  not (_18126_, _18125_);
  nor (_18128_, _18126_, _18121_);
  nor (_18129_, _18128_, _18085_);
  nor (_18130_, _18129_, _02853_);
  and (_18131_, _04703_, _06155_);
  nor (_18132_, _18078_, _05540_);
  not (_18133_, _18132_);
  nor (_18134_, _18133_, _18131_);
  or (_18135_, _18134_, _02579_);
  nor (_18136_, _18135_, _18130_);
  nor (_18137_, _11906_, _08449_);
  nor (_18139_, _18137_, _18078_);
  nor (_18140_, _18139_, _02838_);
  or (_18141_, _18140_, _02802_);
  or (_18142_, _18141_, _18136_);
  and (_18143_, _04703_, _05701_);
  nor (_18144_, _18143_, _18078_);
  nand (_18145_, _18144_, _02802_);
  and (_18146_, _18145_, _18142_);
  and (_18147_, _18146_, _03887_);
  and (_18148_, _11921_, _04703_);
  nor (_18150_, _18148_, _18078_);
  nor (_18151_, _18150_, _03887_);
  or (_18152_, _18151_, _18147_);
  and (_18153_, _18152_, _03128_);
  nor (_18154_, _18153_, _18081_);
  nor (_18155_, _18154_, _02970_);
  nor (_18156_, _18078_, _05130_);
  not (_18157_, _18156_);
  nor (_18158_, _18144_, _03883_);
  and (_18159_, _18158_, _18157_);
  nor (_18161_, _18159_, _18155_);
  nor (_18162_, _18161_, _03135_);
  nor (_18163_, _18097_, _03137_);
  and (_18164_, _18163_, _18157_);
  nor (_18165_, _18164_, _02965_);
  not (_18166_, _18165_);
  nor (_18167_, _18166_, _18162_);
  nor (_18168_, _11919_, _08449_);
  or (_18169_, _18078_, _05783_);
  nor (_18170_, _18169_, _18168_);
  or (_18172_, _18170_, _03123_);
  nor (_18173_, _18172_, _18167_);
  nor (_18174_, _11926_, _08449_);
  nor (_18175_, _18174_, _18078_);
  nor (_18176_, _18175_, _05788_);
  or (_18177_, _18176_, _18173_);
  and (_18178_, _18177_, _03906_);
  nor (_18179_, _18092_, _03906_);
  or (_18180_, _18179_, _18178_);
  and (_18181_, _18180_, _02498_);
  nor (_18183_, _18112_, _02498_);
  or (_18184_, _18183_, _18181_);
  and (_18185_, _18184_, _02890_);
  and (_18186_, _11985_, _04703_);
  nor (_18187_, _18186_, _18078_);
  nor (_18188_, _18187_, _02890_);
  or (_18189_, _18188_, _18185_);
  or (_18190_, _18189_, _42672_);
  or (_18191_, _42668_, \oc8051_golden_model_1.IE [2]);
  and (_18192_, _18191_, _43998_);
  and (_43448_, _18192_, _18190_);
  not (_18194_, \oc8051_golden_model_1.IE [3]);
  nor (_18195_, _04703_, _18194_);
  and (_18196_, _12133_, _04703_);
  nor (_18197_, _18196_, _18195_);
  nor (_18198_, _18197_, _03128_);
  and (_18199_, _04703_, _04241_);
  nor (_18200_, _18199_, _18195_);
  and (_18201_, _18200_, _06770_);
  and (_18202_, _04703_, \oc8051_golden_model_1.ACC [3]);
  nor (_18204_, _18202_, _18195_);
  nor (_18205_, _18204_, _03814_);
  nor (_18206_, _03813_, _18194_);
  or (_18207_, _18206_, _18205_);
  and (_18208_, _18207_, _03810_);
  nor (_18209_, _12017_, _08449_);
  nor (_18210_, _18209_, _18195_);
  nor (_18211_, _18210_, _03810_);
  or (_18212_, _18211_, _18208_);
  and (_18213_, _18212_, _02881_);
  nor (_18215_, _05340_, _18194_);
  and (_18216_, _12021_, _05340_);
  nor (_18217_, _18216_, _18215_);
  nor (_18218_, _18217_, _02881_);
  or (_18219_, _18218_, _03069_);
  or (_18220_, _18219_, _18213_);
  nand (_18221_, _18200_, _03069_);
  and (_18222_, _18221_, _18220_);
  and (_18223_, _18222_, _03084_);
  nor (_18224_, _18204_, _03084_);
  or (_18226_, _18224_, _18223_);
  and (_18227_, _18226_, _02877_);
  and (_18228_, _12005_, _05340_);
  nor (_18229_, _18228_, _18215_);
  nor (_18230_, _18229_, _02877_);
  or (_18231_, _18230_, _02869_);
  or (_18232_, _18231_, _18227_);
  nor (_18233_, _18215_, _12036_);
  nor (_18234_, _18233_, _18217_);
  or (_18235_, _18234_, _02870_);
  and (_18237_, _18235_, _02864_);
  and (_18238_, _18237_, _18232_);
  nor (_18239_, _12054_, _08433_);
  nor (_18240_, _18239_, _18215_);
  nor (_18241_, _18240_, _02864_);
  nor (_18242_, _18241_, _06770_);
  not (_18243_, _18242_);
  nor (_18244_, _18243_, _18238_);
  nor (_18245_, _18244_, _18201_);
  nor (_18246_, _18245_, _02853_);
  and (_18248_, _04703_, _06154_);
  nor (_18249_, _18195_, _05540_);
  not (_18250_, _18249_);
  nor (_18251_, _18250_, _18248_);
  or (_18252_, _18251_, _02579_);
  nor (_18253_, _18252_, _18246_);
  nor (_18254_, _12112_, _08449_);
  nor (_18255_, _18254_, _18195_);
  nor (_18256_, _18255_, _02838_);
  or (_18257_, _18256_, _02802_);
  or (_18259_, _18257_, _18253_);
  and (_18260_, _04703_, _05658_);
  nor (_18261_, _18260_, _18195_);
  nand (_18262_, _18261_, _02802_);
  and (_18263_, _18262_, _18259_);
  and (_18264_, _18263_, _03887_);
  and (_18265_, _12127_, _04703_);
  nor (_18266_, _18265_, _18195_);
  nor (_18267_, _18266_, _03887_);
  or (_18268_, _18267_, _18264_);
  and (_18270_, _18268_, _03128_);
  nor (_18271_, _18270_, _18198_);
  nor (_18272_, _18271_, _02970_);
  nor (_18273_, _18195_, _05079_);
  not (_18274_, _18273_);
  nor (_18275_, _18261_, _03883_);
  and (_18276_, _18275_, _18274_);
  nor (_18277_, _18276_, _18272_);
  nor (_18278_, _18277_, _03135_);
  nor (_18279_, _18204_, _03137_);
  and (_18281_, _18279_, _18274_);
  or (_18282_, _18281_, _18278_);
  and (_18283_, _18282_, _05783_);
  nor (_18284_, _12125_, _08449_);
  nor (_18285_, _18284_, _18195_);
  nor (_18286_, _18285_, _05783_);
  or (_18287_, _18286_, _18283_);
  and (_18288_, _18287_, _05788_);
  nor (_18289_, _12132_, _08449_);
  nor (_18290_, _18289_, _18195_);
  nor (_18292_, _18290_, _05788_);
  or (_18293_, _18292_, _18288_);
  and (_18294_, _18293_, _03906_);
  nor (_18295_, _18210_, _03906_);
  or (_18296_, _18295_, _18294_);
  and (_18297_, _18296_, _02498_);
  nor (_18298_, _18229_, _02498_);
  or (_18299_, _18298_, _18297_);
  and (_18300_, _18299_, _02890_);
  and (_18301_, _12183_, _04703_);
  nor (_18303_, _18301_, _18195_);
  nor (_18304_, _18303_, _02890_);
  or (_18305_, _18304_, _18300_);
  or (_18306_, _18305_, _42672_);
  or (_18307_, _42668_, \oc8051_golden_model_1.IE [3]);
  and (_18308_, _18307_, _43998_);
  and (_43449_, _18308_, _18306_);
  not (_18309_, \oc8051_golden_model_1.IE [4]);
  nor (_18310_, _04703_, _18309_);
  and (_18311_, _12207_, _04703_);
  nor (_18313_, _18311_, _18310_);
  nor (_18314_, _18313_, _03128_);
  and (_18315_, _04703_, _04982_);
  nor (_18316_, _18315_, _18310_);
  and (_18317_, _18316_, _06770_);
  nor (_18318_, _05340_, _18309_);
  and (_18319_, _12213_, _05340_);
  nor (_18320_, _18319_, _18318_);
  nor (_18321_, _18320_, _02877_);
  and (_18322_, _04703_, \oc8051_golden_model_1.ACC [4]);
  nor (_18324_, _18322_, _18310_);
  nor (_18325_, _18324_, _03814_);
  nor (_18326_, _03813_, _18309_);
  or (_18327_, _18326_, _18325_);
  and (_18328_, _18327_, _03810_);
  nor (_18329_, _12217_, _08449_);
  nor (_18330_, _18329_, _18310_);
  nor (_18331_, _18330_, _03810_);
  or (_18332_, _18331_, _18328_);
  and (_18333_, _18332_, _02881_);
  and (_18335_, _12231_, _05340_);
  nor (_18336_, _18335_, _18318_);
  nor (_18337_, _18336_, _02881_);
  or (_18338_, _18337_, _03069_);
  or (_18339_, _18338_, _18333_);
  nand (_18340_, _18316_, _03069_);
  and (_18341_, _18340_, _18339_);
  and (_18342_, _18341_, _03084_);
  nor (_18343_, _18324_, _03084_);
  or (_18344_, _18343_, _18342_);
  and (_18346_, _18344_, _02877_);
  nor (_18347_, _18346_, _18321_);
  nor (_18348_, _18347_, _02869_);
  nor (_18349_, _18318_, _12246_);
  or (_18350_, _18336_, _02870_);
  nor (_18351_, _18350_, _18349_);
  nor (_18352_, _18351_, _18348_);
  nor (_18353_, _18352_, _02863_);
  nor (_18354_, _12264_, _08433_);
  nor (_18355_, _18354_, _18318_);
  nor (_18357_, _18355_, _02864_);
  nor (_18358_, _18357_, _06770_);
  not (_18359_, _18358_);
  nor (_18360_, _18359_, _18353_);
  nor (_18361_, _18360_, _18317_);
  nor (_18362_, _18361_, _02853_);
  and (_18363_, _04703_, _06159_);
  nor (_18364_, _18310_, _05540_);
  not (_18365_, _18364_);
  nor (_18366_, _18365_, _18363_);
  nor (_18368_, _18366_, _02579_);
  not (_18369_, _18368_);
  nor (_18370_, _18369_, _18362_);
  nor (_18371_, _12321_, _08449_);
  nor (_18372_, _18371_, _18310_);
  nor (_18373_, _18372_, _02838_);
  or (_18374_, _18373_, _02802_);
  or (_18375_, _18374_, _18370_);
  and (_18376_, _05666_, _04703_);
  nor (_18377_, _18376_, _18310_);
  nand (_18379_, _18377_, _02802_);
  and (_18380_, _18379_, _18375_);
  and (_18381_, _18380_, _03887_);
  and (_18382_, _12211_, _04703_);
  nor (_18383_, _18382_, _18310_);
  nor (_18384_, _18383_, _03887_);
  or (_18385_, _18384_, _18381_);
  and (_18386_, _18385_, _03128_);
  nor (_18387_, _18386_, _18314_);
  nor (_18388_, _18387_, _02970_);
  nor (_18390_, _18310_, _05031_);
  not (_18391_, _18390_);
  nor (_18392_, _18377_, _03883_);
  and (_18393_, _18392_, _18391_);
  nor (_18394_, _18393_, _18388_);
  nor (_18395_, _18394_, _03135_);
  nor (_18396_, _18324_, _03137_);
  and (_18397_, _18396_, _18391_);
  or (_18398_, _18397_, _18395_);
  and (_18399_, _18398_, _05783_);
  nor (_18401_, _12209_, _08449_);
  nor (_18402_, _18401_, _18310_);
  nor (_18403_, _18402_, _05783_);
  or (_18404_, _18403_, _18399_);
  and (_18405_, _18404_, _05788_);
  nor (_18406_, _12206_, _08449_);
  nor (_18407_, _18406_, _18310_);
  nor (_18408_, _18407_, _05788_);
  or (_18409_, _18408_, _18405_);
  and (_18410_, _18409_, _03906_);
  nor (_18412_, _18330_, _03906_);
  or (_18413_, _18412_, _18410_);
  and (_18414_, _18413_, _02498_);
  nor (_18415_, _18320_, _02498_);
  or (_18416_, _18415_, _18414_);
  and (_18417_, _18416_, _02890_);
  and (_18418_, _12389_, _04703_);
  nor (_18419_, _18418_, _18310_);
  nor (_18420_, _18419_, _02890_);
  or (_18421_, _18420_, _18417_);
  or (_18423_, _18421_, _42672_);
  or (_18424_, _42668_, \oc8051_golden_model_1.IE [4]);
  and (_18425_, _18424_, _43998_);
  and (_43450_, _18425_, _18423_);
  not (_18426_, \oc8051_golden_model_1.IE [5]);
  nor (_18427_, _04703_, _18426_);
  and (_18428_, _12411_, _04703_);
  nor (_18429_, _18428_, _18427_);
  nor (_18430_, _18429_, _03128_);
  and (_18431_, _04703_, _06158_);
  or (_18433_, _18431_, _18427_);
  and (_18434_, _18433_, _02853_);
  nor (_18435_, _12407_, _08449_);
  nor (_18436_, _18435_, _18427_);
  and (_18437_, _18436_, _02974_);
  and (_18438_, _04703_, \oc8051_golden_model_1.ACC [5]);
  nor (_18439_, _18438_, _18427_);
  or (_18440_, _18439_, _03814_);
  or (_18441_, _03813_, _18426_);
  and (_18442_, _18441_, _03810_);
  and (_18444_, _18442_, _18440_);
  or (_18445_, _18444_, _02880_);
  nor (_18446_, _18445_, _18437_);
  nor (_18447_, _05340_, _18426_);
  and (_18448_, _12435_, _05340_);
  nor (_18449_, _18448_, _18447_);
  nor (_18450_, _18449_, _02881_);
  or (_18451_, _18450_, _03069_);
  or (_18452_, _18451_, _18446_);
  and (_18453_, _04703_, _04877_);
  nor (_18455_, _18453_, _18427_);
  nand (_18456_, _18455_, _03069_);
  and (_18457_, _18456_, _18452_);
  and (_18458_, _18457_, _03084_);
  nor (_18459_, _18439_, _03084_);
  or (_18460_, _18459_, _18458_);
  and (_18461_, _18460_, _02877_);
  and (_18462_, _12417_, _05340_);
  nor (_18463_, _18462_, _18447_);
  nor (_18464_, _18463_, _02877_);
  or (_18466_, _18464_, _18461_);
  and (_18467_, _18466_, _02870_);
  nor (_18468_, _18447_, _12450_);
  nor (_18469_, _18468_, _18449_);
  and (_18470_, _18469_, _02869_);
  or (_18471_, _18470_, _18467_);
  and (_18472_, _18471_, _02864_);
  nor (_18473_, _12468_, _08433_);
  nor (_18474_, _18473_, _18447_);
  nor (_18475_, _18474_, _02864_);
  nor (_18477_, _18475_, _06770_);
  not (_18478_, _18477_);
  nor (_18479_, _18478_, _18472_);
  and (_18480_, _18455_, _06770_);
  or (_18481_, _18480_, _02853_);
  nor (_18482_, _18481_, _18479_);
  or (_18483_, _18482_, _18434_);
  and (_18484_, _18483_, _02838_);
  nor (_18485_, _12527_, _08449_);
  nor (_18486_, _18485_, _18427_);
  nor (_18488_, _18486_, _02838_);
  or (_18489_, _18488_, _02802_);
  or (_18490_, _18489_, _18484_);
  and (_18491_, _05614_, _04703_);
  nor (_18492_, _18491_, _18427_);
  nand (_18493_, _18492_, _02802_);
  and (_18494_, _18493_, _18490_);
  and (_18495_, _18494_, _03887_);
  and (_18496_, _12415_, _04703_);
  nor (_18497_, _18496_, _18427_);
  nor (_18499_, _18497_, _03887_);
  or (_18500_, _18499_, _18495_);
  and (_18501_, _18500_, _03128_);
  nor (_18502_, _18501_, _18430_);
  nor (_18503_, _18502_, _02970_);
  nor (_18504_, _18427_, _04924_);
  not (_18505_, _18504_);
  nor (_18506_, _18492_, _03883_);
  and (_18507_, _18506_, _18505_);
  nor (_18508_, _18507_, _18503_);
  nor (_18510_, _18508_, _03135_);
  nor (_18511_, _18439_, _03137_);
  and (_18512_, _18511_, _18505_);
  or (_18513_, _18512_, _18510_);
  and (_18514_, _18513_, _05783_);
  nor (_18515_, _12413_, _08449_);
  nor (_18516_, _18515_, _18427_);
  nor (_18517_, _18516_, _05783_);
  or (_18518_, _18517_, _18514_);
  and (_18519_, _18518_, _05788_);
  nor (_18521_, _12410_, _08449_);
  nor (_18522_, _18521_, _18427_);
  nor (_18523_, _18522_, _05788_);
  or (_18524_, _18523_, _18519_);
  and (_18525_, _18524_, _03906_);
  nor (_18526_, _18436_, _03906_);
  or (_18527_, _18526_, _18525_);
  and (_18528_, _18527_, _02498_);
  nor (_18529_, _18463_, _02498_);
  or (_18530_, _18529_, _18528_);
  and (_18532_, _18530_, _02890_);
  and (_18533_, _12589_, _04703_);
  nor (_18534_, _18533_, _18427_);
  nor (_18535_, _18534_, _02890_);
  or (_18536_, _18535_, _18532_);
  or (_18537_, _18536_, _42672_);
  or (_18538_, _42668_, \oc8051_golden_model_1.IE [5]);
  and (_18539_, _18538_, _43998_);
  and (_43451_, _18539_, _18537_);
  not (_18540_, \oc8051_golden_model_1.IE [6]);
  nor (_18542_, _04703_, _18540_);
  and (_18543_, _12613_, _04703_);
  nor (_18544_, _18543_, _18542_);
  nor (_18545_, _18544_, _03128_);
  and (_18546_, _04703_, _05849_);
  or (_18547_, _18546_, _18542_);
  and (_18548_, _18547_, _02853_);
  and (_18549_, _04703_, \oc8051_golden_model_1.ACC [6]);
  nor (_18550_, _18549_, _18542_);
  nor (_18551_, _18550_, _03814_);
  nor (_18553_, _03813_, _18540_);
  or (_18554_, _18553_, _18551_);
  and (_18555_, _18554_, _03810_);
  nor (_18556_, _12603_, _08449_);
  nor (_18557_, _18556_, _18542_);
  nor (_18558_, _18557_, _03810_);
  or (_18559_, _18558_, _18555_);
  and (_18560_, _18559_, _02881_);
  nor (_18561_, _05340_, _18540_);
  and (_18562_, _12618_, _05340_);
  nor (_18564_, _18562_, _18561_);
  nor (_18565_, _18564_, _02881_);
  or (_18566_, _18565_, _03069_);
  or (_18567_, _18566_, _18560_);
  and (_18568_, _04703_, _04770_);
  nor (_18569_, _18568_, _18542_);
  nand (_18570_, _18569_, _03069_);
  and (_18571_, _18570_, _18567_);
  and (_18572_, _18571_, _03084_);
  nor (_18573_, _18550_, _03084_);
  or (_18575_, _18573_, _18572_);
  and (_18576_, _18575_, _02877_);
  and (_18577_, _12616_, _05340_);
  nor (_18578_, _18577_, _18561_);
  nor (_18579_, _18578_, _02877_);
  or (_18580_, _18579_, _02869_);
  or (_18581_, _18580_, _18576_);
  nor (_18582_, _18561_, _12646_);
  nor (_18583_, _18582_, _18564_);
  or (_18584_, _18583_, _02870_);
  and (_18586_, _18584_, _02864_);
  and (_18587_, _18586_, _18581_);
  nor (_18588_, _12664_, _08433_);
  nor (_18589_, _18588_, _18561_);
  nor (_18590_, _18589_, _02864_);
  nor (_18591_, _18590_, _06770_);
  not (_18592_, _18591_);
  nor (_18593_, _18592_, _18587_);
  and (_18594_, _18569_, _06770_);
  or (_18595_, _18594_, _02853_);
  nor (_18597_, _18595_, _18593_);
  or (_18598_, _18597_, _18548_);
  and (_18599_, _18598_, _02838_);
  nor (_18600_, _12722_, _08449_);
  nor (_18601_, _18600_, _18542_);
  nor (_18602_, _18601_, _02838_);
  or (_18603_, _18602_, _02802_);
  or (_18604_, _18603_, _18599_);
  and (_18605_, _12729_, _04703_);
  nor (_18606_, _18605_, _18542_);
  nand (_18608_, _18606_, _02802_);
  and (_18609_, _18608_, _18604_);
  and (_18610_, _18609_, _03887_);
  and (_18611_, _12739_, _04703_);
  nor (_18612_, _18611_, _18542_);
  nor (_18613_, _18612_, _03887_);
  or (_18614_, _18613_, _18610_);
  and (_18615_, _18614_, _03128_);
  nor (_18616_, _18615_, _18545_);
  nor (_18617_, _18616_, _02970_);
  nor (_18619_, _18542_, _04819_);
  not (_18620_, _18619_);
  nor (_18621_, _18606_, _03883_);
  and (_18622_, _18621_, _18620_);
  nor (_18623_, _18622_, _18617_);
  nor (_18624_, _18623_, _03135_);
  nor (_18625_, _18550_, _03137_);
  and (_18626_, _18625_, _18620_);
  nor (_18627_, _18626_, _02965_);
  not (_18628_, _18627_);
  nor (_18630_, _18628_, _18624_);
  nor (_18631_, _12737_, _08449_);
  or (_18632_, _18542_, _05783_);
  nor (_18633_, _18632_, _18631_);
  or (_18634_, _18633_, _03123_);
  nor (_18635_, _18634_, _18630_);
  nor (_18636_, _12612_, _08449_);
  nor (_18637_, _18636_, _18542_);
  nor (_18638_, _18637_, _05788_);
  or (_18639_, _18638_, _18635_);
  and (_18641_, _18639_, _03906_);
  nor (_18642_, _18557_, _03906_);
  or (_18643_, _18642_, _18641_);
  and (_18644_, _18643_, _02498_);
  nor (_18645_, _18578_, _02498_);
  or (_18646_, _18645_, _18644_);
  and (_18647_, _18646_, _02890_);
  and (_18648_, _12794_, _04703_);
  nor (_18649_, _18648_, _18542_);
  nor (_18650_, _18649_, _02890_);
  or (_18652_, _18650_, _18647_);
  or (_18653_, _18652_, _42672_);
  or (_18654_, _42668_, \oc8051_golden_model_1.IE [6]);
  and (_18655_, _18654_, _43998_);
  and (_43452_, _18655_, _18653_);
  not (_18656_, \oc8051_golden_model_1.IP [0]);
  nor (_18657_, _04693_, _18656_);
  and (_18658_, _11522_, _04693_);
  nor (_18659_, _18658_, _18657_);
  nor (_18660_, _18659_, _03128_);
  and (_18662_, _04693_, _03808_);
  nor (_18663_, _18662_, _18657_);
  and (_18664_, _18663_, _06770_);
  and (_18665_, _04693_, \oc8051_golden_model_1.ACC [0]);
  nor (_18666_, _18665_, _18657_);
  nor (_18667_, _18666_, _03814_);
  nor (_18668_, _03813_, _18656_);
  or (_18669_, _18668_, _18667_);
  and (_18670_, _18669_, _03810_);
  and (_18671_, _05226_, _04693_);
  nor (_18673_, _18671_, _18657_);
  nor (_18674_, _18673_, _03810_);
  or (_18675_, _18674_, _18670_);
  and (_18676_, _18675_, _02881_);
  nor (_18677_, _05328_, _18656_);
  and (_18678_, _11417_, _05328_);
  nor (_18679_, _18678_, _18677_);
  nor (_18680_, _18679_, _02881_);
  nor (_18681_, _18680_, _18676_);
  nor (_18682_, _18681_, _03069_);
  nor (_18684_, _18663_, _03336_);
  or (_18685_, _18684_, _18682_);
  and (_18686_, _18685_, _03084_);
  nor (_18687_, _18666_, _03084_);
  or (_18688_, _18687_, _18686_);
  and (_18689_, _18688_, _02877_);
  and (_18690_, _18657_, _02876_);
  or (_18691_, _18690_, _18689_);
  and (_18692_, _18691_, _02870_);
  nor (_18693_, _18673_, _02870_);
  or (_18695_, _18693_, _18692_);
  and (_18696_, _18695_, _02864_);
  nor (_18697_, _11448_, _08542_);
  nor (_18698_, _18697_, _18677_);
  nor (_18699_, _18698_, _02864_);
  or (_18700_, _18699_, _06770_);
  nor (_18701_, _18700_, _18696_);
  nor (_18702_, _18701_, _18664_);
  nor (_18703_, _18702_, _02853_);
  and (_18704_, _04693_, _06152_);
  nor (_18706_, _18657_, _05540_);
  not (_18707_, _18706_);
  nor (_18708_, _18707_, _18704_);
  or (_18709_, _18708_, _02579_);
  nor (_18710_, _18709_, _18703_);
  nor (_18711_, _11505_, _08558_);
  nor (_18712_, _18711_, _18657_);
  nor (_18713_, _18712_, _02838_);
  or (_18714_, _18713_, _02802_);
  or (_18715_, _18714_, _18710_);
  and (_18717_, _04693_, _05672_);
  nor (_18718_, _18717_, _18657_);
  nand (_18719_, _18718_, _02802_);
  and (_18720_, _18719_, _18715_);
  and (_18721_, _18720_, _03887_);
  and (_18722_, _11399_, _04693_);
  nor (_18723_, _18722_, _18657_);
  nor (_18724_, _18723_, _03887_);
  or (_18725_, _18724_, _18721_);
  and (_18726_, _18725_, _03128_);
  nor (_18728_, _18726_, _18660_);
  nor (_18729_, _18728_, _02970_);
  or (_18730_, _18718_, _03883_);
  nor (_18731_, _18730_, _18671_);
  nor (_18732_, _18731_, _18729_);
  nor (_18733_, _18732_, _03135_);
  nor (_18734_, _18657_, _09409_);
  or (_18735_, _18734_, _03137_);
  nor (_18736_, _18735_, _18666_);
  or (_18737_, _18736_, _18733_);
  and (_18739_, _18737_, _05783_);
  nor (_18740_, _11396_, _08558_);
  nor (_18741_, _18740_, _18657_);
  nor (_18742_, _18741_, _05783_);
  or (_18743_, _18742_, _18739_);
  and (_18744_, _18743_, _05788_);
  nor (_18745_, _11520_, _08558_);
  nor (_18746_, _18745_, _18657_);
  nor (_18747_, _18746_, _05788_);
  or (_18748_, _18747_, _18744_);
  and (_18750_, _18748_, _03906_);
  nor (_18751_, _18673_, _03906_);
  or (_18752_, _18751_, _18750_);
  and (_18753_, _18752_, _02498_);
  and (_18754_, _18657_, _02497_);
  nor (_18755_, _18754_, _02888_);
  not (_18756_, _18755_);
  nor (_18757_, _18756_, _18753_);
  and (_18758_, _18673_, _02888_);
  or (_18759_, _18758_, _18757_);
  nand (_18761_, _18759_, _42668_);
  or (_18762_, _42668_, \oc8051_golden_model_1.IP [0]);
  and (_18763_, _18762_, _43998_);
  and (_43454_, _18763_, _18761_);
  and (_18764_, _04693_, _03698_);
  not (_18765_, _18764_);
  nor (_18766_, _04693_, \oc8051_golden_model_1.IP [1]);
  nor (_18767_, _18766_, _02803_);
  and (_18768_, _18767_, _18765_);
  not (_18769_, \oc8051_golden_model_1.IP [1]);
  nor (_18771_, _04693_, _18769_);
  nor (_18772_, _11695_, _08558_);
  or (_18773_, _18772_, _18771_);
  and (_18774_, _18773_, _02579_);
  and (_18775_, _04693_, _06151_);
  or (_18776_, _18775_, _18771_);
  and (_18777_, _18776_, _02853_);
  and (_18778_, _04693_, _02551_);
  nor (_18779_, _18778_, _18766_);
  and (_18780_, _18779_, _03813_);
  nor (_18782_, _03813_, _18769_);
  or (_18783_, _18782_, _18780_);
  and (_18784_, _18783_, _03810_);
  and (_18785_, _11606_, _04693_);
  nor (_18786_, _18785_, _18766_);
  and (_18787_, _18786_, _02974_);
  or (_18788_, _18787_, _18784_);
  and (_18789_, _18788_, _02881_);
  nor (_18790_, _05328_, _18769_);
  and (_18791_, _11592_, _05328_);
  nor (_18793_, _18791_, _18790_);
  nor (_18794_, _18793_, _02881_);
  or (_18795_, _18794_, _18789_);
  and (_18796_, _18795_, _03336_);
  and (_18797_, _04693_, _04000_);
  nor (_18798_, _18797_, _18771_);
  nor (_18799_, _18798_, _03336_);
  or (_18800_, _18799_, _18796_);
  and (_18801_, _18800_, _03084_);
  and (_18802_, _18779_, _03075_);
  or (_18804_, _18802_, _18801_);
  and (_18805_, _18804_, _02877_);
  and (_18806_, _11595_, _05328_);
  nor (_18807_, _18806_, _18790_);
  nor (_18808_, _18807_, _02877_);
  or (_18809_, _18808_, _18805_);
  and (_18810_, _18809_, _02870_);
  and (_18811_, _18791_, _11591_);
  or (_18812_, _18811_, _18790_);
  and (_18813_, _18812_, _02869_);
  or (_18815_, _18813_, _18810_);
  and (_18816_, _18815_, _02864_);
  nor (_18817_, _11638_, _08542_);
  nor (_18818_, _18790_, _18817_);
  nor (_18819_, _18818_, _02864_);
  or (_18820_, _18819_, _06770_);
  nor (_18821_, _18820_, _18816_);
  and (_18822_, _18798_, _06770_);
  or (_18823_, _18822_, _02853_);
  nor (_18824_, _18823_, _18821_);
  or (_18826_, _18824_, _18777_);
  and (_18827_, _18826_, _02838_);
  nor (_18828_, _18827_, _18774_);
  nor (_18829_, _18828_, _02802_);
  nor (_18830_, _18829_, _18768_);
  nor (_18831_, _18830_, _02980_);
  not (_18832_, _18766_);
  nor (_18833_, _11710_, _08558_);
  nor (_18834_, _18833_, _03887_);
  and (_18835_, _18834_, _18832_);
  nor (_18837_, _18835_, _18831_);
  nor (_18838_, _18837_, _03127_);
  nor (_18839_, _11715_, _08558_);
  nor (_18840_, _18839_, _03128_);
  and (_18841_, _18840_, _18832_);
  nor (_18842_, _18841_, _18838_);
  nor (_18843_, _18842_, _02970_);
  nor (_18844_, _11709_, _08558_);
  nor (_18845_, _18844_, _03883_);
  and (_18846_, _18845_, _18832_);
  nor (_18848_, _18846_, _18843_);
  nor (_18849_, _18848_, _03135_);
  nor (_18850_, _18771_, _13722_);
  nor (_18851_, _18850_, _03137_);
  and (_18852_, _18851_, _18779_);
  nor (_18853_, _18852_, _18849_);
  or (_18854_, _18853_, _17961_);
  and (_18855_, _11714_, _04693_);
  or (_18856_, _18855_, _05788_);
  or (_18857_, _18856_, _18766_);
  and (_18859_, _18857_, _03906_);
  and (_18860_, _18764_, _05178_);
  or (_18861_, _18766_, _05783_);
  or (_18862_, _18861_, _18860_);
  and (_18863_, _18862_, _18859_);
  and (_18864_, _18863_, _18854_);
  nor (_18865_, _18786_, _03906_);
  or (_18866_, _18865_, _02497_);
  nor (_18867_, _18866_, _18864_);
  nor (_18868_, _18807_, _02498_);
  or (_18870_, _18868_, _02888_);
  nor (_18871_, _18870_, _18867_);
  nor (_18872_, _18785_, _18771_);
  and (_18873_, _18872_, _02888_);
  nor (_18874_, _18873_, _18871_);
  or (_18875_, _18874_, _42672_);
  or (_18876_, _42668_, \oc8051_golden_model_1.IP [1]);
  and (_18877_, _18876_, _43998_);
  and (_43455_, _18877_, _18875_);
  not (_18878_, \oc8051_golden_model_1.IP [2]);
  nor (_18880_, _04693_, _18878_);
  and (_18881_, _11927_, _04693_);
  nor (_18882_, _18881_, _18880_);
  nor (_18883_, _18882_, _03128_);
  and (_18884_, _04693_, _04435_);
  nor (_18885_, _18884_, _18880_);
  and (_18886_, _18885_, _06770_);
  and (_18887_, _04693_, \oc8051_golden_model_1.ACC [2]);
  nor (_18888_, _18887_, _18880_);
  nor (_18889_, _18888_, _03814_);
  nor (_18891_, _03813_, _18878_);
  or (_18892_, _18891_, _18889_);
  and (_18893_, _18892_, _03810_);
  nor (_18894_, _11801_, _08558_);
  nor (_18895_, _18894_, _18880_);
  nor (_18896_, _18895_, _03810_);
  or (_18897_, _18896_, _18893_);
  and (_18898_, _18897_, _02881_);
  nor (_18899_, _05328_, _18878_);
  and (_18900_, _11815_, _05328_);
  nor (_18902_, _18900_, _18899_);
  nor (_18903_, _18902_, _02881_);
  or (_18904_, _18903_, _18898_);
  and (_18905_, _18904_, _03336_);
  nor (_18906_, _18885_, _03336_);
  or (_18907_, _18906_, _18905_);
  and (_18908_, _18907_, _03084_);
  nor (_18909_, _18888_, _03084_);
  or (_18910_, _18909_, _18908_);
  and (_18911_, _18910_, _02877_);
  and (_18913_, _11797_, _05328_);
  nor (_18914_, _18913_, _18899_);
  nor (_18915_, _18914_, _02877_);
  or (_18916_, _18915_, _02869_);
  or (_18917_, _18916_, _18911_);
  and (_18918_, _18900_, _11830_);
  or (_18919_, _18899_, _02870_);
  or (_18920_, _18919_, _18918_);
  and (_18921_, _18920_, _02864_);
  and (_18922_, _18921_, _18917_);
  nor (_18924_, _11848_, _08542_);
  nor (_18925_, _18924_, _18899_);
  nor (_18926_, _18925_, _02864_);
  nor (_18927_, _18926_, _06770_);
  not (_18928_, _18927_);
  nor (_18929_, _18928_, _18922_);
  nor (_18930_, _18929_, _18886_);
  nor (_18931_, _18930_, _02853_);
  and (_18932_, _04693_, _06155_);
  nor (_18933_, _18880_, _05540_);
  not (_18935_, _18933_);
  nor (_18936_, _18935_, _18932_);
  or (_18937_, _18936_, _02579_);
  nor (_18938_, _18937_, _18931_);
  nor (_18939_, _11906_, _08558_);
  nor (_18940_, _18939_, _18880_);
  nor (_18941_, _18940_, _02838_);
  or (_18942_, _18941_, _02802_);
  or (_18943_, _18942_, _18938_);
  and (_18944_, _04693_, _05701_);
  nor (_18946_, _18944_, _18880_);
  nand (_18947_, _18946_, _02802_);
  and (_18948_, _18947_, _18943_);
  and (_18949_, _18948_, _03887_);
  and (_18950_, _11921_, _04693_);
  nor (_18951_, _18950_, _18880_);
  nor (_18952_, _18951_, _03887_);
  or (_18953_, _18952_, _18949_);
  and (_18954_, _18953_, _03128_);
  nor (_18955_, _18954_, _18883_);
  nor (_18957_, _18955_, _02970_);
  nor (_18958_, _18880_, _05130_);
  not (_18959_, _18958_);
  nor (_18960_, _18946_, _03883_);
  and (_18961_, _18960_, _18959_);
  nor (_18962_, _18961_, _18957_);
  nor (_18963_, _18962_, _03135_);
  nor (_18964_, _18888_, _03137_);
  and (_18965_, _18964_, _18959_);
  or (_18966_, _18965_, _18963_);
  and (_18968_, _18966_, _05783_);
  nor (_18969_, _11919_, _08558_);
  nor (_18970_, _18969_, _18880_);
  nor (_18971_, _18970_, _05783_);
  or (_18972_, _18971_, _18968_);
  and (_18973_, _18972_, _05788_);
  nor (_18974_, _11926_, _08558_);
  nor (_18975_, _18974_, _18880_);
  nor (_18976_, _18975_, _05788_);
  or (_18977_, _18976_, _18973_);
  and (_18979_, _18977_, _03906_);
  nor (_18980_, _18895_, _03906_);
  or (_18981_, _18980_, _18979_);
  and (_18982_, _18981_, _02498_);
  nor (_18983_, _18914_, _02498_);
  or (_18984_, _18983_, _18982_);
  and (_18985_, _18984_, _02890_);
  and (_18986_, _11985_, _04693_);
  nor (_18987_, _18986_, _18880_);
  nor (_18988_, _18987_, _02890_);
  or (_18990_, _18988_, _18985_);
  or (_18991_, _18990_, _42672_);
  or (_18992_, _42668_, \oc8051_golden_model_1.IP [2]);
  and (_18993_, _18992_, _43998_);
  and (_43456_, _18993_, _18991_);
  not (_18994_, \oc8051_golden_model_1.IP [3]);
  nor (_18995_, _04693_, _18994_);
  and (_18996_, _12133_, _04693_);
  nor (_18997_, _18996_, _18995_);
  nor (_18998_, _18997_, _03128_);
  and (_19000_, _04693_, _04241_);
  nor (_19001_, _19000_, _18995_);
  and (_19002_, _19001_, _06770_);
  and (_19003_, _04693_, \oc8051_golden_model_1.ACC [3]);
  nor (_19004_, _19003_, _18995_);
  nor (_19005_, _19004_, _03814_);
  nor (_19006_, _03813_, _18994_);
  or (_19007_, _19006_, _19005_);
  and (_19008_, _19007_, _03810_);
  nor (_19009_, _12017_, _08558_);
  nor (_19011_, _19009_, _18995_);
  nor (_19012_, _19011_, _03810_);
  or (_19013_, _19012_, _19008_);
  and (_19014_, _19013_, _02881_);
  nor (_19015_, _05328_, _18994_);
  and (_19016_, _12021_, _05328_);
  nor (_19017_, _19016_, _19015_);
  nor (_19018_, _19017_, _02881_);
  or (_19019_, _19018_, _03069_);
  or (_19020_, _19019_, _19014_);
  nand (_19022_, _19001_, _03069_);
  and (_19023_, _19022_, _19020_);
  and (_19024_, _19023_, _03084_);
  nor (_19025_, _19004_, _03084_);
  or (_19026_, _19025_, _19024_);
  and (_19027_, _19026_, _02877_);
  and (_19028_, _12005_, _05328_);
  nor (_19029_, _19028_, _19015_);
  nor (_19030_, _19029_, _02877_);
  or (_19031_, _19030_, _02869_);
  or (_19033_, _19031_, _19027_);
  nor (_19034_, _19015_, _12036_);
  nor (_19035_, _19034_, _19017_);
  or (_19036_, _19035_, _02870_);
  and (_19037_, _19036_, _02864_);
  and (_19038_, _19037_, _19033_);
  nor (_19039_, _12054_, _08542_);
  nor (_19040_, _19039_, _19015_);
  nor (_19041_, _19040_, _02864_);
  nor (_19042_, _19041_, _06770_);
  not (_19044_, _19042_);
  nor (_19045_, _19044_, _19038_);
  nor (_19046_, _19045_, _19002_);
  nor (_19047_, _19046_, _02853_);
  and (_19048_, _04693_, _06154_);
  nor (_19049_, _18995_, _05540_);
  not (_19050_, _19049_);
  nor (_19051_, _19050_, _19048_);
  or (_19052_, _19051_, _02579_);
  nor (_19053_, _19052_, _19047_);
  nor (_19055_, _12112_, _08558_);
  nor (_19056_, _19055_, _18995_);
  nor (_19057_, _19056_, _02838_);
  or (_19058_, _19057_, _02802_);
  or (_19059_, _19058_, _19053_);
  and (_19060_, _04693_, _05658_);
  nor (_19061_, _19060_, _18995_);
  nand (_19062_, _19061_, _02802_);
  and (_19063_, _19062_, _19059_);
  and (_19064_, _19063_, _03887_);
  and (_19066_, _12127_, _04693_);
  nor (_19067_, _19066_, _18995_);
  nor (_19068_, _19067_, _03887_);
  or (_19069_, _19068_, _19064_);
  and (_19070_, _19069_, _03128_);
  nor (_19071_, _19070_, _18998_);
  nor (_19072_, _19071_, _02970_);
  nor (_19073_, _18995_, _05079_);
  not (_19074_, _19073_);
  nor (_19075_, _19061_, _03883_);
  and (_19077_, _19075_, _19074_);
  nor (_19078_, _19077_, _19072_);
  nor (_19079_, _19078_, _03135_);
  nor (_19080_, _19004_, _03137_);
  and (_19081_, _19080_, _19074_);
  or (_19082_, _19081_, _19079_);
  and (_19083_, _19082_, _05783_);
  nor (_19084_, _12125_, _08558_);
  nor (_19085_, _19084_, _18995_);
  nor (_19086_, _19085_, _05783_);
  or (_19088_, _19086_, _19083_);
  and (_19089_, _19088_, _05788_);
  nor (_19090_, _12132_, _08558_);
  nor (_19091_, _19090_, _18995_);
  nor (_19092_, _19091_, _05788_);
  or (_19093_, _19092_, _19089_);
  and (_19094_, _19093_, _03906_);
  nor (_19095_, _19011_, _03906_);
  or (_19096_, _19095_, _19094_);
  and (_19097_, _19096_, _02498_);
  nor (_19099_, _19029_, _02498_);
  or (_19100_, _19099_, _19097_);
  and (_19101_, _19100_, _02890_);
  and (_19102_, _12183_, _04693_);
  nor (_19103_, _19102_, _18995_);
  nor (_19104_, _19103_, _02890_);
  or (_19105_, _19104_, _19101_);
  or (_19106_, _19105_, _42672_);
  or (_19107_, _42668_, \oc8051_golden_model_1.IP [3]);
  and (_19108_, _19107_, _43998_);
  and (_43457_, _19108_, _19106_);
  not (_19110_, \oc8051_golden_model_1.IP [4]);
  nor (_19111_, _04693_, _19110_);
  and (_19112_, _12207_, _04693_);
  nor (_19113_, _19112_, _19111_);
  nor (_19114_, _19113_, _03128_);
  and (_19115_, _04693_, _04982_);
  nor (_19116_, _19115_, _19111_);
  and (_19117_, _19116_, _06770_);
  nor (_19118_, _05328_, _19110_);
  and (_19120_, _12213_, _05328_);
  nor (_19121_, _19120_, _19118_);
  nor (_19122_, _19121_, _02877_);
  and (_19123_, _04693_, \oc8051_golden_model_1.ACC [4]);
  nor (_19124_, _19123_, _19111_);
  nor (_19125_, _19124_, _03814_);
  nor (_19126_, _03813_, _19110_);
  or (_19127_, _19126_, _19125_);
  and (_19128_, _19127_, _03810_);
  nor (_19129_, _12217_, _08558_);
  nor (_19131_, _19129_, _19111_);
  nor (_19132_, _19131_, _03810_);
  or (_19133_, _19132_, _19128_);
  and (_19134_, _19133_, _02881_);
  and (_19135_, _12231_, _05328_);
  nor (_19136_, _19135_, _19118_);
  nor (_19137_, _19136_, _02881_);
  or (_19138_, _19137_, _03069_);
  or (_19139_, _19138_, _19134_);
  nand (_19140_, _19116_, _03069_);
  and (_19142_, _19140_, _19139_);
  and (_19143_, _19142_, _03084_);
  nor (_19144_, _19124_, _03084_);
  or (_19145_, _19144_, _19143_);
  and (_19146_, _19145_, _02877_);
  nor (_19147_, _19146_, _19122_);
  nor (_19148_, _19147_, _02869_);
  and (_19149_, _12247_, _05328_);
  nor (_19150_, _19149_, _19118_);
  nor (_19151_, _19150_, _02870_);
  nor (_19153_, _19151_, _19148_);
  nor (_19154_, _19153_, _02863_);
  nor (_19155_, _12264_, _08542_);
  nor (_19156_, _19155_, _19118_);
  nor (_19157_, _19156_, _02864_);
  nor (_19158_, _19157_, _06770_);
  not (_19159_, _19158_);
  nor (_19160_, _19159_, _19154_);
  nor (_19161_, _19160_, _19117_);
  nor (_19162_, _19161_, _02853_);
  and (_19164_, _04693_, _06159_);
  nor (_19165_, _19111_, _05540_);
  not (_19166_, _19165_);
  nor (_19167_, _19166_, _19164_);
  nor (_19168_, _19167_, _02579_);
  not (_19169_, _19168_);
  nor (_19170_, _19169_, _19162_);
  nor (_19171_, _12321_, _08558_);
  nor (_19172_, _19171_, _19111_);
  nor (_19173_, _19172_, _02838_);
  or (_19175_, _19173_, _02802_);
  or (_19176_, _19175_, _19170_);
  and (_19177_, _05666_, _04693_);
  nor (_19178_, _19177_, _19111_);
  nand (_19179_, _19178_, _02802_);
  and (_19180_, _19179_, _19176_);
  and (_19181_, _19180_, _03887_);
  and (_19182_, _12211_, _04693_);
  nor (_19183_, _19182_, _19111_);
  nor (_19184_, _19183_, _03887_);
  or (_19186_, _19184_, _19181_);
  and (_19187_, _19186_, _03128_);
  nor (_19188_, _19187_, _19114_);
  nor (_19189_, _19188_, _02970_);
  nor (_19190_, _19111_, _05031_);
  not (_19191_, _19190_);
  nor (_19192_, _19178_, _03883_);
  and (_19193_, _19192_, _19191_);
  nor (_19194_, _19193_, _19189_);
  nor (_19195_, _19194_, _03135_);
  nor (_19197_, _19124_, _03137_);
  and (_19198_, _19197_, _19191_);
  or (_19199_, _19198_, _19195_);
  and (_19200_, _19199_, _05783_);
  nor (_19201_, _12209_, _08558_);
  nor (_19202_, _19201_, _19111_);
  nor (_19203_, _19202_, _05783_);
  or (_19204_, _19203_, _19200_);
  and (_19205_, _19204_, _05788_);
  nor (_19206_, _12206_, _08558_);
  nor (_19208_, _19206_, _19111_);
  nor (_19209_, _19208_, _05788_);
  or (_19210_, _19209_, _19205_);
  and (_19211_, _19210_, _03906_);
  nor (_19212_, _19131_, _03906_);
  or (_19213_, _19212_, _19211_);
  and (_19214_, _19213_, _02498_);
  nor (_19215_, _19121_, _02498_);
  or (_19216_, _19215_, _19214_);
  and (_19217_, _19216_, _02890_);
  and (_19219_, _12389_, _04693_);
  nor (_19220_, _19219_, _19111_);
  nor (_19221_, _19220_, _02890_);
  or (_19222_, _19221_, _19217_);
  or (_19223_, _19222_, _42672_);
  or (_19224_, _42668_, \oc8051_golden_model_1.IP [4]);
  and (_19225_, _19224_, _43998_);
  and (_43458_, _19225_, _19223_);
  not (_19226_, \oc8051_golden_model_1.IP [5]);
  nor (_19227_, _04693_, _19226_);
  and (_19229_, _12411_, _04693_);
  nor (_19230_, _19229_, _19227_);
  nor (_19231_, _19230_, _03128_);
  and (_19232_, _04693_, _06158_);
  or (_19233_, _19232_, _19227_);
  and (_19234_, _19233_, _02853_);
  nor (_19235_, _12407_, _08558_);
  nor (_19236_, _19235_, _19227_);
  and (_19237_, _19236_, _02974_);
  and (_19238_, _04693_, \oc8051_golden_model_1.ACC [5]);
  nor (_19240_, _19238_, _19227_);
  or (_19241_, _19240_, _03814_);
  or (_19242_, _03813_, _19226_);
  and (_19243_, _19242_, _03810_);
  and (_19244_, _19243_, _19241_);
  or (_19245_, _19244_, _02880_);
  nor (_19246_, _19245_, _19237_);
  nor (_19247_, _05328_, _19226_);
  and (_19248_, _12435_, _05328_);
  nor (_19249_, _19248_, _19247_);
  nor (_19251_, _19249_, _02881_);
  or (_19252_, _19251_, _03069_);
  or (_19253_, _19252_, _19246_);
  and (_19254_, _04693_, _04877_);
  nor (_19255_, _19254_, _19227_);
  nand (_19256_, _19255_, _03069_);
  and (_19257_, _19256_, _19253_);
  and (_19258_, _19257_, _03084_);
  nor (_19259_, _19240_, _03084_);
  or (_19260_, _19259_, _19258_);
  and (_19262_, _19260_, _02877_);
  and (_19263_, _12417_, _05328_);
  nor (_19264_, _19263_, _19247_);
  nor (_19265_, _19264_, _02877_);
  or (_19266_, _19265_, _19262_);
  and (_19267_, _19266_, _02870_);
  nor (_19268_, _19247_, _12450_);
  nor (_19269_, _19268_, _19249_);
  and (_19270_, _19269_, _02869_);
  or (_19271_, _19270_, _19267_);
  and (_19273_, _19271_, _02864_);
  nor (_19274_, _12468_, _08542_);
  nor (_19275_, _19274_, _19247_);
  nor (_19276_, _19275_, _02864_);
  nor (_19277_, _19276_, _06770_);
  not (_19278_, _19277_);
  nor (_19279_, _19278_, _19273_);
  and (_19280_, _19255_, _06770_);
  or (_19281_, _19280_, _02853_);
  nor (_19282_, _19281_, _19279_);
  or (_19284_, _19282_, _19234_);
  and (_19285_, _19284_, _02838_);
  nor (_19286_, _12527_, _08558_);
  nor (_19287_, _19286_, _19227_);
  nor (_19288_, _19287_, _02838_);
  or (_19289_, _19288_, _02802_);
  or (_19290_, _19289_, _19285_);
  and (_19291_, _05614_, _04693_);
  nor (_19292_, _19291_, _19227_);
  nand (_19293_, _19292_, _02802_);
  and (_19295_, _19293_, _19290_);
  and (_19296_, _19295_, _03887_);
  and (_19297_, _12415_, _04693_);
  nor (_19298_, _19297_, _19227_);
  nor (_19299_, _19298_, _03887_);
  or (_19300_, _19299_, _19296_);
  and (_19301_, _19300_, _03128_);
  nor (_19302_, _19301_, _19231_);
  nor (_19303_, _19302_, _02970_);
  nor (_19304_, _19227_, _04924_);
  not (_19306_, _19304_);
  nor (_19307_, _19292_, _03883_);
  and (_19308_, _19307_, _19306_);
  nor (_19309_, _19308_, _19303_);
  nor (_19310_, _19309_, _03135_);
  nor (_19311_, _19240_, _03137_);
  and (_19312_, _19311_, _19306_);
  nor (_19313_, _19312_, _02965_);
  not (_19314_, _19313_);
  nor (_19315_, _19314_, _19310_);
  nor (_19317_, _12413_, _08558_);
  or (_19318_, _19227_, _05783_);
  nor (_19319_, _19318_, _19317_);
  or (_19320_, _19319_, _03123_);
  nor (_19321_, _19320_, _19315_);
  nor (_19322_, _12410_, _08558_);
  nor (_19323_, _19322_, _19227_);
  nor (_19324_, _19323_, _05788_);
  or (_19325_, _19324_, _19321_);
  and (_19326_, _19325_, _03906_);
  nor (_19328_, _19236_, _03906_);
  or (_19329_, _19328_, _19326_);
  and (_19330_, _19329_, _02498_);
  nor (_19331_, _19264_, _02498_);
  or (_19332_, _19331_, _19330_);
  and (_19333_, _19332_, _02890_);
  and (_19334_, _12589_, _04693_);
  nor (_19335_, _19334_, _19227_);
  nor (_19336_, _19335_, _02890_);
  or (_19337_, _19336_, _19333_);
  or (_19339_, _19337_, _42672_);
  or (_19340_, _42668_, \oc8051_golden_model_1.IP [5]);
  and (_19341_, _19340_, _43998_);
  and (_43459_, _19341_, _19339_);
  not (_19342_, \oc8051_golden_model_1.IP [6]);
  nor (_19343_, _04693_, _19342_);
  and (_19344_, _12613_, _04693_);
  nor (_19345_, _19344_, _19343_);
  nor (_19346_, _19345_, _03128_);
  and (_19347_, _04693_, _05849_);
  or (_19349_, _19347_, _19343_);
  and (_19350_, _19349_, _02853_);
  and (_19351_, _04693_, \oc8051_golden_model_1.ACC [6]);
  nor (_19352_, _19351_, _19343_);
  nor (_19353_, _19352_, _03814_);
  nor (_19354_, _03813_, _19342_);
  or (_19355_, _19354_, _19353_);
  and (_19356_, _19355_, _03810_);
  nor (_19357_, _12603_, _08558_);
  nor (_19358_, _19357_, _19343_);
  nor (_19360_, _19358_, _03810_);
  or (_19361_, _19360_, _19356_);
  and (_19362_, _19361_, _02881_);
  nor (_19363_, _05328_, _19342_);
  and (_19364_, _12618_, _05328_);
  nor (_19365_, _19364_, _19363_);
  nor (_19366_, _19365_, _02881_);
  or (_19367_, _19366_, _03069_);
  or (_19368_, _19367_, _19362_);
  and (_19369_, _04693_, _04770_);
  nor (_19371_, _19369_, _19343_);
  nand (_19372_, _19371_, _03069_);
  and (_19373_, _19372_, _19368_);
  and (_19374_, _19373_, _03084_);
  nor (_19375_, _19352_, _03084_);
  or (_19376_, _19375_, _19374_);
  and (_19377_, _19376_, _02877_);
  and (_19378_, _12616_, _05328_);
  nor (_19379_, _19378_, _19363_);
  nor (_19380_, _19379_, _02877_);
  or (_19382_, _19380_, _02869_);
  or (_19383_, _19382_, _19377_);
  nor (_19384_, _19363_, _12646_);
  nor (_19385_, _19384_, _19365_);
  or (_19386_, _19385_, _02870_);
  and (_19387_, _19386_, _02864_);
  and (_19388_, _19387_, _19383_);
  nor (_19389_, _12664_, _08542_);
  nor (_19390_, _19389_, _19363_);
  nor (_19391_, _19390_, _02864_);
  nor (_19393_, _19391_, _06770_);
  not (_19394_, _19393_);
  nor (_19395_, _19394_, _19388_);
  and (_19396_, _19371_, _06770_);
  or (_19397_, _19396_, _02853_);
  nor (_19398_, _19397_, _19395_);
  or (_19399_, _19398_, _19350_);
  and (_19400_, _19399_, _02838_);
  nor (_19401_, _12722_, _08558_);
  nor (_19402_, _19401_, _19343_);
  nor (_19404_, _19402_, _02838_);
  or (_19405_, _19404_, _02802_);
  or (_19406_, _19405_, _19400_);
  and (_19407_, _12729_, _04693_);
  nor (_19408_, _19407_, _19343_);
  nand (_19409_, _19408_, _02802_);
  and (_19410_, _19409_, _19406_);
  and (_19411_, _19410_, _03887_);
  and (_19412_, _12739_, _04693_);
  nor (_19413_, _19412_, _19343_);
  nor (_19415_, _19413_, _03887_);
  or (_19416_, _19415_, _19411_);
  and (_19417_, _19416_, _03128_);
  nor (_19418_, _19417_, _19346_);
  nor (_19419_, _19418_, _02970_);
  nor (_19420_, _19343_, _04819_);
  not (_19421_, _19420_);
  nor (_19422_, _19408_, _03883_);
  and (_19423_, _19422_, _19421_);
  nor (_19424_, _19423_, _19419_);
  nor (_19426_, _19424_, _03135_);
  nor (_19427_, _19352_, _03137_);
  and (_19428_, _19427_, _19421_);
  or (_19429_, _19428_, _19426_);
  and (_19430_, _19429_, _05783_);
  nor (_19431_, _12737_, _08558_);
  nor (_19432_, _19431_, _19343_);
  nor (_19433_, _19432_, _05783_);
  or (_19434_, _19433_, _19430_);
  and (_19435_, _19434_, _05788_);
  nor (_19437_, _12612_, _08558_);
  nor (_19438_, _19437_, _19343_);
  nor (_19439_, _19438_, _05788_);
  or (_19440_, _19439_, _19435_);
  and (_19441_, _19440_, _03906_);
  nor (_19442_, _19358_, _03906_);
  or (_19443_, _19442_, _19441_);
  and (_19444_, _19443_, _02498_);
  nor (_19445_, _19379_, _02498_);
  or (_19446_, _19445_, _19444_);
  and (_19448_, _19446_, _02890_);
  and (_19449_, _12794_, _04693_);
  nor (_19450_, _19449_, _19343_);
  nor (_19451_, _19450_, _02890_);
  or (_19452_, _19451_, _19448_);
  or (_19453_, _19452_, _42672_);
  or (_19454_, _42668_, \oc8051_golden_model_1.IP [6]);
  and (_19455_, _19454_, _43998_);
  and (_43461_, _19455_, _19453_);
  not (_19456_, \oc8051_golden_model_1.P0 [0]);
  nor (_19458_, _42668_, _19456_);
  or (_19459_, _19458_, rst);
  nor (_19460_, _04628_, _19456_);
  and (_19461_, _11522_, _04628_);
  or (_19462_, _19461_, _19460_);
  and (_19463_, _19462_, _03127_);
  and (_19464_, _04628_, _03808_);
  or (_19465_, _19464_, _19460_);
  or (_19466_, _19465_, _05535_);
  and (_19467_, _05226_, _04628_);
  or (_19469_, _19467_, _19460_);
  or (_19470_, _19469_, _03810_);
  and (_19471_, _04628_, \oc8051_golden_model_1.ACC [0]);
  or (_19472_, _19471_, _19460_);
  and (_19473_, _19472_, _03813_);
  nor (_19474_, _03813_, _19456_);
  or (_19475_, _19474_, _02974_);
  or (_19476_, _19475_, _19473_);
  and (_19477_, _19476_, _02881_);
  and (_19478_, _19477_, _19470_);
  nor (_19480_, _04609_, _19456_);
  and (_19481_, _11417_, _04609_);
  or (_19482_, _19481_, _19480_);
  and (_19483_, _19482_, _02880_);
  or (_19484_, _19483_, _19478_);
  and (_19485_, _19484_, _03336_);
  and (_19486_, _19465_, _03069_);
  or (_19487_, _19486_, _03075_);
  or (_19488_, _19487_, _19485_);
  or (_19489_, _19472_, _03084_);
  and (_19491_, _19489_, _02877_);
  and (_19492_, _19491_, _19488_);
  and (_19493_, _19460_, _02876_);
  or (_19494_, _19493_, _02869_);
  or (_19495_, _19494_, _19492_);
  or (_19496_, _19469_, _02870_);
  and (_19497_, _19496_, _02864_);
  and (_19498_, _19497_, _19495_);
  or (_19499_, _11447_, _11405_);
  and (_19500_, _19499_, _04609_);
  or (_19502_, _19500_, _19480_);
  and (_19503_, _19502_, _02863_);
  or (_19504_, _19503_, _06770_);
  or (_19505_, _19504_, _19498_);
  and (_19506_, _19505_, _19466_);
  or (_19507_, _19506_, _02853_);
  and (_19508_, _04628_, _06152_);
  or (_19509_, _19460_, _05540_);
  or (_19510_, _19509_, _19508_);
  and (_19511_, _19510_, _02838_);
  and (_19513_, _19511_, _19507_);
  and (_19514_, _05710_, \oc8051_golden_model_1.P0 [0]);
  and (_19515_, _05717_, \oc8051_golden_model_1.P1 [0]);
  and (_19516_, _05720_, \oc8051_golden_model_1.P2 [0]);
  and (_19517_, _08669_, \oc8051_golden_model_1.P3 [0]);
  or (_19518_, _19517_, _19516_);
  or (_19519_, _19518_, _19515_);
  nor (_19520_, _19519_, _19514_);
  and (_19521_, _19520_, _11467_);
  and (_19522_, _19521_, _11486_);
  nand (_19523_, _19522_, _11502_);
  or (_19524_, _19523_, _11460_);
  and (_19525_, _19524_, _04628_);
  or (_19526_, _19525_, _19460_);
  and (_19527_, _19526_, _02579_);
  or (_19528_, _19527_, _02802_);
  or (_19529_, _19528_, _19513_);
  and (_19530_, _04628_, _05672_);
  or (_19531_, _19530_, _19460_);
  or (_19532_, _19531_, _02803_);
  and (_19534_, _19532_, _19529_);
  or (_19535_, _19534_, _02980_);
  and (_19536_, _11399_, _04628_);
  or (_19537_, _19460_, _03887_);
  or (_19538_, _19537_, _19536_);
  and (_19539_, _19538_, _03128_);
  and (_19540_, _19539_, _19535_);
  or (_19541_, _19540_, _19463_);
  and (_19542_, _19541_, _03883_);
  nand (_19543_, _19531_, _02970_);
  nor (_19545_, _19543_, _19467_);
  or (_19546_, _19545_, _19542_);
  and (_19547_, _19546_, _03137_);
  or (_19548_, _19460_, _09409_);
  and (_19549_, _19472_, _03135_);
  and (_19550_, _19549_, _19548_);
  or (_19551_, _19550_, _02965_);
  or (_19552_, _19551_, _19547_);
  nor (_19553_, _11396_, _08705_);
  or (_19554_, _19460_, _05783_);
  or (_19556_, _19554_, _19553_);
  and (_19557_, _19556_, _05788_);
  and (_19558_, _19557_, _19552_);
  nor (_19559_, _11520_, _08705_);
  or (_19560_, _19559_, _19460_);
  and (_19561_, _19560_, _03123_);
  or (_19562_, _19561_, _03163_);
  or (_19563_, _19562_, _19558_);
  or (_19564_, _19469_, _03906_);
  and (_19565_, _19564_, _02498_);
  and (_19566_, _19565_, _19563_);
  and (_19567_, _19460_, _02497_);
  or (_19568_, _19567_, _02888_);
  or (_19569_, _19568_, _19566_);
  or (_19570_, _19469_, _02890_);
  and (_19571_, _19570_, _42668_);
  and (_19572_, _19571_, _19569_);
  or (_43462_, _19572_, _19459_);
  not (_19573_, \oc8051_golden_model_1.P0 [1]);
  nor (_19574_, _42668_, _19573_);
  or (_19576_, _19574_, rst);
  nand (_19577_, _04628_, _03698_);
  or (_19578_, _04628_, \oc8051_golden_model_1.P0 [1]);
  and (_19579_, _19578_, _02802_);
  and (_19580_, _19579_, _19577_);
  nor (_19581_, _04628_, _19573_);
  and (_19582_, _04628_, _04000_);
  or (_19583_, _19582_, _19581_);
  or (_19584_, _19583_, _03336_);
  and (_19585_, _11606_, _04628_);
  not (_19586_, _19585_);
  and (_19587_, _19586_, _19578_);
  or (_19588_, _19587_, _03810_);
  nand (_19589_, _04628_, _02551_);
  and (_19590_, _19589_, _19578_);
  and (_19591_, _19590_, _03813_);
  nor (_19592_, _03813_, _19573_);
  or (_19593_, _19592_, _02974_);
  or (_19594_, _19593_, _19591_);
  and (_19595_, _19594_, _02881_);
  and (_19597_, _19595_, _19588_);
  nor (_19598_, _04609_, _19573_);
  and (_19599_, _11592_, _04609_);
  or (_19600_, _19599_, _19598_);
  and (_19601_, _19600_, _02880_);
  or (_19602_, _19601_, _03069_);
  or (_19603_, _19602_, _19597_);
  and (_19604_, _19603_, _19584_);
  or (_19605_, _19604_, _03075_);
  or (_19606_, _19590_, _03084_);
  and (_19608_, _19606_, _02877_);
  and (_19609_, _19608_, _19605_);
  and (_19610_, _11595_, _04609_);
  or (_19611_, _19610_, _19598_);
  and (_19612_, _19611_, _02876_);
  or (_19613_, _19612_, _02869_);
  or (_19614_, _19613_, _19609_);
  and (_19615_, _19599_, _11591_);
  or (_19616_, _19598_, _02870_);
  or (_19617_, _19616_, _19615_);
  and (_19618_, _19617_, _19614_);
  and (_19619_, _19618_, _02864_);
  or (_19620_, _11637_, _11595_);
  and (_19621_, _19620_, _04609_);
  or (_19622_, _19598_, _19621_);
  and (_19623_, _19622_, _02863_);
  or (_19624_, _19623_, _06770_);
  or (_19625_, _19624_, _19619_);
  or (_19626_, _19583_, _05535_);
  and (_19627_, _19626_, _19625_);
  or (_19629_, _19627_, _02853_);
  and (_19630_, _04628_, _06151_);
  or (_19631_, _19581_, _05540_);
  or (_19632_, _19631_, _19630_);
  and (_19633_, _19632_, _02838_);
  and (_19634_, _19633_, _19629_);
  and (_19635_, _05710_, \oc8051_golden_model_1.P0 [1]);
  and (_19636_, _05717_, \oc8051_golden_model_1.P1 [1]);
  and (_19637_, _05720_, \oc8051_golden_model_1.P2 [1]);
  and (_19638_, _08669_, \oc8051_golden_model_1.P3 [1]);
  or (_19640_, _19638_, _19637_);
  or (_19641_, _19640_, _19636_);
  nor (_19642_, _19641_, _19635_);
  and (_19643_, _19642_, _11662_);
  and (_19644_, _19643_, _11676_);
  nand (_19645_, _19644_, _11692_);
  or (_19646_, _19645_, _11650_);
  and (_19647_, _19646_, _04628_);
  or (_19648_, _19647_, _19581_);
  and (_19649_, _19648_, _02579_);
  or (_19650_, _19649_, _19634_);
  and (_19651_, _19650_, _02803_);
  or (_19652_, _19651_, _19580_);
  and (_19653_, _19652_, _03887_);
  or (_19654_, _11710_, _08705_);
  and (_19655_, _19578_, _02980_);
  and (_19656_, _19655_, _19654_);
  or (_19657_, _19656_, _19653_);
  and (_19658_, _19657_, _03128_);
  or (_19659_, _11715_, _08705_);
  and (_19661_, _19578_, _03127_);
  and (_19662_, _19661_, _19659_);
  or (_19663_, _19662_, _19658_);
  and (_19664_, _19663_, _03883_);
  or (_19665_, _11709_, _08705_);
  and (_19666_, _19578_, _02970_);
  and (_19667_, _19666_, _19665_);
  or (_19668_, _19667_, _19664_);
  and (_19669_, _19668_, _03137_);
  or (_19670_, _19581_, _13722_);
  and (_19672_, _19590_, _03135_);
  and (_19673_, _19672_, _19670_);
  or (_19674_, _19673_, _19669_);
  and (_19675_, _19674_, _03124_);
  or (_19676_, _19577_, _13722_);
  and (_19677_, _19578_, _02965_);
  and (_19678_, _19677_, _19676_);
  or (_19679_, _19589_, _13722_);
  and (_19680_, _19578_, _03123_);
  and (_19681_, _19680_, _19679_);
  or (_19682_, _19681_, _03163_);
  or (_19683_, _19682_, _19678_);
  or (_19684_, _19683_, _19675_);
  or (_19685_, _19587_, _03906_);
  and (_19686_, _19685_, _02498_);
  and (_19687_, _19686_, _19684_);
  and (_19688_, _19611_, _02497_);
  or (_19689_, _19688_, _02888_);
  or (_19690_, _19689_, _19687_);
  or (_19691_, _19581_, _02890_);
  or (_19693_, _19691_, _19585_);
  and (_19694_, _19693_, _42668_);
  and (_19695_, _19694_, _19690_);
  or (_43463_, _19695_, _19576_);
  not (_19696_, \oc8051_golden_model_1.P0 [2]);
  nor (_19697_, _42668_, _19696_);
  or (_19698_, _19697_, rst);
  nor (_19699_, _04628_, _19696_);
  and (_19700_, _11927_, _04628_);
  or (_19701_, _19700_, _19699_);
  and (_19703_, _19701_, _03127_);
  and (_19704_, _04628_, _04435_);
  or (_19705_, _19704_, _19699_);
  or (_19706_, _19705_, _05535_);
  and (_19707_, _19705_, _03069_);
  nor (_19708_, _04609_, _19696_);
  and (_19709_, _11815_, _04609_);
  or (_19710_, _19709_, _19708_);
  or (_19711_, _19710_, _02881_);
  nor (_19712_, _11801_, _08705_);
  or (_19713_, _19712_, _19699_);
  and (_19714_, _19713_, _02974_);
  nor (_19715_, _03813_, _19696_);
  and (_19716_, _04628_, \oc8051_golden_model_1.ACC [2]);
  or (_19717_, _19716_, _19699_);
  and (_19718_, _19717_, _03813_);
  or (_19719_, _19718_, _19715_);
  and (_19720_, _19719_, _03810_);
  or (_19721_, _19720_, _02880_);
  or (_19722_, _19721_, _19714_);
  and (_19724_, _19722_, _19711_);
  and (_19725_, _19724_, _03336_);
  or (_19726_, _19725_, _19707_);
  or (_19727_, _19726_, _03075_);
  or (_19728_, _19717_, _03084_);
  and (_19729_, _19728_, _02877_);
  and (_19730_, _19729_, _19727_);
  and (_19731_, _11797_, _04609_);
  or (_19732_, _19731_, _19708_);
  and (_19733_, _19732_, _02876_);
  or (_19735_, _19733_, _02869_);
  or (_19736_, _19735_, _19730_);
  or (_19737_, _19708_, _11830_);
  and (_19738_, _19737_, _19710_);
  or (_19739_, _19738_, _02870_);
  and (_19740_, _19739_, _02864_);
  and (_19741_, _19740_, _19736_);
  or (_19742_, _11847_, _11797_);
  and (_19743_, _19742_, _04609_);
  or (_19744_, _19743_, _19708_);
  and (_19745_, _19744_, _02863_);
  or (_19746_, _19745_, _06770_);
  or (_19747_, _19746_, _19741_);
  and (_19748_, _19747_, _19706_);
  or (_19749_, _19748_, _02853_);
  and (_19750_, _04628_, _06155_);
  or (_19751_, _19699_, _05540_);
  or (_19752_, _19751_, _19750_);
  and (_19753_, _19752_, _02838_);
  and (_19754_, _19753_, _19749_);
  and (_19756_, _05717_, \oc8051_golden_model_1.P1 [2]);
  and (_19757_, _05710_, \oc8051_golden_model_1.P0 [2]);
  and (_19758_, _05720_, \oc8051_golden_model_1.P2 [2]);
  and (_19759_, _08669_, \oc8051_golden_model_1.P3 [2]);
  or (_19760_, _19759_, _19758_);
  or (_19761_, _19760_, _19757_);
  or (_19762_, _19761_, _19756_);
  nor (_19763_, _19762_, _11877_);
  and (_19764_, _19763_, _11903_);
  nand (_19765_, _19764_, _11876_);
  or (_19767_, _19765_, _11860_);
  and (_19768_, _19767_, _04628_);
  or (_19769_, _19768_, _19699_);
  and (_19770_, _19769_, _02579_);
  or (_19771_, _19770_, _02802_);
  or (_19772_, _19771_, _19754_);
  and (_19773_, _04628_, _05701_);
  or (_19774_, _19773_, _19699_);
  or (_19775_, _19774_, _02803_);
  and (_19776_, _19775_, _19772_);
  or (_19777_, _19776_, _02980_);
  and (_19778_, _11921_, _04628_);
  or (_19779_, _19699_, _03887_);
  or (_19780_, _19779_, _19778_);
  and (_19781_, _19780_, _03128_);
  and (_19782_, _19781_, _19777_);
  or (_19783_, _19782_, _19703_);
  and (_19784_, _19783_, _03883_);
  or (_19785_, _19699_, _05130_);
  and (_19786_, _19774_, _02970_);
  and (_19788_, _19786_, _19785_);
  or (_19789_, _19788_, _19784_);
  and (_19790_, _19789_, _03137_);
  and (_19791_, _19717_, _03135_);
  and (_19792_, _19791_, _19785_);
  or (_19793_, _19792_, _02965_);
  or (_19794_, _19793_, _19790_);
  nor (_19795_, _11919_, _08705_);
  or (_19796_, _19699_, _05783_);
  or (_19797_, _19796_, _19795_);
  and (_19799_, _19797_, _05788_);
  and (_19800_, _19799_, _19794_);
  nor (_19801_, _11926_, _08705_);
  or (_19802_, _19801_, _19699_);
  and (_19803_, _19802_, _03123_);
  or (_19804_, _19803_, _03163_);
  or (_19805_, _19804_, _19800_);
  or (_19806_, _19713_, _03906_);
  and (_19807_, _19806_, _02498_);
  and (_19808_, _19807_, _19805_);
  and (_19809_, _19732_, _02497_);
  or (_19810_, _19809_, _02888_);
  or (_19811_, _19810_, _19808_);
  and (_19812_, _11985_, _04628_);
  or (_19813_, _19699_, _02890_);
  or (_19814_, _19813_, _19812_);
  and (_19815_, _19814_, _42668_);
  and (_19816_, _19815_, _19811_);
  or (_43465_, _19816_, _19698_);
  not (_19817_, \oc8051_golden_model_1.P0 [3]);
  nor (_19819_, _42668_, _19817_);
  or (_19820_, _19819_, rst);
  nor (_19821_, _04628_, _19817_);
  and (_19822_, _12133_, _04628_);
  or (_19823_, _19822_, _19821_);
  and (_19824_, _19823_, _03127_);
  and (_19825_, _04628_, _04241_);
  or (_19826_, _19825_, _19821_);
  or (_19827_, _19826_, _05535_);
  nor (_19828_, _12017_, _08705_);
  or (_19830_, _19828_, _19821_);
  or (_19831_, _19830_, _03810_);
  and (_19832_, _04628_, \oc8051_golden_model_1.ACC [3]);
  or (_19833_, _19832_, _19821_);
  and (_19834_, _19833_, _03813_);
  nor (_19835_, _03813_, _19817_);
  or (_19836_, _19835_, _02974_);
  or (_19837_, _19836_, _19834_);
  and (_19838_, _19837_, _02881_);
  and (_19839_, _19838_, _19831_);
  nor (_19840_, _04609_, _19817_);
  and (_19841_, _12021_, _04609_);
  or (_19842_, _19841_, _19840_);
  and (_19843_, _19842_, _02880_);
  or (_19844_, _19843_, _03069_);
  or (_19845_, _19844_, _19839_);
  or (_19846_, _19826_, _03336_);
  and (_19847_, _19846_, _19845_);
  or (_19848_, _19847_, _03075_);
  or (_19849_, _19833_, _03084_);
  and (_19851_, _19849_, _02877_);
  and (_19852_, _19851_, _19848_);
  and (_19853_, _12005_, _04609_);
  or (_19854_, _19853_, _19840_);
  and (_19855_, _19854_, _02876_);
  or (_19856_, _19855_, _02869_);
  or (_19857_, _19856_, _19852_);
  or (_19858_, _19840_, _12036_);
  and (_19859_, _19858_, _19842_);
  or (_19860_, _19859_, _02870_);
  and (_19862_, _19860_, _02864_);
  and (_19863_, _19862_, _19857_);
  or (_19864_, _12005_, _12052_);
  and (_19865_, _19864_, _04609_);
  or (_19866_, _19865_, _19840_);
  and (_19867_, _19866_, _02863_);
  or (_19868_, _19867_, _06770_);
  or (_19869_, _19868_, _19863_);
  and (_19870_, _19869_, _19827_);
  or (_19871_, _19870_, _02853_);
  and (_19872_, _04628_, _06154_);
  or (_19873_, _19821_, _05540_);
  or (_19874_, _19873_, _19872_);
  and (_19875_, _19874_, _02838_);
  and (_19876_, _19875_, _19871_);
  and (_19877_, _05717_, \oc8051_golden_model_1.P1 [3]);
  and (_19878_, _05710_, \oc8051_golden_model_1.P0 [3]);
  and (_19879_, _05720_, \oc8051_golden_model_1.P2 [3]);
  and (_19880_, _08669_, \oc8051_golden_model_1.P3 [3]);
  or (_19881_, _19880_, _19879_);
  or (_19883_, _19881_, _19878_);
  nor (_19884_, _19883_, _19877_);
  and (_19885_, _19884_, _12080_);
  and (_19886_, _19885_, _12094_);
  nand (_19887_, _19886_, _12110_);
  or (_19888_, _19887_, _12067_);
  and (_19889_, _19888_, _04628_);
  or (_19890_, _19889_, _19821_);
  and (_19891_, _19890_, _02579_);
  or (_19892_, _19891_, _02802_);
  or (_19894_, _19892_, _19876_);
  and (_19895_, _04628_, _05658_);
  or (_19896_, _19895_, _19821_);
  or (_19897_, _19896_, _02803_);
  and (_19898_, _19897_, _19894_);
  or (_19899_, _19898_, _02980_);
  and (_19900_, _12127_, _04628_);
  or (_19901_, _19821_, _03887_);
  or (_19902_, _19901_, _19900_);
  and (_19903_, _19902_, _03128_);
  and (_19904_, _19903_, _19899_);
  or (_19905_, _19904_, _19824_);
  and (_19906_, _19905_, _03883_);
  or (_19907_, _19821_, _05079_);
  and (_19908_, _19896_, _02970_);
  and (_19909_, _19908_, _19907_);
  or (_19910_, _19909_, _19906_);
  and (_19911_, _19910_, _03137_);
  and (_19912_, _19833_, _03135_);
  and (_19913_, _19912_, _19907_);
  or (_19915_, _19913_, _02965_);
  or (_19916_, _19915_, _19911_);
  nor (_19917_, _12125_, _08705_);
  or (_19918_, _19821_, _05783_);
  or (_19919_, _19918_, _19917_);
  and (_19920_, _19919_, _05788_);
  and (_19921_, _19920_, _19916_);
  nor (_19922_, _12132_, _08705_);
  or (_19923_, _19922_, _19821_);
  and (_19924_, _19923_, _03123_);
  or (_19926_, _19924_, _03163_);
  or (_19927_, _19926_, _19921_);
  or (_19928_, _19830_, _03906_);
  and (_19929_, _19928_, _02498_);
  and (_19930_, _19929_, _19927_);
  and (_19931_, _19854_, _02497_);
  or (_19932_, _19931_, _02888_);
  or (_19933_, _19932_, _19930_);
  and (_19934_, _12183_, _04628_);
  or (_19935_, _19821_, _02890_);
  or (_19937_, _19935_, _19934_);
  and (_19938_, _19937_, _42668_);
  and (_19939_, _19938_, _19933_);
  or (_43466_, _19939_, _19820_);
  not (_19940_, \oc8051_golden_model_1.P0 [4]);
  nor (_19941_, _42668_, _19940_);
  or (_19942_, _19941_, rst);
  nor (_19943_, _04628_, _19940_);
  and (_19944_, _12207_, _04628_);
  or (_19945_, _19944_, _19943_);
  and (_19946_, _19945_, _03127_);
  and (_19947_, _04628_, _04982_);
  or (_19948_, _19947_, _19943_);
  or (_19949_, _19948_, _05535_);
  nor (_19950_, _04609_, _19940_);
  and (_19951_, _12213_, _04609_);
  or (_19952_, _19951_, _19950_);
  and (_19953_, _19952_, _02876_);
  nor (_19954_, _12217_, _08705_);
  or (_19955_, _19954_, _19943_);
  or (_19957_, _19955_, _03810_);
  and (_19958_, _04628_, \oc8051_golden_model_1.ACC [4]);
  or (_19959_, _19958_, _19943_);
  and (_19960_, _19959_, _03813_);
  nor (_19961_, _03813_, _19940_);
  or (_19962_, _19961_, _02974_);
  or (_19963_, _19962_, _19960_);
  and (_19964_, _19963_, _02881_);
  and (_19965_, _19964_, _19957_);
  and (_19966_, _12231_, _04609_);
  or (_19968_, _19966_, _19950_);
  and (_19969_, _19968_, _02880_);
  or (_19970_, _19969_, _03069_);
  or (_19971_, _19970_, _19965_);
  or (_19972_, _19948_, _03336_);
  and (_19973_, _19972_, _19971_);
  or (_19974_, _19973_, _03075_);
  or (_19975_, _19959_, _03084_);
  and (_19976_, _19975_, _02877_);
  and (_19977_, _19976_, _19974_);
  or (_19978_, _19977_, _19953_);
  and (_19979_, _19978_, _02870_);
  or (_19980_, _19950_, _12246_);
  and (_19981_, _19980_, _02869_);
  and (_19982_, _19981_, _19968_);
  or (_19983_, _19982_, _19979_);
  and (_19984_, _19983_, _02864_);
  or (_19985_, _12263_, _12213_);
  and (_19986_, _19985_, _04609_);
  or (_19987_, _19986_, _19950_);
  and (_19989_, _19987_, _02863_);
  or (_19990_, _19989_, _06770_);
  or (_19991_, _19990_, _19984_);
  and (_19992_, _19991_, _19949_);
  or (_19993_, _19992_, _02853_);
  and (_19994_, _04628_, _06159_);
  or (_19995_, _19943_, _05540_);
  or (_19996_, _19995_, _19994_);
  and (_19997_, _19996_, _02838_);
  and (_19998_, _19997_, _19993_);
  and (_20000_, _05710_, \oc8051_golden_model_1.P0 [4]);
  and (_20001_, _05717_, \oc8051_golden_model_1.P1 [4]);
  and (_20002_, _05720_, \oc8051_golden_model_1.P2 [4]);
  and (_20003_, _08669_, \oc8051_golden_model_1.P3 [4]);
  or (_20004_, _20003_, _20002_);
  or (_20005_, _20004_, _20001_);
  nor (_20006_, _20005_, _20000_);
  and (_20007_, _20006_, _12290_);
  and (_20008_, _20007_, _12285_);
  nand (_20009_, _20008_, _12319_);
  or (_20011_, _20009_, _12277_);
  and (_20012_, _20011_, _04628_);
  or (_20013_, _20012_, _19943_);
  and (_20014_, _20013_, _02579_);
  or (_20015_, _20014_, _02802_);
  or (_20016_, _20015_, _19998_);
  and (_20017_, _05666_, _04628_);
  or (_20018_, _20017_, _19943_);
  or (_20019_, _20018_, _02803_);
  and (_20020_, _20019_, _20016_);
  or (_20021_, _20020_, _02980_);
  and (_20022_, _12211_, _04628_);
  or (_20023_, _19943_, _03887_);
  or (_20024_, _20023_, _20022_);
  and (_20025_, _20024_, _03128_);
  and (_20026_, _20025_, _20021_);
  or (_20027_, _20026_, _19946_);
  and (_20028_, _20027_, _03883_);
  or (_20029_, _19943_, _05031_);
  and (_20030_, _20018_, _02970_);
  and (_20032_, _20030_, _20029_);
  or (_20033_, _20032_, _20028_);
  and (_20034_, _20033_, _03137_);
  and (_20035_, _19959_, _03135_);
  and (_20036_, _20035_, _20029_);
  or (_20037_, _20036_, _02965_);
  or (_20038_, _20037_, _20034_);
  nor (_20039_, _12209_, _08705_);
  or (_20040_, _19943_, _05783_);
  or (_20041_, _20040_, _20039_);
  and (_20043_, _20041_, _05788_);
  and (_20044_, _20043_, _20038_);
  nor (_20045_, _12206_, _08705_);
  or (_20046_, _20045_, _19943_);
  and (_20047_, _20046_, _03123_);
  or (_20048_, _20047_, _03163_);
  or (_20049_, _20048_, _20044_);
  or (_20050_, _19955_, _03906_);
  and (_20051_, _20050_, _02498_);
  and (_20052_, _20051_, _20049_);
  and (_20053_, _19952_, _02497_);
  or (_20054_, _20053_, _02888_);
  or (_20055_, _20054_, _20052_);
  and (_20056_, _12389_, _04628_);
  or (_20057_, _19943_, _02890_);
  or (_20058_, _20057_, _20056_);
  and (_20059_, _20058_, _42668_);
  and (_20060_, _20059_, _20055_);
  or (_43467_, _20060_, _19942_);
  not (_20061_, \oc8051_golden_model_1.P0 [5]);
  nor (_20063_, _42668_, _20061_);
  or (_20064_, _20063_, rst);
  nor (_20065_, _04628_, _20061_);
  and (_20066_, _12411_, _04628_);
  or (_20067_, _20066_, _20065_);
  and (_20068_, _20067_, _03127_);
  nor (_20069_, _12407_, _08705_);
  or (_20070_, _20069_, _20065_);
  or (_20071_, _20070_, _03810_);
  and (_20072_, _04628_, \oc8051_golden_model_1.ACC [5]);
  or (_20074_, _20072_, _20065_);
  and (_20075_, _20074_, _03813_);
  nor (_20076_, _03813_, _20061_);
  or (_20077_, _20076_, _02974_);
  or (_20078_, _20077_, _20075_);
  and (_20079_, _20078_, _02881_);
  and (_20080_, _20079_, _20071_);
  nor (_20081_, _04609_, _20061_);
  and (_20082_, _12435_, _04609_);
  or (_20083_, _20082_, _20081_);
  and (_20085_, _20083_, _02880_);
  or (_20086_, _20085_, _03069_);
  or (_20087_, _20086_, _20080_);
  and (_20088_, _04628_, _04877_);
  or (_20089_, _20088_, _20065_);
  or (_20090_, _20089_, _03336_);
  and (_20091_, _20090_, _20087_);
  or (_20092_, _20091_, _03075_);
  or (_20093_, _20074_, _03084_);
  and (_20094_, _20093_, _02877_);
  and (_20096_, _20094_, _20092_);
  and (_20097_, _12417_, _04609_);
  or (_20098_, _20097_, _20081_);
  and (_20099_, _20098_, _02876_);
  or (_20100_, _20099_, _02869_);
  or (_20101_, _20100_, _20096_);
  or (_20102_, _20081_, _12450_);
  and (_20103_, _20102_, _20083_);
  or (_20104_, _20103_, _02870_);
  and (_20105_, _20104_, _02864_);
  and (_20107_, _20105_, _20101_);
  or (_20108_, _12467_, _12417_);
  and (_20109_, _20108_, _04609_);
  or (_20110_, _20109_, _20081_);
  and (_20111_, _20110_, _02863_);
  or (_20112_, _20111_, _06770_);
  or (_20113_, _20112_, _20107_);
  or (_20114_, _20089_, _05535_);
  and (_20115_, _20114_, _20113_);
  or (_20116_, _20115_, _02853_);
  and (_20118_, _04628_, _06158_);
  or (_20119_, _20065_, _05540_);
  or (_20120_, _20119_, _20118_);
  and (_20121_, _20120_, _02838_);
  and (_20122_, _20121_, _20116_);
  and (_20123_, _05717_, \oc8051_golden_model_1.P1 [5]);
  and (_20124_, _05710_, \oc8051_golden_model_1.P0 [5]);
  and (_20125_, _05720_, \oc8051_golden_model_1.P2 [5]);
  or (_20126_, _20125_, _20124_);
  nor (_20127_, _20126_, _20123_);
  nand (_20129_, _20127_, _12489_);
  not (_20130_, _12494_);
  and (_20131_, _12513_, _20130_);
  nand (_20132_, _20131_, _12509_);
  or (_20133_, _12518_, _12520_);
  and (_20134_, _05714_, \oc8051_golden_model_1.P3 [5]);
  or (_20135_, _20134_, _12491_);
  or (_20136_, _20135_, _20133_);
  nor (_20137_, _12493_, _12490_);
  nand (_20138_, _20137_, _12516_);
  or (_20140_, _20138_, _20136_);
  or (_20141_, _20140_, _20132_);
  or (_20142_, _20141_, _20129_);
  or (_20143_, _20142_, _12481_);
  and (_20144_, _20143_, _04628_);
  or (_20145_, _20144_, _20065_);
  and (_20146_, _20145_, _02579_);
  or (_20147_, _20146_, _02802_);
  or (_20148_, _20147_, _20122_);
  and (_20149_, _05614_, _04628_);
  or (_20151_, _20149_, _20065_);
  or (_20152_, _20151_, _02803_);
  and (_20153_, _20152_, _20148_);
  or (_20154_, _20153_, _02980_);
  and (_20155_, _12415_, _04628_);
  or (_20156_, _20065_, _03887_);
  or (_20157_, _20156_, _20155_);
  and (_20158_, _20157_, _03128_);
  and (_20159_, _20158_, _20154_);
  or (_20160_, _20159_, _20068_);
  and (_20161_, _20160_, _03883_);
  or (_20162_, _20065_, _04924_);
  and (_20163_, _20151_, _02970_);
  and (_20164_, _20163_, _20162_);
  or (_20165_, _20164_, _20161_);
  and (_20166_, _20165_, _03137_);
  and (_20167_, _20074_, _03135_);
  and (_20168_, _20167_, _20162_);
  or (_20169_, _20168_, _02965_);
  or (_20170_, _20169_, _20166_);
  nor (_20171_, _12413_, _08705_);
  or (_20172_, _20065_, _05783_);
  or (_20173_, _20172_, _20171_);
  and (_20174_, _20173_, _05788_);
  and (_20175_, _20174_, _20170_);
  nor (_20176_, _12410_, _08705_);
  or (_20177_, _20176_, _20065_);
  and (_20178_, _20177_, _03123_);
  or (_20179_, _20178_, _03163_);
  or (_20180_, _20179_, _20175_);
  or (_20182_, _20070_, _03906_);
  and (_20183_, _20182_, _02498_);
  and (_20184_, _20183_, _20180_);
  and (_20185_, _20098_, _02497_);
  or (_20186_, _20185_, _02888_);
  or (_20187_, _20186_, _20184_);
  and (_20188_, _12589_, _04628_);
  or (_20189_, _20065_, _02890_);
  or (_20190_, _20189_, _20188_);
  and (_20191_, _20190_, _42668_);
  and (_20193_, _20191_, _20187_);
  or (_43468_, _20193_, _20064_);
  not (_20194_, \oc8051_golden_model_1.P0 [6]);
  nor (_20195_, _42668_, _20194_);
  or (_20196_, _20195_, rst);
  nor (_20197_, _04628_, _20194_);
  and (_20198_, _12613_, _04628_);
  or (_20199_, _20198_, _20197_);
  and (_20200_, _20199_, _03127_);
  nor (_20201_, _12603_, _08705_);
  or (_20203_, _20201_, _20197_);
  or (_20204_, _20203_, _03810_);
  and (_20205_, _04628_, \oc8051_golden_model_1.ACC [6]);
  or (_20206_, _20205_, _20197_);
  and (_20207_, _20206_, _03813_);
  nor (_20208_, _03813_, _20194_);
  or (_20209_, _20208_, _02974_);
  or (_20210_, _20209_, _20207_);
  and (_20211_, _20210_, _02881_);
  and (_20212_, _20211_, _20204_);
  nor (_20214_, _04609_, _20194_);
  and (_20215_, _12618_, _04609_);
  or (_20216_, _20215_, _20214_);
  and (_20217_, _20216_, _02880_);
  or (_20218_, _20217_, _03069_);
  or (_20219_, _20218_, _20212_);
  and (_20220_, _04628_, _04770_);
  or (_20221_, _20220_, _20197_);
  or (_20222_, _20221_, _03336_);
  and (_20223_, _20222_, _20219_);
  or (_20225_, _20223_, _03075_);
  or (_20226_, _20206_, _03084_);
  and (_20227_, _20226_, _02877_);
  and (_20228_, _20227_, _20225_);
  and (_20229_, _12616_, _04609_);
  or (_20230_, _20229_, _20214_);
  and (_20231_, _20230_, _02876_);
  or (_20232_, _20231_, _02869_);
  or (_20233_, _20232_, _20228_);
  or (_20234_, _20214_, _12646_);
  and (_20236_, _20234_, _20216_);
  or (_20237_, _20236_, _02870_);
  and (_20238_, _20237_, _02864_);
  and (_20239_, _20238_, _20233_);
  or (_20240_, _12663_, _12616_);
  and (_20241_, _20240_, _04609_);
  or (_20242_, _20241_, _20214_);
  and (_20243_, _20242_, _02863_);
  or (_20244_, _20243_, _06770_);
  or (_20245_, _20244_, _20239_);
  or (_20247_, _20221_, _05535_);
  and (_20248_, _20247_, _20245_);
  or (_20249_, _20248_, _02853_);
  and (_20250_, _04628_, _05849_);
  or (_20251_, _20197_, _05540_);
  or (_20252_, _20251_, _20250_);
  and (_20253_, _20252_, _02838_);
  and (_20254_, _20253_, _20249_);
  and (_20255_, _05717_, \oc8051_golden_model_1.P1 [6]);
  and (_20256_, _05710_, \oc8051_golden_model_1.P0 [6]);
  and (_20258_, _05720_, \oc8051_golden_model_1.P2 [6]);
  and (_20259_, _08669_, \oc8051_golden_model_1.P3 [6]);
  or (_20260_, _20259_, _20258_);
  or (_20261_, _20260_, _20256_);
  or (_20262_, _20261_, _20255_);
  nor (_20263_, _20262_, _12699_);
  and (_20264_, _20263_, _12718_);
  and (_20265_, _20264_, _12698_);
  nand (_20266_, _20265_, _12691_);
  or (_20267_, _20266_, _12676_);
  and (_20269_, _20267_, _04628_);
  or (_20270_, _20269_, _20197_);
  and (_20271_, _20270_, _02579_);
  or (_20272_, _20271_, _02802_);
  or (_20273_, _20272_, _20254_);
  and (_20274_, _12729_, _04628_);
  or (_20275_, _20274_, _20197_);
  or (_20276_, _20275_, _02803_);
  and (_20277_, _20276_, _20273_);
  or (_20278_, _20277_, _02980_);
  and (_20280_, _12739_, _04628_);
  or (_20281_, _20197_, _03887_);
  or (_20282_, _20281_, _20280_);
  and (_20283_, _20282_, _03128_);
  and (_20284_, _20283_, _20278_);
  or (_20285_, _20284_, _20200_);
  and (_20286_, _20285_, _03883_);
  or (_20287_, _20197_, _04819_);
  and (_20288_, _20275_, _02970_);
  and (_20289_, _20288_, _20287_);
  or (_20291_, _20289_, _20286_);
  and (_20292_, _20291_, _03137_);
  and (_20293_, _20206_, _03135_);
  and (_20294_, _20293_, _20287_);
  or (_20295_, _20294_, _02965_);
  or (_20296_, _20295_, _20292_);
  nor (_20297_, _12737_, _08705_);
  or (_20298_, _20197_, _05783_);
  or (_20299_, _20298_, _20297_);
  and (_20300_, _20299_, _05788_);
  and (_20302_, _20300_, _20296_);
  nor (_20303_, _12612_, _08705_);
  or (_20304_, _20303_, _20197_);
  and (_20305_, _20304_, _03123_);
  or (_20306_, _20305_, _03163_);
  or (_20307_, _20306_, _20302_);
  or (_20308_, _20203_, _03906_);
  and (_20309_, _20308_, _02498_);
  and (_20310_, _20309_, _20307_);
  and (_20311_, _20230_, _02497_);
  or (_20313_, _20311_, _02888_);
  or (_20314_, _20313_, _20310_);
  and (_20315_, _12794_, _04628_);
  or (_20316_, _20197_, _02890_);
  or (_20317_, _20316_, _20315_);
  and (_20318_, _20317_, _42668_);
  and (_20319_, _20318_, _20314_);
  or (_43469_, _20319_, _20196_);
  not (_20320_, \oc8051_golden_model_1.P1 [0]);
  nor (_20321_, _42668_, _20320_);
  or (_20323_, _20321_, rst);
  nor (_20324_, _04634_, _20320_);
  and (_20325_, _11522_, _04634_);
  or (_20326_, _20325_, _20324_);
  and (_20327_, _20326_, _03127_);
  and (_20328_, _04634_, _03808_);
  or (_20329_, _20328_, _20324_);
  or (_20330_, _20329_, _05535_);
  and (_20331_, _05226_, _04634_);
  or (_20332_, _20331_, _20324_);
  and (_20334_, _20332_, _02974_);
  nor (_20335_, _03813_, _20320_);
  and (_20336_, _04634_, \oc8051_golden_model_1.ACC [0]);
  or (_20337_, _20336_, _20324_);
  and (_20338_, _20337_, _03813_);
  or (_20339_, _20338_, _20335_);
  and (_20340_, _20339_, _03810_);
  or (_20341_, _20340_, _02880_);
  or (_20342_, _20341_, _20334_);
  and (_20343_, _11417_, _05344_);
  nor (_20345_, _05344_, _20320_);
  or (_20346_, _20345_, _02881_);
  or (_20347_, _20346_, _20343_);
  and (_20348_, _20347_, _03336_);
  and (_20349_, _20348_, _20342_);
  and (_20350_, _20329_, _03069_);
  or (_20351_, _20350_, _03075_);
  or (_20352_, _20351_, _20349_);
  or (_20353_, _20337_, _03084_);
  and (_20354_, _20353_, _02877_);
  and (_20356_, _20354_, _20352_);
  and (_20357_, _20324_, _02876_);
  or (_20358_, _20357_, _02869_);
  or (_20359_, _20358_, _20356_);
  or (_20360_, _20332_, _02870_);
  and (_20361_, _20360_, _02864_);
  and (_20362_, _20361_, _20359_);
  and (_20363_, _19499_, _05344_);
  or (_20364_, _20363_, _20345_);
  and (_20365_, _20364_, _02863_);
  or (_20367_, _20365_, _06770_);
  or (_20368_, _20367_, _20362_);
  and (_20369_, _20368_, _20330_);
  or (_20370_, _20369_, _02853_);
  and (_20371_, _04634_, _06152_);
  or (_20372_, _20324_, _05540_);
  or (_20373_, _20372_, _20371_);
  and (_20374_, _20373_, _02838_);
  and (_20375_, _20374_, _20370_);
  and (_20376_, _19524_, _04634_);
  or (_20378_, _20376_, _20324_);
  and (_20379_, _20378_, _02579_);
  or (_20380_, _20379_, _02802_);
  or (_20381_, _20380_, _20375_);
  and (_20382_, _04634_, _05672_);
  or (_20383_, _20382_, _20324_);
  or (_20384_, _20383_, _02803_);
  and (_20385_, _20384_, _20381_);
  or (_20386_, _20385_, _02980_);
  and (_20387_, _11399_, _04634_);
  or (_20389_, _20324_, _03887_);
  or (_20390_, _20389_, _20387_);
  and (_20391_, _20390_, _03128_);
  and (_20392_, _20391_, _20386_);
  or (_20393_, _20392_, _20327_);
  and (_20394_, _20393_, _03883_);
  nand (_20395_, _20383_, _02970_);
  nor (_20396_, _20395_, _20331_);
  or (_20397_, _20396_, _20394_);
  and (_20398_, _20397_, _03137_);
  or (_20400_, _20324_, _09409_);
  and (_20401_, _20337_, _03135_);
  and (_20402_, _20401_, _20400_);
  or (_20403_, _20402_, _02965_);
  or (_20404_, _20403_, _20398_);
  nor (_20405_, _11396_, _08808_);
  or (_20406_, _20324_, _05783_);
  or (_20407_, _20406_, _20405_);
  and (_20408_, _20407_, _05788_);
  and (_20409_, _20408_, _20404_);
  nor (_20411_, _11520_, _08808_);
  or (_20412_, _20411_, _20324_);
  and (_20413_, _20412_, _03123_);
  or (_20414_, _20413_, _03163_);
  or (_20415_, _20414_, _20409_);
  or (_20416_, _20332_, _03906_);
  and (_20417_, _20416_, _02498_);
  and (_20418_, _20417_, _20415_);
  and (_20419_, _20324_, _02497_);
  or (_20420_, _20419_, _02888_);
  or (_20422_, _20420_, _20418_);
  or (_20423_, _20332_, _02890_);
  and (_20424_, _20423_, _42668_);
  and (_20425_, _20424_, _20422_);
  or (_43470_, _20425_, _20323_);
  not (_20426_, \oc8051_golden_model_1.P1 [1]);
  nor (_20427_, _42668_, _20426_);
  or (_20428_, _20427_, rst);
  nand (_20429_, _04634_, _03698_);
  or (_20430_, _04634_, \oc8051_golden_model_1.P1 [1]);
  and (_20432_, _20430_, _02802_);
  and (_20433_, _20432_, _20429_);
  or (_20434_, _19646_, _08808_);
  and (_20435_, _20430_, _02579_);
  and (_20436_, _20435_, _20434_);
  nor (_20437_, _04634_, _20426_);
  and (_20438_, _04634_, _04000_);
  or (_20439_, _20438_, _20437_);
  or (_20440_, _20439_, _03336_);
  and (_20441_, _11606_, _04634_);
  not (_20443_, _20441_);
  and (_20444_, _20443_, _20430_);
  or (_20445_, _20444_, _03810_);
  nand (_20446_, _04634_, _02551_);
  and (_20447_, _20446_, _20430_);
  and (_20448_, _20447_, _03813_);
  nor (_20449_, _03813_, _20426_);
  or (_20450_, _20449_, _02974_);
  or (_20451_, _20450_, _20448_);
  and (_20452_, _20451_, _02881_);
  and (_20454_, _20452_, _20445_);
  nor (_20455_, _05344_, _20426_);
  and (_20456_, _11592_, _05344_);
  or (_20457_, _20456_, _20455_);
  and (_20458_, _20457_, _02880_);
  or (_20459_, _20458_, _03069_);
  or (_20460_, _20459_, _20454_);
  and (_20461_, _20460_, _20440_);
  or (_20462_, _20461_, _03075_);
  or (_20463_, _20447_, _03084_);
  and (_20465_, _20463_, _02877_);
  and (_20466_, _20465_, _20462_);
  and (_20467_, _11595_, _05344_);
  or (_20468_, _20467_, _20455_);
  and (_20469_, _20468_, _02876_);
  or (_20470_, _20469_, _02869_);
  or (_20471_, _20470_, _20466_);
  and (_20472_, _20456_, _11591_);
  or (_20473_, _20455_, _02870_);
  or (_20474_, _20473_, _20472_);
  and (_20476_, _20474_, _20471_);
  and (_20477_, _20476_, _02864_);
  and (_20478_, _19620_, _05344_);
  or (_20479_, _20455_, _20478_);
  and (_20480_, _20479_, _02863_);
  or (_20481_, _20480_, _06770_);
  or (_20482_, _20481_, _20477_);
  or (_20483_, _20439_, _05535_);
  and (_20484_, _20483_, _20482_);
  or (_20485_, _20484_, _02853_);
  and (_20487_, _04634_, _06151_);
  or (_20488_, _20437_, _05540_);
  or (_20489_, _20488_, _20487_);
  and (_20490_, _20489_, _02838_);
  and (_20491_, _20490_, _20485_);
  or (_20492_, _20491_, _20436_);
  and (_20493_, _20492_, _02803_);
  or (_20494_, _20493_, _20433_);
  and (_20495_, _20494_, _03887_);
  or (_20496_, _11710_, _08808_);
  and (_20498_, _20430_, _02980_);
  and (_20499_, _20498_, _20496_);
  or (_20500_, _20499_, _20495_);
  and (_20501_, _20500_, _03128_);
  or (_20502_, _11715_, _08808_);
  and (_20503_, _20430_, _03127_);
  and (_20504_, _20503_, _20502_);
  or (_20505_, _20504_, _20501_);
  and (_20506_, _20505_, _03883_);
  or (_20507_, _11709_, _08808_);
  and (_20509_, _20430_, _02970_);
  and (_20510_, _20509_, _20507_);
  or (_20511_, _20510_, _20506_);
  and (_20512_, _20511_, _03137_);
  or (_20513_, _20437_, _13722_);
  and (_20514_, _20447_, _03135_);
  and (_20515_, _20514_, _20513_);
  or (_20516_, _20515_, _20512_);
  and (_20517_, _20516_, _03124_);
  or (_20518_, _20429_, _13722_);
  and (_20520_, _20430_, _02965_);
  and (_20521_, _20520_, _20518_);
  or (_20522_, _20446_, _13722_);
  and (_20523_, _20430_, _03123_);
  and (_20524_, _20523_, _20522_);
  or (_20525_, _20524_, _03163_);
  or (_20526_, _20525_, _20521_);
  or (_20527_, _20526_, _20517_);
  or (_20528_, _20444_, _03906_);
  and (_20529_, _20528_, _02498_);
  and (_20531_, _20529_, _20527_);
  and (_20532_, _20468_, _02497_);
  or (_20533_, _20532_, _02888_);
  or (_20534_, _20533_, _20531_);
  or (_20535_, _20437_, _02890_);
  or (_20536_, _20535_, _20441_);
  and (_20537_, _20536_, _42668_);
  and (_20538_, _20537_, _20534_);
  or (_43471_, _20538_, _20428_);
  not (_20539_, \oc8051_golden_model_1.P1 [2]);
  nor (_20541_, _42668_, _20539_);
  or (_20542_, _20541_, rst);
  nor (_20543_, _04634_, _20539_);
  and (_20544_, _11927_, _04634_);
  or (_20545_, _20544_, _20543_);
  and (_20546_, _20545_, _03127_);
  and (_20547_, _04634_, _04435_);
  or (_20548_, _20547_, _20543_);
  or (_20549_, _20548_, _05535_);
  or (_20550_, _20548_, _03336_);
  nor (_20552_, _11801_, _08808_);
  or (_20553_, _20552_, _20543_);
  or (_20554_, _20553_, _03810_);
  and (_20555_, _04634_, \oc8051_golden_model_1.ACC [2]);
  or (_20556_, _20555_, _20543_);
  and (_20557_, _20556_, _03813_);
  nor (_20558_, _03813_, _20539_);
  or (_20559_, _20558_, _02974_);
  or (_20560_, _20559_, _20557_);
  and (_20561_, _20560_, _02881_);
  and (_20563_, _20561_, _20554_);
  nor (_20564_, _05344_, _20539_);
  and (_20565_, _11815_, _05344_);
  or (_20566_, _20565_, _20564_);
  and (_20567_, _20566_, _02880_);
  or (_20568_, _20567_, _03069_);
  or (_20569_, _20568_, _20563_);
  and (_20570_, _20569_, _20550_);
  or (_20571_, _20570_, _03075_);
  or (_20572_, _20556_, _03084_);
  and (_20574_, _20572_, _02877_);
  and (_20575_, _20574_, _20571_);
  and (_20576_, _11797_, _05344_);
  or (_20577_, _20576_, _20564_);
  and (_20578_, _20577_, _02876_);
  or (_20579_, _20578_, _02869_);
  or (_20580_, _20579_, _20575_);
  and (_20581_, _20565_, _11830_);
  or (_20582_, _20564_, _02870_);
  or (_20583_, _20582_, _20581_);
  and (_20585_, _20583_, _02864_);
  and (_20586_, _20585_, _20580_);
  and (_20587_, _19742_, _05344_);
  or (_20588_, _20587_, _20564_);
  and (_20589_, _20588_, _02863_);
  or (_20590_, _20589_, _06770_);
  or (_20591_, _20590_, _20586_);
  and (_20592_, _20591_, _20549_);
  or (_20593_, _20592_, _02853_);
  and (_20594_, _04634_, _06155_);
  or (_20596_, _20543_, _05540_);
  or (_20597_, _20596_, _20594_);
  and (_20598_, _20597_, _02838_);
  and (_20599_, _20598_, _20593_);
  and (_20600_, _19767_, _04634_);
  or (_20601_, _20600_, _20543_);
  and (_20602_, _20601_, _02579_);
  or (_20603_, _20602_, _02802_);
  or (_20604_, _20603_, _20599_);
  and (_20605_, _04634_, _05701_);
  or (_20607_, _20605_, _20543_);
  or (_20608_, _20607_, _02803_);
  and (_20609_, _20608_, _20604_);
  or (_20610_, _20609_, _02980_);
  and (_20611_, _11921_, _04634_);
  or (_20612_, _20543_, _03887_);
  or (_20613_, _20612_, _20611_);
  and (_20614_, _20613_, _03128_);
  and (_20615_, _20614_, _20610_);
  or (_20616_, _20615_, _20546_);
  and (_20618_, _20616_, _03883_);
  or (_20619_, _20543_, _05130_);
  and (_20620_, _20607_, _02970_);
  and (_20621_, _20620_, _20619_);
  or (_20622_, _20621_, _20618_);
  and (_20623_, _20622_, _03137_);
  and (_20624_, _20556_, _03135_);
  and (_20625_, _20624_, _20619_);
  or (_20626_, _20625_, _02965_);
  or (_20627_, _20626_, _20623_);
  nor (_20629_, _11919_, _08808_);
  or (_20630_, _20543_, _05783_);
  or (_20631_, _20630_, _20629_);
  and (_20632_, _20631_, _05788_);
  and (_20633_, _20632_, _20627_);
  nor (_20634_, _11926_, _08808_);
  or (_20635_, _20634_, _20543_);
  and (_20636_, _20635_, _03123_);
  or (_20637_, _20636_, _03163_);
  or (_20638_, _20637_, _20633_);
  or (_20640_, _20553_, _03906_);
  and (_20641_, _20640_, _02498_);
  and (_20642_, _20641_, _20638_);
  and (_20643_, _20577_, _02497_);
  or (_20644_, _20643_, _02888_);
  or (_20645_, _20644_, _20642_);
  and (_20646_, _11985_, _04634_);
  or (_20647_, _20543_, _02890_);
  or (_20648_, _20647_, _20646_);
  and (_20649_, _20648_, _42668_);
  and (_20651_, _20649_, _20645_);
  or (_43472_, _20651_, _20542_);
  nor (_20652_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_20653_, _20652_, _04182_);
  and (_20654_, _08808_, \oc8051_golden_model_1.P1 [3]);
  and (_20655_, _12133_, _04634_);
  or (_20656_, _20655_, _20654_);
  and (_20657_, _20656_, _03127_);
  and (_20658_, _04634_, _04241_);
  or (_20659_, _20658_, _20654_);
  or (_20661_, _20659_, _05535_);
  nor (_20662_, _12017_, _08808_);
  or (_20663_, _20662_, _20654_);
  or (_20664_, _20663_, _03810_);
  and (_20665_, _04634_, \oc8051_golden_model_1.ACC [3]);
  or (_20666_, _20665_, _20654_);
  and (_20667_, _20666_, _03813_);
  and (_20668_, _03814_, \oc8051_golden_model_1.P1 [3]);
  or (_20669_, _20668_, _02974_);
  or (_20670_, _20669_, _20667_);
  and (_20672_, _20670_, _02881_);
  and (_20673_, _20672_, _20664_);
  not (_20674_, _05344_);
  and (_20675_, _20674_, \oc8051_golden_model_1.P1 [3]);
  and (_20676_, _12021_, _05344_);
  or (_20677_, _20676_, _20675_);
  and (_20678_, _20677_, _02880_);
  or (_20679_, _20678_, _03069_);
  or (_20680_, _20679_, _20673_);
  or (_20681_, _20659_, _03336_);
  and (_20683_, _20681_, _20680_);
  or (_20684_, _20683_, _03075_);
  or (_20685_, _20666_, _03084_);
  and (_20686_, _20685_, _02877_);
  and (_20687_, _20686_, _20684_);
  and (_20688_, _12005_, _05344_);
  or (_20689_, _20688_, _20675_);
  and (_20690_, _20689_, _02876_);
  or (_20691_, _20690_, _02869_);
  or (_20692_, _20691_, _20687_);
  or (_20694_, _20675_, _12036_);
  and (_20695_, _20694_, _20677_);
  or (_20696_, _20695_, _02870_);
  and (_20697_, _20696_, _02864_);
  and (_20698_, _20697_, _20692_);
  and (_20699_, _19864_, _05344_);
  or (_20700_, _20699_, _20675_);
  and (_20701_, _20700_, _02863_);
  or (_20702_, _20701_, _06770_);
  or (_20703_, _20702_, _20698_);
  and (_20705_, _20703_, _20661_);
  or (_20706_, _20705_, _02853_);
  and (_20707_, _04634_, _06154_);
  or (_20708_, _20654_, _05540_);
  or (_20709_, _20708_, _20707_);
  and (_20710_, _20709_, _02838_);
  and (_20711_, _20710_, _20706_);
  and (_20712_, _19888_, _04634_);
  or (_20713_, _20712_, _20654_);
  and (_20714_, _20713_, _02579_);
  or (_20716_, _20714_, _02802_);
  or (_20717_, _20716_, _20711_);
  and (_20718_, _04634_, _05658_);
  or (_20719_, _20718_, _20654_);
  or (_20720_, _20719_, _02803_);
  and (_20721_, _20720_, _20717_);
  or (_20722_, _20721_, _02980_);
  and (_20723_, _12127_, _04634_);
  or (_20724_, _20654_, _03887_);
  or (_20725_, _20724_, _20723_);
  and (_20727_, _20725_, _03128_);
  and (_20728_, _20727_, _20722_);
  or (_20729_, _20728_, _20657_);
  and (_20730_, _20729_, _03883_);
  or (_20731_, _20654_, _05079_);
  and (_20732_, _20719_, _02970_);
  and (_20733_, _20732_, _20731_);
  or (_20734_, _20733_, _20730_);
  and (_20735_, _20734_, _03137_);
  and (_20736_, _20666_, _03135_);
  and (_20738_, _20736_, _20731_);
  or (_20739_, _20738_, _02965_);
  or (_20740_, _20739_, _20735_);
  nor (_20741_, _12125_, _08808_);
  or (_20742_, _20654_, _05783_);
  or (_20743_, _20742_, _20741_);
  and (_20744_, _20743_, _05788_);
  and (_20745_, _20744_, _20740_);
  nor (_20746_, _12132_, _08808_);
  or (_20747_, _20746_, _20654_);
  and (_20749_, _20747_, _03123_);
  or (_20750_, _20749_, _03163_);
  or (_20751_, _20750_, _20745_);
  or (_20752_, _20663_, _03906_);
  and (_20753_, _20752_, _02498_);
  and (_20754_, _20753_, _20751_);
  and (_20755_, _20689_, _02497_);
  or (_20756_, _20755_, _02888_);
  or (_20757_, _20756_, _20754_);
  and (_20758_, _12183_, _04634_);
  or (_20760_, _20654_, _02890_);
  or (_20761_, _20760_, _20758_);
  and (_20762_, _20761_, _42668_);
  and (_20763_, _20762_, _20757_);
  or (_43473_, _20763_, _20653_);
  nor (_20764_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_20765_, _20764_, _04182_);
  and (_20766_, _08808_, \oc8051_golden_model_1.P1 [4]);
  and (_20767_, _12207_, _04634_);
  or (_20768_, _20767_, _20766_);
  and (_20770_, _20768_, _03127_);
  and (_20771_, _04634_, _04982_);
  or (_20772_, _20771_, _20766_);
  or (_20773_, _20772_, _05535_);
  and (_20774_, _20674_, \oc8051_golden_model_1.P1 [4]);
  and (_20775_, _12213_, _05344_);
  or (_20776_, _20775_, _20774_);
  and (_20777_, _20776_, _02876_);
  nor (_20778_, _12217_, _08808_);
  or (_20779_, _20778_, _20766_);
  or (_20781_, _20779_, _03810_);
  and (_20782_, _04634_, \oc8051_golden_model_1.ACC [4]);
  or (_20783_, _20782_, _20766_);
  and (_20784_, _20783_, _03813_);
  and (_20785_, _03814_, \oc8051_golden_model_1.P1 [4]);
  or (_20786_, _20785_, _02974_);
  or (_20787_, _20786_, _20784_);
  and (_20788_, _20787_, _02881_);
  and (_20789_, _20788_, _20781_);
  and (_20790_, _12231_, _05344_);
  or (_20792_, _20790_, _20774_);
  and (_20793_, _20792_, _02880_);
  or (_20794_, _20793_, _03069_);
  or (_20795_, _20794_, _20789_);
  or (_20796_, _20772_, _03336_);
  and (_20797_, _20796_, _20795_);
  or (_20798_, _20797_, _03075_);
  or (_20799_, _20783_, _03084_);
  and (_20800_, _20799_, _02877_);
  and (_20801_, _20800_, _20798_);
  or (_20803_, _20801_, _20777_);
  and (_20804_, _20803_, _02870_);
  and (_20805_, _12247_, _05344_);
  or (_20806_, _20805_, _20774_);
  and (_20807_, _20806_, _02869_);
  or (_20808_, _20807_, _20804_);
  and (_20809_, _20808_, _02864_);
  and (_20810_, _19985_, _05344_);
  or (_20811_, _20810_, _20774_);
  and (_20812_, _20811_, _02863_);
  or (_20814_, _20812_, _06770_);
  or (_20815_, _20814_, _20809_);
  and (_20816_, _20815_, _20773_);
  or (_20817_, _20816_, _02853_);
  and (_20818_, _04634_, _06159_);
  or (_20819_, _20766_, _05540_);
  or (_20820_, _20819_, _20818_);
  and (_20821_, _20820_, _02838_);
  and (_20822_, _20821_, _20817_);
  and (_20823_, _20011_, _04634_);
  or (_20825_, _20823_, _20766_);
  and (_20826_, _20825_, _02579_);
  or (_20827_, _20826_, _02802_);
  or (_20828_, _20827_, _20822_);
  and (_20829_, _05666_, _04634_);
  or (_20830_, _20829_, _20766_);
  or (_20831_, _20830_, _02803_);
  and (_20832_, _20831_, _20828_);
  or (_20833_, _20832_, _02980_);
  and (_20834_, _12211_, _04634_);
  or (_20836_, _20766_, _03887_);
  or (_20837_, _20836_, _20834_);
  and (_20838_, _20837_, _03128_);
  and (_20839_, _20838_, _20833_);
  or (_20840_, _20839_, _20770_);
  and (_20841_, _20840_, _03883_);
  or (_20842_, _20766_, _05031_);
  and (_20843_, _20830_, _02970_);
  and (_20844_, _20843_, _20842_);
  or (_20845_, _20844_, _20841_);
  and (_20847_, _20845_, _03137_);
  and (_20848_, _20783_, _03135_);
  and (_20849_, _20848_, _20842_);
  or (_20850_, _20849_, _02965_);
  or (_20851_, _20850_, _20847_);
  nor (_20852_, _12209_, _08808_);
  or (_20853_, _20766_, _05783_);
  or (_20854_, _20853_, _20852_);
  and (_20855_, _20854_, _05788_);
  and (_20856_, _20855_, _20851_);
  nor (_20858_, _12206_, _08808_);
  or (_20859_, _20858_, _20766_);
  and (_20860_, _20859_, _03123_);
  or (_20861_, _20860_, _03163_);
  or (_20862_, _20861_, _20856_);
  or (_20863_, _20779_, _03906_);
  and (_20864_, _20863_, _02498_);
  and (_20865_, _20864_, _20862_);
  and (_20866_, _20776_, _02497_);
  or (_20867_, _20866_, _02888_);
  or (_20869_, _20867_, _20865_);
  and (_20870_, _12389_, _04634_);
  or (_20871_, _20766_, _02890_);
  or (_20872_, _20871_, _20870_);
  and (_20873_, _20872_, _42668_);
  and (_20874_, _20873_, _20869_);
  or (_43474_, _20874_, _20765_);
  nor (_20875_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_20876_, _20875_, _04182_);
  and (_20877_, _08808_, \oc8051_golden_model_1.P1 [5]);
  and (_20879_, _12411_, _04634_);
  or (_20880_, _20879_, _20877_);
  and (_20881_, _20880_, _03127_);
  nor (_20882_, _12407_, _08808_);
  or (_20883_, _20882_, _20877_);
  or (_20884_, _20883_, _03810_);
  and (_20885_, _04634_, \oc8051_golden_model_1.ACC [5]);
  or (_20886_, _20885_, _20877_);
  and (_20887_, _20886_, _03813_);
  and (_20888_, _03814_, \oc8051_golden_model_1.P1 [5]);
  or (_20890_, _20888_, _02974_);
  or (_20891_, _20890_, _20887_);
  and (_20892_, _20891_, _02881_);
  and (_20893_, _20892_, _20884_);
  and (_20894_, _20674_, \oc8051_golden_model_1.P1 [5]);
  and (_20895_, _12435_, _05344_);
  or (_20896_, _20895_, _20894_);
  and (_20897_, _20896_, _02880_);
  or (_20898_, _20897_, _03069_);
  or (_20899_, _20898_, _20893_);
  and (_20901_, _04634_, _04877_);
  or (_20902_, _20901_, _20877_);
  or (_20903_, _20902_, _03336_);
  and (_20904_, _20903_, _20899_);
  or (_20905_, _20904_, _03075_);
  or (_20906_, _20886_, _03084_);
  and (_20907_, _20906_, _02877_);
  and (_20908_, _20907_, _20905_);
  and (_20909_, _12417_, _05344_);
  or (_20910_, _20909_, _20894_);
  and (_20912_, _20910_, _02876_);
  or (_20913_, _20912_, _02869_);
  or (_20914_, _20913_, _20908_);
  or (_20915_, _20894_, _12450_);
  and (_20916_, _20915_, _20896_);
  or (_20917_, _20916_, _02870_);
  and (_20918_, _20917_, _02864_);
  and (_20919_, _20918_, _20914_);
  and (_20920_, _20108_, _05344_);
  or (_20921_, _20920_, _20894_);
  and (_20923_, _20921_, _02863_);
  or (_20924_, _20923_, _06770_);
  or (_20925_, _20924_, _20919_);
  or (_20926_, _20902_, _05535_);
  and (_20927_, _20926_, _20925_);
  or (_20928_, _20927_, _02853_);
  and (_20929_, _04634_, _06158_);
  or (_20930_, _20877_, _05540_);
  or (_20931_, _20930_, _20929_);
  and (_20932_, _20931_, _02838_);
  and (_20934_, _20932_, _20928_);
  and (_20935_, _20143_, _04634_);
  or (_20936_, _20935_, _20877_);
  and (_20937_, _20936_, _02579_);
  or (_20938_, _20937_, _02802_);
  or (_20939_, _20938_, _20934_);
  and (_20940_, _05614_, _04634_);
  or (_20941_, _20940_, _20877_);
  or (_20942_, _20941_, _02803_);
  and (_20943_, _20942_, _20939_);
  or (_20945_, _20943_, _02980_);
  and (_20946_, _12415_, _04634_);
  or (_20947_, _20877_, _03887_);
  or (_20948_, _20947_, _20946_);
  and (_20949_, _20948_, _03128_);
  and (_20950_, _20949_, _20945_);
  or (_20951_, _20950_, _20881_);
  and (_20952_, _20951_, _03883_);
  or (_20953_, _20877_, _04924_);
  and (_20954_, _20941_, _02970_);
  and (_20956_, _20954_, _20953_);
  or (_20957_, _20956_, _20952_);
  and (_20958_, _20957_, _03137_);
  and (_20959_, _20886_, _03135_);
  and (_20960_, _20959_, _20953_);
  or (_20961_, _20960_, _02965_);
  or (_20962_, _20961_, _20958_);
  nor (_20963_, _12413_, _08808_);
  or (_20964_, _20877_, _05783_);
  or (_20965_, _20964_, _20963_);
  and (_20967_, _20965_, _05788_);
  and (_20968_, _20967_, _20962_);
  nor (_20969_, _12410_, _08808_);
  or (_20970_, _20969_, _20877_);
  and (_20971_, _20970_, _03123_);
  or (_20972_, _20971_, _03163_);
  or (_20973_, _20972_, _20968_);
  or (_20974_, _20883_, _03906_);
  and (_20975_, _20974_, _02498_);
  and (_20976_, _20975_, _20973_);
  and (_20978_, _20910_, _02497_);
  or (_20979_, _20978_, _02888_);
  or (_20980_, _20979_, _20976_);
  and (_20981_, _12589_, _04634_);
  or (_20982_, _20877_, _02890_);
  or (_20983_, _20982_, _20981_);
  and (_20984_, _20983_, _42668_);
  and (_20985_, _20984_, _20980_);
  or (_43475_, _20985_, _20876_);
  not (_20986_, \oc8051_golden_model_1.P1 [6]);
  nor (_20988_, _42668_, _20986_);
  or (_20989_, _20988_, rst);
  nor (_20990_, _04634_, _20986_);
  and (_20991_, _12613_, _04634_);
  or (_20992_, _20991_, _20990_);
  and (_20993_, _20992_, _03127_);
  nor (_20994_, _12603_, _08808_);
  or (_20995_, _20994_, _20990_);
  or (_20996_, _20995_, _03810_);
  and (_20997_, _04634_, \oc8051_golden_model_1.ACC [6]);
  or (_20999_, _20997_, _20990_);
  and (_21000_, _20999_, _03813_);
  nor (_21001_, _03813_, _20986_);
  or (_21002_, _21001_, _02974_);
  or (_21003_, _21002_, _21000_);
  and (_21004_, _21003_, _02881_);
  and (_21005_, _21004_, _20996_);
  nor (_21006_, _05344_, _20986_);
  and (_21007_, _12618_, _05344_);
  or (_21008_, _21007_, _21006_);
  and (_21010_, _21008_, _02880_);
  or (_21011_, _21010_, _03069_);
  or (_21012_, _21011_, _21005_);
  and (_21013_, _04634_, _04770_);
  or (_21014_, _21013_, _20990_);
  or (_21015_, _21014_, _03336_);
  and (_21016_, _21015_, _21012_);
  or (_21017_, _21016_, _03075_);
  or (_21018_, _20999_, _03084_);
  and (_21019_, _21018_, _02877_);
  and (_21021_, _21019_, _21017_);
  and (_21022_, _12616_, _05344_);
  or (_21023_, _21022_, _21006_);
  and (_21024_, _21023_, _02876_);
  or (_21025_, _21024_, _02869_);
  or (_21026_, _21025_, _21021_);
  or (_21027_, _21006_, _12646_);
  and (_21028_, _21027_, _21008_);
  or (_21029_, _21028_, _02870_);
  and (_21030_, _21029_, _02864_);
  and (_21032_, _21030_, _21026_);
  and (_21033_, _20240_, _05344_);
  or (_21034_, _21033_, _21006_);
  and (_21035_, _21034_, _02863_);
  or (_21036_, _21035_, _06770_);
  or (_21037_, _21036_, _21032_);
  or (_21038_, _21014_, _05535_);
  and (_21039_, _21038_, _21037_);
  or (_21040_, _21039_, _02853_);
  and (_21041_, _04634_, _05849_);
  or (_21043_, _20990_, _05540_);
  or (_21044_, _21043_, _21041_);
  and (_21045_, _21044_, _02838_);
  and (_21046_, _21045_, _21040_);
  and (_21047_, _20267_, _04634_);
  or (_21048_, _21047_, _20990_);
  and (_21049_, _21048_, _02579_);
  or (_21050_, _21049_, _02802_);
  or (_21051_, _21050_, _21046_);
  and (_21052_, _12729_, _04634_);
  or (_21054_, _21052_, _20990_);
  or (_21055_, _21054_, _02803_);
  and (_21056_, _21055_, _21051_);
  or (_21057_, _21056_, _02980_);
  and (_21058_, _12739_, _04634_);
  or (_21059_, _20990_, _03887_);
  or (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _03128_);
  and (_21062_, _21061_, _21057_);
  or (_21063_, _21062_, _20993_);
  and (_21065_, _21063_, _03883_);
  or (_21066_, _20990_, _04819_);
  and (_21067_, _21054_, _02970_);
  and (_21068_, _21067_, _21066_);
  or (_21069_, _21068_, _21065_);
  and (_21070_, _21069_, _03137_);
  and (_21071_, _20999_, _03135_);
  and (_21072_, _21071_, _21066_);
  or (_21073_, _21072_, _02965_);
  or (_21074_, _21073_, _21070_);
  nor (_21076_, _12737_, _08808_);
  or (_21077_, _20990_, _05783_);
  or (_21078_, _21077_, _21076_);
  and (_21079_, _21078_, _05788_);
  and (_21080_, _21079_, _21074_);
  nor (_21081_, _12612_, _08808_);
  or (_21082_, _21081_, _20990_);
  and (_21083_, _21082_, _03123_);
  or (_21084_, _21083_, _03163_);
  or (_21085_, _21084_, _21080_);
  or (_21087_, _20995_, _03906_);
  and (_21088_, _21087_, _02498_);
  and (_21089_, _21088_, _21085_);
  and (_21090_, _21023_, _02497_);
  or (_21091_, _21090_, _02888_);
  or (_21092_, _21091_, _21089_);
  and (_21093_, _12794_, _04634_);
  or (_21094_, _20990_, _02890_);
  or (_21095_, _21094_, _21093_);
  and (_21096_, _21095_, _42668_);
  and (_21098_, _21096_, _21092_);
  or (_43476_, _21098_, _20989_);
  not (_21099_, \oc8051_golden_model_1.P2 [0]);
  nor (_21100_, _42668_, _21099_);
  or (_21101_, _21100_, rst);
  nor (_21102_, _04641_, _21099_);
  and (_21103_, _11522_, _04641_);
  or (_21104_, _21103_, _21102_);
  and (_21105_, _21104_, _03127_);
  and (_21106_, _04641_, _03808_);
  or (_21108_, _21106_, _21102_);
  or (_21109_, _21108_, _05535_);
  and (_21110_, _05226_, _04641_);
  or (_21111_, _21110_, _21102_);
  or (_21112_, _21111_, _03810_);
  and (_21113_, _04641_, \oc8051_golden_model_1.ACC [0]);
  or (_21114_, _21113_, _21102_);
  and (_21115_, _21114_, _03813_);
  nor (_21116_, _03813_, _21099_);
  or (_21117_, _21116_, _02974_);
  or (_21119_, _21117_, _21115_);
  and (_21120_, _21119_, _02881_);
  and (_21121_, _21120_, _21112_);
  nor (_21122_, _05347_, _21099_);
  and (_21123_, _11417_, _05347_);
  or (_21124_, _21123_, _21122_);
  and (_21125_, _21124_, _02880_);
  or (_21126_, _21125_, _21121_);
  and (_21127_, _21126_, _03336_);
  and (_21128_, _21108_, _03069_);
  or (_21130_, _21128_, _03075_);
  or (_21131_, _21130_, _21127_);
  or (_21132_, _21114_, _03084_);
  and (_21133_, _21132_, _02877_);
  and (_21134_, _21133_, _21131_);
  and (_21135_, _21102_, _02876_);
  or (_21136_, _21135_, _02869_);
  or (_21137_, _21136_, _21134_);
  or (_21138_, _21111_, _02870_);
  and (_21139_, _21138_, _02864_);
  and (_21141_, _21139_, _21137_);
  and (_21142_, _19499_, _05347_);
  or (_21143_, _21142_, _21122_);
  and (_21144_, _21143_, _02863_);
  or (_21145_, _21144_, _06770_);
  or (_21146_, _21145_, _21141_);
  and (_21147_, _21146_, _21109_);
  or (_21148_, _21147_, _02853_);
  and (_21149_, _04641_, _06152_);
  or (_21150_, _21102_, _05540_);
  or (_21152_, _21150_, _21149_);
  and (_21153_, _21152_, _02838_);
  and (_21154_, _21153_, _21148_);
  and (_21155_, _19524_, _04641_);
  or (_21156_, _21155_, _21102_);
  and (_21157_, _21156_, _02579_);
  or (_21158_, _21157_, _02802_);
  or (_21159_, _21158_, _21154_);
  and (_21160_, _04641_, _05672_);
  or (_21161_, _21160_, _21102_);
  or (_21163_, _21161_, _02803_);
  and (_21164_, _21163_, _21159_);
  or (_21165_, _21164_, _02980_);
  and (_21166_, _11399_, _04641_);
  or (_21167_, _21102_, _03887_);
  or (_21168_, _21167_, _21166_);
  and (_21169_, _21168_, _03128_);
  and (_21170_, _21169_, _21165_);
  or (_21171_, _21170_, _21105_);
  and (_21172_, _21171_, _03883_);
  nand (_21174_, _21161_, _02970_);
  nor (_21175_, _21174_, _21110_);
  or (_21176_, _21175_, _21172_);
  and (_21177_, _21176_, _03137_);
  or (_21178_, _21102_, _09409_);
  and (_21179_, _21114_, _03135_);
  and (_21180_, _21179_, _21178_);
  or (_21181_, _21180_, _02965_);
  or (_21182_, _21181_, _21177_);
  nor (_21183_, _11396_, _08911_);
  or (_21185_, _21102_, _05783_);
  or (_21186_, _21185_, _21183_);
  and (_21187_, _21186_, _05788_);
  and (_21188_, _21187_, _21182_);
  nor (_21189_, _11520_, _08911_);
  or (_21190_, _21189_, _21102_);
  and (_21191_, _21190_, _03123_);
  or (_21192_, _21191_, _03163_);
  or (_21193_, _21192_, _21188_);
  or (_21194_, _21111_, _03906_);
  and (_21196_, _21194_, _02498_);
  and (_21197_, _21196_, _21193_);
  and (_21198_, _21102_, _02497_);
  or (_21199_, _21198_, _02888_);
  or (_21200_, _21199_, _21197_);
  or (_21201_, _21111_, _02890_);
  and (_21202_, _21201_, _42668_);
  and (_21203_, _21202_, _21200_);
  or (_43478_, _21203_, _21101_);
  not (_21204_, \oc8051_golden_model_1.P2 [1]);
  nor (_21206_, _42668_, _21204_);
  or (_21207_, _21206_, rst);
  nand (_21208_, _04641_, _03698_);
  or (_21209_, _04641_, \oc8051_golden_model_1.P2 [1]);
  and (_21210_, _21209_, _02802_);
  and (_21211_, _21210_, _21208_);
  nor (_21212_, _04641_, _21204_);
  and (_21213_, _04641_, _04000_);
  or (_21214_, _21213_, _21212_);
  or (_21215_, _21214_, _03336_);
  and (_21217_, _11606_, _04641_);
  not (_21218_, _21217_);
  and (_21219_, _21218_, _21209_);
  or (_21220_, _21219_, _03810_);
  nand (_21221_, _04641_, _02551_);
  and (_21222_, _21221_, _21209_);
  and (_21223_, _21222_, _03813_);
  nor (_21224_, _03813_, _21204_);
  or (_21225_, _21224_, _02974_);
  or (_21226_, _21225_, _21223_);
  and (_21228_, _21226_, _02881_);
  and (_21229_, _21228_, _21220_);
  nor (_21230_, _05347_, _21204_);
  and (_21231_, _11592_, _05347_);
  or (_21232_, _21231_, _21230_);
  and (_21233_, _21232_, _02880_);
  or (_21234_, _21233_, _03069_);
  or (_21235_, _21234_, _21229_);
  and (_21236_, _21235_, _21215_);
  or (_21237_, _21236_, _03075_);
  or (_21239_, _21222_, _03084_);
  and (_21240_, _21239_, _02877_);
  and (_21241_, _21240_, _21237_);
  and (_21242_, _11595_, _05347_);
  or (_21243_, _21242_, _21230_);
  and (_21244_, _21243_, _02876_);
  or (_21245_, _21244_, _02869_);
  or (_21246_, _21245_, _21241_);
  and (_21247_, _21231_, _11591_);
  or (_21248_, _21230_, _02870_);
  or (_21250_, _21248_, _21247_);
  and (_21251_, _21250_, _21246_);
  and (_21252_, _21251_, _02864_);
  and (_21253_, _19620_, _05347_);
  or (_21254_, _21230_, _21253_);
  and (_21255_, _21254_, _02863_);
  or (_21256_, _21255_, _06770_);
  or (_21257_, _21256_, _21252_);
  or (_21258_, _21214_, _05535_);
  and (_21259_, _21258_, _21257_);
  or (_21261_, _21259_, _02853_);
  and (_21262_, _04641_, _06151_);
  or (_21263_, _21212_, _05540_);
  or (_21264_, _21263_, _21262_);
  and (_21265_, _21264_, _02838_);
  and (_21266_, _21265_, _21261_);
  and (_21267_, _19646_, _04641_);
  or (_21268_, _21267_, _21212_);
  and (_21269_, _21268_, _02579_);
  or (_21270_, _21269_, _21266_);
  and (_21272_, _21270_, _02803_);
  or (_21273_, _21272_, _21211_);
  and (_21274_, _21273_, _03887_);
  or (_21275_, _11710_, _08911_);
  and (_21276_, _21209_, _02980_);
  and (_21277_, _21276_, _21275_);
  or (_21278_, _21277_, _21274_);
  and (_21279_, _21278_, _03128_);
  or (_21280_, _11715_, _08911_);
  and (_21281_, _21209_, _03127_);
  and (_21283_, _21281_, _21280_);
  or (_21284_, _21283_, _21279_);
  and (_21285_, _21284_, _03883_);
  or (_21286_, _11709_, _08911_);
  and (_21287_, _21209_, _02970_);
  and (_21288_, _21287_, _21286_);
  or (_21289_, _21288_, _21285_);
  and (_21290_, _21289_, _03137_);
  or (_21291_, _21212_, _13722_);
  and (_21292_, _21222_, _03135_);
  and (_21294_, _21292_, _21291_);
  or (_21295_, _21294_, _21290_);
  and (_21296_, _21295_, _03124_);
  or (_21297_, _21208_, _13722_);
  and (_21298_, _21209_, _02965_);
  and (_21299_, _21298_, _21297_);
  or (_21300_, _21221_, _13722_);
  and (_21301_, _21209_, _03123_);
  and (_21302_, _21301_, _21300_);
  or (_21303_, _21302_, _03163_);
  or (_21305_, _21303_, _21299_);
  or (_21306_, _21305_, _21296_);
  or (_21307_, _21219_, _03906_);
  and (_21308_, _21307_, _02498_);
  and (_21309_, _21308_, _21306_);
  and (_21310_, _21243_, _02497_);
  or (_21311_, _21310_, _02888_);
  or (_21312_, _21311_, _21309_);
  or (_21313_, _21212_, _02890_);
  or (_21314_, _21313_, _21217_);
  and (_21316_, _21314_, _42668_);
  and (_21317_, _21316_, _21312_);
  or (_43479_, _21317_, _21207_);
  not (_21318_, \oc8051_golden_model_1.P2 [2]);
  nor (_21319_, _42668_, _21318_);
  or (_21320_, _21319_, rst);
  nor (_21321_, _04641_, _21318_);
  and (_21322_, _11927_, _04641_);
  or (_21323_, _21322_, _21321_);
  and (_21324_, _21323_, _03127_);
  and (_21326_, _04641_, _04435_);
  or (_21327_, _21326_, _21321_);
  or (_21328_, _21327_, _05535_);
  and (_21329_, _21327_, _03069_);
  nor (_21330_, _05347_, _21318_);
  and (_21331_, _11815_, _05347_);
  or (_21332_, _21331_, _21330_);
  or (_21333_, _21332_, _02881_);
  nor (_21334_, _11801_, _08911_);
  or (_21335_, _21334_, _21321_);
  and (_21337_, _21335_, _02974_);
  nor (_21338_, _03813_, _21318_);
  and (_21339_, _04641_, \oc8051_golden_model_1.ACC [2]);
  or (_21340_, _21339_, _21321_);
  and (_21341_, _21340_, _03813_);
  or (_21342_, _21341_, _21338_);
  and (_21343_, _21342_, _03810_);
  or (_21344_, _21343_, _02880_);
  or (_21345_, _21344_, _21337_);
  and (_21346_, _21345_, _21333_);
  and (_21348_, _21346_, _03336_);
  or (_21349_, _21348_, _21329_);
  or (_21350_, _21349_, _03075_);
  or (_21351_, _21340_, _03084_);
  and (_21352_, _21351_, _02877_);
  and (_21353_, _21352_, _21350_);
  and (_21354_, _11797_, _05347_);
  or (_21355_, _21354_, _21330_);
  and (_21356_, _21355_, _02876_);
  or (_21357_, _21356_, _02869_);
  or (_21359_, _21357_, _21353_);
  or (_21360_, _21330_, _11830_);
  and (_21361_, _21360_, _21332_);
  or (_21362_, _21361_, _02870_);
  and (_21363_, _21362_, _02864_);
  and (_21364_, _21363_, _21359_);
  and (_21365_, _19742_, _05347_);
  or (_21366_, _21365_, _21330_);
  and (_21367_, _21366_, _02863_);
  or (_21368_, _21367_, _06770_);
  or (_21370_, _21368_, _21364_);
  and (_21371_, _21370_, _21328_);
  or (_21372_, _21371_, _02853_);
  and (_21373_, _04641_, _06155_);
  or (_21374_, _21321_, _05540_);
  or (_21375_, _21374_, _21373_);
  and (_21376_, _21375_, _02838_);
  and (_21377_, _21376_, _21372_);
  and (_21378_, _19767_, _04641_);
  or (_21379_, _21378_, _21321_);
  and (_21381_, _21379_, _02579_);
  or (_21382_, _21381_, _02802_);
  or (_21383_, _21382_, _21377_);
  and (_21384_, _04641_, _05701_);
  or (_21385_, _21384_, _21321_);
  or (_21386_, _21385_, _02803_);
  and (_21387_, _21386_, _21383_);
  or (_21388_, _21387_, _02980_);
  and (_21389_, _11921_, _04641_);
  or (_21390_, _21321_, _03887_);
  or (_21392_, _21390_, _21389_);
  and (_21393_, _21392_, _03128_);
  and (_21394_, _21393_, _21388_);
  or (_21395_, _21394_, _21324_);
  and (_21396_, _21395_, _03883_);
  or (_21397_, _21321_, _05130_);
  and (_21398_, _21385_, _02970_);
  and (_21399_, _21398_, _21397_);
  or (_21400_, _21399_, _21396_);
  and (_21401_, _21400_, _03137_);
  and (_21403_, _21340_, _03135_);
  and (_21404_, _21403_, _21397_);
  or (_21405_, _21404_, _02965_);
  or (_21406_, _21405_, _21401_);
  nor (_21407_, _11919_, _08911_);
  or (_21408_, _21321_, _05783_);
  or (_21409_, _21408_, _21407_);
  and (_21410_, _21409_, _05788_);
  and (_21411_, _21410_, _21406_);
  nor (_21412_, _11926_, _08911_);
  or (_21414_, _21412_, _21321_);
  and (_21415_, _21414_, _03123_);
  or (_21416_, _21415_, _03163_);
  or (_21417_, _21416_, _21411_);
  or (_21418_, _21335_, _03906_);
  and (_21419_, _21418_, _02498_);
  and (_21420_, _21419_, _21417_);
  and (_21421_, _21355_, _02497_);
  or (_21422_, _21421_, _02888_);
  or (_21423_, _21422_, _21420_);
  and (_21425_, _11985_, _04641_);
  or (_21426_, _21321_, _02890_);
  or (_21427_, _21426_, _21425_);
  and (_21428_, _21427_, _42668_);
  and (_21429_, _21428_, _21423_);
  or (_43480_, _21429_, _21320_);
  nor (_21430_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_21431_, _21430_, _04182_);
  and (_21432_, _08911_, \oc8051_golden_model_1.P2 [3]);
  and (_21433_, _12133_, _04641_);
  or (_21435_, _21433_, _21432_);
  and (_21436_, _21435_, _03127_);
  and (_21437_, _04641_, _04241_);
  or (_21438_, _21437_, _21432_);
  or (_21439_, _21438_, _05535_);
  nor (_21440_, _12017_, _08911_);
  or (_21441_, _21440_, _21432_);
  or (_21442_, _21441_, _03810_);
  and (_21443_, _04641_, \oc8051_golden_model_1.ACC [3]);
  or (_21444_, _21443_, _21432_);
  and (_21446_, _21444_, _03813_);
  and (_21447_, _03814_, \oc8051_golden_model_1.P2 [3]);
  or (_21448_, _21447_, _02974_);
  or (_21449_, _21448_, _21446_);
  and (_21450_, _21449_, _02881_);
  and (_21451_, _21450_, _21442_);
  not (_21452_, _05347_);
  and (_21453_, _21452_, \oc8051_golden_model_1.P2 [3]);
  and (_21454_, _12021_, _05347_);
  or (_21455_, _21454_, _21453_);
  and (_21457_, _21455_, _02880_);
  or (_21458_, _21457_, _03069_);
  or (_21459_, _21458_, _21451_);
  or (_21460_, _21438_, _03336_);
  and (_21461_, _21460_, _21459_);
  or (_21462_, _21461_, _03075_);
  or (_21463_, _21444_, _03084_);
  and (_21464_, _21463_, _02877_);
  and (_21465_, _21464_, _21462_);
  and (_21466_, _12005_, _05347_);
  or (_21468_, _21466_, _21453_);
  and (_21469_, _21468_, _02876_);
  or (_21470_, _21469_, _02869_);
  or (_21471_, _21470_, _21465_);
  or (_21472_, _21453_, _12036_);
  and (_21473_, _21472_, _21455_);
  or (_21474_, _21473_, _02870_);
  and (_21475_, _21474_, _02864_);
  and (_21476_, _21475_, _21471_);
  and (_21477_, _19864_, _05347_);
  or (_21479_, _21477_, _21453_);
  and (_21480_, _21479_, _02863_);
  or (_21481_, _21480_, _06770_);
  or (_21482_, _21481_, _21476_);
  and (_21483_, _21482_, _21439_);
  or (_21484_, _21483_, _02853_);
  and (_21485_, _04641_, _06154_);
  or (_21486_, _21432_, _05540_);
  or (_21487_, _21486_, _21485_);
  and (_21488_, _21487_, _02838_);
  and (_21490_, _21488_, _21484_);
  and (_21491_, _19888_, _04641_);
  or (_21492_, _21491_, _21432_);
  and (_21493_, _21492_, _02579_);
  or (_21494_, _21493_, _02802_);
  or (_21495_, _21494_, _21490_);
  and (_21496_, _04641_, _05658_);
  or (_21497_, _21496_, _21432_);
  or (_21498_, _21497_, _02803_);
  and (_21499_, _21498_, _21495_);
  or (_21501_, _21499_, _02980_);
  and (_21502_, _12127_, _04641_);
  or (_21503_, _21432_, _03887_);
  or (_21504_, _21503_, _21502_);
  and (_21505_, _21504_, _03128_);
  and (_21506_, _21505_, _21501_);
  or (_21507_, _21506_, _21436_);
  and (_21508_, _21507_, _03883_);
  or (_21509_, _21432_, _05079_);
  and (_21510_, _21497_, _02970_);
  and (_21512_, _21510_, _21509_);
  or (_21513_, _21512_, _21508_);
  and (_21514_, _21513_, _03137_);
  and (_21515_, _21444_, _03135_);
  and (_21516_, _21515_, _21509_);
  or (_21517_, _21516_, _02965_);
  or (_21518_, _21517_, _21514_);
  nor (_21519_, _12125_, _08911_);
  or (_21520_, _21432_, _05783_);
  or (_21521_, _21520_, _21519_);
  and (_21523_, _21521_, _05788_);
  and (_21524_, _21523_, _21518_);
  nor (_21525_, _12132_, _08911_);
  or (_21526_, _21525_, _21432_);
  and (_21527_, _21526_, _03123_);
  or (_21528_, _21527_, _03163_);
  or (_21529_, _21528_, _21524_);
  or (_21530_, _21441_, _03906_);
  and (_21531_, _21530_, _02498_);
  and (_21532_, _21531_, _21529_);
  and (_21534_, _21468_, _02497_);
  or (_21535_, _21534_, _02888_);
  or (_21536_, _21535_, _21532_);
  and (_21537_, _12183_, _04641_);
  or (_21538_, _21432_, _02890_);
  or (_21539_, _21538_, _21537_);
  and (_21540_, _21539_, _42668_);
  and (_21541_, _21540_, _21536_);
  or (_43481_, _21541_, _21431_);
  nor (_21542_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_21544_, _21542_, _04182_);
  and (_21545_, _08911_, \oc8051_golden_model_1.P2 [4]);
  and (_21546_, _12207_, _04641_);
  or (_21547_, _21546_, _21545_);
  and (_21548_, _21547_, _03127_);
  and (_21549_, _04641_, _04982_);
  or (_21550_, _21549_, _21545_);
  or (_21551_, _21550_, _05535_);
  and (_21552_, _21452_, \oc8051_golden_model_1.P2 [4]);
  and (_21553_, _12213_, _05347_);
  or (_21555_, _21553_, _21552_);
  and (_21556_, _21555_, _02876_);
  nor (_21557_, _12217_, _08911_);
  or (_21558_, _21557_, _21545_);
  or (_21559_, _21558_, _03810_);
  and (_21560_, _04641_, \oc8051_golden_model_1.ACC [4]);
  or (_21561_, _21560_, _21545_);
  and (_21562_, _21561_, _03813_);
  and (_21563_, _03814_, \oc8051_golden_model_1.P2 [4]);
  or (_21564_, _21563_, _02974_);
  or (_21566_, _21564_, _21562_);
  and (_21567_, _21566_, _02881_);
  and (_21568_, _21567_, _21559_);
  and (_21569_, _12231_, _05347_);
  or (_21570_, _21569_, _21552_);
  and (_21571_, _21570_, _02880_);
  or (_21572_, _21571_, _03069_);
  or (_21573_, _21572_, _21568_);
  or (_21574_, _21550_, _03336_);
  and (_21575_, _21574_, _21573_);
  or (_21577_, _21575_, _03075_);
  or (_21578_, _21561_, _03084_);
  and (_21579_, _21578_, _02877_);
  and (_21580_, _21579_, _21577_);
  or (_21581_, _21580_, _21556_);
  and (_21582_, _21581_, _02870_);
  or (_21583_, _21552_, _12246_);
  and (_21584_, _21583_, _02869_);
  and (_21585_, _21584_, _21570_);
  or (_21586_, _21585_, _21582_);
  and (_21588_, _21586_, _02864_);
  and (_21589_, _19985_, _05347_);
  or (_21590_, _21589_, _21552_);
  and (_21591_, _21590_, _02863_);
  or (_21592_, _21591_, _06770_);
  or (_21593_, _21592_, _21588_);
  and (_21594_, _21593_, _21551_);
  or (_21595_, _21594_, _02853_);
  and (_21596_, _04641_, _06159_);
  or (_21597_, _21545_, _05540_);
  or (_21599_, _21597_, _21596_);
  and (_21600_, _21599_, _02838_);
  and (_21601_, _21600_, _21595_);
  and (_21602_, _20011_, _04641_);
  or (_21603_, _21602_, _21545_);
  and (_21604_, _21603_, _02579_);
  or (_21605_, _21604_, _02802_);
  or (_21606_, _21605_, _21601_);
  and (_21607_, _05666_, _04641_);
  or (_21608_, _21607_, _21545_);
  or (_21610_, _21608_, _02803_);
  and (_21611_, _21610_, _21606_);
  or (_21612_, _21611_, _02980_);
  and (_21613_, _12211_, _04641_);
  or (_21614_, _21545_, _03887_);
  or (_21615_, _21614_, _21613_);
  and (_21616_, _21615_, _03128_);
  and (_21617_, _21616_, _21612_);
  or (_21618_, _21617_, _21548_);
  and (_21619_, _21618_, _03883_);
  or (_21622_, _21545_, _05031_);
  and (_21623_, _21608_, _02970_);
  and (_21624_, _21623_, _21622_);
  or (_21625_, _21624_, _21619_);
  and (_21626_, _21625_, _03137_);
  and (_21627_, _21561_, _03135_);
  and (_21628_, _21627_, _21622_);
  or (_21629_, _21628_, _02965_);
  or (_21630_, _21629_, _21626_);
  nor (_21631_, _12209_, _08911_);
  or (_21634_, _21545_, _05783_);
  or (_21635_, _21634_, _21631_);
  and (_21636_, _21635_, _05788_);
  and (_21637_, _21636_, _21630_);
  nor (_21638_, _12206_, _08911_);
  or (_21639_, _21638_, _21545_);
  and (_21640_, _21639_, _03123_);
  or (_21641_, _21640_, _03163_);
  or (_21642_, _21641_, _21637_);
  or (_21643_, _21558_, _03906_);
  and (_21646_, _21643_, _02498_);
  and (_21647_, _21646_, _21642_);
  and (_21648_, _21555_, _02497_);
  or (_21649_, _21648_, _02888_);
  or (_21650_, _21649_, _21647_);
  and (_21651_, _12389_, _04641_);
  or (_21652_, _21545_, _02890_);
  or (_21653_, _21652_, _21651_);
  and (_21654_, _21653_, _42668_);
  and (_21655_, _21654_, _21650_);
  or (_43483_, _21655_, _21544_);
  nor (_21658_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_21659_, _21658_, _04182_);
  and (_21660_, _08911_, \oc8051_golden_model_1.P2 [5]);
  and (_21661_, _12411_, _04641_);
  or (_21662_, _21661_, _21660_);
  and (_21663_, _21662_, _03127_);
  nor (_21664_, _12407_, _08911_);
  or (_21665_, _21664_, _21660_);
  or (_21666_, _21665_, _03810_);
  and (_21669_, _04641_, \oc8051_golden_model_1.ACC [5]);
  or (_21670_, _21669_, _21660_);
  and (_21671_, _21670_, _03813_);
  and (_21672_, _03814_, \oc8051_golden_model_1.P2 [5]);
  or (_21673_, _21672_, _02974_);
  or (_21674_, _21673_, _21671_);
  and (_21675_, _21674_, _02881_);
  and (_21676_, _21675_, _21666_);
  and (_21677_, _21452_, \oc8051_golden_model_1.P2 [5]);
  and (_21678_, _12435_, _05347_);
  or (_21681_, _21678_, _21677_);
  and (_21682_, _21681_, _02880_);
  or (_21683_, _21682_, _03069_);
  or (_21684_, _21683_, _21676_);
  and (_21685_, _04641_, _04877_);
  or (_21686_, _21685_, _21660_);
  or (_21687_, _21686_, _03336_);
  and (_21688_, _21687_, _21684_);
  or (_21689_, _21688_, _03075_);
  or (_21690_, _21670_, _03084_);
  and (_21692_, _21690_, _02877_);
  and (_21693_, _21692_, _21689_);
  and (_21694_, _12417_, _05347_);
  or (_21695_, _21694_, _21677_);
  and (_21696_, _21695_, _02876_);
  or (_21697_, _21696_, _02869_);
  or (_21698_, _21697_, _21693_);
  or (_21699_, _21677_, _12450_);
  and (_21700_, _21699_, _21681_);
  or (_21701_, _21700_, _02870_);
  and (_21703_, _21701_, _02864_);
  and (_21704_, _21703_, _21698_);
  and (_21705_, _20108_, _05347_);
  or (_21706_, _21705_, _21677_);
  and (_21707_, _21706_, _02863_);
  or (_21708_, _21707_, _06770_);
  or (_21709_, _21708_, _21704_);
  or (_21710_, _21686_, _05535_);
  and (_21711_, _21710_, _21709_);
  or (_21712_, _21711_, _02853_);
  and (_21714_, _04641_, _06158_);
  or (_21715_, _21660_, _05540_);
  or (_21716_, _21715_, _21714_);
  and (_21717_, _21716_, _02838_);
  and (_21718_, _21717_, _21712_);
  and (_21719_, _20143_, _04641_);
  or (_21720_, _21719_, _21660_);
  and (_21721_, _21720_, _02579_);
  or (_21722_, _21721_, _02802_);
  or (_21723_, _21722_, _21718_);
  and (_21725_, _05614_, _04641_);
  or (_21726_, _21725_, _21660_);
  or (_21727_, _21726_, _02803_);
  and (_21728_, _21727_, _21723_);
  or (_21729_, _21728_, _02980_);
  and (_21730_, _12415_, _04641_);
  or (_21731_, _21660_, _03887_);
  or (_21732_, _21731_, _21730_);
  and (_21733_, _21732_, _03128_);
  and (_21734_, _21733_, _21729_);
  or (_21736_, _21734_, _21663_);
  and (_21737_, _21736_, _03883_);
  or (_21738_, _21660_, _04924_);
  and (_21739_, _21726_, _02970_);
  and (_21740_, _21739_, _21738_);
  or (_21741_, _21740_, _21737_);
  and (_21742_, _21741_, _03137_);
  and (_21743_, _21670_, _03135_);
  and (_21744_, _21743_, _21738_);
  or (_21745_, _21744_, _02965_);
  or (_21747_, _21745_, _21742_);
  nor (_21748_, _12413_, _08911_);
  or (_21749_, _21660_, _05783_);
  or (_21750_, _21749_, _21748_);
  and (_21751_, _21750_, _05788_);
  and (_21752_, _21751_, _21747_);
  nor (_21753_, _12410_, _08911_);
  or (_21754_, _21753_, _21660_);
  and (_21755_, _21754_, _03123_);
  or (_21756_, _21755_, _03163_);
  or (_21758_, _21756_, _21752_);
  or (_21759_, _21665_, _03906_);
  and (_21760_, _21759_, _02498_);
  and (_21761_, _21760_, _21758_);
  and (_21762_, _21695_, _02497_);
  or (_21763_, _21762_, _02888_);
  or (_21764_, _21763_, _21761_);
  and (_21765_, _12589_, _04641_);
  or (_21766_, _21660_, _02890_);
  or (_21767_, _21766_, _21765_);
  and (_21769_, _21767_, _42668_);
  and (_21770_, _21769_, _21764_);
  or (_43484_, _21770_, _21659_);
  not (_21771_, \oc8051_golden_model_1.P2 [6]);
  nor (_21772_, _42668_, _21771_);
  or (_21773_, _21772_, rst);
  nor (_21774_, _04641_, _21771_);
  and (_21775_, _12613_, _04641_);
  or (_21776_, _21775_, _21774_);
  and (_21777_, _21776_, _03127_);
  nor (_21779_, _12603_, _08911_);
  or (_21780_, _21779_, _21774_);
  or (_21781_, _21780_, _03810_);
  and (_21782_, _04641_, \oc8051_golden_model_1.ACC [6]);
  or (_21783_, _21782_, _21774_);
  and (_21784_, _21783_, _03813_);
  nor (_21785_, _03813_, _21771_);
  or (_21786_, _21785_, _02974_);
  or (_21787_, _21786_, _21784_);
  and (_21788_, _21787_, _02881_);
  and (_21790_, _21788_, _21781_);
  nor (_21791_, _05347_, _21771_);
  and (_21792_, _12618_, _05347_);
  or (_21793_, _21792_, _21791_);
  and (_21794_, _21793_, _02880_);
  or (_21795_, _21794_, _03069_);
  or (_21796_, _21795_, _21790_);
  and (_21797_, _04641_, _04770_);
  or (_21798_, _21797_, _21774_);
  or (_21799_, _21798_, _03336_);
  and (_21801_, _21799_, _21796_);
  or (_21802_, _21801_, _03075_);
  or (_21803_, _21783_, _03084_);
  and (_21804_, _21803_, _02877_);
  and (_21805_, _21804_, _21802_);
  and (_21806_, _12616_, _05347_);
  or (_21807_, _21806_, _21791_);
  and (_21808_, _21807_, _02876_);
  or (_21809_, _21808_, _02869_);
  or (_21810_, _21809_, _21805_);
  or (_21812_, _21791_, _12646_);
  and (_21813_, _21812_, _21793_);
  or (_21814_, _21813_, _02870_);
  and (_21815_, _21814_, _02864_);
  and (_21816_, _21815_, _21810_);
  and (_21817_, _20240_, _05347_);
  or (_21818_, _21817_, _21791_);
  and (_21819_, _21818_, _02863_);
  or (_21820_, _21819_, _06770_);
  or (_21821_, _21820_, _21816_);
  or (_21823_, _21798_, _05535_);
  and (_21824_, _21823_, _21821_);
  or (_21825_, _21824_, _02853_);
  and (_21826_, _04641_, _05849_);
  or (_21827_, _21774_, _05540_);
  or (_21828_, _21827_, _21826_);
  and (_21829_, _21828_, _02838_);
  and (_21830_, _21829_, _21825_);
  and (_21831_, _20267_, _04641_);
  or (_21832_, _21831_, _21774_);
  and (_21834_, _21832_, _02579_);
  or (_21835_, _21834_, _02802_);
  or (_21836_, _21835_, _21830_);
  and (_21837_, _12729_, _04641_);
  or (_21838_, _21837_, _21774_);
  or (_21839_, _21838_, _02803_);
  and (_21840_, _21839_, _21836_);
  or (_21841_, _21840_, _02980_);
  and (_21842_, _12739_, _04641_);
  or (_21843_, _21774_, _03887_);
  or (_21845_, _21843_, _21842_);
  and (_21846_, _21845_, _03128_);
  and (_21847_, _21846_, _21841_);
  or (_21848_, _21847_, _21777_);
  and (_21849_, _21848_, _03883_);
  or (_21850_, _21774_, _04819_);
  and (_21851_, _21838_, _02970_);
  and (_21852_, _21851_, _21850_);
  or (_21853_, _21852_, _21849_);
  and (_21854_, _21853_, _03137_);
  and (_21856_, _21783_, _03135_);
  and (_21857_, _21856_, _21850_);
  or (_21858_, _21857_, _02965_);
  or (_21859_, _21858_, _21854_);
  nor (_21860_, _12737_, _08911_);
  or (_21861_, _21774_, _05783_);
  or (_21862_, _21861_, _21860_);
  and (_21863_, _21862_, _05788_);
  and (_21864_, _21863_, _21859_);
  nor (_21865_, _12612_, _08911_);
  or (_21867_, _21865_, _21774_);
  and (_21868_, _21867_, _03123_);
  or (_21869_, _21868_, _03163_);
  or (_21870_, _21869_, _21864_);
  or (_21871_, _21780_, _03906_);
  and (_21872_, _21871_, _02498_);
  and (_21873_, _21872_, _21870_);
  and (_21874_, _21807_, _02497_);
  or (_21875_, _21874_, _02888_);
  or (_21876_, _21875_, _21873_);
  and (_21878_, _12794_, _04641_);
  or (_21879_, _21774_, _02890_);
  or (_21880_, _21879_, _21878_);
  and (_21881_, _21880_, _42668_);
  and (_21882_, _21881_, _21876_);
  or (_43485_, _21882_, _21773_);
  not (_21883_, \oc8051_golden_model_1.P3 [0]);
  nor (_21884_, _42668_, _21883_);
  or (_21885_, _21884_, rst);
  nor (_21886_, _04645_, _21883_);
  and (_21888_, _11522_, _04645_);
  or (_21889_, _21888_, _21886_);
  and (_21890_, _21889_, _03127_);
  and (_21891_, _04645_, _03808_);
  or (_21892_, _21891_, _21886_);
  or (_21893_, _21892_, _05535_);
  and (_21894_, _05226_, _04645_);
  or (_21895_, _21894_, _21886_);
  or (_21896_, _21895_, _03810_);
  and (_21897_, _04645_, \oc8051_golden_model_1.ACC [0]);
  or (_21899_, _21897_, _21886_);
  and (_21900_, _21899_, _03813_);
  nor (_21901_, _03813_, _21883_);
  or (_21902_, _21901_, _02974_);
  or (_21903_, _21902_, _21900_);
  and (_21904_, _21903_, _02881_);
  and (_21905_, _21904_, _21896_);
  nor (_21906_, _05349_, _21883_);
  and (_21907_, _11417_, _05349_);
  or (_21908_, _21907_, _21906_);
  and (_21910_, _21908_, _02880_);
  or (_21911_, _21910_, _21905_);
  and (_21912_, _21911_, _03336_);
  and (_21913_, _21892_, _03069_);
  or (_21914_, _21913_, _03075_);
  or (_21915_, _21914_, _21912_);
  or (_21916_, _21899_, _03084_);
  and (_21917_, _21916_, _02877_);
  and (_21918_, _21917_, _21915_);
  and (_21919_, _21886_, _02876_);
  or (_21921_, _21919_, _02869_);
  or (_21922_, _21921_, _21918_);
  or (_21923_, _21895_, _02870_);
  and (_21924_, _21923_, _02864_);
  and (_21925_, _21924_, _21922_);
  and (_21926_, _19499_, _05349_);
  or (_21927_, _21926_, _21906_);
  and (_21928_, _21927_, _02863_);
  or (_21929_, _21928_, _06770_);
  or (_21930_, _21929_, _21925_);
  and (_21932_, _21930_, _21893_);
  or (_21933_, _21932_, _02853_);
  and (_21934_, _04645_, _06152_);
  or (_21935_, _21886_, _05540_);
  or (_21936_, _21935_, _21934_);
  and (_21937_, _21936_, _02838_);
  and (_21938_, _21937_, _21933_);
  and (_21939_, _19524_, _04645_);
  or (_21940_, _21939_, _21886_);
  and (_21941_, _21940_, _02579_);
  or (_21943_, _21941_, _02802_);
  or (_21944_, _21943_, _21938_);
  and (_21945_, _04645_, _05672_);
  or (_21946_, _21945_, _21886_);
  or (_21947_, _21946_, _02803_);
  and (_21948_, _21947_, _21944_);
  or (_21949_, _21948_, _02980_);
  and (_21950_, _11399_, _04645_);
  or (_21951_, _21886_, _03887_);
  or (_21952_, _21951_, _21950_);
  and (_21954_, _21952_, _03128_);
  and (_21955_, _21954_, _21949_);
  or (_21956_, _21955_, _21890_);
  and (_21957_, _21956_, _03883_);
  nand (_21958_, _21946_, _02970_);
  nor (_21959_, _21958_, _21894_);
  or (_21960_, _21959_, _21957_);
  and (_21961_, _21960_, _03137_);
  or (_21962_, _21886_, _09409_);
  and (_21963_, _21899_, _03135_);
  and (_21965_, _21963_, _21962_);
  or (_21966_, _21965_, _02965_);
  or (_21967_, _21966_, _21961_);
  nor (_21968_, _11396_, _09020_);
  or (_21969_, _21886_, _05783_);
  or (_21970_, _21969_, _21968_);
  and (_21971_, _21970_, _05788_);
  and (_21972_, _21971_, _21967_);
  nor (_21973_, _11520_, _09020_);
  or (_21974_, _21973_, _21886_);
  and (_21976_, _21974_, _03123_);
  or (_21977_, _21976_, _03163_);
  or (_21978_, _21977_, _21972_);
  or (_21979_, _21895_, _03906_);
  and (_21980_, _21979_, _02498_);
  and (_21981_, _21980_, _21978_);
  and (_21982_, _21886_, _02497_);
  or (_21983_, _21982_, _02888_);
  or (_21984_, _21983_, _21981_);
  or (_21985_, _21895_, _02890_);
  and (_21987_, _21985_, _42668_);
  and (_21988_, _21987_, _21984_);
  or (_43487_, _21988_, _21885_);
  not (_21989_, \oc8051_golden_model_1.P3 [1]);
  nor (_21990_, _42668_, _21989_);
  or (_21991_, _21990_, rst);
  nand (_21992_, _04645_, _03698_);
  or (_21993_, _04645_, \oc8051_golden_model_1.P3 [1]);
  and (_21994_, _21993_, _02802_);
  and (_21995_, _21994_, _21992_);
  or (_21997_, _19646_, _09020_);
  and (_21998_, _21993_, _02579_);
  and (_21999_, _21998_, _21997_);
  nor (_22000_, _04645_, _21989_);
  and (_22001_, _04645_, _04000_);
  or (_22002_, _22001_, _22000_);
  or (_22003_, _22002_, _03336_);
  and (_22004_, _11606_, _04645_);
  not (_22005_, _22004_);
  and (_22006_, _22005_, _21993_);
  or (_22008_, _22006_, _03810_);
  nand (_22009_, _04645_, _02551_);
  and (_22010_, _22009_, _21993_);
  and (_22011_, _22010_, _03813_);
  nor (_22012_, _03813_, _21989_);
  or (_22013_, _22012_, _02974_);
  or (_22014_, _22013_, _22011_);
  and (_22015_, _22014_, _02881_);
  and (_22016_, _22015_, _22008_);
  nor (_22017_, _05349_, _21989_);
  and (_22019_, _11592_, _05349_);
  or (_22020_, _22019_, _22017_);
  and (_22021_, _22020_, _02880_);
  or (_22022_, _22021_, _03069_);
  or (_22023_, _22022_, _22016_);
  and (_22024_, _22023_, _22003_);
  or (_22025_, _22024_, _03075_);
  or (_22026_, _22010_, _03084_);
  and (_22027_, _22026_, _02877_);
  and (_22028_, _22027_, _22025_);
  and (_22030_, _11595_, _05349_);
  or (_22031_, _22030_, _22017_);
  and (_22032_, _22031_, _02876_);
  or (_22033_, _22032_, _02869_);
  or (_22034_, _22033_, _22028_);
  and (_22035_, _22019_, _11591_);
  or (_22036_, _22017_, _02870_);
  or (_22037_, _22036_, _22035_);
  and (_22038_, _22037_, _22034_);
  and (_22039_, _22038_, _02864_);
  and (_22041_, _19620_, _05349_);
  or (_22042_, _22017_, _22041_);
  and (_22043_, _22042_, _02863_);
  or (_22044_, _22043_, _06770_);
  or (_22045_, _22044_, _22039_);
  or (_22046_, _22002_, _05535_);
  and (_22047_, _22046_, _22045_);
  or (_22048_, _22047_, _02853_);
  and (_22049_, _04645_, _06151_);
  or (_22050_, _22000_, _05540_);
  or (_22052_, _22050_, _22049_);
  and (_22053_, _22052_, _02838_);
  and (_22054_, _22053_, _22048_);
  or (_22055_, _22054_, _21999_);
  and (_22056_, _22055_, _02803_);
  or (_22057_, _22056_, _21995_);
  and (_22058_, _22057_, _03887_);
  or (_22059_, _11710_, _09020_);
  and (_22060_, _21993_, _02980_);
  and (_22061_, _22060_, _22059_);
  or (_22063_, _22061_, _22058_);
  and (_22064_, _22063_, _03128_);
  or (_22065_, _11715_, _09020_);
  and (_22066_, _21993_, _03127_);
  and (_22067_, _22066_, _22065_);
  or (_22068_, _22067_, _22064_);
  and (_22069_, _22068_, _03883_);
  or (_22070_, _11709_, _09020_);
  and (_22071_, _21993_, _02970_);
  and (_22072_, _22071_, _22070_);
  or (_22074_, _22072_, _22069_);
  and (_22075_, _22074_, _03137_);
  or (_22076_, _22000_, _13722_);
  and (_22077_, _22010_, _03135_);
  and (_22078_, _22077_, _22076_);
  or (_22079_, _22078_, _22075_);
  and (_22080_, _22079_, _03124_);
  or (_22081_, _22009_, _13722_);
  and (_22082_, _21993_, _03123_);
  and (_22083_, _22082_, _22081_);
  or (_22085_, _22083_, _03163_);
  or (_22086_, _21992_, _13722_);
  and (_22087_, _21993_, _02965_);
  and (_22088_, _22087_, _22086_);
  or (_22089_, _22088_, _22085_);
  or (_22090_, _22089_, _22080_);
  or (_22091_, _22006_, _03906_);
  and (_22092_, _22091_, _02498_);
  and (_22093_, _22092_, _22090_);
  and (_22094_, _22031_, _02497_);
  or (_22096_, _22094_, _02888_);
  or (_22097_, _22096_, _22093_);
  or (_22098_, _22000_, _02890_);
  or (_22099_, _22098_, _22004_);
  and (_22100_, _22099_, _42668_);
  and (_22101_, _22100_, _22097_);
  or (_43488_, _22101_, _21991_);
  not (_22102_, \oc8051_golden_model_1.P3 [2]);
  nor (_22103_, _42668_, _22102_);
  or (_22104_, _22103_, rst);
  nor (_22106_, _04645_, _22102_);
  and (_22107_, _11927_, _04645_);
  or (_22108_, _22107_, _22106_);
  and (_22109_, _22108_, _03127_);
  and (_22110_, _04645_, _04435_);
  or (_22111_, _22110_, _22106_);
  or (_22112_, _22111_, _05535_);
  or (_22113_, _22111_, _03336_);
  nor (_22114_, _11801_, _09020_);
  or (_22115_, _22114_, _22106_);
  or (_22117_, _22115_, _03810_);
  and (_22118_, _04645_, \oc8051_golden_model_1.ACC [2]);
  or (_22119_, _22118_, _22106_);
  and (_22120_, _22119_, _03813_);
  nor (_22121_, _03813_, _22102_);
  or (_22122_, _22121_, _02974_);
  or (_22123_, _22122_, _22120_);
  and (_22124_, _22123_, _02881_);
  and (_22125_, _22124_, _22117_);
  nor (_22126_, _05349_, _22102_);
  and (_22128_, _11815_, _05349_);
  or (_22129_, _22128_, _22126_);
  and (_22130_, _22129_, _02880_);
  or (_22131_, _22130_, _03069_);
  or (_22132_, _22131_, _22125_);
  and (_22133_, _22132_, _22113_);
  or (_22134_, _22133_, _03075_);
  or (_22135_, _22119_, _03084_);
  and (_22136_, _22135_, _02877_);
  and (_22137_, _22136_, _22134_);
  and (_22139_, _11797_, _05349_);
  or (_22140_, _22139_, _22126_);
  and (_22141_, _22140_, _02876_);
  or (_22142_, _22141_, _02869_);
  or (_22143_, _22142_, _22137_);
  and (_22144_, _22128_, _11830_);
  or (_22145_, _22126_, _02870_);
  or (_22146_, _22145_, _22144_);
  and (_22147_, _22146_, _02864_);
  and (_22148_, _22147_, _22143_);
  and (_22150_, _19742_, _05349_);
  or (_22151_, _22150_, _22126_);
  and (_22152_, _22151_, _02863_);
  or (_22153_, _22152_, _06770_);
  or (_22154_, _22153_, _22148_);
  and (_22155_, _22154_, _22112_);
  or (_22156_, _22155_, _02853_);
  and (_22157_, _04645_, _06155_);
  or (_22158_, _22106_, _05540_);
  or (_22159_, _22158_, _22157_);
  and (_22161_, _22159_, _02838_);
  and (_22162_, _22161_, _22156_);
  and (_22163_, _19767_, _04645_);
  or (_22164_, _22163_, _22106_);
  and (_22165_, _22164_, _02579_);
  or (_22166_, _22165_, _02802_);
  or (_22167_, _22166_, _22162_);
  and (_22168_, _04645_, _05701_);
  or (_22169_, _22168_, _22106_);
  or (_22170_, _22169_, _02803_);
  and (_22172_, _22170_, _22167_);
  or (_22173_, _22172_, _02980_);
  and (_22174_, _11921_, _04645_);
  or (_22175_, _22106_, _03887_);
  or (_22176_, _22175_, _22174_);
  and (_22177_, _22176_, _03128_);
  and (_22178_, _22177_, _22173_);
  or (_22179_, _22178_, _22109_);
  and (_22180_, _22179_, _03883_);
  or (_22181_, _22106_, _05130_);
  and (_22182_, _22169_, _02970_);
  and (_22183_, _22182_, _22181_);
  or (_22184_, _22183_, _22180_);
  and (_22185_, _22184_, _03137_);
  and (_22186_, _22119_, _03135_);
  and (_22187_, _22186_, _22181_);
  or (_22188_, _22187_, _02965_);
  or (_22189_, _22188_, _22185_);
  nor (_22190_, _11919_, _09020_);
  or (_22191_, _22106_, _05783_);
  or (_22194_, _22191_, _22190_);
  and (_22195_, _22194_, _05788_);
  and (_22196_, _22195_, _22189_);
  nor (_22197_, _11926_, _09020_);
  or (_22198_, _22197_, _22106_);
  and (_22199_, _22198_, _03123_);
  or (_22200_, _22199_, _03163_);
  or (_22201_, _22200_, _22196_);
  or (_22202_, _22115_, _03906_);
  and (_22203_, _22202_, _02498_);
  and (_22205_, _22203_, _22201_);
  and (_22206_, _22140_, _02497_);
  or (_22207_, _22206_, _02888_);
  or (_22208_, _22207_, _22205_);
  and (_22209_, _11985_, _04645_);
  or (_22210_, _22106_, _02890_);
  or (_22211_, _22210_, _22209_);
  and (_22212_, _22211_, _42668_);
  and (_22213_, _22212_, _22208_);
  or (_43489_, _22213_, _22104_);
  nor (_22215_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_22216_, _22215_, _04182_);
  and (_22217_, _09020_, \oc8051_golden_model_1.P3 [3]);
  and (_22218_, _12133_, _04645_);
  or (_22219_, _22218_, _22217_);
  and (_22220_, _22219_, _03127_);
  and (_22221_, _04645_, _04241_);
  or (_22222_, _22221_, _22217_);
  or (_22223_, _22222_, _05535_);
  nor (_22224_, _12017_, _09020_);
  or (_22226_, _22224_, _22217_);
  or (_22227_, _22226_, _03810_);
  and (_22228_, _04645_, \oc8051_golden_model_1.ACC [3]);
  or (_22229_, _22228_, _22217_);
  and (_22230_, _22229_, _03813_);
  and (_22231_, _03814_, \oc8051_golden_model_1.P3 [3]);
  or (_22232_, _22231_, _02974_);
  or (_22233_, _22232_, _22230_);
  and (_22234_, _22233_, _02881_);
  and (_22235_, _22234_, _22227_);
  not (_22237_, _05349_);
  and (_22238_, _22237_, \oc8051_golden_model_1.P3 [3]);
  and (_22239_, _12021_, _05349_);
  or (_22240_, _22239_, _22238_);
  and (_22241_, _22240_, _02880_);
  or (_22242_, _22241_, _03069_);
  or (_22243_, _22242_, _22235_);
  or (_22244_, _22222_, _03336_);
  and (_22245_, _22244_, _22243_);
  or (_22246_, _22245_, _03075_);
  or (_22248_, _22229_, _03084_);
  and (_22249_, _22248_, _02877_);
  and (_22250_, _22249_, _22246_);
  and (_22251_, _12005_, _05349_);
  or (_22252_, _22251_, _22238_);
  and (_22253_, _22252_, _02876_);
  or (_22254_, _22253_, _02869_);
  or (_22255_, _22254_, _22250_);
  or (_22256_, _22238_, _12036_);
  and (_22257_, _22256_, _22240_);
  or (_22259_, _22257_, _02870_);
  and (_22260_, _22259_, _02864_);
  and (_22261_, _22260_, _22255_);
  and (_22262_, _19864_, _05349_);
  or (_22263_, _22262_, _22238_);
  and (_22264_, _22263_, _02863_);
  or (_22265_, _22264_, _06770_);
  or (_22266_, _22265_, _22261_);
  and (_22267_, _22266_, _22223_);
  or (_22268_, _22267_, _02853_);
  and (_22270_, _04645_, _06154_);
  or (_22271_, _22217_, _05540_);
  or (_22272_, _22271_, _22270_);
  and (_22273_, _22272_, _02838_);
  and (_22274_, _22273_, _22268_);
  and (_22275_, _19888_, _04645_);
  or (_22276_, _22275_, _22217_);
  and (_22277_, _22276_, _02579_);
  or (_22278_, _22277_, _02802_);
  or (_22279_, _22278_, _22274_);
  and (_22281_, _04645_, _05658_);
  or (_22282_, _22281_, _22217_);
  or (_22283_, _22282_, _02803_);
  and (_22284_, _22283_, _22279_);
  or (_22285_, _22284_, _02980_);
  and (_22286_, _12127_, _04645_);
  or (_22287_, _22217_, _03887_);
  or (_22288_, _22287_, _22286_);
  and (_22289_, _22288_, _03128_);
  and (_22290_, _22289_, _22285_);
  or (_22292_, _22290_, _22220_);
  and (_22293_, _22292_, _03883_);
  or (_22294_, _22217_, _05079_);
  and (_22295_, _22282_, _02970_);
  and (_22296_, _22295_, _22294_);
  or (_22297_, _22296_, _22293_);
  and (_22298_, _22297_, _03137_);
  and (_22299_, _22229_, _03135_);
  and (_22300_, _22299_, _22294_);
  or (_22301_, _22300_, _02965_);
  or (_22303_, _22301_, _22298_);
  nor (_22304_, _12125_, _09020_);
  or (_22305_, _22217_, _05783_);
  or (_22306_, _22305_, _22304_);
  and (_22307_, _22306_, _05788_);
  and (_22308_, _22307_, _22303_);
  nor (_22309_, _12132_, _09020_);
  or (_22310_, _22309_, _22217_);
  and (_22311_, _22310_, _03123_);
  or (_22312_, _22311_, _03163_);
  or (_22314_, _22312_, _22308_);
  or (_22315_, _22226_, _03906_);
  and (_22316_, _22315_, _02498_);
  and (_22317_, _22316_, _22314_);
  and (_22318_, _22252_, _02497_);
  or (_22319_, _22318_, _02888_);
  or (_22320_, _22319_, _22317_);
  and (_22321_, _12183_, _04645_);
  or (_22322_, _22217_, _02890_);
  or (_22323_, _22322_, _22321_);
  and (_22325_, _22323_, _42668_);
  and (_22326_, _22325_, _22320_);
  or (_43490_, _22326_, _22216_);
  nor (_22327_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_22328_, _22327_, _04182_);
  and (_22329_, _09020_, \oc8051_golden_model_1.P3 [4]);
  and (_22330_, _12207_, _04645_);
  or (_22331_, _22330_, _22329_);
  and (_22332_, _22331_, _03127_);
  and (_22333_, _04645_, _04982_);
  or (_22335_, _22333_, _22329_);
  or (_22336_, _22335_, _05535_);
  and (_22337_, _22237_, \oc8051_golden_model_1.P3 [4]);
  and (_22338_, _12213_, _05349_);
  or (_22339_, _22338_, _22337_);
  and (_22340_, _22339_, _02876_);
  nor (_22341_, _12217_, _09020_);
  or (_22342_, _22341_, _22329_);
  or (_22343_, _22342_, _03810_);
  and (_22344_, _04645_, \oc8051_golden_model_1.ACC [4]);
  or (_22346_, _22344_, _22329_);
  and (_22347_, _22346_, _03813_);
  and (_22348_, _03814_, \oc8051_golden_model_1.P3 [4]);
  or (_22349_, _22348_, _02974_);
  or (_22350_, _22349_, _22347_);
  and (_22351_, _22350_, _02881_);
  and (_22352_, _22351_, _22343_);
  and (_22353_, _12231_, _05349_);
  or (_22354_, _22353_, _22337_);
  and (_22355_, _22354_, _02880_);
  or (_22356_, _22355_, _03069_);
  or (_22357_, _22356_, _22352_);
  or (_22358_, _22335_, _03336_);
  and (_22359_, _22358_, _22357_);
  or (_22360_, _22359_, _03075_);
  or (_22361_, _22346_, _03084_);
  and (_22362_, _22361_, _02877_);
  and (_22363_, _22362_, _22360_);
  or (_22364_, _22363_, _22340_);
  and (_22365_, _22364_, _02870_);
  or (_22367_, _22337_, _12246_);
  and (_22368_, _22367_, _02869_);
  and (_22369_, _22368_, _22354_);
  or (_22370_, _22369_, _22365_);
  and (_22371_, _22370_, _02864_);
  and (_22372_, _19985_, _05349_);
  or (_22373_, _22372_, _22337_);
  and (_22374_, _22373_, _02863_);
  or (_22375_, _22374_, _06770_);
  or (_22376_, _22375_, _22371_);
  and (_22378_, _22376_, _22336_);
  or (_22379_, _22378_, _02853_);
  and (_22380_, _04645_, _06159_);
  or (_22381_, _22329_, _05540_);
  or (_22382_, _22381_, _22380_);
  and (_22383_, _22382_, _02838_);
  and (_22384_, _22383_, _22379_);
  and (_22385_, _20011_, _04645_);
  or (_22386_, _22385_, _22329_);
  and (_22387_, _22386_, _02579_);
  or (_22388_, _22387_, _02802_);
  or (_22389_, _22388_, _22384_);
  and (_22390_, _05666_, _04645_);
  or (_22391_, _22390_, _22329_);
  or (_22392_, _22391_, _02803_);
  and (_22393_, _22392_, _22389_);
  or (_22394_, _22393_, _02980_);
  and (_22395_, _12211_, _04645_);
  or (_22396_, _22329_, _03887_);
  or (_22397_, _22396_, _22395_);
  and (_22398_, _22397_, _03128_);
  and (_22399_, _22398_, _22394_);
  or (_22400_, _22399_, _22332_);
  and (_22401_, _22400_, _03883_);
  or (_22402_, _22329_, _05031_);
  and (_22403_, _22391_, _02970_);
  and (_22404_, _22403_, _22402_);
  or (_22405_, _22404_, _22401_);
  and (_22406_, _22405_, _03137_);
  and (_22407_, _22346_, _03135_);
  and (_22408_, _22407_, _22402_);
  or (_22409_, _22408_, _02965_);
  or (_22410_, _22409_, _22406_);
  nor (_22411_, _12209_, _09020_);
  or (_22412_, _22329_, _05783_);
  or (_22413_, _22412_, _22411_);
  and (_22414_, _22413_, _05788_);
  and (_22415_, _22414_, _22410_);
  nor (_22416_, _12206_, _09020_);
  or (_22417_, _22416_, _22329_);
  and (_22418_, _22417_, _03123_);
  or (_22419_, _22418_, _03163_);
  or (_22420_, _22419_, _22415_);
  or (_22421_, _22342_, _03906_);
  and (_22422_, _22421_, _02498_);
  and (_22423_, _22422_, _22420_);
  and (_22424_, _22339_, _02497_);
  or (_22425_, _22424_, _02888_);
  or (_22426_, _22425_, _22423_);
  and (_22427_, _12389_, _04645_);
  or (_22428_, _22329_, _02890_);
  or (_22429_, _22428_, _22427_);
  and (_22430_, _22429_, _42668_);
  and (_22431_, _22430_, _22426_);
  or (_43491_, _22431_, _22328_);
  nor (_22432_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_22433_, _22432_, _04182_);
  and (_22434_, _09020_, \oc8051_golden_model_1.P3 [5]);
  and (_22435_, _12411_, _04645_);
  or (_22436_, _22435_, _22434_);
  and (_22438_, _22436_, _03127_);
  nor (_22439_, _12407_, _09020_);
  or (_22440_, _22439_, _22434_);
  or (_22441_, _22440_, _03810_);
  and (_22442_, _04645_, \oc8051_golden_model_1.ACC [5]);
  or (_22443_, _22442_, _22434_);
  and (_22444_, _22443_, _03813_);
  and (_22445_, _03814_, \oc8051_golden_model_1.P3 [5]);
  or (_22446_, _22445_, _02974_);
  or (_22447_, _22446_, _22444_);
  and (_22450_, _22447_, _02881_);
  and (_22451_, _22450_, _22441_);
  and (_22452_, _22237_, \oc8051_golden_model_1.P3 [5]);
  and (_22453_, _12435_, _05349_);
  or (_22454_, _22453_, _22452_);
  and (_22455_, _22454_, _02880_);
  or (_22456_, _22455_, _03069_);
  or (_22457_, _22456_, _22451_);
  and (_22458_, _04645_, _04877_);
  or (_22459_, _22458_, _22434_);
  or (_22460_, _22459_, _03336_);
  and (_22461_, _22460_, _22457_);
  or (_22462_, _22461_, _03075_);
  or (_22463_, _22443_, _03084_);
  and (_22464_, _22463_, _02877_);
  and (_22465_, _22464_, _22462_);
  and (_22466_, _12417_, _05349_);
  or (_22467_, _22466_, _22452_);
  and (_22468_, _22467_, _02876_);
  or (_22469_, _22468_, _02869_);
  or (_22471_, _22469_, _22465_);
  or (_22472_, _22452_, _12450_);
  and (_22473_, _22472_, _22454_);
  or (_22474_, _22473_, _02870_);
  and (_22475_, _22474_, _02864_);
  and (_22476_, _22475_, _22471_);
  and (_22477_, _20108_, _05349_);
  or (_22478_, _22477_, _22452_);
  and (_22479_, _22478_, _02863_);
  or (_22480_, _22479_, _06770_);
  or (_22482_, _22480_, _22476_);
  or (_22483_, _22459_, _05535_);
  and (_22484_, _22483_, _22482_);
  or (_22485_, _22484_, _02853_);
  and (_22486_, _04645_, _06158_);
  or (_22487_, _22434_, _05540_);
  or (_22488_, _22487_, _22486_);
  and (_22489_, _22488_, _02838_);
  and (_22490_, _22489_, _22485_);
  and (_22491_, _20143_, _04645_);
  or (_22493_, _22491_, _22434_);
  and (_22494_, _22493_, _02579_);
  or (_22495_, _22494_, _02802_);
  or (_22496_, _22495_, _22490_);
  and (_22497_, _05614_, _04645_);
  or (_22498_, _22497_, _22434_);
  or (_22499_, _22498_, _02803_);
  and (_22500_, _22499_, _22496_);
  or (_22501_, _22500_, _02980_);
  and (_22502_, _12415_, _04645_);
  or (_22504_, _22434_, _03887_);
  or (_22505_, _22504_, _22502_);
  and (_22506_, _22505_, _03128_);
  and (_22507_, _22506_, _22501_);
  or (_22508_, _22507_, _22438_);
  and (_22509_, _22508_, _03883_);
  or (_22510_, _22434_, _04924_);
  and (_22511_, _22498_, _02970_);
  and (_22512_, _22511_, _22510_);
  or (_22513_, _22512_, _22509_);
  and (_22515_, _22513_, _03137_);
  and (_22516_, _22443_, _03135_);
  and (_22517_, _22516_, _22510_);
  or (_22518_, _22517_, _02965_);
  or (_22519_, _22518_, _22515_);
  nor (_22520_, _12413_, _09020_);
  or (_22521_, _22434_, _05783_);
  or (_22522_, _22521_, _22520_);
  and (_22523_, _22522_, _05788_);
  and (_22524_, _22523_, _22519_);
  nor (_22525_, _12410_, _09020_);
  or (_22526_, _22525_, _22434_);
  and (_22527_, _22526_, _03123_);
  or (_22528_, _22527_, _03163_);
  or (_22529_, _22528_, _22524_);
  or (_22530_, _22440_, _03906_);
  and (_22531_, _22530_, _02498_);
  and (_22532_, _22531_, _22529_);
  and (_22533_, _22467_, _02497_);
  or (_22534_, _22533_, _02888_);
  or (_22536_, _22534_, _22532_);
  and (_22537_, _12589_, _04645_);
  or (_22538_, _22434_, _02890_);
  or (_22539_, _22538_, _22537_);
  and (_22540_, _22539_, _42668_);
  and (_22541_, _22540_, _22536_);
  or (_43492_, _22541_, _22433_);
  not (_22542_, \oc8051_golden_model_1.P3 [6]);
  nor (_22543_, _42668_, _22542_);
  or (_22544_, _22543_, rst);
  nor (_22546_, _04645_, _22542_);
  and (_22547_, _12613_, _04645_);
  or (_22548_, _22547_, _22546_);
  and (_22549_, _22548_, _03127_);
  nor (_22550_, _12603_, _09020_);
  or (_22551_, _22550_, _22546_);
  or (_22552_, _22551_, _03810_);
  and (_22553_, _04645_, \oc8051_golden_model_1.ACC [6]);
  or (_22554_, _22553_, _22546_);
  and (_22555_, _22554_, _03813_);
  nor (_22557_, _03813_, _22542_);
  or (_22558_, _22557_, _02974_);
  or (_22559_, _22558_, _22555_);
  and (_22560_, _22559_, _02881_);
  and (_22561_, _22560_, _22552_);
  nor (_22562_, _05349_, _22542_);
  and (_22563_, _12618_, _05349_);
  or (_22564_, _22563_, _22562_);
  and (_22565_, _22564_, _02880_);
  or (_22566_, _22565_, _03069_);
  or (_22568_, _22566_, _22561_);
  and (_22569_, _04645_, _04770_);
  or (_22570_, _22569_, _22546_);
  or (_22571_, _22570_, _03336_);
  and (_22572_, _22571_, _22568_);
  or (_22573_, _22572_, _03075_);
  or (_22574_, _22554_, _03084_);
  and (_22575_, _22574_, _02877_);
  and (_22576_, _22575_, _22573_);
  and (_22577_, _12616_, _05349_);
  or (_22579_, _22577_, _22562_);
  and (_22580_, _22579_, _02876_);
  or (_22581_, _22580_, _02869_);
  or (_22582_, _22581_, _22576_);
  or (_22583_, _22562_, _12646_);
  and (_22584_, _22583_, _22564_);
  or (_22585_, _22584_, _02870_);
  and (_22586_, _22585_, _02864_);
  and (_22587_, _22586_, _22582_);
  and (_22588_, _20240_, _05349_);
  or (_22589_, _22588_, _22562_);
  and (_22590_, _22589_, _02863_);
  or (_22591_, _22590_, _06770_);
  or (_22592_, _22591_, _22587_);
  or (_22593_, _22570_, _05535_);
  and (_22594_, _22593_, _22592_);
  or (_22595_, _22594_, _02853_);
  and (_22596_, _04645_, _05849_);
  or (_22597_, _22546_, _05540_);
  or (_22598_, _22597_, _22596_);
  and (_22600_, _22598_, _02838_);
  and (_22601_, _22600_, _22595_);
  and (_22602_, _20267_, _04645_);
  or (_22603_, _22602_, _22546_);
  and (_22604_, _22603_, _02579_);
  or (_22605_, _22604_, _02802_);
  or (_22606_, _22605_, _22601_);
  and (_22607_, _12729_, _04645_);
  or (_22608_, _22607_, _22546_);
  or (_22609_, _22608_, _02803_);
  and (_22611_, _22609_, _22606_);
  or (_22612_, _22611_, _02980_);
  and (_22613_, _12739_, _04645_);
  or (_22614_, _22546_, _03887_);
  or (_22615_, _22614_, _22613_);
  and (_22616_, _22615_, _03128_);
  and (_22617_, _22616_, _22612_);
  or (_22618_, _22617_, _22549_);
  and (_22619_, _22618_, _03883_);
  or (_22620_, _22546_, _04819_);
  and (_22622_, _22608_, _02970_);
  and (_22623_, _22622_, _22620_);
  or (_22624_, _22623_, _22619_);
  and (_22625_, _22624_, _03137_);
  and (_22626_, _22554_, _03135_);
  and (_22627_, _22626_, _22620_);
  or (_22628_, _22627_, _02965_);
  or (_22629_, _22628_, _22625_);
  nor (_22630_, _12737_, _09020_);
  or (_22631_, _22546_, _05783_);
  or (_22633_, _22631_, _22630_);
  and (_22634_, _22633_, _05788_);
  and (_22635_, _22634_, _22629_);
  nor (_22636_, _12612_, _09020_);
  or (_22637_, _22636_, _22546_);
  and (_22638_, _22637_, _03123_);
  or (_22639_, _22638_, _03163_);
  or (_22640_, _22639_, _22635_);
  or (_22641_, _22551_, _03906_);
  and (_22642_, _22641_, _02498_);
  and (_22644_, _22642_, _22640_);
  and (_22645_, _22579_, _02497_);
  or (_22646_, _22645_, _02888_);
  or (_22647_, _22646_, _22644_);
  and (_22648_, _12794_, _04645_);
  or (_22649_, _22546_, _02890_);
  or (_22650_, _22649_, _22648_);
  and (_22651_, _22650_, _42668_);
  and (_22652_, _22651_, _22647_);
  or (_43493_, _22652_, _22544_);
  and (_22653_, _09979_, _02244_);
  nor (_22654_, _02937_, _02523_);
  not (_22655_, _22654_);
  and (_22656_, _22655_, _03486_);
  nor (_22657_, _09964_, _09970_);
  nor (_22658_, _22657_, _02244_);
  and (_22659_, _09941_, _09948_);
  nor (_22660_, _22659_, _02244_);
  and (_22661_, _09063_, _08112_);
  nor (_22662_, _22661_, _02244_);
  nor (_22664_, _03486_, _02535_);
  and (_22665_, _09074_, _05783_);
  nor (_22666_, _22665_, _02244_);
  not (_22667_, _09076_);
  nor (_22668_, _07799_, _02244_);
  and (_22669_, _07799_, _02244_);
  nor (_22670_, _22669_, _22668_);
  nor (_22671_, _22670_, _22667_);
  and (_22672_, _09081_, _03883_);
  nor (_22673_, _22672_, _02244_);
  not (_22675_, _09672_);
  and (_22676_, _09657_, _03887_);
  nor (_22677_, _22676_, _02244_);
  not (_22678_, _09083_);
  not (_22679_, _09611_);
  and (_22680_, _02802_, _02244_);
  nor (_22681_, _02981_, _02579_);
  and (_22682_, _22681_, _09200_);
  nor (_22683_, _22682_, _02244_);
  nor (_22684_, _03486_, _02619_);
  nor (_22686_, _09543_, _02244_);
  nor (_22687_, _03486_, _02614_);
  and (_22688_, _09392_, _02244_);
  and (_22689_, _03486_, \oc8051_golden_model_1.PC [0]);
  nor (_22690_, _22689_, _09272_);
  not (_22691_, _22690_);
  nor (_22692_, _22691_, _09392_);
  nor (_22693_, _22692_, _22688_);
  nor (_22694_, _22693_, _09396_);
  nor (_22695_, _03486_, _02621_);
  and (_22697_, _02616_, _02611_);
  or (_22698_, _22697_, _03486_);
  and (_22699_, _09427_, _09426_);
  nor (_22700_, _22699_, _02244_);
  or (_22701_, _22700_, _09425_);
  nor (_22702_, _09430_, _02244_);
  and (_22703_, _09430_, _02244_);
  nor (_22704_, _22703_, _22702_);
  and (_22705_, _22704_, _02611_);
  not (_22706_, _22705_);
  and (_22708_, _22706_, _22699_);
  or (_22709_, _22708_, _22701_);
  and (_22710_, _22709_, _05362_);
  and (_22711_, _22710_, _22698_);
  and (_22712_, _02837_, _02244_);
  nor (_22713_, _22712_, _09143_);
  or (_22714_, _22713_, _09420_);
  nand (_22715_, _09420_, _02244_);
  and (_22716_, _22715_, _22714_);
  nor (_22717_, _22716_, _05362_);
  nor (_22718_, _22717_, _22711_);
  nor (_22719_, _22718_, _02886_);
  and (_22720_, _02886_, \oc8051_golden_model_1.PC [0]);
  nor (_22721_, _22720_, _02974_);
  not (_22722_, _22721_);
  nor (_22723_, _22722_, _22719_);
  not (_22724_, _22723_);
  nor (_22725_, _22690_, _09412_);
  and (_22726_, _09412_, \oc8051_golden_model_1.PC [0]);
  or (_22727_, _22726_, _03810_);
  or (_22729_, _22727_, _22725_);
  and (_22730_, _22729_, _09405_);
  and (_22731_, _22730_, _22724_);
  nor (_22732_, _09405_, _02244_);
  nor (_22733_, _22732_, _04252_);
  not (_22734_, _22733_);
  nor (_22735_, _22734_, _22731_);
  nor (_22736_, _03486_, _02609_);
  and (_22737_, _09470_, _09463_);
  not (_22738_, _22737_);
  nor (_22740_, _22738_, _22736_);
  not (_22741_, _22740_);
  nor (_22742_, _22741_, _22735_);
  nor (_22743_, _22737_, _02244_);
  nor (_22744_, _22743_, _09474_);
  not (_22745_, _22744_);
  nor (_22746_, _22745_, _22742_);
  nor (_22747_, _22746_, _22695_);
  nor (_22748_, _22747_, _09481_);
  nor (_22749_, _22748_, _22694_);
  nor (_22751_, _22749_, _02978_);
  nand (_22752_, _09357_, \oc8051_golden_model_1.PC [0]);
  or (_22753_, _22690_, _09357_);
  and (_22754_, _22753_, _02978_);
  and (_22755_, _22754_, _22752_);
  or (_22756_, _22755_, _22751_);
  and (_22757_, _22756_, _09500_);
  and (_22758_, _09514_, _02244_);
  nor (_22759_, _22691_, _09514_);
  nor (_22760_, _22759_, _22758_);
  nor (_22762_, _22760_, _09500_);
  nor (_22763_, _22762_, _22757_);
  nor (_22764_, _22763_, _02952_);
  and (_22765_, _09528_, \oc8051_golden_model_1.PC [0]);
  nor (_22766_, _22690_, _09528_);
  or (_22767_, _22766_, _09531_);
  nor (_22768_, _22767_, _22765_);
  or (_22769_, _22768_, _22764_);
  and (_22770_, _22769_, _09490_);
  and (_22771_, _09489_, _02244_);
  or (_22773_, _22771_, _22770_);
  and (_22774_, _22773_, _02614_);
  or (_22775_, _22774_, _09544_);
  nor (_22776_, _22775_, _22687_);
  or (_22777_, _22776_, _09551_);
  nor (_22778_, _22777_, _22686_);
  and (_22779_, _09557_, _02605_);
  not (_22780_, _22779_);
  or (_22781_, _22780_, _22778_);
  nor (_22782_, _22781_, _22684_);
  nor (_22783_, _22779_, _02244_);
  nor (_22784_, _22783_, _02581_);
  not (_22785_, _22784_);
  nor (_22786_, _22785_, _22782_);
  nor (_22787_, _03486_, _04251_);
  not (_22788_, _22682_);
  nor (_22789_, _22788_, _22787_);
  not (_22790_, _22789_);
  nor (_22791_, _22790_, _22786_);
  or (_22792_, _22791_, _02518_);
  nor (_22794_, _22792_, _22683_);
  not (_22795_, _02518_);
  nor (_22796_, _03486_, _22795_);
  or (_22797_, _22796_, _09594_);
  nor (_22798_, _22797_, _22794_);
  nor (_22799_, _22713_, _09599_);
  nor (_22800_, _22799_, _22798_);
  and (_22801_, _22800_, _02803_);
  or (_22802_, _22801_, _22680_);
  and (_22803_, _22802_, _22679_);
  and (_22805_, _09611_, _02677_);
  or (_22806_, _22805_, _22803_);
  and (_22807_, _22806_, _04093_);
  nor (_22808_, _03486_, _04093_);
  or (_22809_, _22808_, _22807_);
  and (_22810_, _22809_, _22678_);
  not (_22811_, _22676_);
  and (_22812_, _08165_, \oc8051_golden_model_1.PC [0]);
  and (_22813_, _22713_, _09676_);
  or (_22814_, _22813_, _22812_);
  and (_22816_, _22814_, _09083_);
  nor (_22817_, _22816_, _22811_);
  not (_22818_, _22817_);
  nor (_22819_, _22818_, _22810_);
  nor (_22820_, _22819_, _22677_);
  and (_22821_, _22820_, _02510_);
  nor (_22822_, _03486_, _02510_);
  or (_22823_, _22822_, _22821_);
  and (_22824_, _22823_, _22675_);
  not (_22825_, _22672_);
  nor (_22827_, _22713_, _09676_);
  nor (_22828_, _08165_, \oc8051_golden_model_1.PC [0]);
  nor (_22829_, _22828_, _22675_);
  not (_22830_, _22829_);
  nor (_22831_, _22830_, _22827_);
  nor (_22832_, _22831_, _22825_);
  not (_22833_, _22832_);
  nor (_22834_, _22833_, _22824_);
  nor (_22835_, _22834_, _22673_);
  and (_22836_, _22835_, _02532_);
  nor (_22838_, _03486_, _02532_);
  or (_22839_, _22838_, _22836_);
  and (_22840_, _22839_, _22667_);
  not (_22841_, _22665_);
  or (_22842_, _22841_, _22840_);
  nor (_22843_, _22842_, _22671_);
  or (_22844_, _22843_, _09069_);
  nor (_22845_, _22844_, _22666_);
  nor (_22846_, _22845_, _22664_);
  nor (_22847_, _22846_, _09068_);
  and (_22849_, _07793_, \oc8051_golden_model_1.PC [0]);
  nor (_22850_, _07793_, \oc8051_golden_model_1.PC [0]);
  nor (_22851_, _22850_, _22849_);
  and (_22852_, _22851_, _09068_);
  and (_22853_, _09066_, _07992_);
  not (_22854_, _22853_);
  nor (_22855_, _22854_, _22852_);
  not (_22856_, _22855_);
  nor (_22857_, _22856_, _22847_);
  nor (_22858_, _22853_, _02244_);
  or (_22860_, _22858_, _03145_);
  nor (_22861_, _22860_, _22857_);
  and (_22862_, _06152_, _03145_);
  or (_22863_, _22862_, _22861_);
  and (_22864_, _22863_, _02529_);
  nor (_22865_, _03486_, _02529_);
  or (_22866_, _22865_, _22864_);
  and (_22867_, _22866_, _03561_);
  and (_22868_, _22691_, _09915_);
  nor (_22869_, _09915_, _02244_);
  or (_22870_, _22869_, _03561_);
  or (_22871_, _22870_, _22868_);
  and (_22872_, _22871_, _22661_);
  not (_22873_, _22872_);
  nor (_22874_, _22873_, _22867_);
  nor (_22875_, _22874_, _22662_);
  and (_22876_, _22875_, _02893_);
  and (_22877_, _06152_, _02892_);
  or (_22878_, _22877_, _22876_);
  and (_22879_, _22878_, _02537_);
  nor (_22881_, _03486_, _02537_);
  nor (_22882_, _22881_, _22879_);
  nor (_22883_, _22882_, _02940_);
  not (_22884_, _22659_);
  and (_22885_, _09915_, \oc8051_golden_model_1.PC [0]);
  nor (_22886_, _22690_, _09915_);
  nor (_22887_, _22886_, _22885_);
  and (_22888_, _22887_, _02940_);
  nor (_22889_, _22888_, _22884_);
  not (_22890_, _22889_);
  nor (_22892_, _22890_, _22883_);
  nor (_22893_, _22892_, _22660_);
  nor (_22894_, _22893_, _04337_);
  and (_22895_, _04337_, _03486_);
  nor (_22896_, _22895_, _02497_);
  not (_22897_, _22896_);
  nor (_22898_, _22897_, _22894_);
  not (_22899_, _22657_);
  and (_22900_, _22887_, _02497_);
  nor (_22901_, _22900_, _22899_);
  not (_22903_, _22901_);
  nor (_22904_, _22903_, _22898_);
  nor (_22905_, _22904_, _22658_);
  nor (_22906_, _22655_, _22905_);
  or (_22907_, _22906_, _09979_);
  nor (_22908_, _22907_, _22656_);
  nor (_22909_, _22908_, _22653_);
  nand (_22910_, _22909_, _42668_);
  or (_22911_, _42668_, \oc8051_golden_model_1.PC [0]);
  and (_22912_, _22911_, _43998_);
  and (_43495_, _22912_, _22910_);
  and (_22914_, _09979_, _09270_);
  nand (_22915_, _02888_, _02215_);
  nor (_22916_, _09274_, _09272_);
  nor (_22917_, _22916_, _09275_);
  or (_22918_, _22917_, _09915_);
  nand (_22919_, _09915_, _09270_);
  and (_22920_, _22919_, _22918_);
  and (_22921_, _22920_, _02497_);
  or (_22922_, _09948_, _09270_);
  and (_22924_, _11949_, _05265_);
  or (_22925_, _22924_, _09270_);
  not (_22926_, _02537_);
  nand (_22927_, _07232_, _02552_);
  or (_22928_, _09066_, _09270_);
  or (_22929_, _09074_, _09270_);
  not (_22930_, _09080_);
  or (_22931_, _09081_, _09270_);
  or (_22932_, _07871_, _09270_);
  or (_22933_, _05753_, _02215_);
  or (_22934_, _09557_, _09270_);
  and (_22935_, _02945_, _03299_);
  nor (_22936_, _22935_, _02618_);
  not (_22937_, _22936_);
  nor (_22938_, _03859_, _03062_);
  and (_22939_, _22938_, _04131_);
  and (_22940_, _22939_, _22937_);
  or (_22941_, _22940_, _02215_);
  nand (_22942_, _09489_, _02552_);
  or (_22943_, _22917_, _09392_);
  nand (_22945_, _09392_, _09270_);
  and (_22946_, _22945_, _22943_);
  or (_22947_, _22946_, _09396_);
  nor (_22948_, _03698_, _02621_);
  or (_22949_, _09470_, _09270_);
  nor (_22950_, _03698_, _02611_);
  nor (_22951_, _22702_, _03813_);
  nand (_22952_, _22951_, _02215_);
  or (_22953_, _22951_, _02215_);
  and (_22954_, _22953_, _02611_);
  and (_22956_, _22954_, _22952_);
  or (_22957_, _22956_, _14356_);
  or (_22958_, _22957_, _22950_);
  or (_22959_, _09427_, _09270_);
  and (_22960_, _22959_, _03387_);
  and (_22961_, _22960_, _22958_);
  and (_22962_, _03072_, _02215_);
  or (_22963_, _22962_, _07646_);
  or (_22964_, _22963_, _22961_);
  nand (_22965_, _07646_, _02552_);
  and (_22967_, _22965_, _02616_);
  and (_22968_, _22967_, _22964_);
  nor (_22969_, _03698_, _02616_);
  or (_22970_, _22969_, _05363_);
  or (_22971_, _22970_, _22968_);
  nand (_22972_, _09420_, \oc8051_golden_model_1.PC [1]);
  nor (_22973_, _09145_, _09143_);
  nor (_22974_, _22973_, _09146_);
  or (_22975_, _22974_, _09420_);
  and (_22976_, _22975_, _22972_);
  or (_22978_, _22976_, _05362_);
  and (_22979_, _22978_, _22971_);
  or (_22980_, _22979_, _02886_);
  nand (_22981_, _02886_, _02552_);
  and (_22982_, _22981_, _03810_);
  and (_22983_, _22982_, _22980_);
  nand (_22984_, _09412_, _09270_);
  or (_22985_, _22917_, _09412_);
  and (_22986_, _22985_, _02974_);
  and (_22987_, _22986_, _22984_);
  or (_22989_, _22987_, _09406_);
  or (_22990_, _22989_, _22983_);
  or (_22991_, _09405_, _09270_);
  and (_22992_, _22991_, _02881_);
  and (_22993_, _22992_, _22990_);
  and (_22994_, _02880_, _02215_);
  or (_22995_, _22994_, _04252_);
  or (_22996_, _22995_, _22993_);
  nand (_22997_, _03698_, _04252_);
  and (_22998_, _22997_, _03336_);
  and (_23000_, _22998_, _22996_);
  and (_23001_, _03069_, _02215_);
  or (_23002_, _23001_, _09461_);
  or (_23003_, _23002_, _23000_);
  nand (_23004_, _09461_, _02552_);
  and (_23005_, _23004_, _03084_);
  and (_23006_, _23005_, _23003_);
  nand (_23007_, _03075_, _02215_);
  nand (_23008_, _23007_, _09470_);
  or (_23009_, _23008_, _23006_);
  and (_23011_, _23009_, _22949_);
  or (_23012_, _23011_, _02876_);
  nand (_23013_, _02876_, \oc8051_golden_model_1.PC [1]);
  and (_23014_, _23013_, _02621_);
  and (_23015_, _23014_, _23012_);
  or (_23016_, _23015_, _22948_);
  and (_23017_, _23016_, _03941_);
  nand (_23018_, _02875_, _02215_);
  nand (_23019_, _23018_, _09396_);
  or (_23020_, _23019_, _23017_);
  and (_23022_, _23020_, _22947_);
  or (_23023_, _23022_, _02978_);
  and (_23024_, _09357_, _02552_);
  not (_23025_, _09357_);
  and (_23026_, _22917_, _23025_);
  or (_23027_, _23026_, _02979_);
  or (_23028_, _23027_, _23024_);
  and (_23029_, _23028_, _09500_);
  and (_23030_, _23029_, _23023_);
  not (_23031_, _09514_);
  and (_23033_, _22917_, _23031_);
  and (_23034_, _09514_, _02552_);
  or (_23035_, _23034_, _23033_);
  and (_23036_, _23035_, _02950_);
  or (_23037_, _23036_, _23030_);
  and (_23038_, _23037_, _09531_);
  nand (_23039_, _09528_, _09270_);
  or (_23040_, _22917_, _09528_);
  and (_23041_, _23040_, _02952_);
  and (_23042_, _23041_, _23039_);
  or (_23044_, _23042_, _09489_);
  or (_23045_, _23044_, _23038_);
  and (_23046_, _23045_, _22942_);
  or (_23047_, _23046_, _02869_);
  nand (_23048_, _02869_, \oc8051_golden_model_1.PC [1]);
  and (_23049_, _23048_, _02614_);
  and (_23050_, _23049_, _23047_);
  not (_23051_, _22940_);
  nor (_23052_, _03698_, _02614_);
  or (_23053_, _23052_, _23051_);
  or (_23055_, _23053_, _23050_);
  and (_23056_, _23055_, _22941_);
  or (_23057_, _23056_, _09544_);
  or (_23058_, _09543_, _09270_);
  and (_23059_, _23058_, _09550_);
  and (_23060_, _23059_, _23057_);
  and (_23061_, _03101_, _02215_);
  or (_23062_, _23061_, _09551_);
  or (_23063_, _23062_, _23060_);
  nand (_23064_, _03698_, _09551_);
  and (_23066_, _23064_, _10016_);
  and (_23067_, _23066_, _23063_);
  nand (_23068_, _03100_, _02215_);
  nand (_23069_, _23068_, _09557_);
  or (_23070_, _23069_, _23067_);
  and (_23071_, _23070_, _22934_);
  or (_23072_, _23071_, _09562_);
  or (_23073_, _09561_, _02215_);
  and (_23074_, _23073_, _02605_);
  and (_23075_, _23074_, _23072_);
  and (_23077_, _02583_, _09270_);
  or (_23078_, _23077_, _02863_);
  or (_23079_, _23078_, _23075_);
  nand (_23080_, _02863_, \oc8051_golden_model_1.PC [1]);
  and (_23081_, _23080_, _23079_);
  or (_23082_, _23081_, _02581_);
  nand (_23083_, _03698_, _02581_);
  and (_23084_, _23083_, _08209_);
  and (_23085_, _23084_, _23082_);
  nand (_23086_, _02981_, _02552_);
  nand (_23088_, _23086_, _02857_);
  or (_23089_, _23088_, _23085_);
  or (_23090_, _02857_, _02215_);
  and (_23091_, _23090_, _02838_);
  and (_23092_, _23091_, _23089_);
  nand (_23093_, _02579_, _02552_);
  nand (_23094_, _23093_, _09200_);
  or (_23095_, _23094_, _23092_);
  or (_23096_, _09200_, _09270_);
  and (_23097_, _23096_, _03490_);
  and (_23099_, _23097_, _23095_);
  and (_23100_, _02933_, _02215_);
  or (_23101_, _23100_, _02518_);
  or (_23102_, _23101_, _23099_);
  nand (_23103_, _03698_, _02518_);
  and (_23104_, _23103_, _09599_);
  and (_23105_, _23104_, _23102_);
  and (_23106_, _22974_, _09594_);
  or (_23107_, _23106_, _05754_);
  or (_23108_, _23107_, _23105_);
  and (_23109_, _23108_, _22933_);
  or (_23110_, _23109_, _02802_);
  nand (_23111_, _02802_, _09270_);
  and (_23112_, _23111_, _07860_);
  and (_23113_, _23112_, _23110_);
  and (_23114_, _07859_, _02215_);
  or (_23115_, _23114_, _09611_);
  or (_23116_, _23115_, _23113_);
  or (_23117_, _22679_, _02692_);
  and (_23118_, _23117_, _03496_);
  and (_23121_, _23118_, _23116_);
  and (_23122_, _02932_, _02215_);
  or (_23123_, _23122_, _02514_);
  or (_23124_, _23123_, _23121_);
  nand (_23125_, _03698_, _02514_);
  and (_23126_, _23125_, _22678_);
  and (_23127_, _23126_, _23124_);
  or (_23128_, _22974_, _08165_);
  nand (_23129_, _08165_, \oc8051_golden_model_1.PC [1]);
  and (_23130_, _23129_, _09083_);
  nand (_23132_, _23130_, _23128_);
  nand (_23133_, _23132_, _07871_);
  or (_23134_, _23133_, _23127_);
  nand (_23135_, _23134_, _22932_);
  nor (_23136_, _15733_, _03499_);
  and (_23137_, _23136_, _07873_);
  nand (_23138_, _23137_, _23135_);
  or (_23139_, _23137_, _09270_);
  and (_23140_, _23139_, _15555_);
  and (_23141_, _23140_, _23138_);
  nand (_23142_, _03504_, _09270_);
  nand (_23143_, _23142_, _09660_);
  or (_23144_, _23143_, _23141_);
  or (_23145_, _09660_, _02215_);
  and (_23146_, _23145_, _03887_);
  and (_23147_, _23146_, _23144_);
  and (_23148_, _02980_, _02552_);
  or (_23149_, _23148_, _03127_);
  or (_23150_, _23149_, _23147_);
  nand (_23151_, _03127_, \oc8051_golden_model_1.PC [1]);
  and (_23154_, _23151_, _23150_);
  or (_23155_, _23154_, _02509_);
  nand (_23156_, _03698_, _02509_);
  and (_23157_, _23156_, _22675_);
  and (_23158_, _23157_, _23155_);
  or (_23159_, _22974_, _09676_);
  or (_23160_, _08165_, _02215_);
  and (_23161_, _23160_, _09672_);
  and (_23162_, _23161_, _23159_);
  or (_23163_, _23162_, _09681_);
  or (_23165_, _23163_, _23158_);
  and (_23166_, _23165_, _22931_);
  or (_23167_, _23166_, _22930_);
  or (_23168_, _09080_, _02215_);
  and (_23169_, _23168_, _03883_);
  and (_23170_, _23169_, _23167_);
  and (_23171_, _02970_, _02552_);
  or (_23172_, _23171_, _03135_);
  or (_23173_, _23172_, _23170_);
  nand (_23174_, _03135_, \oc8051_golden_model_1.PC [1]);
  and (_23175_, _23174_, _23173_);
  or (_23176_, _23175_, _03880_);
  nand (_23177_, _03698_, _03880_);
  and (_23178_, _23177_, _22667_);
  and (_23179_, _23178_, _23176_);
  or (_23180_, _22974_, \oc8051_golden_model_1.PSW [7]);
  nand (_23181_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_23182_, _23181_, _09076_);
  and (_23183_, _23182_, _23180_);
  or (_23184_, _23183_, _09694_);
  or (_23187_, _23184_, _23179_);
  and (_23188_, _23187_, _22929_);
  or (_23189_, _23188_, _07944_);
  or (_23190_, _07943_, _02215_);
  and (_23191_, _23190_, _05783_);
  and (_23192_, _23191_, _23189_);
  and (_23193_, _02965_, _02552_);
  or (_23194_, _23193_, _03123_);
  or (_23195_, _23194_, _23192_);
  nand (_23196_, _03123_, \oc8051_golden_model_1.PC [1]);
  and (_23198_, _23196_, _23195_);
  or (_23199_, _23198_, _09069_);
  not (_23200_, _09068_);
  nand (_23201_, _03698_, _09069_);
  and (_23202_, _23201_, _23200_);
  and (_23203_, _23202_, _23199_);
  or (_23204_, _22974_, _07293_);
  or (_23205_, \oc8051_golden_model_1.PSW [7], _02215_);
  and (_23206_, _23205_, _09068_);
  and (_23207_, _23206_, _23204_);
  or (_23208_, _23207_, _09711_);
  or (_23209_, _23208_, _23203_);
  and (_23210_, _23209_, _22928_);
  or (_23211_, _23210_, _10365_);
  or (_23212_, _09065_, _02215_);
  and (_23213_, _23212_, _07992_);
  and (_23214_, _23213_, _23211_);
  and (_23215_, _07991_, _09270_);
  or (_23216_, _23215_, _03145_);
  or (_23217_, _23216_, _23214_);
  or (_23220_, _06151_, _09726_);
  and (_23221_, _23220_, _23217_);
  or (_23222_, _23221_, _03898_);
  nand (_23223_, _03698_, _03898_);
  and (_23224_, _23223_, _03561_);
  and (_23225_, _23224_, _23222_);
  not (_23226_, _09915_);
  or (_23227_, _22917_, _23226_);
  or (_23228_, _09915_, _02552_);
  and (_23229_, _23228_, _02968_);
  and (_23231_, _23229_, _23227_);
  or (_23232_, _23231_, _07232_);
  or (_23233_, _23232_, _23225_);
  nand (_23234_, _23233_, _22927_);
  and (_23235_, _05747_, _02891_);
  nor (_23236_, _23235_, _07229_);
  and (_23237_, _23236_, _07236_);
  nand (_23238_, _23237_, _23234_);
  and (_23239_, _03411_, _02891_);
  nor (_23240_, _23237_, _09270_);
  nor (_23241_, _23240_, _23239_);
  and (_23242_, _23241_, _23238_);
  nand (_23243_, _23239_, _09270_);
  nand (_23244_, _23243_, _08066_);
  or (_23245_, _23244_, _23242_);
  or (_23246_, _08066_, _02215_);
  and (_23247_, _23246_, _08112_);
  and (_23248_, _23247_, _23245_);
  and (_23249_, _08111_, _09270_);
  or (_23250_, _23249_, _02892_);
  or (_23253_, _23250_, _23248_);
  or (_23254_, _06151_, _02893_);
  and (_23255_, _23254_, _23253_);
  or (_23256_, _23255_, _22926_);
  nand (_23257_, _03698_, _22926_);
  and (_23258_, _23257_, _03164_);
  and (_23259_, _23258_, _23256_);
  nand (_23260_, _22920_, _02940_);
  nand (_23261_, _23260_, _22924_);
  or (_23262_, _23261_, _23259_);
  nand (_23264_, _23262_, _22925_);
  not (_23265_, _02367_);
  nor (_23266_, _05748_, _23265_);
  nor (_23267_, _23266_, _03576_);
  nand (_23268_, _23267_, _23264_);
  or (_23269_, _23267_, _09270_);
  and (_23270_, _23269_, _03906_);
  and (_23271_, _23270_, _23268_);
  nand (_23272_, _03163_, _02215_);
  nand (_23273_, _23272_, _09948_);
  or (_23274_, _23273_, _23271_);
  and (_23275_, _23274_, _22922_);
  or (_23276_, _23275_, _04337_);
  nand (_23277_, _04337_, _03698_);
  and (_23278_, _23277_, _02498_);
  and (_23279_, _23278_, _23276_);
  or (_23280_, _23279_, _22921_);
  nand (_23281_, _23280_, _05237_);
  nor (_23282_, _05237_, _02552_);
  nor (_23283_, _23282_, _03920_);
  and (_23286_, _23283_, _23281_);
  and (_23287_, _03920_, _02552_);
  or (_23288_, _23287_, _02888_);
  or (_23289_, _23288_, _23286_);
  and (_23290_, _23289_, _22915_);
  nor (_23291_, _23290_, _09970_);
  nor (_23292_, _09044_, _02552_);
  nor (_23293_, _23292_, _22655_);
  not (_23294_, _23293_);
  nor (_23295_, _23294_, _23291_);
  and (_23297_, _22655_, _03698_);
  or (_23298_, _23297_, _09979_);
  nor (_23299_, _23298_, _23295_);
  or (_23300_, _23299_, _22914_);
  or (_23301_, _23300_, _42672_);
  or (_23302_, _42668_, \oc8051_golden_model_1.PC [1]);
  and (_23303_, _23302_, _43998_);
  and (_43496_, _23303_, _23301_);
  and (_23304_, _09979_, _02549_);
  and (_23305_, _02888_, _02648_);
  nand (_23306_, _03163_, _02648_);
  nor (_23307_, _09063_, _02549_);
  nor (_23308_, _09066_, _02549_);
  nor (_23309_, _09074_, _02549_);
  nor (_23310_, _09081_, _02549_);
  nor (_23311_, _09657_, _02549_);
  nor (_23312_, _09200_, _02549_);
  nor (_23313_, _02851_, _02648_);
  and (_23314_, _02863_, _09140_);
  nor (_23315_, _22940_, _02648_);
  and (_23318_, _09489_, _02995_);
  and (_23319_, _09279_, _09276_);
  nor (_23320_, _23319_, _09280_);
  nor (_23321_, _23320_, _09412_);
  and (_23322_, _09268_, _09412_);
  or (_23323_, _23322_, _23321_);
  and (_23324_, _23323_, _02974_);
  nand (_23325_, _09420_, _02648_);
  and (_23326_, _09150_, _09147_);
  or (_23327_, _23326_, _09151_);
  or (_23329_, _23327_, _09420_);
  and (_23330_, _23329_, _23325_);
  and (_23331_, _23330_, _05363_);
  or (_23332_, _03297_, _02611_);
  nand (_23333_, _09429_, _02549_);
  or (_23334_, _09429_, _02220_);
  and (_23335_, _23334_, _23333_);
  or (_23336_, _23335_, _03813_);
  not (_23337_, _07636_);
  nand (_23338_, _03813_, _02648_);
  and (_23340_, _23338_, _23337_);
  and (_23341_, _23340_, _23336_);
  and (_23342_, _07636_, _02995_);
  or (_23343_, _23342_, _03818_);
  or (_23344_, _23343_, _23341_);
  and (_23345_, _23344_, _09427_);
  and (_23346_, _23345_, _23332_);
  nor (_23347_, _09427_, _02549_);
  or (_23348_, _23347_, _03072_);
  or (_23349_, _23348_, _23346_);
  nand (_23351_, _03072_, _02648_);
  and (_23352_, _23351_, _09426_);
  and (_23353_, _23352_, _23349_);
  and (_23354_, _07646_, _02995_);
  or (_23355_, _23354_, _09425_);
  or (_23356_, _23355_, _23353_);
  or (_23357_, _03297_, _02616_);
  and (_23358_, _23357_, _05362_);
  and (_23359_, _23358_, _23356_);
  or (_23360_, _23359_, _02886_);
  or (_23362_, _23360_, _23331_);
  nand (_23363_, _02886_, _02549_);
  and (_23364_, _23363_, _03810_);
  and (_23365_, _23364_, _23362_);
  or (_23366_, _23365_, _23324_);
  and (_23367_, _23366_, _09405_);
  nor (_23368_, _09405_, _02549_);
  or (_23369_, _23368_, _02880_);
  or (_23370_, _23369_, _23367_);
  nand (_23371_, _02880_, _02648_);
  and (_23373_, _23371_, _02609_);
  and (_23374_, _23373_, _23370_);
  and (_23375_, _03297_, _04252_);
  or (_23376_, _23375_, _03069_);
  or (_23377_, _23376_, _23374_);
  and (_23378_, _03069_, _02648_);
  nor (_23379_, _23378_, _09461_);
  and (_23380_, _23379_, _23377_);
  and (_23381_, _09461_, _02995_);
  or (_23382_, _23381_, _03075_);
  or (_23384_, _23382_, _23380_);
  nand (_23385_, _03075_, _02648_);
  and (_23386_, _23385_, _09470_);
  and (_23387_, _23386_, _23384_);
  nor (_23388_, _09470_, _02549_);
  or (_23389_, _23388_, _02876_);
  or (_23390_, _23389_, _23387_);
  nand (_23391_, _02876_, _02648_);
  and (_23392_, _23391_, _02621_);
  and (_23393_, _23392_, _23390_);
  and (_23395_, _03297_, _09474_);
  or (_23396_, _23395_, _02875_);
  or (_23397_, _23396_, _23393_);
  nand (_23398_, _02875_, _02648_);
  and (_23399_, _23398_, _09396_);
  and (_23400_, _23399_, _23397_);
  nand (_23401_, _09392_, _09267_);
  not (_23402_, _23320_);
  or (_23403_, _23402_, _09392_);
  and (_23404_, _23403_, _23401_);
  and (_23406_, _23404_, _09481_);
  or (_23407_, _23406_, _02978_);
  or (_23408_, _23407_, _23400_);
  nor (_23409_, _23320_, _09357_);
  and (_23410_, _09357_, _09268_);
  or (_23411_, _23410_, _02979_);
  or (_23412_, _23411_, _23409_);
  and (_23413_, _23412_, _09500_);
  and (_23414_, _23413_, _23408_);
  or (_23415_, _23402_, _09514_);
  nand (_23417_, _09514_, _09267_);
  and (_23418_, _23417_, _02950_);
  and (_23419_, _23418_, _23415_);
  or (_23420_, _23419_, _02952_);
  or (_23421_, _23420_, _23414_);
  nor (_23422_, _23320_, _09528_);
  and (_23423_, _09528_, _09268_);
  or (_23424_, _23423_, _09531_);
  or (_23425_, _23424_, _23422_);
  and (_23426_, _23425_, _09490_);
  and (_23428_, _23426_, _23421_);
  or (_23429_, _23428_, _23318_);
  and (_23430_, _23429_, _02870_);
  and (_23431_, _02869_, _09140_);
  or (_23432_, _23431_, _04095_);
  or (_23433_, _23432_, _23430_);
  or (_23434_, _03297_, _02614_);
  and (_23435_, _23434_, _22940_);
  and (_23436_, _23435_, _23433_);
  or (_23437_, _23436_, _23315_);
  and (_23439_, _23437_, _09543_);
  nor (_23440_, _09543_, _02549_);
  or (_23441_, _23440_, _03101_);
  or (_23442_, _23441_, _23439_);
  nand (_23443_, _03101_, _02648_);
  and (_23444_, _23443_, _02619_);
  and (_23445_, _23444_, _23442_);
  and (_23446_, _03297_, _09551_);
  or (_23447_, _23446_, _03100_);
  or (_23448_, _23447_, _23445_);
  nand (_23450_, _03100_, _02648_);
  and (_23451_, _23450_, _09557_);
  and (_23452_, _23451_, _23448_);
  nor (_23453_, _09557_, _02549_);
  or (_23454_, _23453_, _23452_);
  and (_23455_, _23454_, _09561_);
  nor (_23456_, _09561_, _02648_);
  or (_23457_, _23456_, _02583_);
  or (_23458_, _23457_, _23455_);
  nand (_23459_, _02583_, _02549_);
  and (_23461_, _23459_, _02864_);
  and (_23462_, _23461_, _23458_);
  or (_23463_, _23462_, _23314_);
  and (_23464_, _23463_, _04251_);
  and (_23465_, _03297_, _02581_);
  or (_23466_, _23465_, _02981_);
  or (_23467_, _23466_, _23464_);
  nand (_23468_, _09267_, _02981_);
  and (_23469_, _23468_, _02851_);
  and (_23470_, _23469_, _23467_);
  or (_23472_, _23470_, _23313_);
  and (_23473_, _23472_, _02856_);
  nor (_23474_, _02856_, _02648_);
  or (_23475_, _23474_, _02579_);
  or (_23476_, _23475_, _23473_);
  nand (_23477_, _09267_, _02579_);
  and (_23478_, _23477_, _09200_);
  and (_23479_, _23478_, _23476_);
  or (_23480_, _23479_, _23312_);
  and (_23481_, _23480_, _03490_);
  and (_23483_, _02933_, _09140_);
  or (_23484_, _23483_, _02518_);
  or (_23485_, _23484_, _23481_);
  or (_23486_, _03297_, _22795_);
  and (_23487_, _23486_, _09599_);
  and (_23488_, _23487_, _23485_);
  and (_23489_, _23327_, _09594_);
  nor (_23490_, _23489_, _23488_);
  nor (_23491_, _23490_, _04146_);
  and (_23492_, _04146_, _09140_);
  or (_23494_, _23492_, _04145_);
  not (_23495_, _05750_);
  not (_23496_, _04129_);
  or (_23497_, _23496_, _04102_);
  or (_23498_, _23497_, _23495_);
  or (_23499_, _23498_, _23494_);
  or (_23500_, _23499_, _23491_);
  nor (_23501_, _23498_, _04145_);
  or (_23502_, _23501_, _09140_);
  and (_23503_, _23502_, _02803_);
  and (_23505_, _23503_, _23500_);
  and (_23506_, _09268_, _02802_);
  or (_23507_, _23506_, _07859_);
  or (_23508_, _23507_, _23505_);
  nand (_23509_, _07859_, _02648_);
  and (_23510_, _23509_, _22679_);
  and (_23511_, _23510_, _23508_);
  nor (_23512_, _22679_, _02653_);
  or (_23513_, _23512_, _02932_);
  or (_23514_, _23513_, _23511_);
  nand (_23516_, _02932_, _02648_);
  and (_23517_, _23516_, _04093_);
  and (_23518_, _23517_, _23514_);
  and (_23519_, _03297_, _02514_);
  or (_23520_, _23519_, _09083_);
  or (_23521_, _23520_, _23518_);
  and (_23522_, _23327_, _09676_);
  nand (_23523_, _08165_, _09140_);
  nand (_23524_, _23523_, _09083_);
  or (_23525_, _23524_, _23522_);
  and (_23527_, _23525_, _09657_);
  and (_23528_, _23527_, _23521_);
  or (_23529_, _23528_, _23311_);
  and (_23530_, _23529_, _09660_);
  nor (_23531_, _09660_, _02648_);
  or (_23532_, _23531_, _02980_);
  or (_23533_, _23532_, _23530_);
  nand (_23534_, _09267_, _02980_);
  and (_23535_, _23534_, _03128_);
  and (_23536_, _23535_, _23533_);
  and (_23538_, _03127_, _09140_);
  or (_23539_, _23538_, _23536_);
  and (_23540_, _23539_, _02510_);
  and (_23541_, _03297_, _02509_);
  or (_23542_, _23541_, _09672_);
  or (_23543_, _23542_, _23540_);
  and (_23544_, _23327_, _08165_);
  or (_23545_, _08165_, _02648_);
  nand (_23546_, _23545_, _09672_);
  or (_23547_, _23546_, _23544_);
  and (_23549_, _23547_, _09081_);
  and (_23550_, _23549_, _23543_);
  or (_23551_, _23550_, _23310_);
  and (_23552_, _23551_, _09080_);
  nor (_23553_, _09080_, _02648_);
  or (_23554_, _23553_, _02970_);
  or (_23555_, _23554_, _23552_);
  nand (_23556_, _09267_, _02970_);
  and (_23557_, _23556_, _03137_);
  and (_23558_, _23557_, _23555_);
  and (_23560_, _03135_, _09140_);
  or (_23561_, _23560_, _23558_);
  and (_23562_, _23561_, _02532_);
  and (_23563_, _03297_, _03880_);
  or (_23564_, _23563_, _09076_);
  or (_23565_, _23564_, _23562_);
  and (_23566_, _23327_, _07293_);
  or (_23567_, _02648_, _07293_);
  nand (_23568_, _23567_, _09076_);
  or (_23569_, _23568_, _23566_);
  and (_23571_, _23569_, _09074_);
  and (_23572_, _23571_, _23565_);
  or (_23573_, _23572_, _23309_);
  and (_23574_, _23573_, _07943_);
  nor (_23575_, _07943_, _02648_);
  or (_23576_, _23575_, _02965_);
  or (_23577_, _23576_, _23574_);
  nand (_23578_, _09267_, _02965_);
  and (_23579_, _23578_, _05788_);
  and (_23580_, _23579_, _23577_);
  and (_23582_, _03123_, _09140_);
  or (_23583_, _23582_, _23580_);
  and (_23584_, _23583_, _02535_);
  and (_23585_, _03297_, _09069_);
  or (_23586_, _23585_, _09068_);
  or (_23587_, _23586_, _23584_);
  and (_23588_, _23327_, \oc8051_golden_model_1.PSW [7]);
  or (_23589_, _02648_, \oc8051_golden_model_1.PSW [7]);
  nand (_23590_, _23589_, _09068_);
  or (_23591_, _23590_, _23588_);
  and (_23593_, _23591_, _09066_);
  and (_23594_, _23593_, _23587_);
  or (_23595_, _23594_, _23308_);
  and (_23596_, _23595_, _09065_);
  nor (_23597_, _09065_, _02648_);
  or (_23598_, _23597_, _07991_);
  or (_23599_, _23598_, _23596_);
  nand (_23600_, _07991_, _02549_);
  and (_23601_, _23600_, _09726_);
  and (_23602_, _23601_, _23599_);
  and (_23604_, _06031_, _03145_);
  or (_23605_, _23604_, _23602_);
  and (_23606_, _23605_, _02529_);
  and (_23607_, _03297_, _03898_);
  or (_23608_, _23607_, _02968_);
  or (_23609_, _23608_, _23606_);
  nor (_23610_, _09915_, _09267_);
  and (_23611_, _23402_, _09915_);
  or (_23612_, _23611_, _03561_);
  or (_23613_, _23612_, _23610_);
  and (_23615_, _23613_, _09063_);
  and (_23616_, _23615_, _23609_);
  or (_23617_, _23616_, _23307_);
  and (_23618_, _23617_, _08066_);
  nor (_23619_, _08066_, _02648_);
  or (_23620_, _23619_, _08111_);
  or (_23621_, _23620_, _23618_);
  nand (_23622_, _08111_, _02549_);
  and (_23623_, _23622_, _02893_);
  and (_23624_, _23623_, _23621_);
  and (_23626_, _06031_, _02892_);
  or (_23627_, _23626_, _23624_);
  and (_23628_, _23627_, _02537_);
  and (_23629_, _03297_, _22926_);
  or (_23630_, _23629_, _02940_);
  or (_23631_, _23630_, _23628_);
  nor (_23632_, _23320_, _09915_);
  and (_23633_, _09915_, _09268_);
  nor (_23634_, _23633_, _23632_);
  nand (_23635_, _23634_, _02940_);
  and (_23637_, _23635_, _09941_);
  and (_23638_, _23637_, _23631_);
  nor (_23639_, _09941_, _02549_);
  or (_23640_, _23639_, _03163_);
  or (_23641_, _23640_, _23638_);
  and (_23642_, _23641_, _23306_);
  nor (_23643_, _23642_, _09949_);
  nor (_23644_, _09948_, _02995_);
  or (_23645_, _23644_, _04337_);
  or (_23646_, _23645_, _23643_);
  nand (_23648_, _04337_, _03297_);
  and (_23649_, _23648_, _02498_);
  and (_23650_, _23649_, _23646_);
  and (_23651_, _23634_, _02497_);
  or (_23652_, _23651_, _09964_);
  or (_23653_, _23652_, _23650_);
  nand (_23654_, _09964_, _02995_);
  and (_23655_, _23654_, _02890_);
  and (_23656_, _23655_, _23653_);
  or (_23657_, _23656_, _23305_);
  and (_23659_, _23657_, _09044_);
  nor (_23660_, _09044_, _02995_);
  or (_23661_, _23660_, _22655_);
  or (_23662_, _23661_, _23659_);
  nand (_23663_, _22655_, _03297_);
  and (_23664_, _23663_, _09983_);
  and (_23665_, _23664_, _23662_);
  or (_23666_, _23665_, _23304_);
  or (_23667_, _23666_, _42672_);
  or (_23668_, _42668_, \oc8051_golden_model_1.PC [2]);
  and (_23670_, _23668_, _43998_);
  and (_43497_, _23670_, _23667_);
  and (_23671_, _09979_, _02606_);
  and (_23672_, _22655_, _03057_);
  or (_23673_, _23672_, _09979_);
  and (_23674_, _02888_, _02629_);
  and (_23675_, _03163_, _02629_);
  nor (_23676_, _09063_, _02606_);
  nor (_23677_, _09066_, _02606_);
  nor (_23678_, _09074_, _02606_);
  nor (_23680_, _09081_, _02606_);
  nor (_23681_, _09657_, _02606_);
  nor (_23682_, _05753_, _02629_);
  nor (_23683_, _02857_, _02629_);
  or (_23684_, _23683_, _02579_);
  nor (_23685_, _22940_, _02629_);
  and (_23686_, _09489_, _02567_);
  and (_23687_, _09263_, _09412_);
  or (_23688_, _09265_, _09264_);
  and (_23689_, _23688_, _09281_);
  nor (_23691_, _23688_, _09281_);
  nor (_23692_, _23691_, _23689_);
  nor (_23693_, _23692_, _09412_);
  nor (_23694_, _23693_, _23687_);
  or (_23695_, _23694_, _03810_);
  or (_23696_, _09139_, _09138_);
  and (_23697_, _23696_, _09152_);
  nor (_23698_, _23696_, _09152_);
  nor (_23699_, _23698_, _23697_);
  or (_23700_, _23699_, _09420_);
  nand (_23702_, _09420_, _02641_);
  and (_23703_, _23702_, _23700_);
  nor (_23704_, _23703_, _05362_);
  nor (_23705_, _09429_, \oc8051_golden_model_1.PC [3]);
  nor (_23706_, _23705_, _03813_);
  and (_23707_, _03813_, _02629_);
  nor (_23708_, _23707_, _07636_);
  not (_23709_, _23708_);
  nor (_23710_, _23709_, _23706_);
  not (_23711_, _23710_);
  nor (_23713_, _09430_, _02606_);
  nor (_23714_, _23713_, _03818_);
  and (_23715_, _23714_, _23711_);
  nor (_23716_, _03057_, _02611_);
  or (_23717_, _23716_, _14356_);
  nor (_23718_, _23717_, _23715_);
  nor (_23719_, _09427_, _02606_);
  nor (_23720_, _23719_, _03072_);
  not (_23721_, _23720_);
  nor (_23722_, _23721_, _23718_);
  and (_23724_, _03072_, _02629_);
  or (_23725_, _23724_, _23722_);
  and (_23726_, _23725_, _09426_);
  and (_23727_, _07646_, _02606_);
  or (_23728_, _23727_, _23726_);
  and (_23729_, _23728_, _02616_);
  nor (_23730_, _03057_, _02616_);
  nor (_23731_, _23730_, _05363_);
  not (_23732_, _23731_);
  nor (_23733_, _23732_, _23729_);
  or (_23735_, _23733_, _02886_);
  nor (_23736_, _23735_, _23704_);
  and (_23737_, _02886_, _02606_);
  or (_23738_, _23737_, _02974_);
  or (_23739_, _23738_, _23736_);
  and (_23740_, _23739_, _23695_);
  nor (_23741_, _23740_, _09406_);
  nor (_23742_, _09405_, _02606_);
  nor (_23743_, _23742_, _02880_);
  not (_23744_, _23743_);
  nor (_23746_, _23744_, _23741_);
  and (_23747_, _02880_, _02629_);
  nor (_23748_, _23747_, _23746_);
  or (_23749_, _23748_, _04252_);
  or (_23750_, _03057_, _02609_);
  and (_23751_, _23750_, _23749_);
  or (_23752_, _23751_, _03069_);
  and (_23753_, _03069_, _02629_);
  nor (_23754_, _23753_, _09461_);
  nand (_23755_, _23754_, _23752_);
  and (_23757_, _09461_, _02567_);
  nor (_23758_, _23757_, _03075_);
  nand (_23759_, _23758_, _23755_);
  and (_23760_, _03075_, _02629_);
  nor (_23761_, _23760_, _09471_);
  nand (_23762_, _23761_, _23759_);
  nor (_23763_, _09470_, _02606_);
  nor (_23764_, _23763_, _02876_);
  nand (_23765_, _23764_, _23762_);
  and (_23766_, _02876_, _02629_);
  nor (_23768_, _23766_, _09474_);
  nand (_23769_, _23768_, _23765_);
  and (_23770_, _03057_, _09474_);
  nor (_23771_, _23770_, _02875_);
  nand (_23772_, _23771_, _23769_);
  and (_23773_, _02875_, _02629_);
  nor (_23774_, _23773_, _09481_);
  nand (_23775_, _23774_, _23772_);
  and (_23776_, _09392_, _09262_);
  not (_23777_, _23692_);
  nor (_23779_, _23777_, _09392_);
  or (_23780_, _23779_, _23776_);
  nor (_23781_, _23780_, _09396_);
  nor (_23782_, _23781_, _02978_);
  and (_23783_, _23782_, _23775_);
  nor (_23784_, _23692_, _09357_);
  and (_23785_, _09357_, _09263_);
  or (_23786_, _23785_, _02979_);
  nor (_23787_, _23786_, _23784_);
  or (_23788_, _23787_, _02950_);
  or (_23790_, _23788_, _23783_);
  nor (_23791_, _23777_, _09514_);
  and (_23792_, _09514_, _09262_);
  or (_23793_, _23792_, _09500_);
  or (_23794_, _23793_, _23791_);
  and (_23795_, _23794_, _09531_);
  nand (_23796_, _23795_, _23790_);
  nor (_23797_, _23692_, _09528_);
  and (_23798_, _09528_, _09263_);
  or (_23799_, _23798_, _09531_);
  nor (_23801_, _23799_, _23797_);
  nor (_23802_, _23801_, _09489_);
  and (_23803_, _23802_, _23796_);
  or (_23804_, _23803_, _23686_);
  nand (_23805_, _23804_, _02870_);
  and (_23806_, _02869_, _02641_);
  nor (_23807_, _23806_, _04095_);
  nand (_23808_, _23807_, _23805_);
  nor (_23809_, _03057_, _02614_);
  nor (_23810_, _23809_, _23051_);
  and (_23812_, _23810_, _23808_);
  or (_23813_, _23812_, _23685_);
  nand (_23814_, _23813_, _09543_);
  nor (_23815_, _09543_, _02606_);
  nor (_23816_, _23815_, _03101_);
  nand (_23817_, _23816_, _23814_);
  and (_23818_, _03101_, _02629_);
  nor (_23819_, _23818_, _09551_);
  nand (_23820_, _23819_, _23817_);
  and (_23821_, _03057_, _09551_);
  nor (_23823_, _23821_, _03100_);
  nand (_23824_, _23823_, _23820_);
  and (_23825_, _03100_, _02629_);
  nor (_23826_, _23825_, _14649_);
  and (_23827_, _23826_, _23824_);
  nor (_23828_, _09557_, _02606_);
  or (_23829_, _23828_, _23827_);
  nand (_23830_, _23829_, _09561_);
  nor (_23831_, _09561_, _02629_);
  nor (_23832_, _23831_, _02583_);
  and (_23834_, _23832_, _23830_);
  and (_23835_, _02583_, _02606_);
  or (_23836_, _23835_, _02863_);
  nor (_23837_, _23836_, _23834_);
  and (_23838_, _02863_, _02641_);
  or (_23839_, _23838_, _23837_);
  nand (_23840_, _23839_, _04251_);
  and (_23841_, _03057_, _02581_);
  nor (_23842_, _23841_, _02981_);
  nand (_23843_, _23842_, _23840_);
  and (_23845_, _09262_, _02981_);
  nor (_23846_, _23845_, _09582_);
  and (_23847_, _23846_, _23843_);
  or (_23848_, _23847_, _23684_);
  and (_23849_, _09262_, _02579_);
  nor (_23850_, _23849_, _09203_);
  nand (_23851_, _23850_, _23848_);
  nor (_23852_, _09200_, _02606_);
  nor (_23853_, _23852_, _02933_);
  nand (_23854_, _23853_, _23851_);
  and (_23856_, _02933_, _02629_);
  nor (_23857_, _23856_, _02518_);
  nand (_23858_, _23857_, _23854_);
  and (_23859_, _03057_, _02518_);
  nor (_23860_, _23859_, _09594_);
  nand (_23861_, _23860_, _23858_);
  and (_23862_, _23699_, _09594_);
  nor (_23863_, _23862_, _05754_);
  and (_23864_, _23863_, _23861_);
  or (_23865_, _23864_, _23682_);
  nand (_23867_, _23865_, _02803_);
  and (_23868_, _09263_, _02802_);
  nor (_23869_, _23868_, _07859_);
  nand (_23870_, _23869_, _23867_);
  and (_23871_, _07859_, _02629_);
  nor (_23872_, _23871_, _09611_);
  nand (_23873_, _23872_, _23870_);
  nor (_23874_, _22679_, _02602_);
  nor (_23875_, _23874_, _02932_);
  and (_23876_, _23875_, _23873_);
  and (_23878_, _02932_, _02629_);
  or (_23879_, _23878_, _02514_);
  or (_23880_, _23879_, _23876_);
  and (_23881_, _03057_, _02514_);
  nor (_23882_, _23881_, _09083_);
  nand (_23883_, _23882_, _23880_);
  not (_23884_, _09657_);
  and (_23885_, _08165_, _02629_);
  and (_23886_, _23699_, _09676_);
  or (_23887_, _23886_, _23885_);
  and (_23889_, _23887_, _09083_);
  nor (_23890_, _23889_, _23884_);
  and (_23891_, _23890_, _23883_);
  or (_23892_, _23891_, _23681_);
  nand (_23893_, _23892_, _09660_);
  nor (_23894_, _09660_, _02629_);
  nor (_23895_, _23894_, _02980_);
  and (_23896_, _23895_, _23893_);
  and (_23897_, _09262_, _02980_);
  or (_23898_, _23897_, _03127_);
  nor (_23900_, _23898_, _23896_);
  and (_23901_, _03127_, _02641_);
  or (_23902_, _23901_, _23900_);
  nand (_23903_, _23902_, _02510_);
  and (_23904_, _03057_, _02509_);
  nor (_23905_, _23904_, _09672_);
  nand (_23906_, _23905_, _23903_);
  nor (_23907_, _08165_, _02641_);
  and (_23908_, _23699_, _08165_);
  or (_23909_, _23908_, _23907_);
  and (_23911_, _23909_, _09672_);
  nor (_23912_, _23911_, _09681_);
  and (_23913_, _23912_, _23906_);
  or (_23914_, _23913_, _23680_);
  nand (_23915_, _23914_, _09080_);
  nor (_23916_, _09080_, _02629_);
  nor (_23917_, _23916_, _02970_);
  and (_23918_, _23917_, _23915_);
  and (_23919_, _09262_, _02970_);
  or (_23920_, _23919_, _03135_);
  nor (_23922_, _23920_, _23918_);
  and (_23923_, _03135_, _02641_);
  or (_23924_, _23923_, _23922_);
  nand (_23925_, _23924_, _02532_);
  and (_23926_, _03057_, _03880_);
  nor (_23927_, _23926_, _09076_);
  nand (_23928_, _23927_, _23925_);
  nor (_23929_, _23699_, \oc8051_golden_model_1.PSW [7]);
  nor (_23930_, _02629_, _07293_);
  nor (_23931_, _23930_, _22667_);
  not (_23933_, _23931_);
  nor (_23934_, _23933_, _23929_);
  nor (_23935_, _23934_, _09694_);
  and (_23936_, _23935_, _23928_);
  or (_23937_, _23936_, _23678_);
  nand (_23938_, _23937_, _07943_);
  nor (_23939_, _07943_, _02629_);
  nor (_23940_, _23939_, _02965_);
  and (_23941_, _23940_, _23938_);
  and (_23942_, _09262_, _02965_);
  or (_23944_, _23942_, _03123_);
  nor (_23945_, _23944_, _23941_);
  and (_23946_, _03123_, _02641_);
  or (_23947_, _23946_, _23945_);
  nand (_23948_, _23947_, _02535_);
  and (_23949_, _03057_, _09069_);
  nor (_23950_, _23949_, _09068_);
  nand (_23951_, _23950_, _23948_);
  nor (_23952_, _23699_, _07293_);
  nor (_23953_, _02629_, \oc8051_golden_model_1.PSW [7]);
  nor (_23955_, _23953_, _23200_);
  not (_23956_, _23955_);
  nor (_23957_, _23956_, _23952_);
  nor (_23958_, _23957_, _09711_);
  and (_23959_, _23958_, _23951_);
  or (_23960_, _23959_, _23677_);
  nand (_23961_, _23960_, _09065_);
  nor (_23962_, _09065_, _02629_);
  nor (_23963_, _23962_, _07991_);
  and (_23964_, _23963_, _23961_);
  and (_23966_, _07991_, _02606_);
  or (_23967_, _23966_, _03145_);
  nor (_23968_, _23967_, _23964_);
  and (_23969_, _05986_, _03145_);
  or (_23970_, _23969_, _23968_);
  nand (_23971_, _23970_, _02529_);
  and (_23972_, _03057_, _03898_);
  nor (_23973_, _23972_, _02968_);
  nand (_23974_, _23973_, _23971_);
  and (_23975_, _23777_, _09915_);
  nor (_23977_, _09915_, _09262_);
  or (_23978_, _23977_, _03561_);
  or (_23979_, _23978_, _23975_);
  and (_23980_, _23979_, _09063_);
  and (_23981_, _23980_, _23974_);
  or (_23982_, _23981_, _23676_);
  nand (_23983_, _23982_, _08066_);
  nor (_23984_, _08066_, _02629_);
  nor (_23985_, _23984_, _08111_);
  nand (_23986_, _23985_, _23983_);
  and (_23988_, _08111_, _02606_);
  nor (_23989_, _23988_, _02892_);
  and (_23990_, _23989_, _23986_);
  and (_23991_, _05986_, _02892_);
  or (_23992_, _23991_, _23990_);
  nand (_23993_, _23992_, _02537_);
  and (_23994_, _03057_, _22926_);
  nor (_23995_, _23994_, _02940_);
  nand (_23996_, _23995_, _23993_);
  and (_23997_, _09915_, _09263_);
  nor (_23999_, _23692_, _09915_);
  nor (_24000_, _23999_, _23997_);
  and (_24001_, _24000_, _02940_);
  nor (_24002_, _24001_, _09942_);
  nand (_24003_, _24002_, _23996_);
  nor (_24004_, _09941_, _02606_);
  nor (_24005_, _24004_, _03163_);
  and (_24006_, _24005_, _24003_);
  or (_24007_, _24006_, _23675_);
  nand (_24008_, _24007_, _09948_);
  nor (_24010_, _09948_, _02567_);
  nor (_24011_, _24010_, _04337_);
  nand (_24012_, _24011_, _24008_);
  and (_24013_, _04337_, _03057_);
  nor (_24014_, _24013_, _02497_);
  nand (_24015_, _24014_, _24012_);
  and (_24016_, _24000_, _02497_);
  nor (_24017_, _24016_, _09964_);
  nand (_24018_, _24017_, _24015_);
  and (_24019_, _09964_, _02567_);
  nor (_24021_, _24019_, _02888_);
  and (_24022_, _24021_, _24018_);
  or (_24023_, _24022_, _23674_);
  nand (_24024_, _24023_, _09044_);
  nor (_24025_, _09044_, _02567_);
  nor (_24026_, _24025_, _22655_);
  and (_24027_, _24026_, _24024_);
  nor (_24028_, _24027_, _23673_);
  or (_24029_, _24028_, _23671_);
  or (_24030_, _24029_, _42672_);
  or (_24032_, _42668_, \oc8051_golden_model_1.PC [3]);
  and (_24033_, _24032_, _43998_);
  and (_43498_, _24033_, _24030_);
  and (_24034_, _02230_, \oc8051_golden_model_1.PC [4]);
  nor (_24035_, _02230_, \oc8051_golden_model_1.PC [4]);
  nor (_24036_, _24035_, _24034_);
  and (_24037_, _24036_, _09979_);
  and (_24038_, _22655_, _05582_);
  or (_24039_, _24038_, _09979_);
  and (_24040_, _05582_, _04337_);
  and (_24042_, _06123_, _03145_);
  nor (_24043_, _09136_, _08165_);
  and (_24044_, _09157_, _09154_);
  nor (_24045_, _24044_, _09158_);
  and (_24046_, _24045_, _08165_);
  or (_24047_, _24046_, _24043_);
  and (_24048_, _24047_, _09672_);
  nor (_24049_, _09135_, _05753_);
  and (_24050_, _09136_, _02863_);
  nor (_24051_, _22940_, _09135_);
  not (_24053_, _24036_);
  and (_24054_, _24053_, _09489_);
  and (_24055_, _09136_, _02876_);
  nor (_24056_, _24036_, _09456_);
  and (_24057_, _05582_, _03818_);
  and (_24058_, _09136_, _03813_);
  or (_24059_, _24058_, _07636_);
  not (_24060_, \oc8051_golden_model_1.PC [4]);
  or (_24061_, _09429_, _24060_);
  and (_24062_, _24061_, _03814_);
  or (_24064_, _24062_, _24059_);
  or (_24065_, _24053_, _09430_);
  and (_24066_, _24065_, _02611_);
  and (_24067_, _24066_, _24064_);
  or (_24068_, _24067_, _14356_);
  or (_24069_, _24068_, _24057_);
  or (_24070_, _24053_, _09427_);
  and (_24071_, _24070_, _03387_);
  and (_24072_, _24071_, _24069_);
  and (_24073_, _09136_, _03072_);
  or (_24075_, _24073_, _24072_);
  nor (_24076_, _24075_, _07646_);
  and (_24077_, _24036_, _07646_);
  or (_24078_, _24077_, _24076_);
  and (_24079_, _24078_, _02616_);
  nor (_24080_, _05582_, _02616_);
  nor (_24081_, _24080_, _05363_);
  not (_24082_, _24081_);
  nor (_24083_, _24082_, _24079_);
  nand (_24084_, _09420_, _09135_);
  not (_24086_, _09420_);
  and (_24087_, _24045_, _24086_);
  nor (_24088_, _24087_, _05362_);
  and (_24089_, _24088_, _24084_);
  or (_24090_, _24089_, _24083_);
  and (_24091_, _24090_, _09449_);
  and (_24092_, _09286_, _09283_);
  nor (_24093_, _24092_, _09287_);
  not (_24094_, _24093_);
  nor (_24095_, _24094_, _09412_);
  not (_24097_, _24095_);
  nand (_24098_, _09257_, _09412_);
  and (_24099_, _24098_, _02974_);
  and (_24100_, _24099_, _24097_);
  or (_24101_, _24100_, _24091_);
  and (_24102_, _24101_, _09405_);
  or (_24103_, _24102_, _24056_);
  or (_24104_, _24103_, _02880_);
  nand (_24105_, _09135_, _02880_);
  and (_24106_, _24105_, _24104_);
  nor (_24108_, _24106_, _04252_);
  nor (_24109_, _05582_, _02609_);
  or (_24110_, _24109_, _03069_);
  nor (_24111_, _24110_, _24108_);
  and (_24112_, _09136_, _03069_);
  or (_24113_, _24112_, _24111_);
  and (_24114_, _24113_, _09463_);
  and (_24115_, _24053_, _09461_);
  or (_24116_, _24115_, _24114_);
  nand (_24117_, _24116_, _03084_);
  and (_24119_, _09136_, _03075_);
  nor (_24120_, _24119_, _09471_);
  nand (_24121_, _24120_, _24117_);
  nor (_24122_, _24053_, _09470_);
  nor (_24123_, _24122_, _02876_);
  and (_24124_, _24123_, _24121_);
  or (_24125_, _24124_, _24055_);
  nand (_24126_, _24125_, _02621_);
  and (_24127_, _05582_, _09474_);
  nor (_24128_, _24127_, _02875_);
  nand (_24130_, _24128_, _24126_);
  and (_24131_, _09135_, _02875_);
  nor (_24132_, _24131_, _09481_);
  and (_24133_, _24132_, _24130_);
  and (_24134_, _09392_, _09257_);
  nor (_24135_, _24094_, _09392_);
  or (_24136_, _24135_, _24134_);
  nor (_24137_, _24136_, _09396_);
  or (_24138_, _24137_, _24133_);
  nand (_24139_, _24138_, _02979_);
  nor (_24141_, _24094_, _09357_);
  and (_24142_, _09357_, _09257_);
  or (_24143_, _24142_, _24141_);
  or (_24144_, _24143_, _02979_);
  and (_24145_, _24144_, _09500_);
  nand (_24146_, _24145_, _24139_);
  nor (_24147_, _24093_, _09514_);
  and (_24148_, _09514_, _09258_);
  or (_24149_, _24148_, _09500_);
  or (_24150_, _24149_, _24147_);
  nand (_24152_, _24150_, _24146_);
  nand (_24153_, _24152_, _09531_);
  and (_24154_, _09528_, _09257_);
  and (_24155_, _24093_, _09529_);
  or (_24156_, _24155_, _24154_);
  and (_24157_, _24156_, _02952_);
  nor (_24158_, _24157_, _09489_);
  and (_24159_, _24158_, _24153_);
  or (_24160_, _24159_, _24054_);
  nand (_24161_, _24160_, _02870_);
  and (_24163_, _09136_, _02869_);
  nor (_24164_, _24163_, _04095_);
  nand (_24165_, _24164_, _24161_);
  nor (_24166_, _05582_, _02614_);
  nor (_24167_, _24166_, _23051_);
  and (_24168_, _24167_, _24165_);
  or (_24169_, _24168_, _24051_);
  nand (_24170_, _24169_, _09543_);
  nor (_24171_, _24036_, _09543_);
  nor (_24172_, _24171_, _03101_);
  nand (_24174_, _24172_, _24170_);
  and (_24175_, _09135_, _03101_);
  nor (_24176_, _24175_, _09551_);
  nand (_24177_, _24176_, _24174_);
  and (_24178_, _05582_, _09551_);
  nor (_24179_, _24178_, _03100_);
  and (_24180_, _24179_, _24177_);
  and (_24181_, _09135_, _03100_);
  or (_24182_, _24181_, _24180_);
  nand (_24183_, _24182_, _09557_);
  nor (_24185_, _24053_, _09557_);
  nor (_24186_, _24185_, _09562_);
  nand (_24187_, _24186_, _24183_);
  nor (_24188_, _09135_, _09561_);
  nor (_24189_, _24188_, _02583_);
  nand (_24190_, _24189_, _24187_);
  and (_24191_, _24036_, _02583_);
  nor (_24192_, _24191_, _02863_);
  and (_24193_, _24192_, _24190_);
  or (_24194_, _24193_, _24050_);
  nand (_24196_, _24194_, _04251_);
  and (_24197_, _05582_, _02581_);
  nor (_24198_, _24197_, _02981_);
  nand (_24199_, _24198_, _24196_);
  and (_24200_, _09257_, _02981_);
  nor (_24201_, _24200_, _09582_);
  and (_24202_, _24201_, _24199_);
  nor (_24203_, _09135_, _02857_);
  or (_24204_, _24203_, _02579_);
  nor (_24205_, _24204_, _24202_);
  and (_24207_, _09257_, _02579_);
  nor (_24208_, _24207_, _24205_);
  nand (_24209_, _24208_, _09200_);
  nor (_24210_, _24036_, _09200_);
  nor (_24211_, _24210_, _02933_);
  nand (_24212_, _24211_, _24209_);
  and (_24213_, _09135_, _02933_);
  nor (_24214_, _24213_, _02518_);
  nand (_24215_, _24214_, _24212_);
  and (_24216_, _05582_, _02518_);
  nor (_24218_, _24216_, _09594_);
  nand (_24219_, _24218_, _24215_);
  and (_24220_, _24045_, _09594_);
  nor (_24221_, _24220_, _05754_);
  and (_24222_, _24221_, _24219_);
  or (_24223_, _24222_, _24049_);
  nand (_24224_, _24223_, _02803_);
  and (_24225_, _09258_, _02802_);
  nor (_24226_, _24225_, _07859_);
  nand (_24227_, _24226_, _24224_);
  and (_24229_, _09135_, _07859_);
  nor (_24230_, _24229_, _09611_);
  nand (_24231_, _24230_, _24227_);
  and (_24232_, _09628_, _09625_);
  nor (_24233_, _24232_, _09629_);
  nor (_24234_, _24233_, _22679_);
  nor (_24235_, _24234_, _02932_);
  and (_24236_, _24235_, _24231_);
  and (_24237_, _09135_, _02932_);
  or (_24238_, _24237_, _02514_);
  or (_24240_, _24238_, _24236_);
  and (_24241_, _05582_, _02514_);
  nor (_24242_, _24241_, _09083_);
  and (_24243_, _24242_, _24240_);
  and (_24244_, _09135_, _08165_);
  and (_24245_, _24045_, _09676_);
  or (_24246_, _24245_, _24244_);
  and (_24247_, _24246_, _09083_);
  or (_24248_, _24247_, _24243_);
  nand (_24249_, _24248_, _09657_);
  nor (_24251_, _24053_, _09657_);
  nor (_24252_, _24251_, _09661_);
  nand (_24253_, _24252_, _24249_);
  nor (_24254_, _09660_, _09135_);
  nor (_24255_, _24254_, _02980_);
  and (_24256_, _24255_, _24253_);
  and (_24257_, _09257_, _02980_);
  or (_24258_, _24257_, _03127_);
  nor (_24259_, _24258_, _24256_);
  and (_24260_, _09136_, _03127_);
  or (_24262_, _24260_, _24259_);
  nand (_24263_, _24262_, _02510_);
  and (_24264_, _05582_, _02509_);
  nor (_24265_, _24264_, _09672_);
  and (_24266_, _24265_, _24263_);
  or (_24267_, _24266_, _24048_);
  nand (_24268_, _24267_, _09081_);
  nor (_24269_, _24053_, _09081_);
  nor (_24270_, _24269_, _22930_);
  nand (_24271_, _24270_, _24268_);
  nor (_24273_, _09135_, _09080_);
  nor (_24274_, _24273_, _02970_);
  nand (_24275_, _24274_, _24271_);
  and (_24276_, _09257_, _02970_);
  nor (_24277_, _24276_, _03135_);
  and (_24278_, _24277_, _24275_);
  and (_24279_, _09136_, _03135_);
  or (_24280_, _24279_, _24278_);
  nand (_24281_, _24280_, _02532_);
  and (_24282_, _05582_, _03880_);
  nor (_24284_, _24282_, _09076_);
  and (_24285_, _24284_, _24281_);
  and (_24286_, _09135_, \oc8051_golden_model_1.PSW [7]);
  and (_24287_, _24045_, _07293_);
  or (_24288_, _24287_, _24286_);
  and (_24289_, _24288_, _09076_);
  or (_24290_, _24289_, _24285_);
  nand (_24291_, _24290_, _09074_);
  nor (_24292_, _24053_, _09074_);
  nor (_24293_, _24292_, _07944_);
  nand (_24295_, _24293_, _24291_);
  nor (_24296_, _09135_, _07943_);
  nor (_24297_, _24296_, _02965_);
  and (_24298_, _24297_, _24295_);
  and (_24299_, _09257_, _02965_);
  or (_24300_, _24299_, _03123_);
  nor (_24301_, _24300_, _24298_);
  and (_24302_, _09136_, _03123_);
  or (_24303_, _24302_, _24301_);
  nand (_24304_, _24303_, _02535_);
  and (_24306_, _05582_, _09069_);
  nor (_24307_, _24306_, _09068_);
  nand (_24308_, _24307_, _24304_);
  nand (_24309_, _09135_, _07293_);
  nand (_24310_, _24045_, \oc8051_golden_model_1.PSW [7]);
  and (_24311_, _24310_, _24309_);
  or (_24312_, _24311_, _23200_);
  nand (_24313_, _24312_, _24308_);
  nand (_24314_, _24313_, _09066_);
  nor (_24315_, _24053_, _09066_);
  nor (_24318_, _24315_, _10365_);
  nand (_24319_, _24318_, _24314_);
  nor (_24320_, _09135_, _09065_);
  nor (_24321_, _24320_, _07991_);
  nand (_24322_, _24321_, _24319_);
  and (_24323_, _24036_, _07991_);
  nor (_24324_, _24323_, _03145_);
  and (_24325_, _24324_, _24322_);
  or (_24326_, _24325_, _24042_);
  nand (_24327_, _24326_, _02529_);
  and (_24330_, _05582_, _03898_);
  nor (_24331_, _24330_, _02968_);
  and (_24332_, _24331_, _24327_);
  nor (_24333_, _09915_, _09258_);
  and (_24334_, _24093_, _09915_);
  nor (_24335_, _24334_, _24333_);
  nor (_24336_, _24335_, _03561_);
  or (_24337_, _24336_, _24332_);
  nand (_24338_, _24337_, _09063_);
  nor (_24339_, _24053_, _09063_);
  nor (_24342_, _24339_, _08067_);
  nand (_24343_, _24342_, _24338_);
  nor (_24344_, _09135_, _08066_);
  nor (_24345_, _24344_, _08111_);
  nand (_24346_, _24345_, _24343_);
  and (_24347_, _24036_, _08111_);
  nor (_24348_, _24347_, _02892_);
  nand (_24349_, _24348_, _24346_);
  and (_24350_, _06123_, _02892_);
  nor (_24351_, _24350_, _22926_);
  and (_24354_, _24351_, _24349_);
  nor (_24355_, _05582_, _02537_);
  or (_24356_, _24355_, _02940_);
  or (_24357_, _24356_, _24354_);
  and (_24358_, _09915_, _09258_);
  nor (_24359_, _24093_, _09915_);
  nor (_24360_, _24359_, _24358_);
  nor (_24361_, _24360_, _03164_);
  nor (_24362_, _24361_, _09942_);
  nand (_24363_, _24362_, _24357_);
  nor (_24366_, _24053_, _09941_);
  nor (_24367_, _24366_, _03163_);
  nand (_24368_, _24367_, _24363_);
  and (_24369_, _09136_, _03163_);
  nor (_24370_, _24369_, _09949_);
  nand (_24371_, _24370_, _24368_);
  nor (_24372_, _24053_, _09948_);
  nor (_24373_, _24372_, _04337_);
  and (_24374_, _24373_, _24371_);
  or (_24375_, _24374_, _24040_);
  nand (_24378_, _24375_, _02498_);
  nor (_24379_, _24360_, _02498_);
  nor (_24380_, _24379_, _09964_);
  nand (_24381_, _24380_, _24378_);
  and (_24382_, _24036_, _09964_);
  nor (_24383_, _24382_, _02888_);
  nand (_24384_, _24383_, _24381_);
  and (_24385_, _09136_, _02888_);
  nor (_24386_, _24385_, _09970_);
  nand (_24387_, _24386_, _24384_);
  nor (_24390_, _24053_, _09044_);
  nor (_24391_, _24390_, _22655_);
  and (_24392_, _24391_, _24387_);
  nor (_24393_, _24392_, _24039_);
  or (_24394_, _24393_, _24037_);
  or (_24395_, _24394_, _42672_);
  or (_24396_, _42668_, \oc8051_golden_model_1.PC [4]);
  and (_24397_, _24396_, _43998_);
  and (_43499_, _24397_, _24395_);
  nor (_24398_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_24400_, _09130_, _02244_);
  nor (_24401_, _24400_, _24398_);
  and (_24402_, _24401_, _09979_);
  and (_24403_, _22655_, _05613_);
  or (_24404_, _24403_, _09979_);
  and (_24405_, _09130_, _02888_);
  nand (_24406_, _09130_, _03163_);
  nor (_24407_, _24401_, _09063_);
  nor (_24408_, _24401_, _09066_);
  nor (_24409_, _24401_, _09074_);
  nor (_24411_, _24401_, _09081_);
  nor (_24412_, _24401_, _09657_);
  nor (_24413_, _09130_, _05753_);
  and (_24414_, _09131_, _02863_);
  nor (_24415_, _22940_, _09130_);
  not (_24416_, _24401_);
  and (_24417_, _24416_, _09489_);
  nand (_24418_, _09252_, _09412_);
  or (_24419_, _09255_, _09254_);
  and (_24420_, _24419_, _09288_);
  nor (_24422_, _24419_, _09288_);
  or (_24423_, _24422_, _24420_);
  or (_24424_, _24423_, _09412_);
  and (_24425_, _24424_, _24418_);
  and (_24426_, _24425_, _02974_);
  or (_24427_, _09133_, _09132_);
  and (_24428_, _24427_, _09159_);
  nor (_24429_, _24427_, _09159_);
  or (_24430_, _24429_, _24428_);
  or (_24431_, _24430_, _09420_);
  nand (_24433_, _09420_, _09130_);
  and (_24434_, _24433_, _24431_);
  and (_24435_, _24434_, _05363_);
  or (_24436_, _05613_, _02611_);
  nor (_24437_, _09429_, \oc8051_golden_model_1.PC [5]);
  or (_24438_, _24437_, _03813_);
  nand (_24439_, _09130_, _03813_);
  and (_24440_, _24439_, _23337_);
  and (_24441_, _24440_, _24438_);
  nor (_24442_, _24401_, _09430_);
  or (_24444_, _24442_, _03818_);
  or (_24445_, _24444_, _24441_);
  and (_24446_, _24445_, _09427_);
  and (_24447_, _24446_, _24436_);
  nor (_24448_, _24401_, _09427_);
  or (_24449_, _24448_, _03072_);
  or (_24450_, _24449_, _24447_);
  nand (_24451_, _09130_, _03072_);
  and (_24452_, _24451_, _09426_);
  and (_24453_, _24452_, _24450_);
  and (_24455_, _24416_, _07646_);
  or (_24456_, _24455_, _09425_);
  or (_24457_, _24456_, _24453_);
  or (_24458_, _05613_, _02616_);
  and (_24459_, _24458_, _05362_);
  and (_24460_, _24459_, _24457_);
  or (_24461_, _24460_, _02886_);
  or (_24462_, _24461_, _24435_);
  nand (_24463_, _24401_, _02886_);
  and (_24464_, _24463_, _03810_);
  and (_24466_, _24464_, _24462_);
  or (_24467_, _24466_, _24426_);
  and (_24468_, _24467_, _09405_);
  nor (_24469_, _24401_, _09405_);
  or (_24470_, _24469_, _02880_);
  or (_24471_, _24470_, _24468_);
  nand (_24472_, _09130_, _02880_);
  and (_24473_, _24472_, _02609_);
  and (_24474_, _24473_, _24471_);
  and (_24475_, _05613_, _04252_);
  or (_24477_, _24475_, _03069_);
  or (_24478_, _24477_, _24474_);
  and (_24479_, _09130_, _03069_);
  nor (_24480_, _24479_, _09461_);
  and (_24481_, _24480_, _24478_);
  and (_24482_, _24416_, _09461_);
  or (_24483_, _24482_, _03075_);
  or (_24484_, _24483_, _24481_);
  nand (_24485_, _09130_, _03075_);
  and (_24486_, _24485_, _09470_);
  and (_24488_, _24486_, _24484_);
  nor (_24489_, _24401_, _09470_);
  or (_24490_, _24489_, _02876_);
  or (_24491_, _24490_, _24488_);
  nand (_24492_, _09130_, _02876_);
  and (_24493_, _24492_, _02621_);
  and (_24494_, _24493_, _24491_);
  and (_24495_, _05613_, _09474_);
  or (_24496_, _24495_, _02875_);
  or (_24497_, _24496_, _24494_);
  nand (_24499_, _09130_, _02875_);
  and (_24500_, _24499_, _09396_);
  and (_24501_, _24500_, _24497_);
  nand (_24502_, _09392_, _09252_);
  or (_24503_, _24423_, _09392_);
  and (_24504_, _24503_, _24502_);
  and (_24505_, _24504_, _09481_);
  or (_24506_, _24505_, _02978_);
  or (_24507_, _24506_, _24501_);
  and (_24508_, _24423_, _23025_);
  and (_24510_, _09357_, _09253_);
  or (_24511_, _24510_, _02979_);
  or (_24512_, _24511_, _24508_);
  and (_24513_, _24512_, _09500_);
  and (_24514_, _24513_, _24507_);
  or (_24515_, _24423_, _09514_);
  nand (_24516_, _09514_, _09252_);
  and (_24517_, _24516_, _02950_);
  and (_24518_, _24517_, _24515_);
  or (_24519_, _24518_, _02952_);
  or (_24521_, _24519_, _24514_);
  and (_24522_, _24423_, _09529_);
  and (_24523_, _09528_, _09253_);
  or (_24524_, _24523_, _09531_);
  or (_24525_, _24524_, _24522_);
  and (_24526_, _24525_, _09490_);
  and (_24527_, _24526_, _24521_);
  or (_24528_, _24527_, _24417_);
  and (_24529_, _24528_, _02870_);
  and (_24530_, _09131_, _02869_);
  or (_24532_, _24530_, _04095_);
  or (_24533_, _24532_, _24529_);
  or (_24534_, _05613_, _02614_);
  and (_24535_, _24534_, _22940_);
  and (_24536_, _24535_, _24533_);
  or (_24537_, _24536_, _24415_);
  and (_24538_, _24537_, _09543_);
  nor (_24539_, _24401_, _09543_);
  or (_24540_, _24539_, _03101_);
  or (_24541_, _24540_, _24538_);
  nand (_24543_, _09130_, _03101_);
  and (_24544_, _24543_, _02619_);
  and (_24545_, _24544_, _24541_);
  and (_24546_, _05613_, _09551_);
  or (_24547_, _24546_, _03100_);
  or (_24548_, _24547_, _24545_);
  nand (_24549_, _09130_, _03100_);
  and (_24550_, _24549_, _09557_);
  and (_24551_, _24550_, _24548_);
  nor (_24552_, _24401_, _09557_);
  or (_24554_, _24552_, _24551_);
  and (_24555_, _24554_, _09561_);
  nor (_24556_, _09130_, _09561_);
  or (_24557_, _24556_, _02583_);
  or (_24558_, _24557_, _24555_);
  nand (_24559_, _24401_, _02583_);
  and (_24560_, _24559_, _02864_);
  and (_24561_, _24560_, _24558_);
  or (_24562_, _24561_, _24414_);
  and (_24563_, _24562_, _04251_);
  and (_24565_, _05613_, _02581_);
  or (_24566_, _24565_, _02981_);
  or (_24567_, _24566_, _24563_);
  nand (_24568_, _09252_, _02981_);
  and (_24569_, _24568_, _02857_);
  and (_24570_, _24569_, _24567_);
  nor (_24571_, _09130_, _02857_);
  or (_24572_, _24571_, _02579_);
  or (_24573_, _24572_, _24570_);
  nand (_24574_, _09252_, _02579_);
  and (_24576_, _24574_, _09200_);
  and (_24577_, _24576_, _24573_);
  nor (_24578_, _24401_, _09200_);
  or (_24579_, _24578_, _02933_);
  or (_24580_, _24579_, _24577_);
  nand (_24581_, _09130_, _02933_);
  and (_24582_, _24581_, _22795_);
  and (_24583_, _24582_, _24580_);
  and (_24584_, _05613_, _02518_);
  or (_24585_, _24584_, _09594_);
  or (_24587_, _24585_, _24583_);
  or (_24588_, _24430_, _09599_);
  and (_24589_, _24588_, _05753_);
  and (_24590_, _24589_, _24587_);
  or (_24591_, _24590_, _24413_);
  and (_24592_, _24591_, _02803_);
  and (_24593_, _09253_, _02802_);
  or (_24594_, _24593_, _07859_);
  or (_24595_, _24594_, _24592_);
  nand (_24596_, _09130_, _07859_);
  and (_24598_, _24596_, _22679_);
  and (_24599_, _24598_, _24595_);
  and (_24600_, _09630_, _09623_);
  or (_24601_, _24600_, _09631_);
  and (_24602_, _24601_, _09611_);
  or (_24603_, _24602_, _02932_);
  or (_24604_, _24603_, _24599_);
  nand (_24605_, _09130_, _02932_);
  and (_24606_, _24605_, _04093_);
  and (_24607_, _24606_, _24604_);
  and (_24609_, _05613_, _02514_);
  or (_24610_, _24609_, _09083_);
  or (_24611_, _24610_, _24607_);
  and (_24612_, _24430_, _09676_);
  or (_24613_, _09130_, _09676_);
  nand (_24614_, _24613_, _09083_);
  or (_24615_, _24614_, _24612_);
  and (_24616_, _24615_, _09657_);
  and (_24617_, _24616_, _24611_);
  or (_24618_, _24617_, _24412_);
  and (_24620_, _24618_, _09660_);
  nor (_24621_, _09660_, _09130_);
  or (_24622_, _24621_, _02980_);
  or (_24623_, _24622_, _24620_);
  nand (_24624_, _09252_, _02980_);
  and (_24625_, _24624_, _03128_);
  and (_24626_, _24625_, _24623_);
  and (_24627_, _09131_, _03127_);
  or (_24628_, _24627_, _24626_);
  and (_24629_, _24628_, _02510_);
  and (_24631_, _05613_, _02509_);
  or (_24632_, _24631_, _09672_);
  or (_24633_, _24632_, _24629_);
  and (_24634_, _24430_, _08165_);
  or (_24635_, _09130_, _08165_);
  nand (_24636_, _24635_, _09672_);
  or (_24637_, _24636_, _24634_);
  and (_24638_, _24637_, _09081_);
  and (_24639_, _24638_, _24633_);
  or (_24640_, _24639_, _24411_);
  and (_24642_, _24640_, _09080_);
  nor (_24643_, _09130_, _09080_);
  or (_24644_, _24643_, _02970_);
  or (_24645_, _24644_, _24642_);
  nand (_24646_, _09252_, _02970_);
  and (_24647_, _24646_, _03137_);
  and (_24648_, _24647_, _24645_);
  and (_24649_, _09131_, _03135_);
  or (_24650_, _24649_, _24648_);
  and (_24651_, _24650_, _02532_);
  and (_24653_, _05613_, _03880_);
  or (_24654_, _24653_, _09076_);
  or (_24655_, _24654_, _24651_);
  and (_24656_, _24430_, _07293_);
  or (_24657_, _09130_, _07293_);
  nand (_24658_, _24657_, _09076_);
  or (_24659_, _24658_, _24656_);
  and (_24660_, _24659_, _09074_);
  and (_24661_, _24660_, _24655_);
  or (_24662_, _24661_, _24409_);
  and (_24664_, _24662_, _07943_);
  nor (_24665_, _09130_, _07943_);
  or (_24666_, _24665_, _02965_);
  or (_24667_, _24666_, _24664_);
  nand (_24668_, _09252_, _02965_);
  and (_24669_, _24668_, _05788_);
  and (_24670_, _24669_, _24667_);
  and (_24671_, _09131_, _03123_);
  or (_24672_, _24671_, _24670_);
  and (_24673_, _24672_, _02535_);
  and (_24675_, _05613_, _09069_);
  or (_24676_, _24675_, _09068_);
  or (_24677_, _24676_, _24673_);
  and (_24678_, _24430_, \oc8051_golden_model_1.PSW [7]);
  or (_24679_, _09130_, \oc8051_golden_model_1.PSW [7]);
  nand (_24680_, _24679_, _09068_);
  or (_24681_, _24680_, _24678_);
  and (_24682_, _24681_, _09066_);
  and (_24683_, _24682_, _24677_);
  or (_24684_, _24683_, _24408_);
  and (_24686_, _24684_, _09065_);
  nor (_24687_, _09130_, _09065_);
  or (_24688_, _24687_, _07991_);
  or (_24689_, _24688_, _24686_);
  nand (_24690_, _24401_, _07991_);
  and (_24691_, _24690_, _09726_);
  and (_24692_, _24691_, _24689_);
  and (_24693_, _06078_, _03145_);
  or (_24694_, _24693_, _24692_);
  and (_24695_, _24694_, _02529_);
  and (_24697_, _05613_, _03898_);
  or (_24698_, _24697_, _02968_);
  or (_24699_, _24698_, _24695_);
  and (_24700_, _24423_, _09915_);
  nor (_24701_, _09915_, _09252_);
  or (_24702_, _24701_, _03561_);
  or (_24703_, _24702_, _24700_);
  and (_24704_, _24703_, _09063_);
  and (_24705_, _24704_, _24699_);
  or (_24706_, _24705_, _24407_);
  and (_24708_, _24706_, _08066_);
  nor (_24709_, _09130_, _08066_);
  or (_24710_, _24709_, _08111_);
  or (_24711_, _24710_, _24708_);
  nand (_24712_, _24401_, _08111_);
  and (_24713_, _24712_, _02893_);
  and (_24714_, _24713_, _24711_);
  and (_24715_, _06078_, _02892_);
  or (_24716_, _24715_, _24714_);
  and (_24717_, _24716_, _02537_);
  and (_24719_, _05613_, _22926_);
  or (_24720_, _24719_, _02940_);
  or (_24721_, _24720_, _24717_);
  and (_24722_, _09915_, _09252_);
  nor (_24723_, _24423_, _09915_);
  or (_24724_, _24723_, _24722_);
  nand (_24725_, _24724_, _02940_);
  and (_24726_, _24725_, _09941_);
  and (_24727_, _24726_, _24721_);
  nor (_24728_, _24401_, _09941_);
  or (_24730_, _24728_, _03163_);
  or (_24731_, _24730_, _24727_);
  and (_24732_, _24731_, _24406_);
  nor (_24733_, _24732_, _09949_);
  nor (_24734_, _24416_, _09948_);
  nor (_24735_, _24734_, _04337_);
  not (_24736_, _24735_);
  nor (_24737_, _24736_, _24733_);
  and (_24738_, _05613_, _04337_);
  nor (_24739_, _24738_, _02497_);
  not (_24741_, _24739_);
  nor (_24742_, _24741_, _24737_);
  and (_24743_, _24724_, _02497_);
  nor (_24744_, _24743_, _09964_);
  not (_24745_, _24744_);
  nor (_24746_, _24745_, _24742_);
  and (_24747_, _24416_, _09964_);
  nor (_24748_, _24747_, _02888_);
  not (_24749_, _24748_);
  nor (_24750_, _24749_, _24746_);
  nor (_24753_, _24750_, _24405_);
  nor (_24754_, _24753_, _09970_);
  nor (_24755_, _24416_, _09044_);
  nor (_24756_, _24755_, _22655_);
  not (_24757_, _24756_);
  nor (_24758_, _24757_, _24754_);
  nor (_24759_, _24758_, _24404_);
  nor (_24760_, _24759_, _24402_);
  nand (_24761_, _24760_, _42668_);
  or (_24762_, _42668_, \oc8051_golden_model_1.PC [5]);
  and (_24764_, _24762_, _43998_);
  and (_43500_, _24764_, _24761_);
  and (_24765_, _05253_, _02230_);
  nor (_24766_, _24765_, \oc8051_golden_model_1.PC [6]);
  nor (_24767_, _24766_, _09045_);
  and (_24768_, _24767_, _09979_);
  nand (_24769_, _05649_, _04337_);
  not (_24770_, _24767_);
  nand (_24771_, _24770_, _08111_);
  nand (_24772_, _09246_, _02965_);
  nand (_24774_, _09246_, _02970_);
  nand (_24775_, _09246_, _02980_);
  nand (_24776_, _09124_, _02932_);
  nand (_24777_, _24770_, _02583_);
  or (_24778_, _22940_, _09123_);
  nand (_24779_, _24770_, _09489_);
  nor (_24780_, _09291_, _09249_);
  nor (_24781_, _24780_, _09292_);
  or (_24782_, _24781_, _09392_);
  nand (_24783_, _09392_, _09246_);
  and (_24785_, _24783_, _24782_);
  or (_24786_, _24785_, _09396_);
  or (_24787_, _24767_, _09456_);
  and (_24788_, _05649_, _03818_);
  and (_24789_, _09124_, _03813_);
  or (_24790_, _24789_, _07636_);
  not (_24791_, \oc8051_golden_model_1.PC [6]);
  or (_24792_, _09429_, _24791_);
  and (_24793_, _24792_, _03814_);
  or (_24794_, _24793_, _24790_);
  or (_24796_, _24770_, _09430_);
  and (_24797_, _24796_, _02611_);
  and (_24798_, _24797_, _24794_);
  or (_24799_, _24798_, _14356_);
  or (_24800_, _24799_, _24788_);
  or (_24801_, _24770_, _09427_);
  and (_24802_, _24801_, _03387_);
  and (_24803_, _24802_, _24800_);
  and (_24804_, _09124_, _03072_);
  or (_24805_, _24804_, _24803_);
  nand (_24807_, _24805_, _09426_);
  nand (_24808_, _24770_, _07646_);
  and (_24809_, _24808_, _02616_);
  and (_24810_, _24809_, _24807_);
  nor (_24811_, _05649_, _02616_);
  or (_24812_, _24811_, _05363_);
  or (_24813_, _24812_, _24810_);
  nor (_24814_, _09162_, _09127_);
  nor (_24815_, _24814_, _09163_);
  and (_24816_, _24815_, _24086_);
  and (_24818_, _09420_, _09123_);
  or (_24819_, _24818_, _05362_);
  or (_24820_, _24819_, _24816_);
  nand (_24821_, _24820_, _24813_);
  nand (_24822_, _24821_, _09449_);
  not (_24823_, _09412_);
  and (_24824_, _24781_, _24823_);
  and (_24825_, _09245_, _09412_);
  or (_24826_, _24825_, _03810_);
  or (_24827_, _24826_, _24824_);
  and (_24829_, _24827_, _24822_);
  or (_24830_, _24829_, _09406_);
  and (_24831_, _24830_, _24787_);
  or (_24832_, _24831_, _02880_);
  nand (_24833_, _09124_, _02880_);
  and (_24834_, _24833_, _02609_);
  and (_24835_, _24834_, _24832_);
  nor (_24836_, _05649_, _02609_);
  or (_24837_, _24836_, _03069_);
  or (_24838_, _24837_, _24835_);
  nand (_24840_, _09124_, _03069_);
  and (_24841_, _24840_, _24838_);
  and (_24842_, _24841_, _09463_);
  and (_24843_, _24767_, _09461_);
  or (_24844_, _24843_, _03075_);
  or (_24845_, _24844_, _24842_);
  nand (_24846_, _09124_, _03075_);
  and (_24847_, _24846_, _09470_);
  and (_24848_, _24847_, _24845_);
  nor (_24849_, _24770_, _09470_);
  or (_24851_, _24849_, _02876_);
  or (_24852_, _24851_, _24848_);
  nand (_24853_, _09124_, _02876_);
  and (_24854_, _24853_, _24852_);
  or (_24855_, _24854_, _09474_);
  nand (_24856_, _05649_, _09474_);
  and (_24857_, _24856_, _03941_);
  and (_24858_, _24857_, _24855_);
  nand (_24859_, _09123_, _02875_);
  nand (_24860_, _24859_, _09396_);
  or (_24862_, _24860_, _24858_);
  and (_24863_, _24862_, _24786_);
  or (_24864_, _24863_, _02978_);
  and (_24865_, _09357_, _09245_);
  and (_24866_, _24781_, _23025_);
  or (_24867_, _24866_, _02979_);
  or (_24868_, _24867_, _24865_);
  and (_24869_, _24868_, _24864_);
  or (_24870_, _24869_, _02950_);
  and (_24871_, _24781_, _23031_);
  and (_24873_, _09514_, _09245_);
  or (_24874_, _24873_, _09500_);
  or (_24875_, _24874_, _24871_);
  and (_24876_, _24875_, _09531_);
  and (_24877_, _24876_, _24870_);
  or (_24878_, _24781_, _09528_);
  nand (_24879_, _09528_, _09246_);
  and (_24880_, _24879_, _02952_);
  and (_24881_, _24880_, _24878_);
  or (_24882_, _24881_, _09489_);
  or (_24884_, _24882_, _24877_);
  and (_24885_, _24884_, _24779_);
  or (_24886_, _24885_, _02869_);
  nand (_24887_, _09124_, _02869_);
  and (_24888_, _24887_, _02614_);
  and (_24889_, _24888_, _24886_);
  nor (_24890_, _05649_, _02614_);
  or (_24891_, _24890_, _23051_);
  or (_24892_, _24891_, _24889_);
  and (_24893_, _24892_, _24778_);
  or (_24895_, _24893_, _09544_);
  or (_24896_, _24767_, _09543_);
  and (_24897_, _24896_, _09550_);
  and (_24898_, _24897_, _24895_);
  and (_24899_, _09123_, _03101_);
  or (_24900_, _24899_, _09551_);
  or (_24901_, _24900_, _24898_);
  nand (_24902_, _05649_, _09551_);
  and (_24903_, _24902_, _10016_);
  and (_24904_, _24903_, _24901_);
  nand (_24906_, _09123_, _03100_);
  nand (_24907_, _24906_, _09557_);
  or (_24908_, _24907_, _24904_);
  or (_24909_, _24767_, _09557_);
  and (_24910_, _24909_, _09561_);
  and (_24911_, _24910_, _24908_);
  nor (_24912_, _09124_, _09561_);
  or (_24913_, _24912_, _02583_);
  or (_24914_, _24913_, _24911_);
  and (_24915_, _24914_, _24777_);
  or (_24917_, _24915_, _02863_);
  nand (_24918_, _09124_, _02863_);
  and (_24919_, _24918_, _04251_);
  and (_24920_, _24919_, _24917_);
  nor (_24921_, _05649_, _04251_);
  or (_24922_, _24921_, _02981_);
  or (_24923_, _24922_, _24920_);
  nand (_24924_, _09246_, _02981_);
  and (_24925_, _24924_, _24923_);
  or (_24926_, _24925_, _09582_);
  or (_24928_, _09123_, _02857_);
  and (_24929_, _24928_, _24926_);
  or (_24930_, _24929_, _02579_);
  nand (_24931_, _09246_, _02579_);
  and (_24932_, _24931_, _09200_);
  and (_24933_, _24932_, _24930_);
  nor (_24934_, _24770_, _09200_);
  or (_24935_, _24934_, _02933_);
  or (_24936_, _24935_, _24933_);
  nand (_24937_, _09124_, _02933_);
  and (_24939_, _24937_, _22795_);
  and (_24940_, _24939_, _24936_);
  nor (_24941_, _05649_, _22795_);
  or (_24942_, _24941_, _24940_);
  and (_24943_, _24942_, _09599_);
  and (_24944_, _24815_, _09594_);
  or (_24945_, _24944_, _24943_);
  and (_24946_, _24945_, _05753_);
  nor (_24947_, _09124_, _05753_);
  or (_24948_, _24947_, _02802_);
  or (_24950_, _24948_, _24946_);
  nand (_24951_, _09246_, _02802_);
  and (_24952_, _24951_, _07860_);
  and (_24953_, _24952_, _24950_);
  and (_24954_, _09123_, _07859_);
  or (_24955_, _24954_, _09611_);
  or (_24956_, _24955_, _24953_);
  nor (_24957_, _09633_, _09619_);
  nor (_24958_, _24957_, _09634_);
  or (_24959_, _24958_, _22679_);
  and (_24961_, _24959_, _24956_);
  or (_24962_, _24961_, _02932_);
  and (_24963_, _24962_, _24776_);
  or (_24964_, _24963_, _02514_);
  nand (_24965_, _05649_, _02514_);
  and (_24966_, _24965_, _22678_);
  and (_24967_, _24966_, _24964_);
  or (_24968_, _24815_, _08165_);
  or (_24969_, _09123_, _09676_);
  and (_24970_, _24969_, _09083_);
  and (_24972_, _24970_, _24968_);
  or (_24973_, _24972_, _23884_);
  or (_24974_, _24973_, _24967_);
  or (_24975_, _24767_, _09657_);
  and (_24976_, _24975_, _09660_);
  and (_24977_, _24976_, _24974_);
  nor (_24978_, _09660_, _09124_);
  or (_24979_, _24978_, _02980_);
  or (_24980_, _24979_, _24977_);
  and (_24981_, _24980_, _24775_);
  or (_24983_, _24981_, _03127_);
  nand (_24984_, _09124_, _03127_);
  and (_24985_, _24984_, _02510_);
  and (_24986_, _24985_, _24983_);
  nor (_24987_, _05649_, _02510_);
  or (_24988_, _24987_, _24986_);
  and (_24989_, _24988_, _22675_);
  or (_24990_, _24815_, _09676_);
  or (_24991_, _09123_, _08165_);
  and (_24992_, _24991_, _09672_);
  and (_24994_, _24992_, _24990_);
  or (_24995_, _24994_, _09681_);
  or (_24996_, _24995_, _24989_);
  or (_24997_, _24767_, _09081_);
  and (_24998_, _24997_, _09080_);
  and (_24999_, _24998_, _24996_);
  nor (_25000_, _09124_, _09080_);
  or (_25001_, _25000_, _02970_);
  or (_25002_, _25001_, _24999_);
  and (_25003_, _25002_, _24774_);
  or (_25005_, _25003_, _03135_);
  nand (_25006_, _09124_, _03135_);
  and (_25007_, _25006_, _02532_);
  and (_25008_, _25007_, _25005_);
  nor (_25009_, _05649_, _02532_);
  or (_25010_, _25009_, _25008_);
  and (_25011_, _25010_, _22667_);
  or (_25012_, _24815_, \oc8051_golden_model_1.PSW [7]);
  or (_25013_, _09123_, _07293_);
  and (_25014_, _25013_, _09076_);
  and (_25016_, _25014_, _25012_);
  or (_25017_, _25016_, _09694_);
  or (_25018_, _25017_, _25011_);
  or (_25019_, _24767_, _09074_);
  and (_25020_, _25019_, _07943_);
  and (_25021_, _25020_, _25018_);
  nor (_25022_, _09124_, _07943_);
  or (_25023_, _25022_, _02965_);
  or (_25024_, _25023_, _25021_);
  and (_25025_, _25024_, _24772_);
  or (_25027_, _25025_, _03123_);
  nand (_25028_, _09124_, _03123_);
  and (_25029_, _25028_, _02535_);
  and (_25030_, _25029_, _25027_);
  nor (_25031_, _05649_, _02535_);
  or (_25032_, _25031_, _25030_);
  and (_25033_, _25032_, _23200_);
  or (_25034_, _24815_, _07293_);
  or (_25035_, _09123_, \oc8051_golden_model_1.PSW [7]);
  and (_25036_, _25035_, _09068_);
  and (_25038_, _25036_, _25034_);
  or (_25039_, _25038_, _09711_);
  or (_25040_, _25039_, _25033_);
  or (_25041_, _24767_, _09066_);
  and (_25042_, _25041_, _09065_);
  and (_25043_, _25042_, _25040_);
  nor (_25044_, _09124_, _09065_);
  or (_25045_, _25044_, _07991_);
  or (_25046_, _25045_, _25043_);
  nand (_25047_, _24770_, _07991_);
  and (_25049_, _25047_, _09726_);
  and (_25050_, _25049_, _25046_);
  and (_25051_, _05849_, _03145_);
  or (_25052_, _25051_, _03898_);
  or (_25053_, _25052_, _25050_);
  nand (_25054_, _05649_, _03898_);
  and (_25055_, _25054_, _03561_);
  and (_25056_, _25055_, _25053_);
  not (_25057_, _09063_);
  or (_25058_, _09915_, _09245_);
  or (_25060_, _24781_, _23226_);
  and (_25061_, _25060_, _02968_);
  and (_25062_, _25061_, _25058_);
  or (_25063_, _25062_, _25057_);
  or (_25064_, _25063_, _25056_);
  or (_25065_, _24767_, _09063_);
  and (_25066_, _25065_, _08066_);
  and (_25067_, _25066_, _25064_);
  nor (_25068_, _09124_, _08066_);
  or (_25069_, _25068_, _08111_);
  or (_25071_, _25069_, _25067_);
  and (_25072_, _25071_, _24771_);
  or (_25073_, _25072_, _02892_);
  or (_25074_, _05849_, _02893_);
  and (_25075_, _25074_, _02537_);
  and (_25076_, _25075_, _25073_);
  nor (_25077_, _05649_, _02537_);
  or (_25078_, _25077_, _02940_);
  or (_25079_, _25078_, _25076_);
  nand (_25080_, _09915_, _09246_);
  or (_25082_, _24781_, _09915_);
  and (_25083_, _25082_, _25080_);
  or (_25084_, _25083_, _03164_);
  and (_25085_, _25084_, _25079_);
  or (_25086_, _25085_, _09942_);
  or (_25087_, _24767_, _09941_);
  and (_25088_, _25087_, _25086_);
  or (_25089_, _25088_, _03163_);
  nand (_25090_, _09124_, _03163_);
  and (_25091_, _25090_, _09948_);
  and (_25093_, _25091_, _25089_);
  nor (_25094_, _24770_, _09948_);
  or (_25095_, _25094_, _04337_);
  or (_25096_, _25095_, _25093_);
  and (_25097_, _25096_, _24769_);
  or (_25098_, _25097_, _02497_);
  not (_25099_, _09964_);
  or (_25100_, _25083_, _02498_);
  and (_25101_, _25100_, _25099_);
  and (_25102_, _25101_, _25098_);
  and (_25104_, _24767_, _09964_);
  or (_25105_, _25104_, _02888_);
  or (_25106_, _25105_, _25102_);
  nand (_25107_, _09124_, _02888_);
  and (_25108_, _25107_, _09044_);
  and (_25109_, _25108_, _25106_);
  nor (_25110_, _24770_, _09044_);
  or (_25111_, _25110_, _22655_);
  or (_25112_, _25111_, _25109_);
  nand (_25113_, _22655_, _05649_);
  and (_25115_, _25113_, _09983_);
  and (_25116_, _25115_, _25112_);
  or (_25117_, _25116_, _24768_);
  or (_25118_, _25117_, _42672_);
  or (_25119_, _42668_, \oc8051_golden_model_1.PC [6]);
  and (_25120_, _25119_, _43998_);
  and (_43501_, _25120_, _25118_);
  nor (_25121_, _09045_, \oc8051_golden_model_1.PC [7]);
  nor (_25122_, _25121_, _09046_);
  and (_25123_, _25122_, _09979_);
  and (_25125_, _05368_, _02888_);
  or (_25126_, _25122_, _09948_);
  or (_25127_, _25122_, _09063_);
  or (_25128_, _25122_, _09066_);
  or (_25129_, _25122_, _09074_);
  or (_25130_, _25122_, _09081_);
  or (_25131_, _25122_, _09657_);
  or (_25132_, _05753_, _05368_);
  nand (_25133_, _05369_, _02863_);
  or (_25134_, _22940_, _05368_);
  not (_25136_, _25122_);
  nand (_25137_, _25136_, _09489_);
  nand (_25138_, _09412_, _05260_);
  or (_25139_, _09241_, _09242_);
  nand (_25140_, _25139_, _09293_);
  or (_25141_, _25139_, _09293_);
  and (_25142_, _25141_, _25140_);
  or (_25143_, _25142_, _09412_);
  and (_25144_, _25143_, _25138_);
  or (_25145_, _25144_, _03810_);
  or (_25147_, _09119_, _09120_);
  nand (_25148_, _25147_, _09164_);
  or (_25149_, _25147_, _09164_);
  and (_25150_, _25149_, _25148_);
  or (_25151_, _25150_, _09420_);
  nand (_25152_, _09420_, _05369_);
  and (_25153_, _25152_, _25151_);
  or (_25154_, _25153_, _05362_);
  nor (_25155_, _05311_, _02611_);
  or (_25156_, _09429_, \oc8051_golden_model_1.PC [7]);
  and (_25158_, _25156_, _03814_);
  and (_25159_, _05368_, _03813_);
  or (_25160_, _25159_, _07636_);
  or (_25161_, _25160_, _25158_);
  or (_25162_, _25122_, _09430_);
  and (_25163_, _25162_, _02611_);
  and (_25164_, _25163_, _25161_);
  or (_25165_, _25164_, _14356_);
  or (_25166_, _25165_, _25155_);
  or (_25167_, _25122_, _09427_);
  and (_25169_, _25167_, _03387_);
  and (_25170_, _25169_, _25166_);
  and (_25171_, _05368_, _03072_);
  or (_25172_, _25171_, _07646_);
  or (_25173_, _25172_, _25170_);
  nand (_25174_, _25136_, _07646_);
  and (_25175_, _25174_, _02616_);
  and (_25176_, _25175_, _25173_);
  nor (_25177_, _05311_, _02616_);
  or (_25178_, _25177_, _05363_);
  or (_25180_, _25178_, _25176_);
  and (_25181_, _25180_, _04265_);
  and (_25182_, _25181_, _25154_);
  and (_25183_, _25122_, _02886_);
  or (_25184_, _25183_, _02974_);
  or (_25185_, _25184_, _25182_);
  and (_25186_, _25185_, _25145_);
  or (_25187_, _25186_, _09406_);
  or (_25188_, _25122_, _09405_);
  and (_25189_, _25188_, _02881_);
  and (_25191_, _25189_, _25187_);
  and (_25192_, _05368_, _02880_);
  or (_25193_, _25192_, _04252_);
  or (_25194_, _25193_, _25191_);
  nand (_25195_, _05311_, _04252_);
  and (_25196_, _25195_, _03336_);
  and (_25197_, _25196_, _25194_);
  and (_25198_, _05368_, _03069_);
  or (_25199_, _25198_, _09461_);
  or (_25200_, _25199_, _25197_);
  nand (_25202_, _25136_, _09461_);
  and (_25203_, _25202_, _03084_);
  and (_25204_, _25203_, _25200_);
  nand (_25205_, _05368_, _03075_);
  nand (_25206_, _25205_, _09470_);
  or (_25207_, _25206_, _25204_);
  or (_25208_, _25122_, _09470_);
  and (_25209_, _25208_, _02877_);
  and (_25210_, _25209_, _25207_);
  and (_25211_, _05368_, _02876_);
  or (_25213_, _25211_, _09474_);
  or (_25214_, _25213_, _25210_);
  nand (_25215_, _05311_, _09474_);
  and (_25216_, _25215_, _03941_);
  and (_25217_, _25216_, _25214_);
  nand (_25218_, _05368_, _02875_);
  nand (_25219_, _25218_, _09396_);
  or (_25220_, _25219_, _25217_);
  or (_25221_, _25142_, _09392_);
  nand (_25222_, _09392_, _05260_);
  and (_25224_, _25222_, _25221_);
  or (_25225_, _25224_, _09396_);
  and (_25226_, _25225_, _02979_);
  and (_25227_, _25226_, _25220_);
  or (_25228_, _25142_, _09357_);
  nand (_25229_, _09357_, _05260_);
  and (_25230_, _25229_, _02978_);
  and (_25231_, _25230_, _25228_);
  or (_25232_, _25231_, _02950_);
  or (_25233_, _25232_, _25227_);
  and (_25234_, _25142_, _23031_);
  and (_25235_, _09514_, _05259_);
  or (_25236_, _25235_, _09500_);
  or (_25237_, _25236_, _25234_);
  and (_25238_, _25237_, _09531_);
  and (_25239_, _25238_, _25233_);
  or (_25240_, _25142_, _09528_);
  nand (_25241_, _09528_, _05260_);
  and (_25242_, _25241_, _02952_);
  and (_25243_, _25242_, _25240_);
  or (_25246_, _25243_, _09489_);
  or (_25247_, _25246_, _25239_);
  and (_25248_, _25247_, _25137_);
  or (_25249_, _25248_, _02869_);
  nand (_25250_, _05369_, _02869_);
  and (_25251_, _25250_, _02614_);
  and (_25252_, _25251_, _25249_);
  nor (_25253_, _05311_, _02614_);
  or (_25254_, _25253_, _23051_);
  or (_25255_, _25254_, _25252_);
  and (_25257_, _25255_, _25134_);
  or (_25258_, _25257_, _09544_);
  or (_25259_, _25122_, _09543_);
  and (_25260_, _25259_, _09550_);
  and (_25261_, _25260_, _25258_);
  and (_25262_, _05368_, _03101_);
  or (_25263_, _25262_, _09551_);
  or (_25264_, _25263_, _25261_);
  nand (_25265_, _05311_, _09551_);
  and (_25266_, _25265_, _10016_);
  and (_25268_, _25266_, _25264_);
  nand (_25269_, _05368_, _03100_);
  nand (_25270_, _25269_, _09557_);
  or (_25271_, _25270_, _25268_);
  or (_25272_, _25122_, _09557_);
  and (_25273_, _25272_, _25271_);
  or (_25274_, _25273_, _09562_);
  or (_25275_, _09561_, _05368_);
  and (_25276_, _25275_, _02605_);
  and (_25277_, _25276_, _25274_);
  and (_25278_, _25122_, _02583_);
  or (_25279_, _25278_, _02863_);
  or (_25280_, _25279_, _25277_);
  and (_25281_, _25280_, _25133_);
  or (_25282_, _25281_, _02581_);
  nand (_25283_, _05311_, _02581_);
  and (_25284_, _25283_, _08209_);
  and (_25285_, _25284_, _25282_);
  nand (_25286_, _05259_, _02981_);
  nand (_25287_, _25286_, _02857_);
  or (_25290_, _25287_, _25285_);
  or (_25291_, _05368_, _02857_);
  and (_25292_, _25291_, _02838_);
  and (_25293_, _25292_, _25290_);
  nand (_25294_, _05259_, _02579_);
  nand (_25295_, _25294_, _09200_);
  or (_25296_, _25295_, _25293_);
  or (_25297_, _25122_, _09200_);
  and (_25298_, _25297_, _03490_);
  and (_25299_, _25298_, _25296_);
  and (_25301_, _05368_, _02933_);
  or (_25302_, _25301_, _02518_);
  or (_25303_, _25302_, _25299_);
  nand (_25304_, _05311_, _02518_);
  and (_25305_, _25304_, _09599_);
  and (_25306_, _25305_, _25303_);
  and (_25307_, _25150_, _09594_);
  or (_25308_, _25307_, _05754_);
  or (_25309_, _25308_, _25306_);
  and (_25310_, _25309_, _25132_);
  or (_25311_, _25310_, _02802_);
  nand (_25312_, _05260_, _02802_);
  and (_25313_, _25312_, _07860_);
  and (_25314_, _25313_, _25311_);
  and (_25315_, _07859_, _05368_);
  or (_25316_, _25315_, _09611_);
  or (_25317_, _25316_, _25314_);
  or (_25318_, _09615_, _09616_);
  nand (_25319_, _25318_, _09635_);
  or (_25320_, _25318_, _09635_);
  and (_25323_, _25320_, _25319_);
  or (_25324_, _25323_, _22679_);
  and (_25325_, _25324_, _03496_);
  and (_25326_, _25325_, _25317_);
  and (_25327_, _05368_, _02932_);
  or (_25328_, _25327_, _02514_);
  or (_25329_, _25328_, _25326_);
  nand (_25330_, _05311_, _02514_);
  and (_25331_, _25330_, _22678_);
  and (_25332_, _25331_, _25329_);
  or (_25334_, _25150_, _08165_);
  or (_25335_, _09676_, _05368_);
  and (_25336_, _25335_, _09083_);
  and (_25337_, _25336_, _25334_);
  or (_25338_, _25337_, _23884_);
  or (_25339_, _25338_, _25332_);
  and (_25340_, _25339_, _25131_);
  or (_25341_, _25340_, _09661_);
  or (_25342_, _09660_, _05368_);
  and (_25343_, _25342_, _03887_);
  and (_25345_, _25343_, _25341_);
  and (_25346_, _05259_, _02980_);
  or (_25347_, _25346_, _03127_);
  or (_25348_, _25347_, _25345_);
  nand (_25349_, _05369_, _03127_);
  and (_25350_, _25349_, _25348_);
  or (_25351_, _25350_, _02509_);
  nand (_25352_, _05311_, _02509_);
  and (_25353_, _25352_, _22675_);
  and (_25354_, _25353_, _25351_);
  or (_25356_, _25150_, _09676_);
  or (_25357_, _08165_, _05368_);
  and (_25358_, _25357_, _09672_);
  and (_25359_, _25358_, _25356_);
  or (_25360_, _25359_, _09681_);
  or (_25361_, _25360_, _25354_);
  and (_25362_, _25361_, _25130_);
  or (_25363_, _25362_, _22930_);
  or (_25364_, _09080_, _05368_);
  and (_25365_, _25364_, _03883_);
  and (_25366_, _25365_, _25363_);
  and (_25367_, _05259_, _02970_);
  or (_25368_, _25367_, _03135_);
  or (_25369_, _25368_, _25366_);
  nand (_25370_, _05369_, _03135_);
  and (_25371_, _25370_, _25369_);
  or (_25372_, _25371_, _03880_);
  nand (_25373_, _05311_, _03880_);
  and (_25374_, _25373_, _22667_);
  and (_25375_, _25374_, _25372_);
  or (_25378_, _25150_, \oc8051_golden_model_1.PSW [7]);
  or (_25379_, _05368_, _07293_);
  and (_25380_, _25379_, _09076_);
  and (_25381_, _25380_, _25378_);
  or (_25382_, _25381_, _09694_);
  or (_25383_, _25382_, _25375_);
  and (_25384_, _25383_, _25129_);
  or (_25385_, _25384_, _07944_);
  or (_25386_, _07943_, _05368_);
  and (_25387_, _25386_, _05783_);
  and (_25389_, _25387_, _25385_);
  and (_25390_, _05259_, _02965_);
  or (_25391_, _25390_, _03123_);
  or (_25392_, _25391_, _25389_);
  nand (_25393_, _05369_, _03123_);
  and (_25394_, _25393_, _25392_);
  or (_25395_, _25394_, _09069_);
  nand (_25396_, _05311_, _09069_);
  and (_25397_, _25396_, _23200_);
  and (_25398_, _25397_, _25395_);
  or (_25400_, _25150_, _07293_);
  or (_25401_, _05368_, \oc8051_golden_model_1.PSW [7]);
  and (_25402_, _25401_, _09068_);
  and (_25403_, _25402_, _25400_);
  or (_25404_, _25403_, _09711_);
  or (_25405_, _25404_, _25398_);
  and (_25406_, _25405_, _25128_);
  or (_25407_, _25406_, _10365_);
  or (_25408_, _09065_, _05368_);
  and (_25409_, _25408_, _07992_);
  and (_25411_, _25409_, _25407_);
  and (_25412_, _25122_, _07991_);
  or (_25413_, _25412_, _03145_);
  or (_25414_, _25413_, _25411_);
  or (_25415_, _05462_, _09726_);
  and (_25416_, _25415_, _25414_);
  or (_25417_, _25416_, _03898_);
  nand (_25418_, _05311_, _03898_);
  and (_25419_, _25418_, _03561_);
  and (_25420_, _25419_, _25417_);
  or (_25422_, _25142_, _23226_);
  or (_25423_, _09915_, _05259_);
  and (_25424_, _25423_, _02968_);
  and (_25425_, _25424_, _25422_);
  or (_25426_, _25425_, _25057_);
  or (_25427_, _25426_, _25420_);
  and (_25428_, _25427_, _25127_);
  or (_25429_, _25428_, _08067_);
  or (_25430_, _08066_, _05368_);
  and (_25431_, _25430_, _08112_);
  and (_25433_, _25431_, _25429_);
  and (_25434_, _25122_, _08111_);
  or (_25435_, _25434_, _02892_);
  or (_25436_, _25435_, _25433_);
  or (_25437_, _05462_, _02893_);
  and (_25438_, _25437_, _25436_);
  or (_25439_, _25438_, _22926_);
  nand (_25440_, _05311_, _22926_);
  and (_25441_, _25440_, _03164_);
  and (_25442_, _25441_, _25439_);
  nand (_25444_, _09915_, _05260_);
  or (_25445_, _25142_, _09915_);
  and (_25446_, _25445_, _25444_);
  and (_25447_, _25446_, _02940_);
  or (_25448_, _25447_, _09942_);
  or (_25449_, _25448_, _25442_);
  or (_25450_, _25122_, _09941_);
  and (_25451_, _25450_, _03906_);
  and (_25452_, _25451_, _25449_);
  nand (_25453_, _05368_, _03163_);
  nand (_25455_, _25453_, _09948_);
  or (_25456_, _25455_, _25452_);
  and (_25457_, _25456_, _25126_);
  or (_25458_, _25457_, _04337_);
  nand (_25459_, _05311_, _04337_);
  and (_25460_, _25459_, _02498_);
  and (_25461_, _25460_, _25458_);
  and (_25462_, _25446_, _02497_);
  or (_25463_, _25462_, _09964_);
  or (_25464_, _25463_, _25461_);
  nand (_25466_, _25136_, _09964_);
  and (_25467_, _25466_, _02890_);
  and (_25468_, _25467_, _25464_);
  or (_25469_, _25468_, _25125_);
  and (_25470_, _25469_, _09044_);
  nor (_25471_, _25136_, _09044_);
  or (_25472_, _25471_, _22655_);
  or (_25473_, _25472_, _25470_);
  nand (_25474_, _22655_, _05311_);
  and (_25475_, _25474_, _09983_);
  and (_25477_, _25475_, _25473_);
  or (_25478_, _25477_, _25123_);
  or (_25479_, _25478_, _42672_);
  or (_25480_, _42668_, \oc8051_golden_model_1.PC [7]);
  and (_25481_, _25480_, _43998_);
  and (_43502_, _25481_, _25479_);
  nor (_25482_, _09979_, _02523_);
  and (_25483_, _02835_, _02937_);
  and (_25484_, _02835_, _02939_);
  nor (_25485_, _09046_, \oc8051_golden_model_1.PC [8]);
  nor (_25487_, _25485_, _09053_);
  and (_25488_, _25487_, _08111_);
  nor (_25489_, _25487_, _09063_);
  nor (_25490_, _25487_, _09066_);
  nor (_25491_, _25487_, _09074_);
  nor (_25492_, _25487_, _09081_);
  and (_25493_, _09297_, _02980_);
  nor (_25494_, _25487_, _09657_);
  nor (_25495_, _09168_, _05753_);
  nor (_25496_, _09594_, _02518_);
  and (_25497_, _09168_, _02933_);
  nor (_25498_, _22940_, _09168_);
  not (_25499_, _09475_);
  and (_25500_, _09168_, _02876_);
  and (_25501_, _09168_, _03069_);
  and (_25502_, _09168_, _02880_);
  nor (_25503_, _09301_, _09295_);
  nor (_25504_, _25503_, _09302_);
  nor (_25505_, _25504_, _09412_);
  and (_25506_, _09298_, _09412_);
  nor (_25509_, _25506_, _25505_);
  or (_25510_, _25509_, _03810_);
  nor (_25511_, _09171_, _09166_);
  nor (_25512_, _25511_, _09172_);
  or (_25513_, _25512_, _09420_);
  not (_25514_, _09168_);
  nand (_25515_, _09420_, _25514_);
  and (_25516_, _25515_, _25513_);
  nor (_25517_, _25516_, _05362_);
  nor (_25518_, _03813_, _03072_);
  nor (_25520_, _25518_, _25514_);
  not (_25521_, _25487_);
  nor (_25522_, _25521_, _09430_);
  not (_25523_, _25522_);
  and (_25524_, _09427_, _02611_);
  not (_25525_, _25524_);
  and (_25526_, _03814_, \oc8051_golden_model_1.PC [8]);
  and (_25527_, _25526_, _09430_);
  nor (_25528_, _25527_, _25525_);
  and (_25529_, _25528_, _25523_);
  nor (_25531_, _25529_, _03072_);
  nor (_25532_, _25531_, _25520_);
  nor (_25533_, _25487_, _09427_);
  nor (_25534_, _25533_, _07646_);
  not (_25535_, _25534_);
  nor (_25536_, _25535_, _25532_);
  and (_25537_, _25487_, _07646_);
  and (_25538_, _05362_, _02616_);
  not (_25539_, _25538_);
  nor (_25540_, _25539_, _25537_);
  not (_25542_, _25540_);
  nor (_25543_, _25542_, _25536_);
  or (_25544_, _25543_, _02886_);
  nor (_25545_, _25544_, _25517_);
  and (_25546_, _25487_, _02886_);
  or (_25547_, _25546_, _02974_);
  or (_25548_, _25547_, _25545_);
  and (_25549_, _25548_, _25510_);
  nor (_25550_, _25549_, _09406_);
  nor (_25551_, _25487_, _09405_);
  nor (_25553_, _25551_, _02880_);
  not (_25554_, _25553_);
  nor (_25555_, _25554_, _25550_);
  nor (_25556_, _25555_, _25502_);
  nor (_25557_, _25556_, _04252_);
  and (_25558_, _25557_, _03336_);
  or (_25559_, _25558_, _09461_);
  nor (_25560_, _25559_, _25501_);
  and (_25561_, _25521_, _09461_);
  nor (_25562_, _25561_, _03075_);
  not (_25564_, _25562_);
  nor (_25565_, _25564_, _25560_);
  and (_25566_, _09168_, _03075_);
  nor (_25567_, _25566_, _09471_);
  not (_25568_, _25567_);
  nor (_25569_, _25568_, _25565_);
  nor (_25570_, _25487_, _09470_);
  nor (_25571_, _25570_, _02876_);
  not (_25572_, _25571_);
  nor (_25573_, _25572_, _25569_);
  nor (_25575_, _25573_, _25500_);
  nor (_25576_, _25575_, _25499_);
  and (_25577_, _09168_, _02875_);
  nor (_25578_, _25577_, _09481_);
  not (_25579_, _25578_);
  nor (_25580_, _25579_, _25576_);
  and (_25581_, _09392_, _09297_);
  not (_25582_, _25504_);
  nor (_25583_, _25582_, _09392_);
  or (_25584_, _25583_, _25581_);
  nor (_25586_, _25584_, _09396_);
  nor (_25587_, _25586_, _25580_);
  nor (_25588_, _25587_, _02978_);
  and (_25589_, _09357_, _09298_);
  nor (_25590_, _25504_, _09357_);
  nor (_25591_, _25590_, _25589_);
  nor (_25592_, _25591_, _02979_);
  or (_25593_, _25592_, _02950_);
  nor (_25594_, _25593_, _25588_);
  and (_25595_, _09514_, _09297_);
  nor (_25597_, _25582_, _09514_);
  nor (_25598_, _25597_, _25595_);
  nor (_25599_, _25598_, _09500_);
  nor (_25600_, _25599_, _25594_);
  nor (_25601_, _25600_, _02952_);
  and (_25602_, _09528_, _09297_);
  and (_25603_, _25504_, _09529_);
  or (_25604_, _25603_, _25602_);
  and (_25605_, _25604_, _02952_);
  nor (_25606_, _25605_, _25601_);
  or (_25608_, _25606_, _09489_);
  nand (_25609_, _25487_, _09489_);
  and (_25610_, _25609_, _25608_);
  or (_25611_, _25610_, _02869_);
  and (_25612_, _09168_, _02869_);
  not (_25613_, _25612_);
  and (_25614_, _22940_, _02614_);
  and (_25615_, _25614_, _25613_);
  and (_25616_, _25615_, _25611_);
  or (_25617_, _25616_, _25498_);
  nand (_25619_, _25617_, _09543_);
  nor (_25620_, _25487_, _09543_);
  nor (_25621_, _25620_, _03101_);
  nand (_25622_, _25621_, _25619_);
  and (_25623_, _09168_, _03101_);
  nor (_25624_, _25623_, _09551_);
  nand (_25625_, _25624_, _25622_);
  nand (_25626_, _25625_, _10016_);
  and (_25627_, _09168_, _03100_);
  nor (_25628_, _25627_, _14649_);
  and (_25630_, _25628_, _25626_);
  nor (_25631_, _25487_, _09557_);
  or (_25632_, _25631_, _25630_);
  nand (_25633_, _25632_, _09561_);
  nor (_25634_, _09168_, _09561_);
  nor (_25635_, _25634_, _02583_);
  nand (_25636_, _25635_, _25633_);
  and (_25637_, _25487_, _02583_);
  nor (_25638_, _25637_, _02863_);
  nand (_25639_, _25638_, _25636_);
  and (_25641_, _25514_, _02863_);
  nor (_25642_, _02981_, _02581_);
  not (_25643_, _25642_);
  nor (_25644_, _25643_, _25641_);
  nand (_25645_, _25644_, _25639_);
  and (_25646_, _09297_, _02981_);
  nor (_25647_, _25646_, _09582_);
  and (_25648_, _25647_, _25645_);
  nor (_25649_, _09168_, _02857_);
  or (_25650_, _25649_, _02579_);
  or (_25652_, _25650_, _25648_);
  and (_25653_, _09297_, _02579_);
  nor (_25654_, _25653_, _09203_);
  nand (_25655_, _25654_, _25652_);
  nor (_25656_, _25487_, _09200_);
  nor (_25657_, _25656_, _02933_);
  and (_25658_, _25657_, _25655_);
  or (_25659_, _25658_, _25497_);
  nand (_25660_, _25659_, _25496_);
  and (_25661_, _25512_, _09594_);
  nor (_25663_, _25661_, _05754_);
  and (_25664_, _25663_, _25660_);
  or (_25665_, _25664_, _25495_);
  nand (_25666_, _25665_, _02803_);
  and (_25667_, _09298_, _02802_);
  nor (_25668_, _25667_, _07859_);
  nand (_25669_, _25668_, _25666_);
  and (_25670_, _09168_, _07859_);
  nor (_25671_, _25670_, _09611_);
  nand (_25672_, _25671_, _25669_);
  nor (_25673_, _09637_, \oc8051_golden_model_1.DPH [0]);
  nor (_25674_, _25673_, _09638_);
  nor (_25675_, _25674_, _22679_);
  nor (_25676_, _25675_, _02932_);
  nand (_25677_, _25676_, _25672_);
  and (_25678_, _09168_, _02932_);
  nor (_25679_, _25678_, _02514_);
  nand (_25680_, _25679_, _25677_);
  nand (_25681_, _25680_, _22678_);
  nor (_25682_, _25512_, _08165_);
  nor (_25685_, _09168_, _09676_);
  nor (_25686_, _25685_, _22678_);
  not (_25687_, _25686_);
  nor (_25688_, _25687_, _25682_);
  nor (_25689_, _25688_, _23884_);
  and (_25690_, _25689_, _25681_);
  or (_25691_, _25690_, _25494_);
  nand (_25692_, _25691_, _09660_);
  nor (_25693_, _09660_, _09168_);
  nor (_25694_, _25693_, _02980_);
  and (_25696_, _25694_, _25692_);
  or (_25697_, _25696_, _25493_);
  nand (_25698_, _25697_, _03128_);
  and (_25699_, _09168_, _03127_);
  nor (_25700_, _25699_, _02509_);
  nand (_25701_, _25700_, _25698_);
  nand (_25702_, _25701_, _22675_);
  and (_25703_, _09168_, _09676_);
  and (_25704_, _25512_, _08165_);
  or (_25705_, _25704_, _25703_);
  and (_25707_, _25705_, _09672_);
  nor (_25708_, _25707_, _09681_);
  and (_25709_, _25708_, _25702_);
  or (_25710_, _25709_, _25492_);
  nand (_25711_, _25710_, _09080_);
  nor (_25712_, _09168_, _09080_);
  nor (_25713_, _25712_, _02970_);
  nand (_25714_, _25713_, _25711_);
  and (_25715_, _09297_, _02970_);
  nor (_25716_, _25715_, _03135_);
  nand (_25718_, _25716_, _25714_);
  nor (_25719_, _09076_, _03880_);
  not (_25720_, _25719_);
  and (_25721_, _25514_, _03135_);
  nor (_25722_, _25721_, _25720_);
  nand (_25723_, _25722_, _25718_);
  nor (_25724_, _25512_, \oc8051_golden_model_1.PSW [7]);
  nor (_25725_, _09168_, _07293_);
  nor (_25726_, _25725_, _22667_);
  not (_25727_, _25726_);
  nor (_25729_, _25727_, _25724_);
  nor (_25730_, _25729_, _09694_);
  and (_25731_, _25730_, _25723_);
  or (_25732_, _25731_, _25491_);
  nand (_25733_, _25732_, _07943_);
  nor (_25734_, _09168_, _07943_);
  nor (_25735_, _25734_, _02965_);
  and (_25736_, _25735_, _25733_);
  and (_25737_, _09297_, _02965_);
  or (_25738_, _25737_, _03123_);
  or (_25740_, _25738_, _25736_);
  nor (_25741_, _09068_, _09069_);
  not (_25742_, _25741_);
  and (_25743_, _25514_, _03123_);
  nor (_25744_, _25743_, _25742_);
  nand (_25745_, _25744_, _25740_);
  nor (_25746_, _25512_, _07293_);
  nor (_25747_, _09168_, \oc8051_golden_model_1.PSW [7]);
  nor (_25748_, _25747_, _23200_);
  not (_25749_, _25748_);
  nor (_25751_, _25749_, _25746_);
  nor (_25752_, _25751_, _09711_);
  and (_25753_, _25752_, _25745_);
  or (_25754_, _25753_, _25490_);
  nand (_25755_, _25754_, _09065_);
  nor (_25756_, _09168_, _09065_);
  nor (_25757_, _25756_, _07991_);
  and (_25758_, _25757_, _25755_);
  and (_25759_, _25487_, _07991_);
  or (_25760_, _25759_, _25758_);
  nand (_25762_, _25760_, _09726_);
  and (_25763_, _03808_, _03145_);
  nor (_25764_, _25763_, _03898_);
  nand (_25765_, _25764_, _25762_);
  nand (_25766_, _25765_, _03561_);
  nor (_25767_, _09915_, _09297_);
  and (_25768_, _25582_, _09915_);
  or (_25769_, _25768_, _03561_);
  or (_25770_, _25769_, _25767_);
  and (_25771_, _25770_, _09063_);
  and (_25773_, _25771_, _25766_);
  or (_25774_, _25773_, _25489_);
  nand (_25775_, _25774_, _08066_);
  nor (_25776_, _09168_, _08066_);
  nor (_25777_, _25776_, _08111_);
  and (_25778_, _25777_, _25775_);
  or (_25779_, _25778_, _25488_);
  nand (_25780_, _25779_, _02893_);
  and (_25781_, _03808_, _02892_);
  nor (_25782_, _25781_, _22926_);
  nand (_25784_, _25782_, _25780_);
  nand (_25785_, _25784_, _03164_);
  and (_25786_, _09915_, _09298_);
  nor (_25787_, _25504_, _09915_);
  nor (_25788_, _25787_, _25786_);
  and (_25789_, _25788_, _02940_);
  nor (_25790_, _25789_, _09942_);
  nand (_25791_, _25790_, _25785_);
  nor (_25792_, _25487_, _09941_);
  nor (_25793_, _25792_, _03163_);
  nand (_25795_, _25793_, _25791_);
  and (_25796_, _09168_, _03163_);
  nor (_25797_, _25796_, _09949_);
  nand (_25798_, _25797_, _25795_);
  nor (_25799_, _25487_, _09948_);
  nor (_25800_, _25799_, _02939_);
  and (_25801_, _25800_, _25798_);
  or (_25802_, _25801_, _25484_);
  nor (_25803_, _02497_, _02525_);
  nand (_25804_, _25803_, _25802_);
  and (_25806_, _25788_, _02497_);
  nor (_25807_, _25806_, _09964_);
  nand (_25808_, _25807_, _25804_);
  and (_25809_, _25521_, _09964_);
  nor (_25810_, _25809_, _02888_);
  nand (_25811_, _25810_, _25808_);
  and (_25812_, _09168_, _02888_);
  nor (_25813_, _25812_, _09970_);
  nand (_25814_, _25813_, _25811_);
  nor (_25815_, _25487_, _09044_);
  nor (_25817_, _25815_, _02937_);
  and (_25818_, _25817_, _25814_);
  or (_25819_, _25818_, _25483_);
  and (_25820_, _25819_, _25482_);
  and (_25821_, _25487_, _09979_);
  or (_25822_, _25821_, _25820_);
  or (_25823_, _25822_, _42672_);
  or (_25824_, _42668_, \oc8051_golden_model_1.PC [8]);
  and (_25825_, _25824_, _43998_);
  and (_43504_, _25825_, _25823_);
  nor (_25827_, _09043_, _03665_);
  nor (_25828_, _06173_, _03665_);
  nor (_25829_, _09053_, \oc8051_golden_model_1.PC [9]);
  nor (_25830_, _25829_, _09054_);
  nor (_25831_, _25830_, _09063_);
  and (_25832_, _09236_, _02965_);
  nor (_25833_, _25830_, _09074_);
  and (_25834_, _09236_, _02970_);
  nor (_25835_, _25830_, _09081_);
  and (_25836_, _09236_, _02980_);
  nor (_25838_, _25830_, _09657_);
  nor (_25839_, _09115_, _05753_);
  and (_25840_, _09115_, _02933_);
  and (_25841_, _09115_, _03100_);
  and (_25842_, _09115_, _03101_);
  and (_25843_, _09115_, _03069_);
  nand (_25844_, _09430_, _09426_);
  and (_25845_, _25844_, _25830_);
  and (_25846_, _03814_, \oc8051_golden_model_1.PC [9]);
  and (_25847_, _25846_, _09430_);
  not (_25849_, _09115_);
  or (_25850_, _25518_, _25849_);
  nand (_25851_, _25850_, _25524_);
  or (_25852_, _25851_, _25847_);
  or (_25853_, _25852_, _25845_);
  or (_25854_, _25830_, _22699_);
  nand (_25855_, _25849_, _03072_);
  and (_25856_, _25855_, _25854_);
  and (_25857_, _25856_, _25853_);
  nor (_25858_, _25857_, _25539_);
  and (_25860_, _09420_, _09115_);
  nor (_25861_, _09172_, _09169_);
  and (_25862_, _25861_, _09118_);
  nor (_25863_, _25861_, _09118_);
  nor (_25864_, _25863_, _25862_);
  nor (_25865_, _25864_, _09420_);
  or (_25866_, _25865_, _25860_);
  nor (_25867_, _25866_, _05362_);
  nor (_25868_, _25867_, _25858_);
  nor (_25869_, _25868_, _02886_);
  not (_25870_, _25830_);
  and (_25871_, _25870_, _02886_);
  or (_25872_, _25871_, _02974_);
  nor (_25873_, _25872_, _25869_);
  and (_25874_, _09237_, _09412_);
  nor (_25875_, _09302_, _09299_);
  and (_25876_, _25875_, _09240_);
  nor (_25877_, _25875_, _09240_);
  nor (_25878_, _25877_, _25876_);
  not (_25879_, _25878_);
  nor (_25882_, _25879_, _09412_);
  or (_25883_, _25882_, _03810_);
  nor (_25884_, _25883_, _25874_);
  or (_25885_, _25884_, _09406_);
  nor (_25886_, _25885_, _25873_);
  nor (_25887_, _25830_, _09405_);
  nor (_25888_, _25887_, _02880_);
  not (_25889_, _25888_);
  nor (_25890_, _25889_, _25886_);
  and (_25891_, _09115_, _02880_);
  or (_25893_, _25891_, _04252_);
  nor (_25894_, _25893_, _25890_);
  nor (_25895_, _25894_, _03069_);
  or (_25896_, _25895_, _09461_);
  nor (_25897_, _25896_, _25843_);
  and (_25898_, _25870_, _09461_);
  nor (_25899_, _25898_, _03075_);
  not (_25900_, _25899_);
  nor (_25901_, _25900_, _25897_);
  and (_25902_, _09115_, _03075_);
  nor (_25904_, _25902_, _09471_);
  not (_25905_, _25904_);
  nor (_25906_, _25905_, _25901_);
  nor (_25907_, _25830_, _09470_);
  nor (_25908_, _25907_, _02876_);
  not (_25909_, _25908_);
  nor (_25910_, _25909_, _25906_);
  and (_25911_, _09115_, _02876_);
  or (_25912_, _25911_, _09474_);
  nor (_25913_, _25912_, _25910_);
  nor (_25915_, _25913_, _02875_);
  and (_25916_, _09115_, _02875_);
  nor (_25917_, _25916_, _09481_);
  not (_25918_, _25917_);
  nor (_25919_, _25918_, _25915_);
  and (_25920_, _09392_, _09236_);
  nor (_25921_, _25878_, _09392_);
  or (_25922_, _25921_, _25920_);
  nor (_25923_, _25922_, _09396_);
  nor (_25924_, _25923_, _25919_);
  nor (_25926_, _25924_, _02978_);
  nor (_25927_, _25878_, _09357_);
  and (_25928_, _09357_, _09236_);
  or (_25929_, _25928_, _25927_);
  nor (_25930_, _25929_, _02979_);
  or (_25931_, _25930_, _02950_);
  nor (_25932_, _25931_, _25926_);
  nor (_25933_, _25878_, _09514_);
  and (_25934_, _09514_, _09236_);
  nor (_25935_, _25934_, _25933_);
  nor (_25937_, _25935_, _09500_);
  nor (_25938_, _25937_, _25932_);
  nor (_25939_, _25938_, _02952_);
  and (_25940_, _09528_, _09236_);
  nor (_25941_, _25878_, _09528_);
  or (_25942_, _25941_, _25940_);
  and (_25943_, _25942_, _02952_);
  or (_25944_, _25943_, _25939_);
  and (_25945_, _25944_, _09490_);
  and (_25946_, _25830_, _09489_);
  or (_25948_, _25946_, _25945_);
  nor (_25949_, _25948_, _02869_);
  and (_25950_, _25849_, _02869_);
  not (_25951_, _25950_);
  and (_25952_, _25951_, _25614_);
  not (_25953_, _25952_);
  nor (_25954_, _25953_, _25949_);
  nor (_25955_, _22940_, _25849_);
  nor (_25956_, _25955_, _09544_);
  not (_25957_, _25956_);
  nor (_25959_, _25957_, _25954_);
  nor (_25960_, _25830_, _09543_);
  nor (_25961_, _25960_, _03101_);
  not (_25962_, _25961_);
  nor (_25963_, _25962_, _25959_);
  or (_25964_, _25963_, _25842_);
  and (_25965_, _25964_, _09552_);
  or (_25966_, _25965_, _14649_);
  nor (_25967_, _25966_, _25841_);
  nor (_25968_, _25830_, _09557_);
  or (_25970_, _25968_, _25967_);
  nand (_25971_, _25970_, _09561_);
  nor (_25972_, _09115_, _09561_);
  nor (_25973_, _25972_, _02583_);
  nand (_25974_, _25973_, _25971_);
  and (_25975_, _25830_, _02583_);
  nor (_25976_, _25975_, _02863_);
  nand (_25977_, _25976_, _25974_);
  and (_25978_, _25849_, _02863_);
  nor (_25979_, _25978_, _25643_);
  nand (_25981_, _25979_, _25977_);
  and (_25982_, _09236_, _02981_);
  nor (_25983_, _25982_, _09582_);
  and (_25984_, _25983_, _25981_);
  nor (_25985_, _09115_, _02857_);
  or (_25986_, _25985_, _02579_);
  or (_25987_, _25986_, _25984_);
  and (_25988_, _09236_, _02579_);
  nor (_25989_, _25988_, _09203_);
  nand (_25990_, _25989_, _25987_);
  nor (_25992_, _25830_, _09200_);
  nor (_25993_, _25992_, _02933_);
  and (_25994_, _25993_, _25990_);
  or (_25995_, _25994_, _25840_);
  nand (_25996_, _25995_, _25496_);
  nor (_25997_, _25864_, _09599_);
  nor (_25998_, _25997_, _05754_);
  and (_25999_, _25998_, _25996_);
  or (_26000_, _25999_, _25839_);
  nand (_26001_, _26000_, _02803_);
  and (_26003_, _09237_, _02802_);
  nor (_26004_, _26003_, _07859_);
  nand (_26005_, _26004_, _26001_);
  and (_26006_, _09115_, _07859_);
  nor (_26007_, _26006_, _09611_);
  nand (_26008_, _26007_, _26005_);
  nor (_26009_, _09638_, \oc8051_golden_model_1.DPH [1]);
  nor (_26010_, _26009_, _09639_);
  nor (_26011_, _26010_, _22679_);
  nor (_26012_, _26011_, _02932_);
  nand (_26014_, _26012_, _26008_);
  and (_26015_, _09115_, _02932_);
  nor (_26016_, _26015_, _02514_);
  nand (_26017_, _26016_, _26014_);
  nand (_26018_, _26017_, _22678_);
  and (_26019_, _09115_, _08165_);
  nor (_26020_, _25864_, _08165_);
  or (_26021_, _26020_, _26019_);
  and (_26022_, _26021_, _09083_);
  nor (_26023_, _26022_, _23884_);
  and (_26025_, _26023_, _26018_);
  or (_26026_, _26025_, _25838_);
  nand (_26027_, _26026_, _09660_);
  nor (_26028_, _09660_, _09115_);
  nor (_26029_, _26028_, _02980_);
  and (_26030_, _26029_, _26027_);
  or (_26031_, _26030_, _25836_);
  nand (_26032_, _26031_, _03128_);
  and (_26033_, _09115_, _03127_);
  nor (_26034_, _26033_, _02509_);
  nand (_26036_, _26034_, _26032_);
  nand (_26037_, _26036_, _22675_);
  and (_26038_, _25864_, _08165_);
  nor (_26039_, _09115_, _08165_);
  nor (_26040_, _26039_, _22675_);
  not (_26041_, _26040_);
  nor (_26042_, _26041_, _26038_);
  nor (_26043_, _26042_, _09681_);
  and (_26044_, _26043_, _26037_);
  or (_26045_, _26044_, _25835_);
  nand (_26047_, _26045_, _09080_);
  nor (_26048_, _09115_, _09080_);
  nor (_26049_, _26048_, _02970_);
  and (_26050_, _26049_, _26047_);
  or (_26051_, _26050_, _25834_);
  nand (_26052_, _26051_, _03137_);
  and (_26053_, _09115_, _03135_);
  nor (_26054_, _26053_, _03880_);
  nand (_26055_, _26054_, _26052_);
  nand (_26056_, _26055_, _22667_);
  and (_26058_, _09115_, \oc8051_golden_model_1.PSW [7]);
  nor (_26059_, _25864_, \oc8051_golden_model_1.PSW [7]);
  or (_26060_, _26059_, _26058_);
  and (_26061_, _26060_, _09076_);
  nor (_26062_, _26061_, _09694_);
  and (_26063_, _26062_, _26056_);
  or (_26064_, _26063_, _25833_);
  nand (_26065_, _26064_, _07943_);
  nor (_26066_, _09115_, _07943_);
  nor (_26067_, _26066_, _02965_);
  and (_26069_, _26067_, _26065_);
  or (_26070_, _26069_, _25832_);
  nand (_26071_, _26070_, _05788_);
  and (_26072_, _09115_, _03123_);
  nor (_26073_, _26072_, _09069_);
  nand (_26074_, _26073_, _26071_);
  and (_26075_, _26074_, _23200_);
  and (_26076_, _09115_, _07293_);
  nor (_26077_, _25864_, _07293_);
  or (_26078_, _26077_, _26076_);
  and (_26080_, _26078_, _09068_);
  or (_26081_, _26080_, _26075_);
  nand (_26082_, _26081_, _09066_);
  nor (_26083_, _25870_, _09066_);
  nor (_26084_, _26083_, _10365_);
  nand (_26085_, _26084_, _26082_);
  nor (_26086_, _09115_, _09065_);
  nor (_26087_, _26086_, _07991_);
  nand (_26088_, _26087_, _26085_);
  and (_26089_, _25830_, _07991_);
  nor (_26091_, _26089_, _03145_);
  nand (_26092_, _26091_, _26088_);
  nor (_26093_, _02968_, _03898_);
  not (_26094_, _26093_);
  nor (_26095_, _04000_, _09726_);
  nor (_26096_, _26095_, _26094_);
  nand (_26097_, _26096_, _26092_);
  and (_26098_, _25878_, _09915_);
  nor (_26099_, _09915_, _09236_);
  or (_26100_, _26099_, _03561_);
  or (_26102_, _26100_, _26098_);
  and (_26103_, _26102_, _09063_);
  and (_26104_, _26103_, _26097_);
  or (_26105_, _26104_, _25831_);
  nand (_26106_, _26105_, _08066_);
  nor (_26107_, _09115_, _08066_);
  nor (_26108_, _26107_, _08111_);
  nand (_26109_, _26108_, _26106_);
  and (_26110_, _25830_, _08111_);
  nor (_26111_, _26110_, _02892_);
  nand (_26113_, _26111_, _26109_);
  nor (_26114_, _04000_, _02893_);
  nor (_26115_, _02940_, _22926_);
  not (_26116_, _26115_);
  nor (_26117_, _26116_, _26114_);
  nand (_26118_, _26117_, _26113_);
  and (_26119_, _09915_, _09237_);
  nor (_26120_, _25879_, _09915_);
  nor (_26121_, _26120_, _26119_);
  and (_26122_, _26121_, _02940_);
  nor (_26124_, _26122_, _09942_);
  nand (_26125_, _26124_, _26118_);
  nor (_26126_, _25830_, _09941_);
  nor (_26127_, _26126_, _03163_);
  nand (_26128_, _26127_, _26125_);
  and (_26129_, _09115_, _03163_);
  nor (_26130_, _26129_, _09949_);
  nand (_26131_, _26130_, _26128_);
  nor (_26132_, _25830_, _09948_);
  nor (_26133_, _26132_, _02939_);
  and (_26135_, _26133_, _26131_);
  or (_26136_, _26135_, _25828_);
  nand (_26137_, _26136_, _25803_);
  and (_26138_, _26121_, _02497_);
  nor (_26139_, _26138_, _09964_);
  nand (_26140_, _26139_, _26137_);
  and (_26141_, _25870_, _09964_);
  nor (_26142_, _26141_, _02888_);
  nand (_26143_, _26142_, _26140_);
  and (_26144_, _09115_, _02888_);
  nor (_26146_, _26144_, _09970_);
  nand (_26147_, _26146_, _26143_);
  nor (_26148_, _25830_, _09044_);
  nor (_26149_, _26148_, _02937_);
  and (_26150_, _26149_, _26147_);
  or (_26151_, _26150_, _25827_);
  and (_26152_, _26151_, _25482_);
  and (_26153_, _25830_, _09979_);
  or (_26154_, _26153_, _26152_);
  or (_26155_, _26154_, _42672_);
  or (_26157_, _42668_, \oc8051_golden_model_1.PC [9]);
  and (_26158_, _26157_, _43998_);
  and (_43505_, _26158_, _26155_);
  and (_26159_, _03256_, _02939_);
  nor (_26160_, _09054_, \oc8051_golden_model_1.PC [10]);
  nor (_26161_, _26160_, _09047_);
  nor (_26162_, _26161_, _09941_);
  not (_26163_, _26161_);
  and (_26164_, _26163_, _07991_);
  and (_26165_, _09229_, _02965_);
  and (_26167_, _09229_, _02970_);
  and (_26168_, _09229_, _02980_);
  not (_26169_, _09109_);
  and (_26170_, _26169_, _03100_);
  and (_26171_, _09109_, _02876_);
  and (_26172_, _26163_, _09461_);
  not (_26173_, _09232_);
  nor (_26174_, _09306_, _09303_);
  nor (_26175_, _26174_, _26173_);
  and (_26176_, _26174_, _26173_);
  nor (_26178_, _26176_, _26175_);
  nor (_26179_, _26178_, _09412_);
  and (_26180_, _09229_, _09412_);
  nor (_26181_, _26180_, _26179_);
  or (_26182_, _26181_, _03810_);
  not (_26183_, _09112_);
  nor (_26184_, _09176_, _09173_);
  nor (_26185_, _26184_, _26183_);
  and (_26186_, _26184_, _26183_);
  nor (_26187_, _26186_, _26185_);
  nor (_26189_, _26187_, _09420_);
  and (_26190_, _09420_, _26169_);
  nor (_26191_, _26190_, _26189_);
  nor (_26192_, _26191_, _05362_);
  nor (_26193_, _26161_, _09431_);
  nor (_26194_, _03813_, \oc8051_golden_model_1.PC [10]);
  and (_26195_, _26194_, _09430_);
  and (_26196_, _26195_, _25524_);
  nor (_26197_, _26196_, _26193_);
  nor (_26198_, _26197_, _03072_);
  nor (_26200_, _25518_, _09109_);
  nor (_26201_, _26200_, _07646_);
  not (_26202_, _26201_);
  nor (_26203_, _26202_, _26198_);
  and (_26204_, _26161_, _07646_);
  nor (_26205_, _26204_, _25539_);
  not (_26206_, _26205_);
  nor (_26207_, _26206_, _26203_);
  or (_26208_, _26207_, _02886_);
  nor (_26209_, _26208_, _26192_);
  and (_26211_, _26161_, _02886_);
  or (_26212_, _26211_, _02974_);
  or (_26213_, _26212_, _26209_);
  and (_26214_, _26213_, _26182_);
  nor (_26215_, _26214_, _09406_);
  nor (_26216_, _26161_, _09405_);
  nor (_26217_, _26216_, _02880_);
  not (_26218_, _26217_);
  nor (_26219_, _26218_, _26215_);
  nor (_26220_, _26219_, _04252_);
  nor (_26221_, _26220_, _03069_);
  nor (_26222_, _26169_, _03076_);
  nor (_26223_, _26222_, _09461_);
  not (_26224_, _26223_);
  nor (_26225_, _26224_, _26221_);
  nor (_26226_, _26225_, _26172_);
  nor (_26227_, _26226_, _03075_);
  and (_26228_, _26169_, _03075_);
  nor (_26229_, _26228_, _09471_);
  not (_26230_, _26229_);
  nor (_26233_, _26230_, _26227_);
  nor (_26234_, _26163_, _09470_);
  nor (_26235_, _26234_, _26233_);
  nor (_26236_, _26235_, _02876_);
  or (_26237_, _26236_, _09474_);
  nor (_26238_, _26237_, _26171_);
  nor (_26239_, _26238_, _02875_);
  and (_26240_, _09109_, _02875_);
  nor (_26241_, _26240_, _09481_);
  not (_26242_, _26241_);
  nor (_26244_, _26242_, _26239_);
  and (_26245_, _09392_, _09228_);
  not (_26246_, _26178_);
  nor (_26247_, _26246_, _09392_);
  or (_26248_, _26247_, _26245_);
  nor (_26249_, _26248_, _09396_);
  nor (_26250_, _26249_, _26244_);
  nor (_26251_, _26250_, _02978_);
  nor (_26252_, _26246_, _09357_);
  and (_26253_, _09357_, _09228_);
  nor (_26255_, _26253_, _26252_);
  and (_26256_, _26255_, _02978_);
  or (_26257_, _26256_, _02950_);
  nor (_26258_, _26257_, _26251_);
  and (_26259_, _09514_, _09228_);
  nor (_26260_, _26246_, _09514_);
  nor (_26261_, _26260_, _26259_);
  nor (_26262_, _26261_, _09500_);
  nor (_26263_, _26262_, _26258_);
  nor (_26264_, _26263_, _02952_);
  and (_26266_, _09528_, _09228_);
  and (_26267_, _26178_, _09529_);
  or (_26268_, _26267_, _26266_);
  and (_26269_, _26268_, _02952_);
  nor (_26270_, _26269_, _26264_);
  or (_26271_, _26270_, _09489_);
  nand (_26272_, _26161_, _09489_);
  and (_26273_, _26272_, _26271_);
  or (_26274_, _26273_, _02869_);
  nand (_26275_, _26274_, _02614_);
  nand (_26277_, _26275_, _22940_);
  and (_26278_, _22940_, _02870_);
  nor (_26279_, _26278_, _26169_);
  nor (_26280_, _26279_, _09544_);
  nand (_26281_, _26280_, _26277_);
  nor (_26282_, _26161_, _09543_);
  nor (_26283_, _26282_, _03101_);
  and (_26284_, _26283_, _26281_);
  and (_26285_, _09109_, _03101_);
  nor (_26286_, _26285_, _26284_);
  and (_26288_, _26286_, _09552_);
  or (_26289_, _26288_, _26170_);
  nand (_26290_, _26289_, _09557_);
  nor (_26291_, _26161_, _09557_);
  nor (_26292_, _26291_, _09562_);
  nand (_26293_, _26292_, _26290_);
  nor (_26294_, _26169_, _09561_);
  nor (_26295_, _26294_, _02583_);
  nand (_26296_, _26295_, _26293_);
  and (_26297_, _26163_, _02583_);
  nor (_26299_, _26297_, _02863_);
  and (_26300_, _26299_, _26296_);
  and (_26301_, _09109_, _02863_);
  nor (_26302_, _26301_, _26300_);
  and (_26303_, _26302_, _25642_);
  and (_26304_, _09229_, _02981_);
  or (_26305_, _26304_, _26303_);
  and (_26306_, _26305_, _02857_);
  nor (_26307_, _09109_, _02857_);
  or (_26308_, _26307_, _26306_);
  nand (_26310_, _26308_, _02838_);
  and (_26311_, _09229_, _02579_);
  nor (_26312_, _26311_, _09203_);
  and (_26313_, _26312_, _26310_);
  nor (_26314_, _26163_, _09200_);
  or (_26315_, _26314_, _26313_);
  nand (_26316_, _26315_, _03490_);
  and (_26317_, _09109_, _02933_);
  not (_26318_, _26317_);
  and (_26319_, _26318_, _25496_);
  nand (_26321_, _26319_, _26316_);
  nor (_26322_, _26187_, _09599_);
  nor (_26323_, _26322_, _05754_);
  and (_26324_, _26323_, _26321_);
  nor (_26325_, _26169_, _05753_);
  or (_26326_, _26325_, _02802_);
  or (_26327_, _26326_, _26324_);
  and (_26328_, _09229_, _02802_);
  nor (_26329_, _26328_, _07859_);
  nand (_26330_, _26329_, _26327_);
  and (_26331_, _09109_, _07859_);
  nor (_26332_, _26331_, _09611_);
  and (_26333_, _26332_, _26330_);
  nor (_26334_, _09639_, \oc8051_golden_model_1.DPH [2]);
  nor (_26335_, _26334_, _09640_);
  nor (_26336_, _26335_, _22679_);
  or (_26337_, _26336_, _26333_);
  or (_26338_, _26337_, _02932_);
  nand (_26339_, _09109_, _02932_);
  and (_26340_, _26339_, _26338_);
  or (_26343_, _26340_, _02514_);
  or (_26344_, _26343_, _09083_);
  and (_26345_, _09109_, _08165_);
  and (_26346_, _26187_, _09676_);
  or (_26347_, _26346_, _26345_);
  and (_26348_, _26347_, _09083_);
  nor (_26349_, _26348_, _23884_);
  nand (_26350_, _26349_, _26344_);
  nor (_26351_, _26161_, _09657_);
  nor (_26352_, _26351_, _09661_);
  nand (_26354_, _26352_, _26350_);
  nor (_26355_, _09660_, _26169_);
  nor (_26356_, _26355_, _02980_);
  and (_26357_, _26356_, _26354_);
  or (_26358_, _26357_, _26168_);
  nand (_26359_, _26358_, _03128_);
  and (_26360_, _26169_, _03127_);
  nor (_26361_, _09672_, _02509_);
  not (_26362_, _26361_);
  nor (_26363_, _26362_, _26360_);
  nand (_26365_, _26363_, _26359_);
  and (_26366_, _09109_, _09676_);
  and (_26367_, _26187_, _08165_);
  or (_26368_, _26367_, _26366_);
  and (_26369_, _26368_, _09672_);
  nor (_26370_, _26369_, _09681_);
  nand (_26371_, _26370_, _26365_);
  nor (_26372_, _26161_, _09081_);
  nor (_26373_, _26372_, _22930_);
  nand (_26374_, _26373_, _26371_);
  nor (_26376_, _26169_, _09080_);
  nor (_26377_, _26376_, _02970_);
  and (_26378_, _26377_, _26374_);
  or (_26379_, _26378_, _26167_);
  nand (_26380_, _26379_, _03137_);
  and (_26381_, _26169_, _03135_);
  nor (_26382_, _26381_, _25720_);
  nand (_26383_, _26382_, _26380_);
  and (_26384_, _09109_, \oc8051_golden_model_1.PSW [7]);
  and (_26385_, _26187_, _07293_);
  or (_26387_, _26385_, _26384_);
  and (_26388_, _26387_, _09076_);
  nor (_26389_, _26388_, _09694_);
  nand (_26390_, _26389_, _26383_);
  nor (_26391_, _26161_, _09074_);
  nor (_26392_, _26391_, _07944_);
  nand (_26393_, _26392_, _26390_);
  nor (_26394_, _26169_, _07943_);
  nor (_26395_, _26394_, _02965_);
  and (_26396_, _26395_, _26393_);
  or (_26398_, _26396_, _26165_);
  nand (_26399_, _26398_, _05788_);
  and (_26400_, _26169_, _03123_);
  nor (_26401_, _26400_, _25742_);
  nand (_26402_, _26401_, _26399_);
  and (_26403_, _09109_, _07293_);
  and (_26404_, _26187_, \oc8051_golden_model_1.PSW [7]);
  or (_26405_, _26404_, _26403_);
  and (_26406_, _26405_, _09068_);
  nor (_26407_, _26406_, _09711_);
  nand (_26409_, _26407_, _26402_);
  nor (_26410_, _26161_, _09066_);
  nor (_26411_, _26410_, _10365_);
  nand (_26412_, _26411_, _26409_);
  nor (_26413_, _26169_, _09065_);
  nor (_26414_, _26413_, _07991_);
  and (_26415_, _26414_, _26412_);
  or (_26416_, _26415_, _26164_);
  nand (_26417_, _26416_, _09726_);
  nor (_26418_, _04435_, _09726_);
  nor (_26420_, _26418_, _26094_);
  nand (_26421_, _26420_, _26417_);
  and (_26422_, _26246_, _09915_);
  nor (_26423_, _09915_, _09228_);
  or (_26424_, _26423_, _03561_);
  or (_26425_, _26424_, _26422_);
  and (_26426_, _26425_, _09063_);
  nand (_26427_, _26426_, _26421_);
  nor (_26428_, _26161_, _09063_);
  nor (_26429_, _26428_, _08067_);
  nand (_26431_, _26429_, _26427_);
  nor (_26432_, _26169_, _08066_);
  nor (_26433_, _26432_, _08111_);
  and (_26434_, _26433_, _26431_);
  and (_26435_, _26163_, _08111_);
  or (_26436_, _26435_, _26434_);
  nand (_26437_, _26436_, _02893_);
  nor (_26438_, _04435_, _02893_);
  nor (_26439_, _26438_, _26116_);
  nand (_26440_, _26439_, _26437_);
  and (_26442_, _09915_, _09229_);
  nor (_26443_, _26178_, _09915_);
  nor (_26444_, _26443_, _26442_);
  and (_26445_, _26444_, _02940_);
  nor (_26446_, _26445_, _09942_);
  and (_26447_, _26446_, _26440_);
  or (_26448_, _26447_, _26162_);
  nand (_26449_, _26448_, _03906_);
  and (_26450_, _26169_, _03163_);
  nor (_26451_, _26450_, _09949_);
  nand (_26453_, _26451_, _26449_);
  nor (_26454_, _26163_, _09948_);
  nor (_26455_, _26454_, _02939_);
  nand (_26456_, _26455_, _26453_);
  nand (_26457_, _26456_, _25803_);
  or (_26458_, _26457_, _26159_);
  and (_26459_, _26444_, _02497_);
  nor (_26460_, _26459_, _09964_);
  and (_26461_, _26460_, _26458_);
  and (_26462_, _26163_, _09964_);
  or (_26464_, _26462_, _26461_);
  nand (_26465_, _26464_, _02890_);
  and (_26466_, _26169_, _02888_);
  nor (_26467_, _26466_, _09970_);
  nand (_26468_, _26467_, _26465_);
  nor (_26469_, _26163_, _09044_);
  nor (_26470_, _26469_, _02937_);
  nand (_26471_, _26470_, _26468_);
  not (_26472_, _25482_);
  and (_26473_, _03256_, _02937_);
  nor (_26475_, _26473_, _26472_);
  and (_26476_, _26475_, _26471_);
  and (_26477_, _26161_, _09979_);
  or (_26478_, _26477_, _26476_);
  or (_26479_, _26478_, _42672_);
  or (_26480_, _42668_, \oc8051_golden_model_1.PC [10]);
  and (_26481_, _26480_, _43998_);
  and (_43506_, _26481_, _26479_);
  nor (_26482_, _09047_, _09219_);
  and (_26483_, _09047_, _09219_);
  or (_26485_, _26483_, _26482_);
  or (_26486_, _26485_, _09063_);
  or (_26487_, _26485_, _09066_);
  or (_26488_, _09104_, _09070_);
  and (_26489_, _26488_, _23200_);
  or (_26490_, _26485_, _09074_);
  or (_26491_, _09104_, _09077_);
  and (_26492_, _26491_, _22667_);
  or (_26493_, _26485_, _09081_);
  nor (_26494_, _26185_, _09110_);
  and (_26496_, _26494_, _09107_);
  nor (_26497_, _26494_, _09107_);
  or (_26498_, _26497_, _26496_);
  or (_26499_, _26498_, _08165_);
  or (_26500_, _09104_, _09676_);
  and (_26501_, _26500_, _09083_);
  and (_26502_, _26501_, _26499_);
  or (_26503_, _09104_, _05753_);
  and (_26504_, _09222_, _02579_);
  or (_26505_, _09104_, _02857_);
  and (_26507_, _26505_, _02838_);
  nor (_26508_, _26175_, _09230_);
  and (_26509_, _26508_, _09226_);
  nor (_26510_, _26508_, _09226_);
  or (_26511_, _26510_, _26509_);
  or (_26512_, _26511_, _09528_);
  nand (_26513_, _09528_, _09223_);
  and (_26514_, _26513_, _02952_);
  and (_26515_, _26514_, _26512_);
  nand (_26516_, _09392_, _09223_);
  or (_26518_, _26511_, _09392_);
  and (_26519_, _26518_, _09481_);
  and (_26520_, _26519_, _26516_);
  and (_26521_, _09104_, _03075_);
  or (_26522_, _09402_, _09104_);
  nand (_26523_, _09223_, _09412_);
  or (_26524_, _26511_, _09412_);
  and (_26525_, _26524_, _02974_);
  and (_26526_, _26525_, _26523_);
  and (_26527_, _26498_, _24086_);
  and (_26529_, _09420_, _09104_);
  or (_26530_, _26529_, _05362_);
  or (_26531_, _26530_, _26527_);
  and (_26532_, _09104_, _03072_);
  not (_26533_, _09104_);
  nor (_26534_, _09434_, _26533_);
  and (_26535_, _02611_, \oc8051_golden_model_1.PC [11]);
  and (_26536_, _26535_, _25518_);
  and (_26537_, _26536_, _09430_);
  or (_26538_, _26537_, _26534_);
  and (_26540_, _26538_, _09427_);
  or (_26541_, _26540_, _26532_);
  and (_26542_, _26541_, _09426_);
  not (_26543_, _26485_);
  nor (_26544_, _26543_, _09432_);
  or (_26545_, _26544_, _26542_);
  and (_26546_, _26545_, _02616_);
  or (_26547_, _26533_, _02616_);
  nand (_26548_, _26547_, _05362_);
  or (_26549_, _26548_, _26546_);
  and (_26551_, _26549_, _09449_);
  and (_26552_, _26551_, _26531_);
  or (_26553_, _26552_, _26526_);
  and (_26554_, _26553_, _09405_);
  not (_26555_, _09402_);
  nor (_26556_, _26543_, _09456_);
  or (_26557_, _26556_, _26555_);
  or (_26558_, _26557_, _26554_);
  and (_26559_, _26558_, _26522_);
  or (_26560_, _26559_, _09461_);
  nand (_26562_, _26543_, _09461_);
  and (_26563_, _26562_, _03084_);
  and (_26564_, _26563_, _26560_);
  or (_26565_, _26564_, _26521_);
  and (_26566_, _26565_, _09470_);
  or (_26567_, _26543_, _09470_);
  nand (_26568_, _26567_, _09476_);
  or (_26569_, _26568_, _26566_);
  or (_26570_, _09476_, _09104_);
  and (_26571_, _26570_, _09396_);
  and (_26573_, _26571_, _26569_);
  or (_26574_, _26573_, _26520_);
  and (_26575_, _26574_, _02979_);
  nand (_26576_, _09357_, _09223_);
  or (_26577_, _26511_, _09357_);
  and (_26578_, _26577_, _02978_);
  and (_26579_, _26578_, _26576_);
  or (_26580_, _26579_, _02950_);
  or (_26581_, _26580_, _26575_);
  and (_26582_, _09514_, _09222_);
  and (_26584_, _26511_, _23031_);
  or (_26585_, _26584_, _09500_);
  or (_26586_, _26585_, _26582_);
  and (_26587_, _26586_, _09531_);
  and (_26588_, _26587_, _26581_);
  or (_26589_, _26588_, _26515_);
  and (_26590_, _26589_, _09490_);
  nand (_26591_, _26485_, _09489_);
  nand (_26592_, _26591_, _09498_);
  or (_26593_, _26592_, _26590_);
  or (_26595_, _09498_, _09104_);
  and (_26596_, _26595_, _09543_);
  and (_26597_, _26596_, _26593_);
  nor (_26598_, _26543_, _09543_);
  or (_26599_, _26598_, _09554_);
  or (_26600_, _26599_, _26597_);
  or (_26601_, _09553_, _09104_);
  and (_26602_, _26601_, _09557_);
  and (_26603_, _26602_, _26600_);
  nor (_26604_, _26543_, _09557_);
  or (_26606_, _26604_, _09562_);
  or (_26607_, _26606_, _26603_);
  or (_26608_, _09104_, _09561_);
  and (_26609_, _26608_, _02605_);
  and (_26610_, _26609_, _26607_);
  nand (_26611_, _26485_, _02583_);
  nand (_26612_, _26611_, _09572_);
  or (_26613_, _26612_, _26610_);
  or (_26614_, _09572_, _09104_);
  and (_26615_, _26614_, _08209_);
  and (_26617_, _26615_, _26613_);
  nand (_26618_, _09222_, _02981_);
  nand (_26619_, _26618_, _02857_);
  or (_26620_, _26619_, _26617_);
  and (_26621_, _26620_, _26507_);
  or (_26622_, _26621_, _26504_);
  and (_26623_, _26622_, _09200_);
  nor (_26624_, _26543_, _09200_);
  or (_26625_, _26624_, _09592_);
  or (_26626_, _26625_, _26623_);
  or (_26628_, _09591_, _09104_);
  and (_26629_, _26628_, _09599_);
  and (_26630_, _26629_, _26626_);
  and (_26631_, _26498_, _09594_);
  or (_26632_, _26631_, _05754_);
  or (_26633_, _26632_, _26630_);
  and (_26634_, _26633_, _26503_);
  or (_26635_, _26634_, _02802_);
  nand (_26636_, _09223_, _02802_);
  and (_26637_, _26636_, _07860_);
  and (_26639_, _26637_, _26635_);
  and (_26640_, _09104_, _07859_);
  or (_26641_, _26640_, _26639_);
  and (_26642_, _26641_, _22679_);
  nor (_26643_, _09640_, \oc8051_golden_model_1.DPH [3]);
  nor (_26644_, _26643_, _09641_);
  and (_26645_, _26644_, _09611_);
  or (_26646_, _26645_, _09650_);
  or (_26647_, _26646_, _26642_);
  or (_26648_, _09649_, _09104_);
  and (_26650_, _26648_, _22678_);
  and (_26651_, _26650_, _26647_);
  or (_26652_, _26651_, _26502_);
  and (_26653_, _26652_, _09657_);
  nor (_26654_, _26543_, _09657_);
  or (_26655_, _26654_, _09661_);
  or (_26656_, _26655_, _26653_);
  or (_26657_, _09660_, _09104_);
  and (_26658_, _26657_, _03887_);
  and (_26659_, _26658_, _26656_);
  nand (_26661_, _09222_, _02980_);
  nand (_26662_, _26661_, _09668_);
  or (_26663_, _26662_, _26659_);
  or (_26664_, _09668_, _09104_);
  and (_26665_, _26664_, _22675_);
  and (_26666_, _26665_, _26663_);
  or (_26667_, _26498_, _09676_);
  or (_26668_, _09104_, _08165_);
  and (_26669_, _26668_, _09672_);
  and (_26670_, _26669_, _26667_);
  or (_26672_, _26670_, _09681_);
  or (_26673_, _26672_, _26666_);
  and (_26674_, _26673_, _26493_);
  or (_26675_, _26674_, _22930_);
  or (_26676_, _09104_, _09080_);
  and (_26677_, _26676_, _03883_);
  and (_26678_, _26677_, _26675_);
  nand (_26679_, _09222_, _02970_);
  nand (_26680_, _26679_, _09077_);
  or (_26681_, _26680_, _26678_);
  and (_26683_, _26681_, _26492_);
  or (_26684_, _26498_, \oc8051_golden_model_1.PSW [7]);
  or (_26685_, _09104_, _07293_);
  and (_26686_, _26685_, _09076_);
  and (_26687_, _26686_, _26684_);
  or (_26688_, _26687_, _09694_);
  or (_26689_, _26688_, _26683_);
  and (_26690_, _26689_, _26490_);
  or (_26691_, _26690_, _07944_);
  or (_26692_, _09104_, _07943_);
  and (_26694_, _26692_, _05783_);
  and (_26695_, _26694_, _26691_);
  nand (_26696_, _09222_, _02965_);
  nand (_26697_, _26696_, _09070_);
  or (_26698_, _26697_, _26695_);
  and (_26699_, _26698_, _26489_);
  or (_26700_, _26498_, _07293_);
  or (_26701_, _09104_, \oc8051_golden_model_1.PSW [7]);
  and (_26702_, _26701_, _09068_);
  and (_26703_, _26702_, _26700_);
  or (_26705_, _26703_, _09711_);
  or (_26706_, _26705_, _26699_);
  and (_26707_, _26706_, _26487_);
  or (_26708_, _26707_, _10365_);
  or (_26709_, _09104_, _09065_);
  and (_26710_, _26709_, _07992_);
  and (_26711_, _26710_, _26708_);
  and (_26712_, _26485_, _07991_);
  or (_26713_, _26712_, _03145_);
  or (_26714_, _26713_, _26711_);
  or (_26716_, _04241_, _09726_);
  and (_26717_, _26716_, _26714_);
  or (_26718_, _26717_, _03898_);
  nor (_26719_, _09104_, _02529_);
  nor (_26720_, _26719_, _02968_);
  and (_26721_, _26720_, _26718_);
  or (_26722_, _26511_, _23226_);
  or (_26723_, _09915_, _09222_);
  and (_26724_, _26723_, _02968_);
  and (_26725_, _26724_, _26722_);
  or (_26727_, _26725_, _25057_);
  or (_26728_, _26727_, _26721_);
  and (_26729_, _26728_, _26486_);
  or (_26730_, _26729_, _08067_);
  or (_26731_, _09104_, _08066_);
  and (_26732_, _26731_, _08112_);
  and (_26733_, _26732_, _26730_);
  and (_26734_, _26485_, _08111_);
  or (_26735_, _26734_, _02892_);
  or (_26736_, _26735_, _26733_);
  or (_26738_, _04241_, _02893_);
  and (_26739_, _26738_, _26736_);
  or (_26740_, _26739_, _22926_);
  nor (_26741_, _09104_, _02537_);
  nor (_26742_, _26741_, _02940_);
  and (_26743_, _26742_, _26740_);
  or (_26744_, _26511_, _09915_);
  nand (_26745_, _09915_, _09223_);
  and (_26746_, _26745_, _26744_);
  and (_26747_, _26746_, _02940_);
  or (_26749_, _26747_, _09942_);
  or (_26750_, _26749_, _26743_);
  or (_26751_, _26485_, _09941_);
  and (_26752_, _26751_, _03906_);
  and (_26753_, _26752_, _26750_);
  nand (_26754_, _09104_, _03163_);
  nand (_26755_, _26754_, _09948_);
  or (_26756_, _26755_, _26753_);
  or (_26757_, _26485_, _09948_);
  and (_26758_, _26757_, _06173_);
  and (_26760_, _26758_, _26756_);
  nor (_26761_, _06173_, _02794_);
  or (_26762_, _26761_, _02525_);
  or (_26763_, _26762_, _26760_);
  nand (_26764_, _26533_, _02525_);
  and (_26765_, _26764_, _02498_);
  and (_26766_, _26765_, _26763_);
  and (_26767_, _26746_, _02497_);
  or (_26768_, _26767_, _09964_);
  or (_26769_, _26768_, _26766_);
  nand (_26771_, _26543_, _09964_);
  and (_26772_, _26771_, _02890_);
  and (_26773_, _26772_, _26769_);
  nand (_26774_, _09104_, _02888_);
  nand (_26775_, _26774_, _09044_);
  or (_26776_, _26775_, _26773_);
  or (_26777_, _26485_, _09044_);
  and (_26778_, _26777_, _09043_);
  and (_26779_, _26778_, _26776_);
  nor (_26780_, _09043_, _02794_);
  or (_26781_, _26780_, _02523_);
  or (_26782_, _26781_, _26779_);
  nand (_26783_, _26533_, _02523_);
  and (_26784_, _26783_, _09983_);
  and (_26785_, _26784_, _26782_);
  and (_26786_, _26485_, _09979_);
  or (_26787_, _26786_, _26785_);
  or (_26788_, _26787_, _42672_);
  or (_26789_, _42668_, \oc8051_golden_model_1.PC [11]);
  and (_26790_, _26789_, _43998_);
  and (_43507_, _26790_, _26788_);
  nor (_26793_, _09048_, \oc8051_golden_model_1.PC [12]);
  nor (_26794_, _26793_, _09049_);
  not (_26795_, _26794_);
  nand (_26796_, _26795_, _09979_);
  nand (_26797_, _26795_, _08111_);
  nor (_26798_, _12395_, _09070_);
  nor (_26799_, _12395_, _09077_);
  nor (_26800_, _09668_, _12395_);
  nor (_26801_, _09649_, _12395_);
  or (_26803_, _09101_, _05753_);
  nor (_26804_, _12395_, _02857_);
  or (_26805_, _26804_, _02579_);
  nor (_26806_, _09313_, _09311_);
  nor (_26807_, _26806_, _09314_);
  and (_26808_, _26807_, _23025_);
  and (_26809_, _09357_, _09217_);
  or (_26810_, _26809_, _26808_);
  and (_26811_, _26810_, _02978_);
  nor (_26812_, _26795_, _09470_);
  nand (_26814_, _26795_, _09461_);
  and (_26815_, _26807_, _24823_);
  and (_26816_, _09217_, _09412_);
  or (_26817_, _26816_, _03810_);
  or (_26818_, _26817_, _26815_);
  nor (_26819_, _09183_, _09181_);
  nor (_26820_, _26819_, _09184_);
  and (_26821_, _26820_, _24086_);
  and (_26822_, _09420_, _09101_);
  or (_26823_, _26822_, _05362_);
  or (_26825_, _26823_, _26821_);
  or (_26826_, _26794_, _09427_);
  nor (_26827_, _09434_, _12395_);
  nor (_26828_, _26795_, _09431_);
  not (_26829_, \oc8051_golden_model_1.PC [12]);
  nor (_26830_, _03813_, _26829_);
  and (_26831_, _26830_, _09430_);
  or (_26832_, _26831_, _26828_);
  and (_26833_, _26832_, _02611_);
  or (_26834_, _26833_, _26827_);
  and (_26836_, _26834_, _26826_);
  or (_26837_, _26836_, _03072_);
  nand (_26838_, _12395_, _03072_);
  and (_26839_, _26838_, _09426_);
  and (_26840_, _26839_, _26837_);
  and (_26841_, _26794_, _07646_);
  or (_26842_, _26841_, _26840_);
  and (_26843_, _26842_, _02616_);
  or (_26844_, _12395_, _02616_);
  nand (_26845_, _26844_, _05362_);
  or (_26847_, _26845_, _26843_);
  and (_26848_, _26847_, _04265_);
  and (_26849_, _26848_, _26825_);
  and (_26850_, _26794_, _02886_);
  or (_26851_, _26850_, _02974_);
  or (_26852_, _26851_, _26849_);
  and (_26853_, _26852_, _26818_);
  or (_26854_, _26853_, _09406_);
  or (_26855_, _26794_, _09405_);
  and (_26856_, _26855_, _09402_);
  and (_26858_, _26856_, _26854_);
  nor (_26859_, _09402_, _12395_);
  or (_26860_, _26859_, _09461_);
  or (_26861_, _26860_, _26858_);
  and (_26862_, _26861_, _26814_);
  or (_26863_, _26862_, _03075_);
  nand (_26864_, _12395_, _03075_);
  and (_26865_, _26864_, _09470_);
  and (_26866_, _26865_, _26863_);
  or (_26867_, _26866_, _26812_);
  and (_26869_, _26867_, _09476_);
  or (_26870_, _09476_, _12395_);
  nand (_26871_, _26870_, _09396_);
  or (_26872_, _26871_, _26869_);
  and (_26873_, _09392_, _09217_);
  not (_26874_, _09392_);
  and (_26875_, _26807_, _26874_);
  or (_26876_, _26875_, _26873_);
  or (_26877_, _26876_, _09396_);
  and (_26878_, _26877_, _02979_);
  and (_26880_, _26878_, _26872_);
  or (_26881_, _26880_, _02950_);
  or (_26882_, _26881_, _26811_);
  and (_26883_, _26807_, _23031_);
  and (_26884_, _09514_, _09217_);
  or (_26885_, _26884_, _09500_);
  or (_26886_, _26885_, _26883_);
  and (_26887_, _26886_, _09531_);
  and (_26888_, _26887_, _26882_);
  or (_26889_, _26807_, _09528_);
  or (_26891_, _09529_, _09217_);
  and (_26892_, _26891_, _02952_);
  and (_26893_, _26892_, _26889_);
  or (_26894_, _26893_, _09489_);
  or (_26895_, _26894_, _26888_);
  nand (_26896_, _26795_, _09489_);
  and (_26897_, _26896_, _09498_);
  and (_26898_, _26897_, _26895_);
  nor (_26899_, _09498_, _12395_);
  or (_26900_, _26899_, _09544_);
  or (_26902_, _26900_, _26898_);
  or (_26903_, _26794_, _09543_);
  and (_26904_, _26903_, _09553_);
  and (_26905_, _26904_, _26902_);
  or (_26906_, _09553_, _12395_);
  nand (_26907_, _26906_, _09557_);
  or (_26908_, _26907_, _26905_);
  nor (_26909_, _26794_, _09557_);
  nor (_26910_, _26909_, _09562_);
  and (_26911_, _26910_, _26908_);
  nor (_26913_, _12395_, _09561_);
  or (_26914_, _26913_, _02583_);
  or (_26915_, _26914_, _26911_);
  nand (_26916_, _26795_, _02583_);
  and (_26917_, _26916_, _09572_);
  and (_26918_, _26917_, _26915_);
  nor (_26919_, _09572_, _12395_);
  or (_26920_, _26919_, _02981_);
  or (_26921_, _26920_, _26918_);
  or (_26922_, _09217_, _08209_);
  and (_26924_, _26922_, _02857_);
  and (_26925_, _26924_, _26921_);
  or (_26926_, _26925_, _26805_);
  or (_26927_, _09217_, _02838_);
  and (_26928_, _26927_, _09200_);
  and (_26929_, _26928_, _26926_);
  nor (_26930_, _26795_, _09200_);
  or (_26931_, _26930_, _09592_);
  or (_26932_, _26931_, _26929_);
  or (_26933_, _09591_, _09101_);
  and (_26935_, _26933_, _09599_);
  and (_26936_, _26935_, _26932_);
  and (_26937_, _26820_, _09594_);
  or (_26938_, _26937_, _05754_);
  or (_26939_, _26938_, _26936_);
  and (_26940_, _26939_, _26803_);
  or (_26941_, _26940_, _02802_);
  or (_26942_, _09217_, _02803_);
  and (_26943_, _26942_, _07860_);
  and (_26944_, _26943_, _26941_);
  and (_26947_, _09101_, _07859_);
  or (_26948_, _26947_, _09611_);
  or (_26949_, _26948_, _26944_);
  nor (_26950_, _09641_, \oc8051_golden_model_1.DPH [4]);
  nor (_26951_, _26950_, _09642_);
  or (_26952_, _26951_, _22679_);
  and (_26953_, _26952_, _09649_);
  and (_26954_, _26953_, _26949_);
  or (_26955_, _26954_, _26801_);
  and (_26956_, _26955_, _22678_);
  or (_26958_, _26820_, _08165_);
  or (_26959_, _09101_, _09676_);
  and (_26960_, _26959_, _09083_);
  and (_26961_, _26960_, _26958_);
  or (_26962_, _26961_, _23884_);
  or (_26963_, _26962_, _26956_);
  or (_26964_, _26794_, _09657_);
  and (_26965_, _26964_, _09660_);
  and (_26966_, _26965_, _26963_);
  nor (_26967_, _09660_, _12395_);
  or (_26969_, _26967_, _02980_);
  or (_26970_, _26969_, _26966_);
  or (_26971_, _09217_, _03887_);
  and (_26972_, _26971_, _09668_);
  and (_26973_, _26972_, _26970_);
  or (_26974_, _26973_, _26800_);
  and (_26975_, _26974_, _22675_);
  or (_26976_, _26820_, _09676_);
  or (_26977_, _09101_, _08165_);
  and (_26978_, _26977_, _09672_);
  and (_26980_, _26978_, _26976_);
  or (_26981_, _26980_, _09681_);
  or (_26982_, _26981_, _26975_);
  or (_26983_, _26794_, _09081_);
  and (_26984_, _26983_, _09080_);
  and (_26985_, _26984_, _26982_);
  nor (_26986_, _12395_, _09080_);
  or (_26987_, _26986_, _02970_);
  or (_26988_, _26987_, _26985_);
  or (_26989_, _09217_, _03883_);
  and (_26991_, _26989_, _09077_);
  and (_26992_, _26991_, _26988_);
  or (_26993_, _26992_, _26799_);
  and (_26994_, _26993_, _22667_);
  or (_26995_, _26820_, \oc8051_golden_model_1.PSW [7]);
  or (_26996_, _09101_, _07293_);
  and (_26997_, _26996_, _09076_);
  and (_26998_, _26997_, _26995_);
  or (_26999_, _26998_, _09694_);
  or (_27000_, _26999_, _26994_);
  or (_27002_, _26794_, _09074_);
  and (_27003_, _27002_, _07943_);
  and (_27004_, _27003_, _27000_);
  nor (_27005_, _12395_, _07943_);
  or (_27006_, _27005_, _02965_);
  or (_27007_, _27006_, _27004_);
  or (_27008_, _09217_, _05783_);
  and (_27009_, _27008_, _09070_);
  and (_27010_, _27009_, _27007_);
  or (_27011_, _27010_, _26798_);
  and (_27013_, _27011_, _23200_);
  or (_27014_, _26820_, _07293_);
  or (_27015_, _09101_, \oc8051_golden_model_1.PSW [7]);
  and (_27016_, _27015_, _09068_);
  and (_27017_, _27016_, _27014_);
  or (_27018_, _27017_, _09711_);
  or (_27019_, _27018_, _27013_);
  or (_27020_, _26794_, _09066_);
  and (_27021_, _27020_, _09065_);
  and (_27022_, _27021_, _27019_);
  nor (_27024_, _12395_, _09065_);
  or (_27025_, _27024_, _07991_);
  or (_27026_, _27025_, _27022_);
  nand (_27027_, _26795_, _07991_);
  and (_27028_, _27027_, _09726_);
  and (_27029_, _27028_, _27026_);
  and (_27030_, _04982_, _03145_);
  or (_27031_, _27030_, _03898_);
  or (_27032_, _27031_, _27029_);
  nor (_27033_, _09101_, _02529_);
  nor (_27035_, _27033_, _02968_);
  and (_27036_, _27035_, _27032_);
  or (_27037_, _09915_, _09217_);
  or (_27038_, _26807_, _23226_);
  and (_27039_, _27038_, _02968_);
  and (_27040_, _27039_, _27037_);
  or (_27041_, _27040_, _25057_);
  or (_27042_, _27041_, _27036_);
  or (_27043_, _26794_, _09063_);
  and (_27044_, _27043_, _08066_);
  and (_27046_, _27044_, _27042_);
  nor (_27047_, _12395_, _08066_);
  or (_27048_, _27047_, _08111_);
  or (_27049_, _27048_, _27046_);
  and (_27050_, _27049_, _26797_);
  or (_27051_, _27050_, _02892_);
  or (_27052_, _04982_, _02893_);
  and (_27053_, _27052_, _02537_);
  and (_27054_, _27053_, _27051_);
  nor (_27055_, _12395_, _02537_);
  or (_27057_, _27055_, _02940_);
  or (_27058_, _27057_, _27054_);
  or (_27059_, _23226_, _09217_);
  or (_27060_, _26807_, _09915_);
  and (_27061_, _27060_, _27059_);
  or (_27062_, _27061_, _03164_);
  and (_27063_, _27062_, _27058_);
  or (_27064_, _27063_, _09942_);
  or (_27065_, _26794_, _09941_);
  and (_27066_, _27065_, _27064_);
  or (_27068_, _27066_, _03163_);
  nand (_27069_, _12395_, _03163_);
  and (_27070_, _27069_, _09948_);
  and (_27071_, _27070_, _27068_);
  nor (_27072_, _26795_, _09948_);
  or (_27073_, _27072_, _02939_);
  or (_27074_, _27073_, _27071_);
  nand (_27075_, _02939_, _03629_);
  and (_27076_, _27075_, _02526_);
  and (_27077_, _27076_, _27074_);
  and (_27078_, _09101_, _02525_);
  or (_27079_, _27078_, _02497_);
  or (_27080_, _27079_, _27077_);
  or (_27081_, _27061_, _02498_);
  and (_27082_, _27081_, _25099_);
  and (_27083_, _27082_, _27080_);
  and (_27084_, _26794_, _09964_);
  or (_27085_, _27084_, _02888_);
  or (_27086_, _27085_, _27083_);
  nand (_27087_, _12395_, _02888_);
  and (_27090_, _27087_, _09044_);
  and (_27091_, _27090_, _27086_);
  nor (_27092_, _26795_, _09044_);
  or (_27093_, _27092_, _02937_);
  or (_27094_, _27093_, _27091_);
  nand (_27095_, _02937_, _03629_);
  and (_27096_, _27095_, _02524_);
  and (_27097_, _27096_, _27094_);
  and (_27098_, _09101_, _02523_);
  or (_27099_, _27098_, _09979_);
  or (_27101_, _27099_, _27097_);
  and (_27102_, _27101_, _26796_);
  or (_27103_, _27102_, _42672_);
  or (_27104_, _42668_, \oc8051_golden_model_1.PC [12]);
  and (_27105_, _27104_, _43998_);
  and (_43508_, _27105_, _27103_);
  and (_27106_, _09046_, _09092_);
  and (_27107_, _27106_, \oc8051_golden_model_1.PC [12]);
  nor (_27108_, _27107_, _09090_);
  and (_27109_, _27107_, _09090_);
  or (_27111_, _27109_, _27108_);
  or (_27112_, _27111_, _09063_);
  or (_27113_, _27111_, _09066_);
  or (_27114_, _09097_, _09070_);
  and (_27115_, _27114_, _23200_);
  or (_27116_, _27111_, _09074_);
  or (_27117_, _09097_, _09077_);
  and (_27118_, _27117_, _22667_);
  or (_27119_, _27111_, _09081_);
  or (_27120_, _27111_, _09657_);
  or (_27122_, _09097_, _05753_);
  or (_27123_, _27111_, _09200_);
  or (_27124_, _09097_, _02857_);
  and (_27125_, _27124_, _02838_);
  or (_27126_, _09215_, _09214_);
  nand (_27127_, _27126_, _09315_);
  or (_27128_, _27126_, _09315_);
  and (_27129_, _27128_, _27127_);
  or (_27130_, _27129_, _09528_);
  nand (_27131_, _09528_, _09213_);
  and (_27133_, _27131_, _02952_);
  and (_27134_, _27133_, _27130_);
  nand (_27135_, _09392_, _09213_);
  or (_27136_, _27129_, _09392_);
  and (_27137_, _27136_, _09481_);
  and (_27138_, _27137_, _27135_);
  and (_27139_, _09097_, _03075_);
  or (_27140_, _09402_, _09097_);
  nand (_27141_, _09213_, _09412_);
  or (_27142_, _27129_, _09412_);
  and (_27144_, _27142_, _02974_);
  and (_27145_, _27144_, _27141_);
  or (_27146_, _09099_, _09098_);
  nand (_27147_, _27146_, _09185_);
  or (_27148_, _27146_, _09185_);
  and (_27149_, _27148_, _27147_);
  and (_27150_, _27149_, _24086_);
  and (_27151_, _09420_, _09097_);
  or (_27152_, _27151_, _05362_);
  or (_27153_, _27152_, _27150_);
  or (_27155_, _27111_, _09432_);
  or (_27156_, _09444_, _09097_);
  or (_27157_, _03072_, \oc8051_golden_model_1.PC [13]);
  nor (_27158_, _27157_, _09435_);
  nand (_27159_, _27158_, _09430_);
  and (_27160_, _27159_, _27156_);
  or (_27161_, _27160_, _07646_);
  and (_27162_, _27161_, _02616_);
  and (_27163_, _27162_, _27155_);
  not (_27164_, _09097_);
  or (_27166_, _27164_, _02616_);
  nand (_27167_, _27166_, _05362_);
  or (_27168_, _27167_, _27163_);
  and (_27169_, _27168_, _09449_);
  and (_27170_, _27169_, _27153_);
  or (_27171_, _27170_, _27145_);
  and (_27172_, _27171_, _09405_);
  not (_27173_, _27111_);
  nor (_27174_, _27173_, _09456_);
  or (_27175_, _27174_, _26555_);
  or (_27177_, _27175_, _27172_);
  and (_27178_, _27177_, _27140_);
  or (_27179_, _27178_, _09461_);
  nand (_27180_, _27173_, _09461_);
  and (_27181_, _27180_, _03084_);
  and (_27182_, _27181_, _27179_);
  or (_27183_, _27182_, _27139_);
  and (_27184_, _27183_, _09470_);
  or (_27185_, _27173_, _09470_);
  nand (_27186_, _27185_, _09476_);
  or (_27187_, _27186_, _27184_);
  or (_27188_, _09476_, _09097_);
  and (_27189_, _27188_, _09396_);
  and (_27190_, _27189_, _27187_);
  or (_27191_, _27190_, _27138_);
  and (_27192_, _27191_, _02979_);
  nand (_27193_, _09357_, _09213_);
  or (_27194_, _27129_, _09357_);
  and (_27195_, _27194_, _02978_);
  and (_27196_, _27195_, _27193_);
  or (_27199_, _27196_, _02950_);
  or (_27200_, _27199_, _27192_);
  and (_27201_, _09514_, _09212_);
  and (_27202_, _27129_, _23031_);
  or (_27203_, _27202_, _09500_);
  or (_27204_, _27203_, _27201_);
  and (_27205_, _27204_, _09531_);
  and (_27206_, _27205_, _27200_);
  or (_27207_, _27206_, _27134_);
  and (_27208_, _27207_, _09490_);
  nand (_27210_, _27111_, _09489_);
  nand (_27211_, _27210_, _09498_);
  or (_27212_, _27211_, _27208_);
  or (_27213_, _09498_, _09097_);
  and (_27214_, _27213_, _09543_);
  and (_27215_, _27214_, _27212_);
  nor (_27216_, _27173_, _09543_);
  or (_27217_, _27216_, _09554_);
  or (_27218_, _27217_, _27215_);
  or (_27219_, _09553_, _09097_);
  and (_27221_, _27219_, _09557_);
  and (_27222_, _27221_, _27218_);
  nor (_27223_, _27173_, _09557_);
  or (_27224_, _27223_, _09562_);
  or (_27225_, _27224_, _27222_);
  or (_27226_, _09097_, _09561_);
  and (_27227_, _27226_, _02605_);
  and (_27228_, _27227_, _27225_);
  nand (_27229_, _27111_, _02583_);
  nand (_27230_, _27229_, _09572_);
  or (_27232_, _27230_, _27228_);
  or (_27233_, _09572_, _09097_);
  and (_27234_, _27233_, _08209_);
  and (_27235_, _27234_, _27232_);
  nand (_27236_, _09212_, _02981_);
  nand (_27237_, _27236_, _02857_);
  or (_27238_, _27237_, _27235_);
  and (_27239_, _27238_, _27125_);
  nand (_27240_, _09212_, _02579_);
  nand (_27241_, _27240_, _09200_);
  or (_27243_, _27241_, _27239_);
  and (_27244_, _27243_, _27123_);
  or (_27245_, _27244_, _09592_);
  or (_27246_, _09591_, _09097_);
  and (_27247_, _27246_, _09599_);
  and (_27248_, _27247_, _27245_);
  and (_27249_, _27149_, _09594_);
  or (_27250_, _27249_, _05754_);
  or (_27251_, _27250_, _27248_);
  and (_27252_, _27251_, _27122_);
  or (_27254_, _27252_, _02802_);
  nand (_27255_, _09213_, _02802_);
  and (_27256_, _27255_, _07860_);
  and (_27257_, _27256_, _27254_);
  and (_27258_, _09097_, _07859_);
  or (_27259_, _27258_, _27257_);
  and (_27260_, _27259_, _22679_);
  nor (_27261_, _09642_, \oc8051_golden_model_1.DPH [5]);
  nor (_27262_, _27261_, _09643_);
  and (_27263_, _27262_, _09611_);
  or (_27265_, _27263_, _09650_);
  or (_27266_, _27265_, _27260_);
  or (_27267_, _09649_, _09097_);
  and (_27268_, _27267_, _22678_);
  and (_27269_, _27268_, _27266_);
  or (_27270_, _27149_, _08165_);
  or (_27271_, _09097_, _09676_);
  and (_27272_, _27271_, _09083_);
  and (_27273_, _27272_, _27270_);
  or (_27274_, _27273_, _23884_);
  or (_27276_, _27274_, _27269_);
  and (_27277_, _27276_, _27120_);
  or (_27278_, _27277_, _09661_);
  or (_27279_, _09660_, _09097_);
  and (_27280_, _27279_, _03887_);
  and (_27281_, _27280_, _27278_);
  nand (_27282_, _09212_, _02980_);
  nand (_27283_, _27282_, _09668_);
  or (_27284_, _27283_, _27281_);
  or (_27285_, _09668_, _09097_);
  and (_27287_, _27285_, _22675_);
  and (_27288_, _27287_, _27284_);
  or (_27289_, _27149_, _09676_);
  or (_27290_, _09097_, _08165_);
  and (_27291_, _27290_, _09672_);
  and (_27292_, _27291_, _27289_);
  or (_27293_, _27292_, _09681_);
  or (_27294_, _27293_, _27288_);
  and (_27295_, _27294_, _27119_);
  or (_27296_, _27295_, _22930_);
  or (_27298_, _09097_, _09080_);
  and (_27299_, _27298_, _03883_);
  and (_27300_, _27299_, _27296_);
  nand (_27301_, _09212_, _02970_);
  nand (_27302_, _27301_, _09077_);
  or (_27303_, _27302_, _27300_);
  and (_27304_, _27303_, _27118_);
  or (_27305_, _27149_, \oc8051_golden_model_1.PSW [7]);
  or (_27306_, _09097_, _07293_);
  and (_27307_, _27306_, _09076_);
  and (_27309_, _27307_, _27305_);
  or (_27310_, _27309_, _09694_);
  or (_27311_, _27310_, _27304_);
  and (_27312_, _27311_, _27116_);
  or (_27313_, _27312_, _07944_);
  or (_27314_, _09097_, _07943_);
  and (_27315_, _27314_, _05783_);
  and (_27316_, _27315_, _27313_);
  nand (_27317_, _09212_, _02965_);
  nand (_27318_, _27317_, _09070_);
  or (_27320_, _27318_, _27316_);
  and (_27321_, _27320_, _27115_);
  or (_27322_, _27149_, _07293_);
  or (_27323_, _09097_, \oc8051_golden_model_1.PSW [7]);
  and (_27324_, _27323_, _09068_);
  and (_27325_, _27324_, _27322_);
  or (_27326_, _27325_, _09711_);
  or (_27327_, _27326_, _27321_);
  and (_27328_, _27327_, _27113_);
  or (_27329_, _27328_, _10365_);
  or (_27331_, _09097_, _09065_);
  and (_27332_, _27331_, _07992_);
  and (_27333_, _27332_, _27329_);
  and (_27334_, _27111_, _07991_);
  or (_27335_, _27334_, _03145_);
  or (_27336_, _27335_, _27333_);
  or (_27337_, _04877_, _09726_);
  and (_27338_, _27337_, _27336_);
  or (_27339_, _27338_, _03898_);
  nor (_27340_, _09097_, _02529_);
  nor (_27342_, _27340_, _02968_);
  and (_27343_, _27342_, _27339_);
  or (_27344_, _27129_, _23226_);
  or (_27345_, _09915_, _09212_);
  and (_27346_, _27345_, _02968_);
  and (_27347_, _27346_, _27344_);
  or (_27348_, _27347_, _25057_);
  or (_27349_, _27348_, _27343_);
  and (_27350_, _27349_, _27112_);
  or (_27351_, _27350_, _08067_);
  or (_27353_, _09097_, _08066_);
  and (_27354_, _27353_, _08112_);
  and (_27355_, _27354_, _27351_);
  and (_27356_, _27111_, _08111_);
  or (_27357_, _27356_, _02892_);
  or (_27358_, _27357_, _27355_);
  or (_27359_, _04877_, _02893_);
  and (_27360_, _27359_, _27358_);
  or (_27361_, _27360_, _22926_);
  nor (_27362_, _09097_, _02537_);
  nor (_27364_, _27362_, _02940_);
  and (_27365_, _27364_, _27361_);
  or (_27366_, _27129_, _09915_);
  nand (_27367_, _09915_, _09213_);
  and (_27368_, _27367_, _27366_);
  and (_27369_, _27368_, _02940_);
  or (_27370_, _27369_, _09942_);
  or (_27371_, _27370_, _27365_);
  or (_27372_, _27111_, _09941_);
  and (_27373_, _27372_, _03906_);
  and (_27375_, _27373_, _27371_);
  nand (_27376_, _09097_, _03163_);
  nand (_27377_, _27376_, _09948_);
  or (_27378_, _27377_, _27375_);
  or (_27379_, _27111_, _09948_);
  and (_27380_, _27379_, _06173_);
  and (_27381_, _27380_, _27378_);
  nor (_27382_, _03211_, _06173_);
  or (_27383_, _27382_, _02525_);
  or (_27384_, _27383_, _27381_);
  nand (_27386_, _27164_, _02525_);
  and (_27387_, _27386_, _02498_);
  and (_27388_, _27387_, _27384_);
  and (_27389_, _27368_, _02497_);
  or (_27390_, _27389_, _09964_);
  or (_27391_, _27390_, _27388_);
  nand (_27392_, _27173_, _09964_);
  and (_27393_, _27392_, _02890_);
  and (_27394_, _27393_, _27391_);
  nand (_27395_, _09097_, _02888_);
  nand (_27397_, _27395_, _09044_);
  or (_27398_, _27397_, _27394_);
  or (_27399_, _27111_, _09044_);
  and (_27400_, _27399_, _09043_);
  and (_27401_, _27400_, _27398_);
  nand (_27402_, _03211_, _02524_);
  and (_27403_, _27402_, _22655_);
  or (_27404_, _27403_, _27401_);
  nand (_27405_, _27164_, _02523_);
  and (_27406_, _27405_, _09983_);
  and (_27407_, _27406_, _27404_);
  and (_27408_, _27111_, _09979_);
  or (_27409_, _27408_, _27407_);
  or (_27410_, _27409_, _42672_);
  or (_27411_, _42668_, \oc8051_golden_model_1.PC [13]);
  and (_27412_, _27411_, _43998_);
  and (_43509_, _27412_, _27410_);
  nor (_27413_, _09050_, \oc8051_golden_model_1.PC [14]);
  nor (_27414_, _27413_, _09051_);
  not (_27415_, _27414_);
  nand (_27418_, _27415_, _08111_);
  nor (_27419_, _12800_, _09070_);
  nor (_27420_, _12800_, _09077_);
  nor (_27421_, _09668_, _12800_);
  nor (_27422_, _09649_, _12800_);
  or (_27423_, _09086_, _05753_);
  nor (_27424_, _09318_, _09210_);
  nor (_27425_, _27424_, _09319_);
  and (_27426_, _27425_, _23025_);
  and (_27427_, _09357_, _09207_);
  or (_27429_, _27427_, _27426_);
  and (_27430_, _27429_, _02978_);
  nor (_27431_, _27415_, _09470_);
  nand (_27432_, _27415_, _09461_);
  and (_27433_, _27425_, _24823_);
  and (_27434_, _09207_, _09412_);
  or (_27435_, _27434_, _03810_);
  or (_27436_, _27435_, _27433_);
  nor (_27437_, _09188_, _09089_);
  nor (_27438_, _27437_, _09189_);
  and (_27440_, _27438_, _24086_);
  and (_27441_, _09420_, _09086_);
  or (_27442_, _27441_, _05362_);
  or (_27443_, _27442_, _27440_);
  nor (_27444_, _27415_, _09432_);
  and (_27445_, _03387_, \oc8051_golden_model_1.PC [14]);
  and (_27446_, _27445_, _09434_);
  and (_27447_, _27446_, _22699_);
  and (_27448_, _27447_, _09430_);
  or (_27449_, _27448_, _27444_);
  and (_27451_, _27449_, _02616_);
  and (_27452_, _09445_, _09086_);
  or (_27453_, _27452_, _05363_);
  or (_27454_, _27453_, _27451_);
  and (_27455_, _27454_, _04265_);
  and (_27456_, _27455_, _27443_);
  and (_27457_, _27414_, _02886_);
  or (_27458_, _27457_, _02974_);
  or (_27459_, _27458_, _27456_);
  and (_27460_, _27459_, _27436_);
  or (_27462_, _27460_, _09406_);
  or (_27463_, _27414_, _09405_);
  and (_27464_, _27463_, _09402_);
  and (_27465_, _27464_, _27462_);
  nor (_27466_, _09402_, _12800_);
  or (_27467_, _27466_, _09461_);
  or (_27468_, _27467_, _27465_);
  and (_27469_, _27468_, _27432_);
  or (_27470_, _27469_, _03075_);
  nand (_27471_, _12800_, _03075_);
  and (_27473_, _27471_, _09470_);
  and (_27474_, _27473_, _27470_);
  or (_27475_, _27474_, _27431_);
  and (_27476_, _27475_, _09476_);
  or (_27477_, _09476_, _12800_);
  nand (_27478_, _27477_, _09396_);
  or (_27479_, _27478_, _27476_);
  and (_27480_, _09392_, _09207_);
  and (_27481_, _27425_, _26874_);
  or (_27482_, _27481_, _27480_);
  or (_27484_, _27482_, _09396_);
  and (_27485_, _27484_, _02979_);
  and (_27486_, _27485_, _27479_);
  or (_27487_, _27486_, _02950_);
  or (_27488_, _27487_, _27430_);
  and (_27489_, _27425_, _23031_);
  and (_27490_, _09514_, _09207_);
  or (_27491_, _27490_, _09500_);
  or (_27492_, _27491_, _27489_);
  and (_27493_, _27492_, _09531_);
  and (_27495_, _27493_, _27488_);
  or (_27496_, _27425_, _09528_);
  or (_27497_, _09529_, _09207_);
  and (_27498_, _27497_, _02952_);
  and (_27499_, _27498_, _27496_);
  or (_27500_, _27499_, _09489_);
  or (_27501_, _27500_, _27495_);
  nand (_27502_, _27415_, _09489_);
  and (_27503_, _27502_, _09498_);
  and (_27504_, _27503_, _27501_);
  nor (_27506_, _09498_, _12800_);
  or (_27507_, _27506_, _09544_);
  or (_27508_, _27507_, _27504_);
  or (_27509_, _27414_, _09543_);
  and (_27510_, _27509_, _09553_);
  and (_27511_, _27510_, _27508_);
  or (_27512_, _09553_, _12800_);
  nand (_27513_, _27512_, _09557_);
  or (_27514_, _27513_, _27511_);
  or (_27515_, _27414_, _09557_);
  and (_27517_, _27515_, _09561_);
  and (_27518_, _27517_, _27514_);
  nor (_27519_, _12800_, _09561_);
  or (_27520_, _27519_, _02583_);
  or (_27521_, _27520_, _27518_);
  nand (_27522_, _27415_, _02583_);
  and (_27523_, _27522_, _09572_);
  and (_27524_, _27523_, _27521_);
  nor (_27525_, _09572_, _12800_);
  or (_27526_, _27525_, _02981_);
  or (_27528_, _27526_, _27524_);
  or (_27529_, _09207_, _08209_);
  and (_27530_, _27529_, _02857_);
  and (_27531_, _27530_, _27528_);
  nor (_27532_, _12800_, _02857_);
  or (_27533_, _27532_, _02579_);
  or (_27534_, _27533_, _27531_);
  or (_27535_, _09207_, _02838_);
  and (_27536_, _27535_, _09200_);
  and (_27537_, _27536_, _27534_);
  nor (_27539_, _27415_, _09200_);
  or (_27540_, _27539_, _09592_);
  or (_27541_, _27540_, _27537_);
  or (_27542_, _09591_, _09086_);
  and (_27543_, _27542_, _09599_);
  and (_27544_, _27543_, _27541_);
  and (_27545_, _27438_, _09594_);
  or (_27546_, _27545_, _05754_);
  or (_27547_, _27546_, _27544_);
  and (_27548_, _27547_, _27423_);
  or (_27550_, _27548_, _02802_);
  or (_27551_, _09207_, _02803_);
  and (_27552_, _27551_, _07860_);
  and (_27553_, _27552_, _27550_);
  and (_27554_, _09086_, _07859_);
  or (_27555_, _27554_, _09611_);
  or (_27556_, _27555_, _27553_);
  nor (_27557_, _09643_, \oc8051_golden_model_1.DPH [6]);
  nor (_27558_, _27557_, _09644_);
  or (_27559_, _27558_, _22679_);
  and (_27561_, _27559_, _09649_);
  and (_27562_, _27561_, _27556_);
  or (_27563_, _27562_, _27422_);
  and (_27564_, _27563_, _22678_);
  or (_27565_, _27438_, _08165_);
  or (_27566_, _09086_, _09676_);
  and (_27567_, _27566_, _09083_);
  and (_27568_, _27567_, _27565_);
  or (_27569_, _27568_, _23884_);
  or (_27570_, _27569_, _27564_);
  or (_27572_, _27414_, _09657_);
  and (_27573_, _27572_, _09660_);
  and (_27574_, _27573_, _27570_);
  nor (_27575_, _09660_, _12800_);
  or (_27576_, _27575_, _02980_);
  or (_27577_, _27576_, _27574_);
  or (_27578_, _09207_, _03887_);
  and (_27579_, _27578_, _09668_);
  and (_27580_, _27579_, _27577_);
  or (_27581_, _27580_, _27421_);
  and (_27583_, _27581_, _22675_);
  or (_27584_, _27438_, _09676_);
  or (_27585_, _09086_, _08165_);
  and (_27586_, _27585_, _09672_);
  and (_27587_, _27586_, _27584_);
  or (_27588_, _27587_, _09681_);
  or (_27589_, _27588_, _27583_);
  or (_27590_, _27414_, _09081_);
  and (_27591_, _27590_, _09080_);
  and (_27592_, _27591_, _27589_);
  nor (_27594_, _12800_, _09080_);
  or (_27595_, _27594_, _02970_);
  or (_27596_, _27595_, _27592_);
  or (_27597_, _09207_, _03883_);
  and (_27598_, _27597_, _09077_);
  and (_27599_, _27598_, _27596_);
  or (_27600_, _27599_, _27420_);
  and (_27601_, _27600_, _22667_);
  or (_27602_, _27438_, \oc8051_golden_model_1.PSW [7]);
  or (_27603_, _09086_, _07293_);
  and (_27605_, _27603_, _09076_);
  and (_27606_, _27605_, _27602_);
  or (_27607_, _27606_, _09694_);
  or (_27608_, _27607_, _27601_);
  or (_27609_, _27414_, _09074_);
  and (_27610_, _27609_, _07943_);
  and (_27611_, _27610_, _27608_);
  nor (_27612_, _12800_, _07943_);
  or (_27613_, _27612_, _02965_);
  or (_27614_, _27613_, _27611_);
  or (_27616_, _09207_, _05783_);
  and (_27617_, _27616_, _09070_);
  and (_27618_, _27617_, _27614_);
  or (_27619_, _27618_, _27419_);
  and (_27620_, _27619_, _23200_);
  or (_27621_, _27438_, _07293_);
  or (_27622_, _09086_, \oc8051_golden_model_1.PSW [7]);
  and (_27623_, _27622_, _09068_);
  and (_27624_, _27623_, _27621_);
  or (_27625_, _27624_, _09711_);
  or (_27627_, _27625_, _27620_);
  or (_27628_, _27414_, _09066_);
  and (_27629_, _27628_, _09065_);
  and (_27630_, _27629_, _27627_);
  nor (_27631_, _12800_, _09065_);
  or (_27632_, _27631_, _07991_);
  or (_27633_, _27632_, _27630_);
  nand (_27634_, _27415_, _07991_);
  and (_27635_, _27634_, _09726_);
  and (_27636_, _27635_, _27633_);
  and (_27638_, _04770_, _03145_);
  or (_27639_, _27638_, _03898_);
  or (_27640_, _27639_, _27636_);
  nor (_27641_, _09086_, _02529_);
  nor (_27642_, _27641_, _02968_);
  and (_27643_, _27642_, _27640_);
  or (_27644_, _09915_, _09207_);
  or (_27645_, _27425_, _23226_);
  and (_27646_, _27645_, _02968_);
  and (_27647_, _27646_, _27644_);
  or (_27649_, _27647_, _25057_);
  or (_27650_, _27649_, _27643_);
  or (_27651_, _27414_, _09063_);
  and (_27652_, _27651_, _08066_);
  and (_27653_, _27652_, _27650_);
  nor (_27654_, _12800_, _08066_);
  or (_27655_, _27654_, _08111_);
  or (_27656_, _27655_, _27653_);
  and (_27657_, _27656_, _27418_);
  or (_27658_, _27657_, _02892_);
  or (_27660_, _04770_, _02893_);
  and (_27661_, _27660_, _02537_);
  and (_27662_, _27661_, _27658_);
  nor (_27663_, _12800_, _02537_);
  or (_27664_, _27663_, _02940_);
  or (_27665_, _27664_, _27662_);
  or (_27666_, _23226_, _09207_);
  or (_27667_, _27425_, _09915_);
  and (_27668_, _27667_, _27666_);
  or (_27669_, _27668_, _03164_);
  and (_27670_, _27669_, _27665_);
  or (_27671_, _27670_, _09942_);
  or (_27672_, _27414_, _09941_);
  and (_27673_, _27672_, _27671_);
  or (_27674_, _27673_, _03163_);
  nand (_27675_, _12800_, _03163_);
  and (_27676_, _27675_, _09948_);
  and (_27677_, _27676_, _27674_);
  nor (_27678_, _27415_, _09948_);
  or (_27679_, _27678_, _02939_);
  or (_27682_, _27679_, _27677_);
  nand (_27683_, _02939_, _02927_);
  and (_27684_, _27683_, _02526_);
  and (_27685_, _27684_, _27682_);
  and (_27686_, _09086_, _02525_);
  or (_27687_, _27686_, _02497_);
  or (_27688_, _27687_, _27685_);
  or (_27689_, _27668_, _02498_);
  and (_27690_, _27689_, _25099_);
  and (_27691_, _27690_, _27688_);
  and (_27693_, _27414_, _09964_);
  or (_27694_, _27693_, _02888_);
  or (_27695_, _27694_, _27691_);
  nand (_27696_, _12800_, _02888_);
  and (_27697_, _27696_, _09044_);
  and (_27698_, _27697_, _27695_);
  nor (_27699_, _27415_, _09044_);
  or (_27700_, _27699_, _02937_);
  or (_27701_, _27700_, _27698_);
  nand (_27702_, _02937_, _02927_);
  and (_27704_, _27702_, _27701_);
  or (_27705_, _27704_, _02523_);
  nand (_27706_, _12800_, _02523_);
  and (_27707_, _27706_, _09983_);
  and (_27708_, _27707_, _27705_);
  and (_27709_, _27414_, _09979_);
  or (_27710_, _27709_, _27708_);
  or (_27711_, _27710_, _42672_);
  or (_27712_, _42668_, \oc8051_golden_model_1.PC [14]);
  and (_27713_, _27712_, _43998_);
  and (_43510_, _27713_, _27711_);
  not (_27715_, \oc8051_golden_model_1.PSW [0]);
  nor (_27716_, _42668_, _27715_);
  not (_27717_, _09522_);
  nor (_27718_, _27717_, _08131_);
  and (_27719_, _14825_, _27717_);
  nor (_27720_, _27719_, _27718_);
  nor (_27721_, _27720_, _15160_);
  and (_27722_, _27720_, _15160_);
  or (_27723_, _27722_, _27721_);
  nor (_27725_, _27723_, _15502_);
  and (_27726_, _27723_, _15502_);
  nor (_27727_, _27726_, _27725_);
  nor (_27728_, _27727_, _15836_);
  and (_27729_, _27727_, _15836_);
  or (_27730_, _27729_, _27728_);
  or (_27731_, _27730_, _16171_);
  nand (_27732_, _27730_, _16171_);
  and (_27733_, _27732_, _27731_);
  nor (_27734_, _27733_, _16506_);
  and (_27736_, _27733_, _16506_);
  nor (_27737_, _27736_, _27734_);
  and (_27738_, _27737_, _08147_);
  nor (_27739_, _27737_, _08147_);
  or (_27740_, _27739_, _27738_);
  and (_27741_, _27740_, _08065_);
  nor (_27742_, _07578_, _07577_);
  nor (_27743_, _14897_, \oc8051_golden_model_1.ACC [3]);
  and (_27744_, _14897_, \oc8051_golden_model_1.ACC [3]);
  nor (_27745_, _27744_, _27743_);
  nor (_27747_, _06826_, _06824_);
  nor (_27748_, _27747_, \oc8051_golden_model_1.ACC [6]);
  and (_27749_, _27747_, \oc8051_golden_model_1.ACC [6]);
  nor (_27750_, _27749_, _27748_);
  and (_27751_, _27750_, _27745_);
  nor (_27752_, _27750_, _27745_);
  nor (_27753_, _27752_, _27751_);
  nor (_27754_, _27753_, _27742_);
  and (_27755_, _27753_, _27742_);
  or (_27756_, _27755_, _27754_);
  and (_27758_, _27756_, _07991_);
  nor (_27759_, _06906_, _06905_);
  nor (_27760_, _27759_, _06806_);
  and (_27761_, _27759_, _06806_);
  nor (_27762_, _27761_, _27760_);
  nor (_27763_, _27747_, _14835_);
  and (_27764_, _27747_, _14835_);
  nor (_27765_, _27764_, _27763_);
  and (_27766_, _27765_, _27762_);
  nor (_27767_, _27765_, _27762_);
  nor (_27769_, _27767_, _27766_);
  nor (_27770_, _27769_, _05771_);
  and (_27771_, _27769_, _05771_);
  nor (_27772_, _27771_, _27770_);
  nor (_27773_, _03062_, _04095_);
  or (_27774_, _27773_, _27772_);
  not (_27775_, _27772_);
  nor (_27776_, _27775_, _09470_);
  or (_27777_, _06032_, _06156_);
  nand (_27778_, _27777_, _11770_);
  or (_27780_, _27777_, _11770_);
  nand (_27781_, _27780_, _27778_);
  nor (_27782_, _06124_, _06160_);
  nand (_27783_, _27782_, _05849_);
  or (_27784_, _27782_, _05849_);
  nand (_27785_, _27784_, _27783_);
  nand (_27786_, _27785_, _27781_);
  or (_27787_, _27785_, _27781_);
  and (_27788_, _27787_, _27786_);
  nor (_27789_, _27788_, _05462_);
  and (_27791_, _27788_, _05462_);
  or (_27792_, _27791_, _27789_);
  or (_27793_, _27792_, _03840_);
  and (_27794_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_27795_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_27796_, _27795_, _27794_);
  and (_27797_, _27796_, _14608_);
  nor (_27798_, _27796_, _14608_);
  nor (_27799_, _27798_, _27797_);
  and (_27800_, _15584_, _15270_);
  and (_27802_, _15583_, _15271_);
  nor (_27803_, _27802_, _27800_);
  nor (_27804_, _27803_, _27799_);
  and (_27805_, _27803_, _27799_);
  nor (_27806_, _27805_, _27804_);
  and (_27807_, _27806_, _15949_);
  nor (_27808_, _27806_, _15949_);
  or (_27809_, _27808_, _27807_);
  nor (_27810_, _16280_, _07673_);
  and (_27811_, _16280_, _07673_);
  nor (_27813_, _27811_, _27810_);
  nor (_27814_, _27813_, _27809_);
  and (_27815_, _27813_, _27809_);
  nor (_27816_, _27815_, _27814_);
  and (_27817_, _27816_, _07649_);
  nor (_27818_, _27817_, _09404_);
  not (_27819_, _16272_);
  not (_27820_, _14370_);
  nor (_27821_, _14602_, _27820_);
  and (_27822_, _14602_, _27820_);
  nor (_27824_, _27822_, _27821_);
  and (_27825_, _27824_, _14890_);
  nor (_27826_, _27824_, _14890_);
  nor (_27827_, _27826_, _27825_);
  and (_27828_, _27827_, _15942_);
  nor (_27829_, _27827_, _15942_);
  or (_27830_, _27829_, _27828_);
  nor (_27831_, _15577_, _15262_);
  and (_27832_, _15577_, _15262_);
  nor (_27833_, _27832_, _27831_);
  and (_27835_, _27833_, _27830_);
  nor (_27836_, _27833_, _27830_);
  nor (_27837_, _27836_, _27835_);
  nor (_27838_, _27837_, _27819_);
  and (_27839_, _27837_, _27819_);
  or (_27840_, _27839_, _27838_);
  and (_27841_, _27840_, _07651_);
  nor (_27842_, _27840_, _07651_);
  or (_27843_, _27842_, _27841_);
  or (_27844_, _27843_, _03810_);
  nor (_27846_, _11584_, _04982_);
  and (_27847_, _11584_, _04982_);
  nor (_27848_, _27847_, _27846_);
  nor (_27849_, _05272_, _05240_);
  and (_27850_, _05246_, _12421_);
  nor (_27851_, _05246_, _12421_);
  nor (_27852_, _27851_, _27850_);
  nor (_27853_, _27852_, _27849_);
  and (_27854_, _27852_, _27849_);
  or (_27855_, _27854_, _27853_);
  nand (_27857_, _27855_, _27848_);
  or (_27858_, _27855_, _27848_);
  and (_27859_, _27858_, _27857_);
  and (_27860_, _27859_, _07633_);
  and (_27861_, _09434_, _09430_);
  nor (_27862_, _27861_, _27772_);
  and (_27863_, _27861_, _27715_);
  nor (_27864_, _27863_, _27862_);
  or (_27865_, _27864_, _03363_);
  and (_27866_, _27865_, _07635_);
  or (_27868_, _27866_, _27860_);
  or (_27869_, _27792_, _07631_);
  and (_27870_, _27869_, _27868_);
  or (_27871_, _27870_, _03072_);
  and (_27872_, _07517_, _07504_);
  nor (_27873_, _27872_, _07518_);
  and (_27874_, _27873_, _07442_);
  nor (_27875_, _27873_, _07442_);
  nor (_27876_, _27875_, _27874_);
  nor (_27877_, _07481_, _07424_);
  and (_27879_, _07481_, _07424_);
  nor (_27880_, _27879_, _27877_);
  not (_27881_, _27880_);
  and (_27882_, _07468_, _07453_);
  and (_27883_, _07467_, _07454_);
  nor (_27884_, _27883_, _27882_);
  and (_27885_, _27884_, _27881_);
  nor (_27886_, _27884_, _27881_);
  nor (_27887_, _27886_, _27885_);
  nor (_27888_, _27887_, _27876_);
  and (_27890_, _27887_, _27876_);
  nor (_27891_, _27890_, _27888_);
  nor (_27892_, _27891_, _10005_);
  and (_27893_, _27891_, _10005_);
  or (_27894_, _27893_, _27892_);
  or (_27895_, _27894_, _03387_);
  and (_27896_, _27895_, _09426_);
  and (_27897_, _27896_, _27871_);
  or (_27898_, _27897_, _25539_);
  or (_27899_, _27772_, _25538_);
  and (_27901_, _27899_, _04265_);
  and (_27902_, _27901_, _27898_);
  nor (_27903_, _27750_, \oc8051_golden_model_1.ACC [7]);
  and (_27904_, _27750_, \oc8051_golden_model_1.ACC [7]);
  nor (_27905_, _27904_, _27903_);
  or (_27906_, _27905_, _27781_);
  nand (_27907_, _27905_, _27781_);
  and (_27908_, _27907_, _27906_);
  and (_27909_, _27908_, _02886_);
  or (_27910_, _27909_, _02974_);
  or (_27912_, _27910_, _27902_);
  and (_27913_, _27912_, _27844_);
  or (_27914_, _27913_, _07649_);
  and (_27915_, _27914_, _27818_);
  and (_27916_, _27772_, _09404_);
  or (_27917_, _27916_, _27915_);
  and (_27918_, _27917_, _02881_);
  and (_27919_, _14615_, _14376_);
  nor (_27920_, _14615_, _14376_);
  or (_27921_, _27920_, _27919_);
  nor (_27923_, _16287_, _15590_);
  and (_27924_, _16287_, _15590_);
  nor (_27925_, _27924_, _27923_);
  nor (_27926_, _27925_, _27921_);
  and (_27927_, _27925_, _27921_);
  or (_27928_, _27927_, _27926_);
  not (_27929_, _15953_);
  nor (_27930_, _15276_, _14906_);
  and (_27931_, _15276_, _14906_);
  nor (_27932_, _27931_, _27930_);
  nor (_27934_, _27932_, _27929_);
  and (_27935_, _27932_, _27929_);
  nor (_27936_, _27935_, _27934_);
  and (_27937_, _27936_, _27928_);
  nor (_27938_, _27936_, _27928_);
  nor (_27939_, _27938_, _27937_);
  and (_27940_, _27939_, _07680_);
  nor (_27941_, _27939_, _07680_);
  or (_27942_, _27941_, _27940_);
  and (_27943_, _27942_, _02880_);
  or (_27945_, _27943_, _04252_);
  or (_27946_, _27945_, _27918_);
  or (_27947_, _27772_, _02609_);
  and (_27948_, _27947_, _27946_);
  or (_27949_, _27948_, _03069_);
  and (_27950_, _14577_, _14348_);
  nor (_27951_, _14577_, _14348_);
  nor (_27952_, _27951_, _27950_);
  not (_27953_, _27952_);
  not (_27954_, _15219_);
  and (_27955_, _27954_, _14871_);
  nor (_27956_, _27954_, _14871_);
  nor (_27957_, _27956_, _27955_);
  and (_27958_, _27957_, _27953_);
  nor (_27959_, _27957_, _27953_);
  nor (_27960_, _27959_, _27958_);
  and (_27961_, _27960_, _15558_);
  nor (_27962_, _27960_, _15558_);
  or (_27963_, _27962_, _27961_);
  and (_27964_, _27963_, _15887_);
  nor (_27966_, _27963_, _15887_);
  or (_27967_, _27966_, _27964_);
  and (_27968_, _27967_, _16223_);
  nor (_27969_, _27967_, _16223_);
  or (_27970_, _27969_, _27968_);
  and (_27971_, _27970_, _07402_);
  nor (_27972_, _27970_, _07402_);
  or (_27973_, _27972_, _27971_);
  or (_27974_, _27973_, _03336_);
  and (_27975_, _27974_, _07628_);
  and (_27977_, _27975_, _27949_);
  and (_27978_, _27859_, _07682_);
  or (_27979_, _27978_, _03399_);
  or (_27980_, _27979_, _27977_);
  and (_27981_, _27980_, _27793_);
  or (_27982_, _27981_, _03075_);
  or (_27983_, _27894_, _03084_);
  and (_27984_, _27983_, _09470_);
  and (_27985_, _27984_, _27982_);
  or (_27986_, _27985_, _27776_);
  and (_27988_, _27986_, _02877_);
  nor (_27989_, _14634_, _14346_);
  and (_27990_, _14634_, _14346_);
  nor (_27991_, _27990_, _27989_);
  nor (_27992_, _16307_, _07700_);
  and (_27993_, _16307_, _07700_);
  nor (_27994_, _27993_, _27992_);
  nor (_27995_, _27994_, _27991_);
  and (_27996_, _27994_, _27991_);
  nor (_27997_, _27996_, _27995_);
  not (_27999_, _15296_);
  and (_28000_, _27999_, _14926_);
  nor (_28001_, _27999_, _14926_);
  nor (_28002_, _28001_, _28000_);
  nor (_28003_, _15973_, _15610_);
  and (_28004_, _15973_, _15610_);
  nor (_28005_, _28004_, _28003_);
  nor (_28006_, _28005_, _28002_);
  and (_28007_, _28005_, _28002_);
  or (_28008_, _28007_, _28006_);
  nor (_28010_, _28008_, _27997_);
  and (_28011_, _28008_, _27997_);
  or (_28012_, _28011_, _28010_);
  nand (_28013_, _28012_, _02876_);
  nor (_28014_, _25499_, _02976_);
  nand (_28015_, _28014_, _28013_);
  or (_28016_, _28015_, _27988_);
  or (_28017_, _28014_, _27772_);
  nand (_28018_, _28017_, _28016_);
  and (_28019_, _02963_, _02949_);
  nand (_28021_, _28019_, _28018_);
  or (_28022_, _28019_, _27772_);
  nor (_28023_, _02978_, _02954_);
  and (_28024_, _28023_, _28022_);
  and (_28025_, _28024_, _28021_);
  or (_28026_, _28023_, _27775_);
  nand (_28027_, _28026_, _09491_);
  or (_28028_, _28027_, _28025_);
  or (_28029_, _27772_, _09491_);
  and (_28030_, _28029_, _02870_);
  and (_28032_, _28030_, _28028_);
  not (_28033_, _14931_);
  and (_28034_, _28033_, _14639_);
  nor (_28035_, _28033_, _14639_);
  nor (_28036_, _28035_, _28034_);
  and (_28037_, _28036_, _15924_);
  nor (_28038_, _28036_, _15924_);
  or (_28039_, _28038_, _28037_);
  nor (_28040_, _15243_, _27820_);
  and (_28041_, _15243_, _27820_);
  nor (_28043_, _28041_, _28040_);
  and (_28044_, _28043_, _15616_);
  nor (_28045_, _28043_, _15616_);
  nor (_28046_, _28045_, _28044_);
  nor (_28047_, _28046_, _28039_);
  and (_28048_, _28046_, _28039_);
  nor (_28049_, _28048_, _28047_);
  not (_28050_, _16312_);
  and (_28051_, _28050_, _07705_);
  nor (_28052_, _28050_, _07705_);
  nor (_28054_, _28052_, _28051_);
  nand (_28055_, _28054_, _28049_);
  or (_28056_, _28054_, _28049_);
  and (_28057_, _28056_, _02869_);
  nand (_28058_, _28057_, _28055_);
  nand (_28059_, _28058_, _27773_);
  or (_28060_, _28059_, _28032_);
  nand (_28061_, _28060_, _27774_);
  nor (_28062_, _03859_, _03059_);
  and (_28063_, _28062_, _09541_);
  nand (_28065_, _28063_, _28061_);
  or (_28066_, _28063_, _27772_);
  and (_28067_, _28066_, _06253_);
  and (_28068_, _28067_, _28065_);
  nor (_28069_, _03101_, _09551_);
  and (_28070_, _28069_, _08225_);
  nor (_28071_, _14645_, _14400_);
  and (_28072_, _14645_, _14400_);
  or (_28073_, _28072_, _28071_);
  nor (_28074_, _28073_, _14936_);
  and (_28076_, _28073_, _14936_);
  nor (_28077_, _28076_, _28074_);
  nor (_28078_, _28077_, _15304_);
  and (_28079_, _28077_, _15304_);
  or (_28080_, _28079_, _28078_);
  nor (_28081_, _28080_, _15621_);
  and (_28082_, _28080_, _15621_);
  or (_28083_, _28082_, _28081_);
  nor (_28084_, _28083_, _15981_);
  and (_28085_, _28083_, _15981_);
  or (_28087_, _28085_, _28084_);
  nor (_28088_, _28087_, _16318_);
  and (_28089_, _28087_, _16318_);
  or (_28090_, _28089_, _28088_);
  or (_28091_, _28090_, _07710_);
  nand (_28092_, _28090_, _07710_);
  and (_28093_, _28092_, _06247_);
  nand (_28094_, _28093_, _28091_);
  nand (_28095_, _28094_, _28070_);
  or (_28096_, _28095_, _28068_);
  or (_28098_, _28070_, _27772_);
  and (_28099_, _28098_, _10016_);
  and (_28100_, _28099_, _28096_);
  and (_28101_, _27772_, _03100_);
  or (_28102_, _28101_, _07716_);
  or (_28103_, _28102_, _28100_);
  not (_28104_, _15640_);
  not (_28105_, _07737_);
  and (_28106_, _14654_, _28105_);
  or (_28107_, _28106_, _07738_);
  nor (_28109_, _28107_, _14956_);
  and (_28110_, _28107_, _14956_);
  or (_28111_, _28110_, _28109_);
  nor (_28112_, _28111_, _15320_);
  and (_28113_, _28111_, _15320_);
  or (_28114_, _28113_, _28112_);
  and (_28115_, _28114_, _28104_);
  nor (_28116_, _28114_, _28104_);
  nor (_28117_, _28116_, _28115_);
  nor (_28118_, _28117_, _15998_);
  and (_28120_, _28117_, _15998_);
  nor (_28121_, _28120_, _28118_);
  nor (_28122_, _28121_, _16334_);
  and (_28123_, _28121_, _16334_);
  or (_28124_, _28123_, _28122_);
  and (_28125_, _28124_, _07747_);
  nor (_28126_, _28124_, _07747_);
  or (_28127_, _28126_, _28125_);
  nor (_28128_, _03711_, _03433_);
  and (_28129_, _28128_, _28127_);
  or (_28131_, _28129_, _07718_);
  and (_28132_, _28131_, _28103_);
  not (_28133_, _28128_);
  and (_28134_, _28133_, _28127_);
  or (_28135_, _28134_, _03434_);
  or (_28136_, _28135_, _28132_);
  not (_28137_, _07614_);
  and (_28138_, _14662_, _28137_);
  nor (_28139_, _28138_, _07615_);
  and (_28140_, _28139_, _14974_);
  nor (_28142_, _28139_, _14974_);
  or (_28143_, _28142_, _28140_);
  nor (_28144_, _28143_, _15237_);
  and (_28145_, _28143_, _15237_);
  nor (_28146_, _28145_, _28144_);
  or (_28147_, _28146_, _15658_);
  nand (_28148_, _28146_, _15658_);
  and (_28149_, _28148_, _28147_);
  or (_28150_, _28149_, _15918_);
  nand (_28151_, _28149_, _15918_);
  and (_28153_, _28151_, _28150_);
  nor (_28154_, _28153_, _16255_);
  and (_28155_, _28153_, _16255_);
  nor (_28156_, _28155_, _28154_);
  nor (_28157_, _28156_, _07624_);
  and (_28158_, _28156_, _07624_);
  or (_28159_, _28158_, _28157_);
  or (_28160_, _28159_, _07626_);
  and (_28161_, _28160_, _03111_);
  and (_28162_, _28161_, _28136_);
  or (_28164_, _07583_, _07573_);
  and (_28165_, _28164_, _07584_);
  and (_28166_, _28165_, _14988_);
  nor (_28167_, _28165_, _14988_);
  nor (_28168_, _28167_, _28166_);
  nor (_28169_, _28168_, _15334_);
  and (_28170_, _28168_, _15334_);
  or (_28171_, _28170_, _28169_);
  nor (_28172_, _28171_, _15671_);
  and (_28173_, _28171_, _15671_);
  or (_28175_, _28173_, _28172_);
  and (_28176_, _28175_, _16019_);
  nor (_28177_, _28175_, _16019_);
  or (_28178_, _28177_, _28176_);
  nor (_28179_, _28178_, _16239_);
  and (_28180_, _28178_, _16239_);
  or (_28181_, _28180_, _28179_);
  nor (_28182_, _28181_, _07596_);
  and (_28183_, _28181_, _07596_);
  or (_28184_, _28183_, _28182_);
  and (_28186_, _28184_, _03106_);
  or (_28187_, _28186_, _07404_);
  or (_28188_, _28187_, _28162_);
  not (_28189_, _15687_);
  not (_28190_, _07804_);
  and (_28191_, _14584_, _28190_);
  nor (_28192_, _14584_, _28190_);
  nor (_28193_, _28192_, _28191_);
  not (_28194_, _28193_);
  nor (_28195_, _28194_, _15004_);
  and (_28197_, _28194_, _15004_);
  nor (_28198_, _28197_, _28195_);
  and (_28199_, _28198_, _15350_);
  nor (_28200_, _28198_, _15350_);
  nor (_28201_, _28200_, _28199_);
  nand (_28202_, _28201_, _28189_);
  or (_28203_, _28201_, _28189_);
  and (_28204_, _28203_, _28202_);
  or (_28205_, _28204_, _15903_);
  nand (_28206_, _28204_, _15903_);
  and (_28208_, _28206_, _28205_);
  nor (_28209_, _28208_, _16352_);
  and (_28210_, _28208_, _16352_);
  nor (_28211_, _28210_, _28209_);
  and (_28212_, _28211_, _07826_);
  nor (_28213_, _28211_, _07826_);
  or (_28214_, _28213_, _28212_);
  or (_28215_, _28214_, _07405_);
  and (_28216_, _28215_, _28188_);
  or (_28217_, _28216_, _02583_);
  nor (_28219_, _04606_, _02928_);
  nor (_28220_, _04639_, _04632_);
  nor (_28221_, _04653_, _04619_);
  nor (_28222_, _04658_, _04626_);
  nor (_28223_, _28222_, _28221_);
  and (_28224_, _28222_, _28221_);
  nor (_28225_, _28224_, _28223_);
  nor (_28226_, _28225_, _28220_);
  and (_28227_, _28225_, _28220_);
  nor (_28228_, _28227_, _28226_);
  not (_28230_, _28228_);
  nor (_28231_, _28230_, _28219_);
  and (_28232_, _28230_, _28219_);
  or (_28233_, _28232_, _28231_);
  or (_28234_, _28233_, _02605_);
  and (_28235_, _28234_, _02864_);
  and (_28236_, _28235_, _28217_);
  not (_28237_, _07835_);
  and (_28238_, _14676_, _14421_);
  nor (_28239_, _14676_, _14421_);
  or (_28241_, _28239_, _28238_);
  nor (_28242_, _16360_, _15696_);
  and (_28243_, _16360_, _15696_);
  nor (_28244_, _28243_, _28242_);
  nor (_28245_, _28244_, _28241_);
  and (_28246_, _28244_, _28241_);
  or (_28247_, _28246_, _28245_);
  not (_28248_, _16030_);
  nor (_28249_, _15359_, _15013_);
  and (_28250_, _15359_, _15013_);
  nor (_28252_, _28250_, _28249_);
  nor (_28253_, _28252_, _28248_);
  and (_28254_, _28252_, _28248_);
  nor (_28255_, _28254_, _28253_);
  and (_28256_, _28255_, _28247_);
  nor (_28257_, _28255_, _28247_);
  nor (_28258_, _28257_, _28256_);
  nand (_28259_, _28258_, _28237_);
  or (_28260_, _28258_, _28237_);
  and (_28261_, _28260_, _02863_);
  and (_28263_, _28261_, _28259_);
  or (_28264_, _28263_, _25643_);
  or (_28265_, _28264_, _28236_);
  or (_28266_, _27772_, _25642_);
  nand (_28267_, _28266_, _28265_);
  and (_28268_, _04009_, _02517_);
  not (_28269_, _28268_);
  and (_28270_, _28269_, _02851_);
  nand (_28271_, _28270_, _28267_);
  nand (_28272_, _02855_, _02462_);
  or (_28274_, _28270_, _27973_);
  and (_28275_, _28274_, _28272_);
  and (_28276_, _28275_, _28271_);
  and (_28277_, _27973_, _03450_);
  or (_28278_, _28277_, _02853_);
  or (_28279_, _28278_, _28276_);
  and (_28280_, _14683_, _14428_);
  nor (_28281_, _14683_, _14428_);
  nor (_28282_, _28281_, _28280_);
  not (_28283_, _28282_);
  not (_28285_, _15367_);
  and (_28286_, _28285_, _15020_);
  nor (_28287_, _28285_, _15020_);
  nor (_28288_, _28287_, _28286_);
  and (_28289_, _28288_, _28283_);
  nor (_28290_, _28288_, _28283_);
  nor (_28291_, _28290_, _28289_);
  not (_28292_, _16038_);
  and (_28293_, _28292_, _15704_);
  nor (_28294_, _28292_, _15704_);
  nor (_28296_, _28294_, _28293_);
  nand (_28297_, _28296_, _16368_);
  or (_28298_, _28296_, _16368_);
  and (_28299_, _28298_, _28297_);
  nor (_28300_, _28299_, _28291_);
  and (_28301_, _28299_, _28291_);
  or (_28302_, _28301_, _28300_);
  nor (_28303_, _28302_, _07842_);
  and (_28304_, _28302_, _07842_);
  or (_28305_, _28304_, _05540_);
  or (_28307_, _28305_, _28303_);
  and (_28308_, _28307_, _02838_);
  and (_28309_, _28308_, _28279_);
  and (_28310_, _14689_, _14433_);
  nor (_28311_, _14689_, _14433_);
  nor (_28312_, _28311_, _28310_);
  not (_28313_, _15372_);
  and (_28314_, _28313_, _15026_);
  nor (_28315_, _28313_, _15026_);
  nor (_28316_, _28315_, _28314_);
  nor (_28318_, _28316_, _28312_);
  and (_28319_, _28316_, _28312_);
  or (_28320_, _28319_, _28318_);
  not (_28321_, _16044_);
  and (_28322_, _28321_, _15709_);
  nor (_28323_, _28321_, _15709_);
  nor (_28324_, _28323_, _28322_);
  not (_28325_, _16374_);
  and (_28326_, _28325_, _07848_);
  nor (_28327_, _28325_, _07848_);
  nor (_28329_, _28327_, _28326_);
  nor (_28330_, _28329_, _28324_);
  and (_28331_, _28329_, _28324_);
  nor (_28332_, _28331_, _28330_);
  or (_28333_, _28332_, _28320_);
  nand (_28334_, _28332_, _28320_);
  and (_28335_, _28334_, _02579_);
  and (_28336_, _28335_, _28333_);
  or (_28337_, _28336_, _06784_);
  or (_28338_, _28337_, _28309_);
  nor (_28340_, _06928_, _06877_);
  and (_28341_, _06928_, _06877_);
  nor (_28342_, _28341_, _28340_);
  not (_28343_, _28342_);
  and (_28344_, _28343_, _06984_);
  nor (_28345_, _28343_, _06984_);
  nor (_28346_, _28345_, _28344_);
  nor (_28347_, _28346_, _16380_);
  and (_28348_, _28346_, _16380_);
  nor (_28349_, _28348_, _28347_);
  nor (_28351_, _06844_, _07852_);
  and (_28352_, _06844_, _07852_);
  nor (_28353_, _28352_, _28351_);
  and (_28354_, _28353_, _28349_);
  nor (_28355_, _28353_, _28349_);
  or (_28356_, _28355_, _28354_);
  and (_28357_, _28356_, _07059_);
  nor (_28358_, _28356_, _07059_);
  nor (_28359_, _28358_, _28357_);
  not (_28360_, _28359_);
  nor (_28362_, _28360_, _07138_);
  and (_28363_, _28360_, _07138_);
  or (_28364_, _28363_, _06791_);
  or (_28365_, _28364_, _28362_);
  and (_28366_, _28365_, _02635_);
  and (_28367_, _28366_, _28338_);
  nand (_28368_, _28233_, _02546_);
  nor (_28369_, _09594_, _04146_);
  and (_28370_, _28369_, _09591_);
  nand (_28371_, _28370_, _28368_);
  or (_28373_, _28371_, _28367_);
  nor (_28374_, _28370_, _27772_);
  nor (_28375_, _28374_, _04145_);
  and (_28376_, _28375_, _28373_);
  nand (_28377_, _27772_, _04145_);
  nand (_28378_, _28377_, _04129_);
  or (_28379_, _28378_, _28376_);
  nor (_28380_, _27772_, _04129_);
  nor (_28381_, _28380_, _04102_);
  and (_28382_, _28381_, _28379_);
  nand (_28384_, _27772_, _04102_);
  nand (_28385_, _28384_, _05750_);
  or (_28386_, _28385_, _28382_);
  or (_28387_, _27772_, _05750_);
  and (_28388_, _28387_, _02803_);
  and (_28389_, _28388_, _28386_);
  nor (_28390_, _15384_, _15038_);
  and (_28391_, _15384_, _15038_);
  nor (_28392_, _28391_, _28390_);
  nor (_28393_, _14701_, _14444_);
  and (_28394_, _14701_, _14444_);
  or (_28395_, _28394_, _28393_);
  nor (_28396_, _28395_, _28392_);
  and (_28397_, _28395_, _28392_);
  nor (_28398_, _28397_, _28396_);
  not (_28399_, _16389_);
  nor (_28400_, _16056_, _15548_);
  and (_28401_, _16056_, _15548_);
  nor (_28402_, _28401_, _28400_);
  nor (_28403_, _28402_, _28399_);
  and (_28406_, _28402_, _28399_);
  nor (_28407_, _28406_, _28403_);
  nor (_28408_, _28407_, _28398_);
  and (_28409_, _28407_, _28398_);
  or (_28410_, _28409_, _28408_);
  nand (_28411_, _28410_, _07862_);
  or (_28412_, _28410_, _07862_);
  and (_28413_, _28412_, _02802_);
  and (_28414_, _28413_, _28411_);
  or (_28415_, _28414_, _28389_);
  and (_28417_, _28415_, _07860_);
  nand (_28418_, _28233_, _07859_);
  and (_28419_, _09649_, _22679_);
  nand (_28420_, _28419_, _28418_);
  or (_28421_, _28420_, _28417_);
  or (_28422_, _28419_, _27772_);
  and (_28423_, _28422_, _22678_);
  and (_28424_, _28423_, _28421_);
  and (_28425_, _27772_, _09083_);
  or (_28426_, _28425_, _07869_);
  or (_28428_, _28426_, _28424_);
  not (_28429_, _07194_);
  and (_28430_, _28429_, _07191_);
  nor (_28431_, _28429_, _07191_);
  nor (_28432_, _28431_, _28430_);
  and (_28433_, _14339_, _07212_);
  nor (_28434_, _28433_, _14949_);
  and (_28435_, _15201_, _07208_);
  nor (_28436_, _15201_, _07208_);
  nor (_28437_, _28436_, _28435_);
  nor (_28439_, _28437_, _28434_);
  and (_28440_, _28437_, _28434_);
  nor (_28441_, _28440_, _28439_);
  and (_28442_, _07201_, _07197_);
  nor (_28443_, _07201_, _07197_);
  nor (_28444_, _28443_, _28442_);
  nor (_28445_, _28444_, _28441_);
  and (_28446_, _28444_, _28441_);
  nor (_28447_, _28446_, _28445_);
  nor (_28448_, _28447_, _28432_);
  and (_28450_, _28447_, _28432_);
  or (_28451_, _28450_, _28448_);
  or (_28452_, _28451_, _07870_);
  and (_28453_, _28452_, _07868_);
  and (_28454_, _28453_, _28428_);
  not (_28455_, _07868_);
  nand (_28456_, _28451_, _28455_);
  nand (_28457_, _28456_, _07874_);
  or (_28458_, _28457_, _28454_);
  or (_28459_, _28451_, _07874_);
  and (_28461_, _28459_, _16401_);
  and (_28462_, _28461_, _28458_);
  not (_28463_, _08027_);
  and (_28464_, _28463_, _07886_);
  nor (_28465_, _28463_, _07886_);
  nor (_28466_, _28465_, _28464_);
  and (_28467_, _14455_, _08045_);
  nor (_28468_, _28467_, _14969_);
  nor (_28469_, _15227_, _08041_);
  and (_28470_, _15227_, _08041_);
  nor (_28472_, _28470_, _28469_);
  nor (_28473_, _28472_, _28468_);
  and (_28474_, _28472_, _28468_);
  nor (_28475_, _28474_, _28473_);
  nor (_28476_, _08030_, _08034_);
  and (_28477_, _08030_, _08034_);
  nor (_28478_, _28477_, _28476_);
  nor (_28479_, _28478_, _28475_);
  and (_28480_, _28478_, _28475_);
  nor (_28481_, _28480_, _28479_);
  nor (_28483_, _28481_, _28466_);
  and (_28484_, _28481_, _28466_);
  or (_28485_, _28484_, _28483_);
  and (_28486_, _28485_, _16400_);
  or (_28487_, _28486_, _03504_);
  or (_28488_, _28487_, _28462_);
  or (_28489_, _28485_, _15555_);
  and (_28490_, _28489_, _07890_);
  and (_28491_, _28490_, _28488_);
  not (_28492_, _12613_);
  and (_28494_, _28492_, _05774_);
  nor (_28495_, _28492_, _05774_);
  nor (_28496_, _28495_, _28494_);
  nor (_28497_, _11715_, _11522_);
  and (_28498_, _11715_, _11522_);
  nor (_28499_, _28498_, _28497_);
  not (_28500_, _11927_);
  nor (_28501_, _12133_, _28500_);
  and (_28502_, _12133_, _28500_);
  nor (_28503_, _28502_, _28501_);
  nor (_28505_, _28503_, _28499_);
  and (_28506_, _28503_, _28499_);
  nor (_28507_, _28506_, _28505_);
  or (_28508_, _28507_, _12207_);
  nand (_28509_, _28507_, _12207_);
  and (_28510_, _28509_, _28508_);
  nor (_28511_, _28510_, _12411_);
  and (_28512_, _28510_, _12411_);
  or (_28513_, _28512_, _28511_);
  and (_28514_, _28513_, _28496_);
  nor (_28516_, _28513_, _28496_);
  or (_28517_, _28516_, _28514_);
  and (_28518_, _28517_, _03129_);
  or (_28519_, _28518_, _07399_);
  or (_28520_, _28519_, _28491_);
  and (_28521_, _08116_, _07896_);
  nor (_28522_, _28521_, _09526_);
  and (_28523_, _27717_, _08131_);
  nor (_28524_, _28523_, _27718_);
  nor (_28525_, _28524_, _14996_);
  and (_28526_, _28524_, _14996_);
  nor (_28527_, _28526_, _28525_);
  and (_28528_, _08123_, _09519_);
  nor (_28529_, _08123_, _09519_);
  or (_28530_, _28529_, _28528_);
  nor (_28531_, _28530_, _08120_);
  and (_28532_, _28530_, _08120_);
  nor (_28533_, _28532_, _28531_);
  nor (_28534_, _28533_, _28527_);
  and (_28535_, _28533_, _28527_);
  nor (_28537_, _28535_, _28534_);
  or (_28538_, _28537_, _28522_);
  nand (_28539_, _28537_, _28522_);
  and (_28540_, _28539_, _28538_);
  or (_28541_, _28540_, _07897_);
  and (_28542_, _28541_, _03887_);
  and (_28543_, _28542_, _28520_);
  and (_28544_, _14734_, _14466_);
  nor (_28545_, _14734_, _14466_);
  nor (_28546_, _28545_, _28544_);
  not (_28548_, _28546_);
  not (_28549_, _15216_);
  and (_28550_, _28549_, _15066_);
  nor (_28551_, _28549_, _15066_);
  nor (_28552_, _28551_, _28550_);
  and (_28553_, _28552_, _28548_);
  nor (_28554_, _28552_, _28548_);
  or (_28555_, _28554_, _28553_);
  nor (_28556_, _16219_, _15883_);
  and (_28557_, _16219_, _15883_);
  nor (_28559_, _28557_, _28556_);
  not (_28560_, _15553_);
  and (_28561_, _28560_, _07902_);
  nor (_28562_, _28560_, _07902_);
  nor (_28563_, _28562_, _28561_);
  nor (_28564_, _28563_, _28559_);
  and (_28565_, _28563_, _28559_);
  nor (_28566_, _28565_, _28564_);
  nand (_28567_, _28566_, _28555_);
  or (_28568_, _28566_, _28555_);
  and (_28570_, _28568_, _02980_);
  and (_28571_, _28570_, _28567_);
  or (_28572_, _28571_, _28543_);
  and (_28573_, _28572_, _03128_);
  nand (_28574_, _27772_, _03127_);
  nor (_28575_, _28574_, _04706_);
  or (_28576_, _28575_, _26362_);
  or (_28577_, _28576_, _28573_);
  not (_28578_, _14470_);
  and (_28579_, _14477_, _28578_);
  or (_28580_, _27772_, _26361_);
  and (_28581_, _28580_, _28579_);
  and (_28582_, _28581_, _28577_);
  not (_28583_, _28579_);
  or (_28584_, _07213_, _07210_);
  nand (_28585_, _07213_, _07210_);
  and (_28586_, _28585_, _28584_);
  and (_28587_, _14862_, _07204_);
  and (_28588_, _07206_, _07205_);
  nor (_28589_, _28588_, _28587_);
  and (_28592_, _28589_, _28586_);
  nor (_28593_, _28589_, _28586_);
  nor (_28594_, _28593_, _28592_);
  not (_28595_, _07195_);
  nor (_28596_, _07199_, _07192_);
  and (_28597_, _07199_, _07192_);
  nor (_28598_, _28597_, _28596_);
  nor (_28599_, _28598_, _28595_);
  and (_28600_, _28598_, _28595_);
  nor (_28601_, _28600_, _28599_);
  and (_28603_, _28601_, _28594_);
  nor (_28604_, _28601_, _28594_);
  or (_28605_, _28604_, _28603_);
  and (_28606_, _28605_, _07190_);
  nor (_28607_, _28605_, _07190_);
  or (_28608_, _28607_, _28606_);
  nand (_28609_, _28608_, _28583_);
  nand (_28610_, _28609_, _14475_);
  or (_28611_, _28610_, _28582_);
  or (_28612_, _28608_, _14475_);
  and (_28614_, _28612_, _07912_);
  and (_28615_, _28614_, _28611_);
  or (_28616_, _08046_, _08043_);
  nand (_28617_, _08046_, _08043_);
  and (_28618_, _28617_, _28616_);
  and (_28619_, _08038_, _08039_);
  nor (_28620_, _08038_, _08039_);
  nor (_28621_, _28620_, _28619_);
  not (_28622_, _28621_);
  and (_28623_, _28622_, _28618_);
  nor (_28625_, _28622_, _28618_);
  nor (_28626_, _28625_, _28623_);
  not (_28627_, _08028_);
  nor (_28628_, _08032_, _08025_);
  and (_28629_, _08032_, _08025_);
  nor (_28630_, _28629_, _28628_);
  nor (_28631_, _28630_, _28627_);
  and (_28632_, _28630_, _28627_);
  nor (_28633_, _28632_, _28631_);
  not (_28634_, _28633_);
  nor (_28636_, _28634_, _28626_);
  and (_28637_, _28634_, _28626_);
  or (_28638_, _28637_, _28636_);
  and (_28639_, _28638_, _07885_);
  nor (_28640_, _28638_, _07885_);
  or (_28641_, _28640_, _28639_);
  and (_28642_, _28641_, _07911_);
  or (_28643_, _28642_, _03138_);
  or (_28644_, _28643_, _28615_);
  nor (_28645_, _11587_, _11521_);
  and (_28647_, _11587_, _11521_);
  nor (_28648_, _28647_, _28645_);
  not (_28649_, _12131_);
  and (_28650_, _28649_, _11925_);
  nor (_28651_, _28649_, _11925_);
  nor (_28652_, _28651_, _28650_);
  and (_28653_, _28652_, _28648_);
  nor (_28654_, _28652_, _28648_);
  nor (_28655_, _28654_, _28653_);
  not (_28656_, _12611_);
  nor (_28658_, _12409_, _12205_);
  and (_28659_, _12409_, _12205_);
  nor (_28660_, _28659_, _28658_);
  nor (_28661_, _28660_, _28656_);
  and (_28662_, _28660_, _28656_);
  nor (_28663_, _28662_, _28661_);
  and (_28664_, _28663_, _28655_);
  nor (_28665_, _28663_, _28655_);
  or (_28666_, _28665_, _28664_);
  nor (_28667_, _28666_, _05772_);
  and (_28669_, _28666_, _05772_);
  or (_28670_, _28669_, _28667_);
  or (_28671_, _28670_, _07396_);
  and (_28672_, _28671_, _07395_);
  and (_28673_, _28672_, _28644_);
  not (_28674_, _08126_);
  or (_28675_, _08132_, _08129_);
  nand (_28676_, _08132_, _08129_);
  and (_28677_, _28676_, _28675_);
  nand (_28678_, _28677_, _28674_);
  or (_28680_, _28677_, _28674_);
  and (_28681_, _28680_, _28678_);
  nor (_28682_, _28681_, _08124_);
  and (_28683_, _28681_, _08124_);
  or (_28684_, _28683_, _28682_);
  and (_28685_, _08114_, _07895_);
  nor (_28686_, _28685_, _10404_);
  nor (_28687_, _08117_, _08121_);
  and (_28688_, _08117_, _08121_);
  nor (_28689_, _28688_, _28687_);
  nor (_28691_, _28689_, _28686_);
  and (_28692_, _28689_, _28686_);
  or (_28693_, _28692_, _28691_);
  nor (_28694_, _28693_, _28684_);
  and (_28695_, _28693_, _28684_);
  or (_28696_, _28695_, _28694_);
  and (_28697_, _28696_, _07394_);
  or (_28698_, _28697_, _28673_);
  and (_28699_, _28698_, _03883_);
  and (_28700_, _09077_, _22667_);
  nor (_28702_, _15088_, _14494_);
  and (_28703_, _15088_, _14494_);
  nor (_28704_, _28703_, _28702_);
  nor (_28705_, _16437_, _15550_);
  and (_28706_, _16437_, _15550_);
  nor (_28707_, _28706_, _28705_);
  and (_28708_, _28707_, _28704_);
  nor (_28709_, _28707_, _28704_);
  nor (_28710_, _28709_, _28708_);
  nor (_28711_, _15430_, _14755_);
  and (_28713_, _15430_, _14755_);
  nor (_28714_, _28713_, _28711_);
  nor (_28715_, _16096_, _07923_);
  and (_28716_, _16096_, _07923_);
  nor (_28717_, _28716_, _28715_);
  and (_28718_, _28717_, _28714_);
  nor (_28719_, _28717_, _28714_);
  nor (_28720_, _28719_, _28718_);
  not (_28721_, _28720_);
  nand (_28722_, _28721_, _28710_);
  or (_28724_, _28721_, _28710_);
  and (_28725_, _28724_, _02970_);
  nand (_28726_, _28725_, _28722_);
  nand (_28727_, _28726_, _28700_);
  or (_28728_, _28727_, _28699_);
  or (_28729_, _27772_, _28700_);
  and (_28730_, _16102_, _15211_);
  and (_28731_, _28730_, _28729_);
  and (_28732_, _28731_, _28728_);
  nor (_28733_, _14338_, _07211_);
  and (_28735_, _14338_, _07211_);
  nor (_28736_, _28735_, _28733_);
  not (_28737_, _28736_);
  nor (_28738_, _07207_, _07203_);
  and (_28739_, _07207_, _07203_);
  nor (_28740_, _28739_, _28738_);
  nor (_28741_, _28740_, _28737_);
  and (_28742_, _28740_, _28737_);
  nor (_28743_, _28742_, _28741_);
  not (_28744_, _07196_);
  nor (_28746_, _07200_, _07193_);
  and (_28747_, _07200_, _07193_);
  nor (_28748_, _28747_, _28746_);
  nor (_28749_, _28748_, _28744_);
  and (_28750_, _28748_, _28744_);
  nor (_28751_, _28750_, _28749_);
  not (_28752_, _28751_);
  nor (_28753_, _28752_, _28743_);
  and (_28754_, _28752_, _28743_);
  or (_28755_, _28754_, _28753_);
  and (_28757_, _28755_, _07189_);
  nor (_28758_, _28755_, _07189_);
  nor (_28759_, _28758_, _28757_);
  nor (_28760_, _28759_, _28730_);
  or (_28761_, _28760_, _07935_);
  or (_28762_, _28761_, _28732_);
  nor (_28763_, _14454_, _08044_);
  and (_28764_, _14454_, _08044_);
  nor (_28765_, _28764_, _28763_);
  not (_28766_, _28765_);
  and (_28768_, _08036_, _08040_);
  nor (_28769_, _08036_, _08040_);
  nor (_28770_, _28769_, _28768_);
  nor (_28771_, _28770_, _28766_);
  and (_28772_, _28770_, _28766_);
  nor (_28773_, _28772_, _28771_);
  not (_28774_, _08029_);
  nor (_28775_, _08033_, _08026_);
  and (_28776_, _08033_, _08026_);
  nor (_28777_, _28776_, _28775_);
  nor (_28779_, _28777_, _28774_);
  and (_28780_, _28777_, _28774_);
  nor (_28781_, _28780_, _28779_);
  nor (_28782_, _28781_, _28773_);
  and (_28783_, _28781_, _28773_);
  nor (_28784_, _28783_, _28782_);
  and (_28785_, _28784_, _07884_);
  nor (_28786_, _28784_, _07884_);
  or (_28787_, _28786_, _28785_);
  or (_28788_, _28787_, _15441_);
  and (_28790_, _28788_, _03122_);
  and (_28791_, _28790_, _28762_);
  nor (_28792_, _11714_, _11520_);
  and (_28793_, _11714_, _11520_);
  nor (_28794_, _28793_, _28792_);
  and (_28795_, _28794_, _11926_);
  nor (_28796_, _28794_, _11926_);
  or (_28797_, _28796_, _28795_);
  nand (_28798_, _28797_, _12132_);
  or (_28799_, _28797_, _12132_);
  and (_28801_, _28799_, _28798_);
  nor (_28802_, _12410_, _12206_);
  and (_28803_, _12410_, _12206_);
  nor (_28804_, _28803_, _28802_);
  nor (_28805_, _28804_, _12612_);
  and (_28806_, _28804_, _12612_);
  nor (_28807_, _28806_, _28805_);
  not (_28808_, _28807_);
  nor (_28809_, _28808_, _28801_);
  and (_28810_, _28808_, _28801_);
  nor (_28813_, _28810_, _28809_);
  or (_28815_, _28813_, _05773_);
  nand (_28817_, _28813_, _05773_);
  and (_28819_, _28817_, _03121_);
  and (_28821_, _28819_, _28815_);
  or (_28823_, _28821_, _07942_);
  or (_28825_, _28823_, _28791_);
  nor (_28827_, _09521_, _08130_);
  and (_28829_, _09521_, _08130_);
  nor (_28831_, _28829_, _28827_);
  and (_28834_, _28831_, _08127_);
  nor (_28835_, _28831_, _08127_);
  or (_28836_, _28835_, _28834_);
  and (_28837_, _28836_, _08125_);
  nor (_28838_, _28836_, _08125_);
  or (_28839_, _28838_, _28837_);
  and (_28840_, _28839_, _08122_);
  nor (_28841_, _28839_, _08122_);
  or (_28842_, _28841_, _28840_);
  and (_28843_, _28842_, _08118_);
  nor (_28845_, _28842_, _08118_);
  or (_28846_, _28845_, _28843_);
  and (_28847_, _28846_, _08115_);
  nor (_28848_, _28846_, _08115_);
  or (_28849_, _28848_, _28847_);
  and (_28850_, _28849_, _07894_);
  nor (_28851_, _28849_, _07894_);
  or (_28852_, _28851_, _28850_);
  or (_28853_, _28852_, _07945_);
  and (_28854_, _28853_, _05783_);
  and (_28856_, _28854_, _28825_);
  and (_28857_, _09070_, _23200_);
  not (_28858_, _16462_);
  and (_28859_, _28858_, _07953_);
  nor (_28860_, _28858_, _07953_);
  nor (_28861_, _28860_, _28859_);
  not (_28862_, _16119_);
  and (_28863_, _28862_, _15792_);
  nor (_28864_, _28862_, _15792_);
  nor (_28865_, _28864_, _28863_);
  not (_28867_, _28865_);
  nor (_28868_, _14781_, _14515_);
  and (_28869_, _14781_, _14515_);
  or (_28870_, _28869_, _28868_);
  and (_28871_, _28870_, _15113_);
  nor (_28872_, _28870_, _15113_);
  or (_28873_, _28872_, _28871_);
  nand (_28874_, _28873_, _15456_);
  or (_28875_, _28873_, _15456_);
  and (_28876_, _28875_, _28874_);
  nor (_28878_, _28876_, _28867_);
  and (_28879_, _28876_, _28867_);
  nor (_28880_, _28879_, _28878_);
  nand (_28881_, _28880_, _28861_);
  or (_28882_, _28880_, _28861_);
  and (_28883_, _28882_, _02965_);
  nand (_28884_, _28883_, _28881_);
  nand (_28885_, _28884_, _28857_);
  or (_28886_, _28885_, _28856_);
  or (_28887_, _27772_, _28857_);
  and (_28889_, _28887_, _07320_);
  and (_28890_, _28889_, _28886_);
  not (_28891_, _07320_);
  nor (_28892_, _07737_, _07372_);
  nor (_28893_, _14787_, _28105_);
  nor (_28894_, _28893_, _28892_);
  nor (_28895_, _28894_, _15118_);
  and (_28896_, _28894_, _15118_);
  nor (_28897_, _28896_, _28895_);
  nor (_28898_, _28897_, _15465_);
  and (_28900_, _28897_, _15465_);
  or (_28901_, _28900_, _28898_);
  nor (_28902_, _28901_, _15797_);
  and (_28903_, _28901_, _15797_);
  or (_28904_, _28903_, _28902_);
  nor (_28905_, _28904_, _16129_);
  and (_28906_, _28904_, _16129_);
  or (_28907_, _28906_, _28905_);
  nor (_28908_, _28907_, _16467_);
  and (_28909_, _28907_, _16467_);
  or (_28911_, _28909_, _28908_);
  nand (_28912_, _28911_, _07391_);
  or (_28913_, _28911_, _07391_);
  and (_28914_, _28913_, _28912_);
  and (_28915_, _28914_, _28891_);
  or (_28916_, _28915_, _03543_);
  or (_28917_, _28916_, _28890_);
  or (_28918_, _28914_, _07317_);
  and (_28919_, _28918_, _16123_);
  and (_28920_, _28919_, _28917_);
  and (_28922_, _28914_, _16122_);
  or (_28923_, _28922_, _03546_);
  or (_28924_, _28923_, _28920_);
  or (_28925_, _28914_, _16127_);
  and (_28926_, _28925_, _28924_);
  or (_28927_, _28926_, _07240_);
  not (_28928_, _03549_);
  nor (_28929_, _07614_, _07292_);
  nor (_28930_, _14792_, _28137_);
  nor (_28931_, _28930_, _28929_);
  nor (_28933_, _28931_, _15124_);
  and (_28934_, _28931_, _15124_);
  nor (_28935_, _28934_, _28933_);
  nor (_28936_, _28935_, _15461_);
  and (_28937_, _28935_, _15461_);
  or (_28938_, _28937_, _28936_);
  nor (_28939_, _28938_, _15803_);
  and (_28940_, _28938_, _15803_);
  or (_28941_, _28940_, _28939_);
  nor (_28942_, _28941_, _16138_);
  and (_28944_, _28941_, _16138_);
  or (_28945_, _28944_, _28942_);
  nor (_28946_, _28945_, _16473_);
  and (_28947_, _28945_, _16473_);
  or (_28948_, _28947_, _28946_);
  nand (_28949_, _28948_, _07312_);
  or (_28950_, _28948_, _07312_);
  and (_28951_, _28950_, _28949_);
  or (_28952_, _28951_, _28928_);
  and (_28953_, _28952_, _03134_);
  nand (_28955_, _07240_, _02543_);
  or (_28956_, _28955_, _28951_);
  and (_28957_, _28956_, _28953_);
  and (_28958_, _28957_, _28927_);
  not (_28959_, _07987_);
  and (_28960_, _14798_, _07573_);
  nor (_28961_, _14798_, _07573_);
  nor (_28962_, _28961_, _28960_);
  nor (_28963_, _28962_, _15129_);
  and (_28964_, _28962_, _15129_);
  nor (_28966_, _28964_, _28963_);
  and (_28967_, _28966_, _15471_);
  nor (_28968_, _28966_, _15471_);
  or (_28969_, _28968_, _28967_);
  nor (_28970_, _28969_, _15808_);
  and (_28971_, _28969_, _15808_);
  or (_28972_, _28971_, _28970_);
  nor (_28973_, _28972_, _16144_);
  and (_28974_, _28972_, _16144_);
  or (_28975_, _28974_, _28973_);
  and (_28977_, _28975_, _16478_);
  nor (_28978_, _28975_, _16478_);
  nor (_28979_, _28978_, _28977_);
  nor (_28980_, _28979_, _28959_);
  and (_28981_, _28979_, _28959_);
  or (_28982_, _28981_, _07962_);
  or (_28983_, _28982_, _28980_);
  and (_28984_, _28983_, _10365_);
  or (_28985_, _28984_, _28958_);
  nor (_28986_, _07804_, _07798_);
  nor (_28988_, _14803_, _28190_);
  nor (_28989_, _28988_, _28986_);
  nor (_28990_, _28989_, _15135_);
  and (_28991_, _28989_, _15135_);
  nor (_28992_, _28991_, _28990_);
  nor (_28993_, _28992_, _15477_);
  and (_28994_, _28992_, _15477_);
  or (_28995_, _28994_, _28993_);
  nor (_28996_, _28995_, _15544_);
  and (_28997_, _28995_, _15544_);
  or (_28999_, _28997_, _28996_);
  nor (_29000_, _28999_, _16149_);
  and (_29001_, _28999_, _16149_);
  or (_29002_, _29001_, _29000_);
  nor (_29003_, _29002_, _16213_);
  and (_29004_, _29002_, _16213_);
  or (_29005_, _29004_, _29003_);
  nand (_29006_, _29005_, _08015_);
  or (_29007_, _29005_, _08015_);
  and (_29008_, _29007_, _29006_);
  or (_29010_, _29008_, _07993_);
  and (_29011_, _29010_, _07992_);
  and (_29012_, _29011_, _28985_);
  or (_29013_, _29012_, _27758_);
  nor (_29014_, _03145_, _03898_);
  and (_29015_, _29014_, _03561_);
  and (_29016_, _29015_, _29013_);
  or (_29017_, _29015_, _27775_);
  nand (_29018_, _29017_, _07238_);
  or (_29019_, _29018_, _29016_);
  not (_29021_, _14338_);
  and (_29022_, _29021_, _07212_);
  nor (_29023_, _29021_, _07212_);
  nor (_29024_, _29023_, _29022_);
  and (_29025_, _29024_, _15143_);
  nor (_29026_, _29024_, _15143_);
  nor (_29027_, _29026_, _29025_);
  and (_29028_, _29027_, _15204_);
  nor (_29029_, _29027_, _15204_);
  nor (_29030_, _29029_, _29028_);
  and (_29032_, _29030_, _15819_);
  nor (_29033_, _29030_, _15819_);
  nor (_29034_, _29033_, _29032_);
  nor (_29035_, _29034_, _15877_);
  and (_29036_, _29034_, _15877_);
  or (_29037_, _29036_, _29035_);
  nor (_29038_, _29037_, _16489_);
  and (_29039_, _29037_, _16489_);
  or (_29040_, _29039_, _29038_);
  nor (_29041_, _29040_, _07228_);
  and (_29043_, _29040_, _07228_);
  or (_29044_, _29043_, _29041_);
  or (_29045_, _29044_, _07238_);
  and (_29046_, _29045_, _08024_);
  and (_29047_, _29046_, _29019_);
  and (_29048_, _07188_, _02543_);
  not (_29049_, _14454_);
  and (_29050_, _29049_, _08045_);
  nor (_29051_, _29049_, _08045_);
  nor (_29052_, _29051_, _29050_);
  and (_29054_, _29052_, _15149_);
  nor (_29055_, _29052_, _15149_);
  nor (_29056_, _29055_, _29054_);
  and (_29057_, _29056_, _15489_);
  nor (_29058_, _29056_, _15489_);
  nor (_29059_, _29058_, _29057_);
  and (_29060_, _29059_, _15825_);
  nor (_29061_, _29059_, _15825_);
  nor (_29062_, _29061_, _29060_);
  nor (_29063_, _29062_, _16160_);
  and (_29065_, _29062_, _16160_);
  or (_29066_, _29065_, _29063_);
  and (_29067_, _29066_, _16495_);
  nor (_29068_, _29066_, _16495_);
  or (_29069_, _29068_, _29067_);
  and (_29070_, _29069_, _08061_);
  nor (_29071_, _29069_, _08061_);
  or (_29072_, _29071_, _29070_);
  and (_29073_, _29072_, _29048_);
  and (_29074_, _29072_, _23239_);
  or (_29076_, _29074_, _02894_);
  or (_29077_, _29076_, _29073_);
  or (_29078_, _29077_, _29047_);
  not (_29079_, _08107_);
  nor (_29080_, _09507_, _10193_);
  and (_29081_, _14820_, _09507_);
  nor (_29082_, _29081_, _29080_);
  nor (_29083_, _29082_, _15154_);
  and (_29084_, _29082_, _15154_);
  nor (_29085_, _29084_, _29083_);
  and (_29087_, _29085_, _15496_);
  nor (_29088_, _29085_, _15496_);
  nor (_29089_, _29088_, _29087_);
  nor (_29090_, _29089_, _15830_);
  and (_29091_, _29089_, _15830_);
  or (_29092_, _29091_, _29090_);
  nor (_29093_, _29092_, _16166_);
  and (_29094_, _29092_, _16166_);
  or (_29095_, _29094_, _29093_);
  nor (_29096_, _29095_, _16500_);
  and (_29098_, _29095_, _16500_);
  or (_29099_, _29098_, _29096_);
  nor (_29100_, _29099_, _29079_);
  and (_29101_, _29099_, _29079_);
  or (_29102_, _29101_, _29100_);
  or (_29103_, _29102_, _02896_);
  and (_29104_, _29103_, _08113_);
  and (_29105_, _29104_, _29078_);
  or (_29106_, _29105_, _27741_);
  nor (_29107_, _08111_, _02892_);
  and (_29109_, _26115_, _29107_);
  and (_29110_, _29109_, _29106_);
  or (_29111_, _29109_, _27775_);
  nand (_29112_, _29111_, _09941_);
  or (_29113_, _29112_, _29110_);
  or (_29114_, _27772_, _09941_);
  and (_29115_, _29114_, _03906_);
  and (_29116_, _29115_, _29113_);
  and (_29117_, _27843_, _03163_);
  or (_29118_, _29117_, _08154_);
  or (_29120_, _29118_, _29116_);
  not (_29121_, _08160_);
  and (_29122_, _14897_, _29121_);
  and (_29123_, _29122_, \oc8051_golden_model_1.ACC [3]);
  nor (_29124_, _29122_, \oc8051_golden_model_1.ACC [3]);
  nor (_29125_, _29124_, _29123_);
  and (_29126_, _29125_, _15849_);
  nor (_29127_, _29125_, _15849_);
  nor (_29128_, _29127_, _29126_);
  and (_29129_, _16182_, _06806_);
  nor (_29130_, _16182_, _06806_);
  nor (_29131_, _29130_, _29129_);
  nor (_29132_, _29131_, _29128_);
  and (_29133_, _29131_, _29128_);
  or (_29134_, _29133_, _29132_);
  nor (_29135_, _29134_, _08166_);
  and (_29136_, _29134_, _08166_);
  nor (_29137_, _29136_, _29135_);
  and (_29138_, _29137_, _08154_);
  nor (_29139_, _29138_, _08159_);
  and (_29142_, _29139_, _29120_);
  and (_29143_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_29144_, _29143_, _07670_);
  nand (_29145_, _29144_, _27753_);
  or (_29146_, _29144_, _27753_);
  and (_29147_, _29146_, _29145_);
  nand (_29148_, _29147_, _08159_);
  nand (_29149_, _29148_, _03915_);
  or (_29150_, _29149_, _29142_);
  or (_29151_, _27772_, _03915_);
  and (_29153_, _29151_, _02498_);
  and (_29154_, _29153_, _29150_);
  and (_29155_, _28012_, _02497_);
  or (_29156_, _29155_, _06142_);
  or (_29157_, _29156_, _29154_);
  nor (_29158_, _27772_, _06141_);
  nor (_29159_, _29158_, _04120_);
  and (_29160_, _29159_, _29157_);
  and (_29161_, _27772_, _04120_);
  or (_29162_, _29161_, _04118_);
  or (_29164_, _29162_, _29160_);
  or (_29165_, _27772_, _04117_);
  and (_29166_, _29165_, _02890_);
  and (_29167_, _29166_, _29164_);
  nor (_29168_, _14847_, _14370_);
  and (_29169_, _14847_, _14370_);
  nor (_29170_, _29169_, _29168_);
  and (_29171_, _29170_, _15184_);
  nor (_29172_, _29170_, _15184_);
  or (_29173_, _29172_, _29171_);
  and (_29175_, _29173_, _15526_);
  nor (_29176_, _29173_, _15526_);
  or (_29177_, _29176_, _29175_);
  and (_29178_, _29177_, _15861_);
  nor (_29179_, _29177_, _15861_);
  or (_29180_, _29179_, _29178_);
  and (_29181_, _29180_, _16195_);
  nor (_29182_, _29180_, _16195_);
  or (_29183_, _29182_, _29181_);
  and (_29184_, _29183_, _16529_);
  nor (_29186_, _29183_, _16529_);
  or (_29187_, _29186_, _29184_);
  and (_29188_, _29187_, _08179_);
  nor (_29189_, _29187_, _08179_);
  or (_29190_, _29189_, _29188_);
  and (_29191_, _29190_, _02888_);
  or (_29192_, _29191_, _08176_);
  or (_29193_, _29192_, _29167_);
  not (_29194_, _08184_);
  and (_29195_, _14897_, _29194_);
  and (_29197_, _29195_, _02564_);
  nor (_29198_, _29195_, _02564_);
  nor (_29199_, _29198_, _29197_);
  nor (_29200_, _29199_, _15866_);
  and (_29201_, _29199_, _15866_);
  or (_29202_, _29201_, _29200_);
  nor (_29203_, _29202_, _16534_);
  and (_29204_, _29202_, _16534_);
  or (_29205_, _29204_, _29203_);
  nor (_29206_, _16201_, _08191_);
  and (_29208_, _16201_, _08191_);
  nor (_29209_, _29208_, _29206_);
  nand (_29210_, _29209_, _29205_);
  or (_29211_, _29209_, _29205_);
  nand (_29212_, _29211_, _29210_);
  and (_29213_, _29212_, _08176_);
  nor (_29214_, _29213_, _08183_);
  and (_29215_, _29214_, _29193_);
  and (_29216_, _22654_, _09983_);
  nand (_29217_, _27772_, _08183_);
  nand (_29219_, _29217_, _29216_);
  or (_29220_, _29219_, _29215_);
  or (_29221_, _27772_, _29216_);
  and (_29222_, _29221_, _42668_);
  and (_29223_, _29222_, _29220_);
  or (_29224_, _29223_, _27716_);
  and (_43512_, _29224_, _43998_);
  nand (_29225_, _04690_, _03698_);
  or (_29226_, _04690_, \oc8051_golden_model_1.PSW [1]);
  and (_29227_, _29226_, _02802_);
  and (_29229_, _29227_, _29225_);
  nand (_29230_, _11695_, _04690_);
  and (_29231_, _29226_, _02579_);
  and (_29232_, _29231_, _29230_);
  not (_29233_, \oc8051_golden_model_1.PSW [1]);
  nor (_29234_, _04690_, _29233_);
  and (_29235_, _04690_, _04000_);
  or (_29236_, _29235_, _29234_);
  or (_29237_, _29236_, _03336_);
  and (_29238_, _11606_, _04690_);
  not (_29240_, _29238_);
  and (_29241_, _29240_, _29226_);
  or (_29242_, _29241_, _03810_);
  nand (_29243_, _04690_, _02551_);
  and (_29244_, _29243_, _29226_);
  and (_29245_, _29244_, _03813_);
  nor (_29246_, _03813_, _29233_);
  or (_29247_, _29246_, _02974_);
  or (_29248_, _29247_, _29245_);
  and (_29249_, _29248_, _02881_);
  and (_29251_, _29249_, _29242_);
  nor (_29252_, _05331_, _29233_);
  and (_29253_, _11592_, _05331_);
  or (_29254_, _29253_, _29252_);
  and (_29255_, _29254_, _02880_);
  or (_29256_, _29255_, _03069_);
  or (_29257_, _29256_, _29251_);
  and (_29258_, _29257_, _29237_);
  or (_29259_, _29258_, _03075_);
  or (_29260_, _29244_, _03084_);
  and (_29261_, _29260_, _02877_);
  and (_29262_, _29261_, _29259_);
  and (_29263_, _11595_, _05331_);
  or (_29264_, _29263_, _29252_);
  and (_29265_, _29264_, _02876_);
  or (_29266_, _29265_, _02869_);
  or (_29267_, _29266_, _29262_);
  and (_29268_, _29253_, _11591_);
  or (_29269_, _29252_, _02870_);
  or (_29270_, _29269_, _29268_);
  and (_29272_, _29270_, _29267_);
  and (_29273_, _29272_, _02864_);
  not (_29274_, _05331_);
  nor (_29275_, _11638_, _29274_);
  or (_29276_, _29252_, _29275_);
  and (_29277_, _29276_, _02863_);
  or (_29278_, _29277_, _06770_);
  or (_29279_, _29278_, _29273_);
  or (_29280_, _29236_, _05535_);
  and (_29281_, _29280_, _29279_);
  or (_29283_, _29281_, _02853_);
  and (_29284_, _04690_, _06151_);
  or (_29285_, _29234_, _05540_);
  or (_29286_, _29285_, _29284_);
  and (_29287_, _29286_, _02838_);
  and (_29288_, _29287_, _29283_);
  or (_29289_, _29288_, _29232_);
  and (_29290_, _29289_, _02803_);
  or (_29291_, _29290_, _29229_);
  and (_29292_, _29291_, _03887_);
  or (_29294_, _11710_, _09998_);
  and (_29295_, _29226_, _02980_);
  and (_29296_, _29295_, _29294_);
  or (_29297_, _29296_, _29292_);
  and (_29298_, _29297_, _03128_);
  or (_29299_, _11715_, _09998_);
  and (_29300_, _29226_, _03127_);
  and (_29301_, _29300_, _29299_);
  or (_29302_, _29301_, _29298_);
  and (_29303_, _29302_, _03883_);
  or (_29305_, _11709_, _09998_);
  and (_29306_, _29226_, _02970_);
  and (_29307_, _29306_, _29305_);
  or (_29308_, _29307_, _29303_);
  and (_29309_, _29308_, _03137_);
  or (_29310_, _29234_, _13722_);
  and (_29311_, _29244_, _03135_);
  and (_29312_, _29311_, _29310_);
  or (_29313_, _29312_, _29309_);
  and (_29314_, _29313_, _03124_);
  or (_29316_, _29225_, _13722_);
  and (_29317_, _29226_, _02965_);
  and (_29318_, _29317_, _29316_);
  or (_29319_, _29243_, _13722_);
  and (_29320_, _29226_, _03123_);
  and (_29321_, _29320_, _29319_);
  or (_29322_, _29321_, _03163_);
  or (_29323_, _29322_, _29318_);
  or (_29324_, _29323_, _29314_);
  or (_29325_, _29241_, _03906_);
  and (_29327_, _29325_, _02498_);
  and (_29328_, _29327_, _29324_);
  and (_29329_, _29264_, _02497_);
  or (_29330_, _29329_, _02888_);
  or (_29331_, _29330_, _29328_);
  or (_29332_, _29234_, _02890_);
  or (_29333_, _29332_, _29238_);
  and (_29334_, _29333_, _29331_);
  or (_29335_, _29334_, _42672_);
  or (_29336_, _42668_, \oc8051_golden_model_1.PSW [1]);
  and (_29338_, _29336_, _43998_);
  and (_43513_, _29338_, _29335_);
  and (_29339_, _07243_, \oc8051_golden_model_1.ACC [7]);
  nor (_29340_, _07243_, \oc8051_golden_model_1.ACC [7]);
  nor (_29341_, _29340_, _10359_);
  nor (_29342_, _29341_, _29339_);
  or (_29343_, _29342_, _07241_);
  nand (_29344_, _29343_, _07314_);
  and (_29345_, _29339_, _03134_);
  nand (_29346_, _29345_, _07309_);
  and (_29348_, _29346_, _29344_);
  not (_29349_, \oc8051_golden_model_1.PSW [2]);
  nor (_29350_, _04690_, _29349_);
  not (_29351_, _29350_);
  nand (_29352_, _11927_, _04690_);
  and (_29353_, _29352_, _29351_);
  or (_29354_, _29353_, _03128_);
  nand (_29355_, _04690_, _04435_);
  and (_29356_, _29355_, _29351_);
  and (_29357_, _29356_, _06770_);
  not (_29359_, _07747_);
  nor (_29360_, _07325_, \oc8051_golden_model_1.ACC [7]);
  and (_29361_, _07325_, \oc8051_golden_model_1.ACC [7]);
  nor (_29362_, _29361_, _29360_);
  and (_29363_, _29362_, _10265_);
  nor (_29364_, _29362_, _10265_);
  or (_29365_, _29364_, _29363_);
  nand (_29366_, _29365_, _29359_);
  or (_29367_, _29365_, _29359_);
  and (_29368_, _29367_, _10106_);
  and (_29370_, _29368_, _29366_);
  nor (_29371_, _05331_, _29349_);
  not (_29372_, _29371_);
  nand (_29373_, _11815_, _05331_);
  and (_29374_, _29373_, _29372_);
  and (_29375_, _29372_, _10028_);
  or (_29376_, _29375_, _02870_);
  or (_29377_, _29376_, _29374_);
  and (_29378_, _11797_, _05331_);
  nor (_29379_, _29378_, _29371_);
  or (_29381_, _29379_, _02877_);
  and (_29382_, _29356_, _03069_);
  nor (_29383_, _11801_, _09998_);
  nor (_29384_, _29383_, _29350_);
  and (_29385_, _29384_, _02974_);
  and (_29386_, _04690_, \oc8051_golden_model_1.ACC [2]);
  nor (_29387_, _29386_, _29350_);
  or (_29388_, _29387_, _03814_);
  or (_29389_, _03813_, _29349_);
  and (_29390_, _29389_, _03810_);
  and (_29392_, _29390_, _29388_);
  or (_29393_, _29392_, _02880_);
  or (_29394_, _29393_, _29385_);
  or (_29395_, _29374_, _02881_);
  and (_29396_, _29395_, _03336_);
  and (_29397_, _29396_, _29394_);
  or (_29398_, _29397_, _29382_);
  and (_29399_, _29398_, _03084_);
  and (_29400_, _29387_, _03075_);
  or (_29401_, _29400_, _02876_);
  or (_29403_, _29401_, _29399_);
  and (_29404_, _29403_, _29381_);
  or (_29405_, _29404_, _02869_);
  and (_29406_, _29405_, _29377_);
  or (_29407_, _29406_, _06247_);
  or (_29408_, _13672_, _13551_);
  or (_29409_, _29408_, _13793_);
  or (_29410_, _29409_, _13913_);
  or (_29411_, _29410_, _14030_);
  or (_29412_, _29411_, _14150_);
  or (_29414_, _29412_, _06766_);
  nor (_29415_, _29414_, _14267_);
  or (_29416_, _29415_, _06253_);
  and (_29417_, _29416_, _07718_);
  and (_29418_, _29417_, _29407_);
  or (_29419_, _29418_, _03434_);
  or (_29420_, _29419_, _29370_);
  not (_29421_, _07244_);
  and (_29422_, _10276_, _29421_);
  nor (_29423_, _10276_, _29421_);
  nor (_29425_, _29423_, _29422_);
  nor (_29426_, _29425_, _07621_);
  and (_29427_, _29425_, _07621_);
  or (_29428_, _29427_, _07626_);
  or (_29429_, _29428_, _29426_);
  and (_29430_, _29429_, _29420_);
  or (_29431_, _29430_, _03106_);
  nor (_29432_, _07521_, \oc8051_golden_model_1.ACC [7]);
  nor (_29433_, _07520_, _10397_);
  nor (_29434_, _29433_, _29432_);
  nor (_29436_, _29434_, _07526_);
  nor (_29437_, _10013_, _07522_);
  or (_29438_, _29437_, _29436_);
  and (_29439_, _29438_, _07593_);
  nor (_29440_, _29438_, _07593_);
  or (_29441_, _29440_, _03111_);
  or (_29442_, _29441_, _29439_);
  and (_29443_, _29442_, _07405_);
  and (_29444_, _29443_, _29431_);
  not (_29445_, _07759_);
  and (_29447_, _07823_, _29445_);
  nand (_29448_, _29447_, _10296_);
  or (_29449_, _29447_, _10296_);
  and (_29450_, _29449_, _29448_);
  and (_29451_, _29450_, _07404_);
  or (_29452_, _29451_, _02863_);
  or (_29453_, _29452_, _29444_);
  or (_29454_, _11848_, _29274_);
  and (_29455_, _29454_, _29372_);
  or (_29456_, _29455_, _02864_);
  and (_29458_, _29456_, _05535_);
  and (_29459_, _29458_, _29453_);
  or (_29460_, _29459_, _29357_);
  and (_29461_, _29460_, _05540_);
  or (_29462_, _09998_, _06031_);
  nor (_29463_, _29350_, _05540_);
  and (_29464_, _29463_, _29462_);
  or (_29465_, _29464_, _02579_);
  or (_29466_, _29465_, _29461_);
  or (_29467_, _11906_, _09998_);
  and (_29469_, _29467_, _29351_);
  or (_29470_, _29469_, _02838_);
  and (_29471_, _29470_, _06791_);
  and (_29472_, _29471_, _29466_);
  nand (_29473_, _06802_, _06825_);
  and (_29474_, _29473_, _06784_);
  or (_29475_, _29474_, _29472_);
  or (_29476_, _29475_, _02802_);
  and (_29477_, _04690_, _05701_);
  nor (_29478_, _29477_, _29350_);
  or (_29480_, _29478_, _02803_);
  and (_29481_, _29480_, _03887_);
  and (_29482_, _29481_, _29476_);
  nand (_29483_, _11921_, _04690_);
  nor (_29484_, _29350_, _03887_);
  and (_29485_, _29484_, _29483_);
  or (_29486_, _29485_, _03127_);
  or (_29487_, _29486_, _29482_);
  and (_29488_, _29487_, _29354_);
  or (_29489_, _29488_, _02970_);
  and (_29491_, _29351_, _05129_);
  or (_29492_, _29478_, _03883_);
  or (_29493_, _29492_, _29491_);
  and (_29494_, _29493_, _29489_);
  or (_29495_, _29494_, _03135_);
  or (_29496_, _29387_, _03137_);
  or (_29497_, _29496_, _29491_);
  and (_29498_, _29497_, _05783_);
  and (_29499_, _29498_, _29495_);
  or (_29500_, _11919_, _09998_);
  and (_29502_, _29500_, _29351_);
  and (_29503_, _29502_, _02965_);
  or (_29504_, _29503_, _29499_);
  and (_29505_, _29504_, _05788_);
  or (_29506_, _11926_, _09998_);
  nor (_29507_, _29350_, _05788_);
  nand (_29508_, _29507_, _29506_);
  nand (_29509_, _29508_, _07319_);
  or (_29510_, _29509_, _29505_);
  nor (_29511_, _29360_, _09991_);
  nor (_29513_, _29511_, _29361_);
  nand (_29514_, _29513_, _07391_);
  nand (_29515_, _29361_, _07388_);
  and (_29516_, _29515_, _29514_);
  or (_29517_, _29516_, _07319_);
  and (_29518_, _29517_, _07318_);
  and (_29519_, _29518_, _29510_);
  and (_29520_, _29516_, _03726_);
  or (_29521_, _29520_, _29519_);
  and (_29522_, _29521_, _07317_);
  and (_29524_, _29516_, _03543_);
  or (_29525_, _29524_, _29522_);
  and (_29526_, _29525_, _16123_);
  and (_29527_, _29516_, _16122_);
  or (_29528_, _29527_, _03546_);
  or (_29529_, _29528_, _29526_);
  or (_29530_, _29516_, _16127_);
  and (_29531_, _29530_, _07241_);
  and (_29532_, _29531_, _29529_);
  or (_29533_, _29532_, _29348_);
  nand (_29535_, _29433_, _07984_);
  nor (_29536_, _10366_, _07985_);
  and (_29537_, _29434_, _29536_);
  or (_29538_, _29433_, _28959_);
  or (_29539_, _29538_, _29537_);
  and (_29540_, _29539_, _29535_);
  or (_29541_, _29540_, _03134_);
  and (_29542_, _29541_, _29533_);
  and (_29543_, _29542_, _07993_);
  and (_29544_, _07758_, \oc8051_golden_model_1.ACC [7]);
  or (_29546_, _07758_, \oc8051_golden_model_1.ACC [7]);
  and (_29547_, _29546_, _10373_);
  or (_29548_, _29547_, _29544_);
  nor (_29549_, _29548_, _08015_);
  and (_29550_, _29548_, _08015_);
  or (_29551_, _29550_, _29549_);
  and (_29552_, _29551_, _07962_);
  or (_29553_, _29552_, _10378_);
  or (_29554_, _29553_, _29543_);
  nor (_29555_, _07225_, _07189_);
  not (_29557_, _10383_);
  or (_29558_, _29557_, _07224_);
  nand (_29559_, _29558_, _10378_);
  or (_29560_, _29559_, _29555_);
  and (_29561_, _29560_, _08024_);
  nand (_29562_, _29561_, _29554_);
  not (_29563_, _07884_);
  nor (_29564_, _08058_, _29563_);
  and (_29565_, _08058_, _07885_);
  or (_29566_, _29565_, _08024_);
  or (_29568_, _29566_, _29564_);
  and (_29569_, _29568_, _08066_);
  and (_29570_, _29569_, _29562_);
  nor (_29571_, _10398_, _02896_);
  or (_29572_, _08104_, _08068_);
  and (_29573_, _29572_, _29571_);
  or (_29574_, _08144_, _07894_);
  and (_29575_, _10406_, _08065_);
  and (_29576_, _29575_, _29574_);
  or (_29577_, _29576_, _03163_);
  or (_29579_, _29577_, _29573_);
  or (_29580_, _29579_, _29570_);
  nand (_29581_, _29384_, _03163_);
  and (_29582_, _29581_, _02498_);
  and (_29583_, _29582_, _29580_);
  nor (_29584_, _29379_, _02498_);
  or (_29585_, _29584_, _02888_);
  or (_29586_, _29585_, _29583_);
  and (_29587_, _11985_, _04690_);
  or (_29588_, _29350_, _02890_);
  or (_29590_, _29588_, _29587_);
  and (_29591_, _29590_, _29586_);
  or (_29592_, _29591_, _42672_);
  or (_29593_, _42668_, \oc8051_golden_model_1.PSW [2]);
  and (_29594_, _29593_, _43998_);
  and (_43514_, _29594_, _29592_);
  not (_29595_, \oc8051_golden_model_1.PSW [3]);
  nor (_29596_, _04690_, _29595_);
  and (_29597_, _12133_, _04690_);
  or (_29598_, _29597_, _29596_);
  and (_29600_, _29598_, _03127_);
  and (_29601_, _04690_, _04241_);
  or (_29602_, _29601_, _29596_);
  or (_29603_, _29602_, _05535_);
  nor (_29604_, _12017_, _09998_);
  or (_29605_, _29604_, _29596_);
  or (_29606_, _29605_, _03810_);
  and (_29607_, _04690_, \oc8051_golden_model_1.ACC [3]);
  or (_29608_, _29607_, _29596_);
  and (_29609_, _29608_, _03813_);
  nor (_29611_, _03813_, _29595_);
  or (_29612_, _29611_, _02974_);
  or (_29613_, _29612_, _29609_);
  and (_29614_, _29613_, _02881_);
  and (_29615_, _29614_, _29606_);
  nor (_29616_, _05331_, _29595_);
  and (_29617_, _12021_, _05331_);
  or (_29618_, _29617_, _29616_);
  and (_29619_, _29618_, _02880_);
  or (_29620_, _29619_, _03069_);
  or (_29622_, _29620_, _29615_);
  or (_29623_, _29602_, _03336_);
  and (_29624_, _29623_, _29622_);
  or (_29625_, _29624_, _03075_);
  or (_29626_, _29608_, _03084_);
  and (_29627_, _29626_, _02877_);
  and (_29628_, _29627_, _29625_);
  and (_29629_, _12005_, _05331_);
  or (_29630_, _29629_, _29616_);
  and (_29631_, _29630_, _02876_);
  or (_29633_, _29631_, _02869_);
  or (_29634_, _29633_, _29628_);
  or (_29635_, _29616_, _12036_);
  and (_29636_, _29635_, _29618_);
  or (_29637_, _29636_, _02870_);
  and (_29638_, _29637_, _02864_);
  and (_29639_, _29638_, _29634_);
  nor (_29640_, _12054_, _29274_);
  or (_29641_, _29640_, _29616_);
  and (_29642_, _29641_, _02863_);
  or (_29644_, _29642_, _06770_);
  or (_29645_, _29644_, _29639_);
  and (_29646_, _29645_, _29603_);
  or (_29647_, _29646_, _02853_);
  and (_29648_, _04690_, _06154_);
  or (_29649_, _29596_, _05540_);
  or (_29650_, _29649_, _29648_);
  and (_29651_, _29650_, _02838_);
  and (_29652_, _29651_, _29647_);
  nor (_29653_, _12112_, _09998_);
  or (_29655_, _29653_, _29596_);
  and (_29656_, _29655_, _02579_);
  or (_29657_, _29656_, _02802_);
  or (_29658_, _29657_, _29652_);
  and (_29659_, _04690_, _05658_);
  or (_29660_, _29659_, _29596_);
  or (_29661_, _29660_, _02803_);
  and (_29662_, _29661_, _29658_);
  or (_29663_, _29662_, _02980_);
  and (_29664_, _12127_, _04690_);
  or (_29666_, _29596_, _03887_);
  or (_29667_, _29666_, _29664_);
  and (_29668_, _29667_, _03128_);
  and (_29669_, _29668_, _29663_);
  or (_29670_, _29669_, _29600_);
  and (_29671_, _29670_, _03883_);
  or (_29672_, _29596_, _05079_);
  and (_29673_, _29660_, _02970_);
  and (_29674_, _29673_, _29672_);
  or (_29675_, _29674_, _29671_);
  and (_29676_, _29675_, _03137_);
  and (_29677_, _29608_, _03135_);
  and (_29678_, _29677_, _29672_);
  or (_29679_, _29678_, _02965_);
  or (_29680_, _29679_, _29676_);
  nor (_29681_, _12125_, _09998_);
  or (_29682_, _29596_, _05783_);
  or (_29683_, _29682_, _29681_);
  and (_29684_, _29683_, _05788_);
  and (_29685_, _29684_, _29680_);
  nor (_29688_, _12132_, _09998_);
  or (_29689_, _29688_, _29596_);
  and (_29690_, _29689_, _03123_);
  or (_29691_, _29690_, _03163_);
  or (_29692_, _29691_, _29685_);
  or (_29693_, _29605_, _03906_);
  and (_29694_, _29693_, _02498_);
  and (_29695_, _29694_, _29692_);
  and (_29696_, _29630_, _02497_);
  or (_29697_, _29696_, _02888_);
  or (_29699_, _29697_, _29695_);
  and (_29700_, _12183_, _04690_);
  or (_29701_, _29596_, _02890_);
  or (_29702_, _29701_, _29700_);
  and (_29703_, _29702_, _29699_);
  or (_29704_, _29703_, _42672_);
  or (_29705_, _42668_, \oc8051_golden_model_1.PSW [3]);
  and (_29706_, _29705_, _43998_);
  and (_43515_, _29706_, _29704_);
  not (_29707_, \oc8051_golden_model_1.PSW [4]);
  nor (_29709_, _04690_, _29707_);
  and (_29710_, _12207_, _04690_);
  nor (_29711_, _29710_, _29709_);
  nor (_29712_, _29711_, _03128_);
  and (_29713_, _04690_, _04982_);
  nor (_29714_, _29713_, _29709_);
  and (_29715_, _29714_, _06770_);
  nor (_29716_, _05331_, _29707_);
  and (_29717_, _12213_, _05331_);
  nor (_29718_, _29717_, _29716_);
  nor (_29720_, _29718_, _02877_);
  and (_29721_, _04690_, \oc8051_golden_model_1.ACC [4]);
  nor (_29722_, _29721_, _29709_);
  nor (_29723_, _29722_, _03814_);
  nor (_29724_, _03813_, _29707_);
  or (_29725_, _29724_, _29723_);
  and (_29726_, _29725_, _03810_);
  nor (_29727_, _12217_, _09998_);
  nor (_29728_, _29727_, _29709_);
  nor (_29729_, _29728_, _03810_);
  or (_29731_, _29729_, _29726_);
  and (_29732_, _29731_, _02881_);
  and (_29733_, _12231_, _05331_);
  nor (_29734_, _29733_, _29716_);
  nor (_29735_, _29734_, _02881_);
  or (_29736_, _29735_, _03069_);
  or (_29737_, _29736_, _29732_);
  nand (_29738_, _29714_, _03069_);
  and (_29739_, _29738_, _29737_);
  and (_29740_, _29739_, _03084_);
  nor (_29742_, _29722_, _03084_);
  or (_29743_, _29742_, _29740_);
  and (_29744_, _29743_, _02877_);
  nor (_29745_, _29744_, _29720_);
  nor (_29746_, _29745_, _02869_);
  and (_29747_, _12247_, _05331_);
  nor (_29748_, _29747_, _29716_);
  nor (_29749_, _29748_, _02870_);
  nor (_29750_, _29749_, _29746_);
  nor (_29751_, _29750_, _02863_);
  nor (_29753_, _12264_, _29274_);
  nor (_29754_, _29753_, _29716_);
  nor (_29755_, _29754_, _02864_);
  nor (_29756_, _29755_, _06770_);
  not (_29757_, _29756_);
  nor (_29758_, _29757_, _29751_);
  nor (_29759_, _29758_, _29715_);
  nor (_29760_, _29759_, _02853_);
  and (_29761_, _04690_, _06159_);
  nor (_29762_, _29709_, _05540_);
  not (_29764_, _29762_);
  nor (_29765_, _29764_, _29761_);
  nor (_29766_, _29765_, _02579_);
  not (_29767_, _29766_);
  nor (_29768_, _29767_, _29760_);
  nor (_29769_, _12321_, _09998_);
  nor (_29770_, _29769_, _29709_);
  nor (_29771_, _29770_, _02838_);
  or (_29772_, _29771_, _02802_);
  or (_29773_, _29772_, _29768_);
  and (_29775_, _05666_, _04690_);
  nor (_29776_, _29775_, _29709_);
  nand (_29777_, _29776_, _02802_);
  and (_29778_, _29777_, _29773_);
  and (_29779_, _29778_, _03887_);
  and (_29780_, _12211_, _04690_);
  nor (_29781_, _29780_, _29709_);
  nor (_29782_, _29781_, _03887_);
  or (_29783_, _29782_, _29779_);
  and (_29784_, _29783_, _03128_);
  nor (_29786_, _29784_, _29712_);
  nor (_29787_, _29786_, _02970_);
  nor (_29788_, _29709_, _05031_);
  not (_29789_, _29788_);
  nor (_29790_, _29776_, _03883_);
  and (_29791_, _29790_, _29789_);
  nor (_29792_, _29791_, _29787_);
  nor (_29793_, _29792_, _03135_);
  nor (_29794_, _29722_, _03137_);
  and (_29795_, _29794_, _29789_);
  or (_29797_, _29795_, _29793_);
  and (_29798_, _29797_, _05783_);
  nor (_29799_, _12209_, _09998_);
  nor (_29800_, _29799_, _29709_);
  nor (_29801_, _29800_, _05783_);
  or (_29802_, _29801_, _29798_);
  and (_29803_, _29802_, _05788_);
  nor (_29804_, _12206_, _09998_);
  nor (_29805_, _29804_, _29709_);
  nor (_29806_, _29805_, _05788_);
  or (_29808_, _29806_, _29803_);
  and (_29809_, _29808_, _03906_);
  nor (_29810_, _29728_, _03906_);
  or (_29811_, _29810_, _29809_);
  and (_29812_, _29811_, _02498_);
  nor (_29813_, _29718_, _02498_);
  or (_29814_, _29813_, _29812_);
  and (_29815_, _29814_, _02890_);
  and (_29816_, _12389_, _04690_);
  nor (_29817_, _29816_, _29709_);
  nor (_29819_, _29817_, _02890_);
  or (_29820_, _29819_, _29815_);
  or (_29821_, _29820_, _42672_);
  or (_29822_, _42668_, \oc8051_golden_model_1.PSW [4]);
  and (_29823_, _29822_, _43998_);
  and (_43516_, _29823_, _29821_);
  not (_29824_, \oc8051_golden_model_1.PSW [5]);
  nor (_29825_, _04690_, _29824_);
  and (_29826_, _12411_, _04690_);
  nor (_29827_, _29826_, _29825_);
  nor (_29829_, _29827_, _03128_);
  and (_29830_, _04690_, _06158_);
  or (_29831_, _29830_, _29825_);
  and (_29832_, _29831_, _02853_);
  nor (_29833_, _12407_, _09998_);
  nor (_29834_, _29833_, _29825_);
  and (_29835_, _29834_, _02974_);
  and (_29836_, _04690_, \oc8051_golden_model_1.ACC [5]);
  nor (_29837_, _29836_, _29825_);
  or (_29838_, _29837_, _03814_);
  or (_29840_, _03813_, _29824_);
  and (_29841_, _29840_, _03810_);
  and (_29842_, _29841_, _29838_);
  or (_29843_, _29842_, _02880_);
  nor (_29844_, _29843_, _29835_);
  nor (_29845_, _05331_, _29824_);
  and (_29846_, _12435_, _05331_);
  nor (_29847_, _29846_, _29845_);
  nor (_29848_, _29847_, _02881_);
  or (_29849_, _29848_, _03069_);
  or (_29851_, _29849_, _29844_);
  and (_29852_, _04690_, _04877_);
  nor (_29853_, _29852_, _29825_);
  nand (_29854_, _29853_, _03069_);
  and (_29855_, _29854_, _29851_);
  and (_29856_, _29855_, _03084_);
  nor (_29857_, _29837_, _03084_);
  or (_29858_, _29857_, _29856_);
  and (_29859_, _29858_, _02877_);
  and (_29860_, _12417_, _05331_);
  nor (_29862_, _29860_, _29845_);
  nor (_29863_, _29862_, _02877_);
  or (_29864_, _29863_, _02869_);
  or (_29865_, _29864_, _29859_);
  nor (_29866_, _29845_, _12450_);
  nor (_29867_, _29866_, _29847_);
  or (_29868_, _29867_, _02870_);
  and (_29869_, _29868_, _02864_);
  and (_29870_, _29869_, _29865_);
  nor (_29871_, _12468_, _29274_);
  nor (_29873_, _29871_, _29845_);
  nor (_29874_, _29873_, _02864_);
  nor (_29875_, _29874_, _06770_);
  not (_29876_, _29875_);
  nor (_29877_, _29876_, _29870_);
  and (_29878_, _29853_, _06770_);
  or (_29879_, _29878_, _02853_);
  nor (_29880_, _29879_, _29877_);
  or (_29881_, _29880_, _29832_);
  and (_29882_, _29881_, _02838_);
  nor (_29884_, _12527_, _09998_);
  nor (_29885_, _29884_, _29825_);
  nor (_29886_, _29885_, _02838_);
  or (_29887_, _29886_, _02802_);
  or (_29888_, _29887_, _29882_);
  and (_29889_, _05614_, _04690_);
  nor (_29890_, _29889_, _29825_);
  nand (_29891_, _29890_, _02802_);
  and (_29892_, _29891_, _29888_);
  and (_29893_, _29892_, _03887_);
  and (_29895_, _12415_, _04690_);
  nor (_29896_, _29895_, _29825_);
  nor (_29897_, _29896_, _03887_);
  or (_29898_, _29897_, _29893_);
  and (_29899_, _29898_, _03128_);
  nor (_29900_, _29899_, _29829_);
  nor (_29901_, _29900_, _02970_);
  nor (_29902_, _29825_, _04924_);
  not (_29903_, _29902_);
  nor (_29904_, _29890_, _03883_);
  and (_29906_, _29904_, _29903_);
  nor (_29907_, _29906_, _29901_);
  nor (_29908_, _29907_, _03135_);
  nor (_29909_, _29837_, _03137_);
  and (_29910_, _29909_, _29903_);
  or (_29911_, _29910_, _29908_);
  and (_29912_, _29911_, _05783_);
  nor (_29913_, _12413_, _09998_);
  nor (_29914_, _29913_, _29825_);
  nor (_29915_, _29914_, _05783_);
  or (_29917_, _29915_, _29912_);
  and (_29918_, _29917_, _05788_);
  nor (_29919_, _12410_, _09998_);
  nor (_29920_, _29919_, _29825_);
  nor (_29921_, _29920_, _05788_);
  or (_29922_, _29921_, _29918_);
  and (_29923_, _29922_, _03906_);
  nor (_29924_, _29834_, _03906_);
  or (_29925_, _29924_, _29923_);
  and (_29926_, _29925_, _02498_);
  nor (_29928_, _29862_, _02498_);
  or (_29929_, _29928_, _29926_);
  and (_29930_, _29929_, _02890_);
  and (_29931_, _12589_, _04690_);
  nor (_29932_, _29931_, _29825_);
  nor (_29933_, _29932_, _02890_);
  or (_29934_, _29933_, _29930_);
  or (_29935_, _29934_, _42672_);
  or (_29936_, _42668_, \oc8051_golden_model_1.PSW [5]);
  and (_29937_, _29936_, _43998_);
  and (_43517_, _29937_, _29935_);
  nor (_29938_, _07265_, _07241_);
  and (_29939_, _29938_, _07303_);
  nor (_29940_, _04690_, _15267_);
  not (_29941_, _29940_);
  nand (_29942_, _12613_, _04690_);
  and (_29943_, _29942_, _29941_);
  or (_29944_, _29943_, _03128_);
  nand (_29945_, _04690_, _04770_);
  and (_29946_, _29945_, _29941_);
  and (_29949_, _29946_, _06770_);
  nor (_29950_, _07816_, _07755_);
  or (_29951_, _29950_, _07405_);
  nor (_29952_, _07617_, _07265_);
  or (_29953_, _29952_, _07626_);
  nor (_29954_, _05331_, _15267_);
  and (_29955_, _12616_, _05331_);
  nor (_29956_, _29955_, _29954_);
  or (_29957_, _29956_, _02877_);
  nor (_29958_, _12603_, _09998_);
  nor (_29960_, _29958_, _29940_);
  and (_29961_, _29960_, _02974_);
  and (_29962_, _04690_, \oc8051_golden_model_1.ACC [6]);
  nor (_29963_, _29962_, _29940_);
  or (_29964_, _29963_, _03814_);
  or (_29965_, _03813_, _15267_);
  and (_29966_, _29965_, _03810_);
  and (_29967_, _29966_, _29964_);
  or (_29968_, _29967_, _02880_);
  or (_29969_, _29968_, _29961_);
  not (_29971_, _29954_);
  nand (_29972_, _12618_, _05331_);
  and (_29973_, _29972_, _29971_);
  or (_29974_, _29973_, _02881_);
  and (_29975_, _29974_, _03336_);
  and (_29976_, _29975_, _29969_);
  and (_29977_, _29946_, _03069_);
  or (_29978_, _29977_, _29976_);
  and (_29979_, _29978_, _03084_);
  and (_29980_, _29963_, _03075_);
  or (_29982_, _29980_, _02876_);
  or (_29983_, _29982_, _29979_);
  and (_29984_, _29983_, _29957_);
  or (_29985_, _29984_, _02869_);
  and (_29986_, _29971_, _10076_);
  or (_29987_, _29986_, _02870_);
  or (_29988_, _29987_, _29973_);
  and (_29989_, _29988_, _07718_);
  and (_29990_, _29989_, _29985_);
  or (_29991_, _07718_, _07345_);
  nor (_29993_, _29991_, _07740_);
  or (_29994_, _29993_, _03434_);
  or (_29995_, _29994_, _29990_);
  and (_29996_, _29995_, _03111_);
  and (_29997_, _29996_, _29953_);
  or (_29998_, _07485_, _03111_);
  nor (_29999_, _29998_, _07586_);
  or (_30000_, _29999_, _07404_);
  or (_30001_, _30000_, _29997_);
  and (_30002_, _30001_, _29951_);
  or (_30004_, _30002_, _02863_);
  or (_30005_, _12664_, _29274_);
  and (_30006_, _30005_, _29971_);
  or (_30007_, _30006_, _02864_);
  and (_30008_, _30007_, _05535_);
  and (_30009_, _30008_, _30004_);
  or (_30010_, _30009_, _29949_);
  and (_30011_, _30010_, _05540_);
  nand (_30012_, _04690_, _05849_);
  nor (_30013_, _29940_, _05540_);
  and (_30014_, _30013_, _30012_);
  or (_30015_, _30014_, _02579_);
  or (_30016_, _30015_, _30011_);
  or (_30017_, _12722_, _09998_);
  and (_30018_, _30017_, _29941_);
  or (_30019_, _30018_, _02838_);
  and (_30020_, _30019_, _02803_);
  and (_30021_, _30020_, _30016_);
  and (_30022_, _12729_, _04690_);
  nor (_30023_, _30022_, _29940_);
  and (_30025_, _30023_, _02802_);
  or (_30026_, _30025_, _30021_);
  and (_30027_, _30026_, _03887_);
  nand (_30028_, _12739_, _04690_);
  nor (_30029_, _29940_, _03887_);
  and (_30030_, _30029_, _30028_);
  or (_30031_, _30030_, _03127_);
  or (_30032_, _30031_, _30027_);
  and (_30033_, _30032_, _29944_);
  or (_30034_, _30033_, _02970_);
  and (_30036_, _29941_, _04818_);
  or (_30037_, _30023_, _03883_);
  or (_30038_, _30037_, _30036_);
  and (_30039_, _30038_, _30034_);
  or (_30040_, _30039_, _03135_);
  or (_30041_, _29963_, _03137_);
  or (_30042_, _30041_, _30036_);
  and (_30043_, _30042_, _05783_);
  and (_30044_, _30043_, _30040_);
  or (_30045_, _12737_, _09998_);
  and (_30047_, _30045_, _29941_);
  and (_30048_, _30047_, _02965_);
  or (_30049_, _30048_, _30044_);
  and (_30050_, _30049_, _05788_);
  or (_30051_, _12612_, _09998_);
  nor (_30052_, _29940_, _05788_);
  and (_30053_, _30052_, _30051_);
  or (_30054_, _30053_, _03312_);
  or (_30055_, _30054_, _30050_);
  and (_30056_, _02846_, _02967_);
  not (_30058_, _03312_);
  not (_30059_, _07345_);
  and (_30060_, _07382_, _30059_);
  nor (_30061_, _30060_, _30058_);
  nor (_30062_, _30061_, _30056_);
  and (_30063_, _30062_, _30055_);
  and (_30064_, _30060_, _30056_);
  or (_30065_, _30064_, _30063_);
  or (_30066_, _30065_, _03548_);
  not (_30067_, _03548_);
  or (_30069_, _30060_, _30067_);
  and (_30070_, _30069_, _30066_);
  or (_30071_, _30070_, _03726_);
  or (_30072_, _30060_, _07318_);
  and (_30073_, _30072_, _07317_);
  and (_30074_, _30073_, _30071_);
  and (_30075_, _30060_, _03543_);
  or (_30076_, _30075_, _07315_);
  or (_30077_, _30076_, _30074_);
  or (_30078_, _30060_, _07316_);
  and (_30080_, _30078_, _07241_);
  and (_30081_, _30080_, _30077_);
  or (_30082_, _30081_, _29939_);
  and (_30083_, _30082_, _03134_);
  nor (_30084_, _07485_, _03134_);
  and (_30085_, _30084_, _07978_);
  or (_30086_, _30085_, _07962_);
  or (_30087_, _30086_, _30083_);
  not (_30088_, _07755_);
  and (_30089_, _08006_, _30088_);
  or (_30091_, _30089_, _07993_);
  and (_30092_, _30091_, _07238_);
  and (_30093_, _30092_, _30087_);
  nor (_30094_, _07238_, _07219_);
  or (_30095_, _30094_, _07188_);
  or (_30096_, _30095_, _30093_);
  nand (_30097_, _08052_, _07188_);
  and (_30098_, _30097_, _02896_);
  and (_30099_, _30098_, _30096_);
  nor (_30100_, _08098_, _02896_);
  or (_30102_, _30100_, _08065_);
  nor (_30103_, _30102_, _30099_);
  and (_30104_, _08138_, _08065_);
  or (_30105_, _30104_, _30103_);
  and (_30106_, _30105_, _03906_);
  nor (_30107_, _29960_, _03906_);
  or (_30108_, _30107_, _30106_);
  and (_30109_, _30108_, _02498_);
  nor (_30110_, _29956_, _02498_);
  or (_30111_, _30110_, _30109_);
  and (_30113_, _30111_, _02890_);
  and (_30114_, _12794_, _04690_);
  nor (_30115_, _30114_, _29940_);
  nor (_30116_, _30115_, _02890_);
  or (_30117_, _30116_, _30113_);
  or (_30118_, _30117_, _42672_);
  or (_30119_, _42668_, \oc8051_golden_model_1.PSW [6]);
  and (_30120_, _30119_, _43998_);
  and (_43518_, _30120_, _30118_);
  not (_30121_, \oc8051_golden_model_1.PCON [0]);
  nor (_30123_, _04685_, _30121_);
  and (_30124_, _05226_, _04685_);
  nor (_30125_, _30124_, _30123_);
  and (_30126_, _30125_, _16625_);
  and (_30127_, _04685_, \oc8051_golden_model_1.ACC [0]);
  nor (_30128_, _30127_, _30123_);
  nor (_30129_, _30128_, _03084_);
  nor (_30130_, _30129_, _06770_);
  nor (_30131_, _30125_, _03810_);
  nor (_30132_, _03813_, _30121_);
  nor (_30134_, _30128_, _03814_);
  nor (_30135_, _30134_, _30132_);
  nor (_30136_, _30135_, _02974_);
  or (_30137_, _30136_, _03069_);
  nor (_30138_, _30137_, _30131_);
  or (_30139_, _30138_, _03075_);
  and (_30140_, _30139_, _30130_);
  and (_30141_, _04685_, _03808_);
  and (_30142_, _05535_, _03336_);
  or (_30143_, _30142_, _30123_);
  nor (_30145_, _30143_, _30141_);
  nor (_30146_, _30145_, _30140_);
  nor (_30147_, _30146_, _02853_);
  and (_30148_, _04685_, _06152_);
  nor (_30149_, _30123_, _05540_);
  not (_30150_, _30149_);
  nor (_30151_, _30150_, _30148_);
  nor (_30152_, _30151_, _30147_);
  and (_30153_, _30152_, _02838_);
  nor (_30154_, _11505_, _10462_);
  nor (_30156_, _30154_, _30123_);
  nor (_30157_, _30156_, _02838_);
  or (_30158_, _30157_, _30153_);
  and (_30159_, _30158_, _02803_);
  and (_30160_, _04685_, _05672_);
  nor (_30161_, _30160_, _30123_);
  nor (_30162_, _30161_, _02803_);
  or (_30163_, _30162_, _30159_);
  and (_30164_, _30163_, _03887_);
  and (_30165_, _11399_, _04685_);
  nor (_30167_, _30165_, _30123_);
  nor (_30168_, _30167_, _03887_);
  or (_30169_, _30168_, _30164_);
  and (_30170_, _30169_, _03128_);
  and (_30171_, _11522_, _04685_);
  nor (_30172_, _30171_, _30123_);
  nor (_30173_, _30172_, _03128_);
  or (_30174_, _30173_, _30170_);
  and (_30175_, _30174_, _03883_);
  or (_30176_, _30161_, _03883_);
  nor (_30178_, _30176_, _30124_);
  nor (_30179_, _30178_, _30175_);
  nor (_30180_, _30179_, _03135_);
  and (_30181_, _11521_, _04685_);
  or (_30182_, _30181_, _30123_);
  and (_30183_, _30182_, _03135_);
  or (_30184_, _30183_, _30180_);
  and (_30185_, _30184_, _05783_);
  nor (_30186_, _11396_, _10462_);
  nor (_30187_, _30186_, _30123_);
  nor (_30189_, _30187_, _05783_);
  or (_30190_, _30189_, _30185_);
  and (_30191_, _30190_, _05788_);
  nor (_30192_, _11520_, _10462_);
  nor (_30193_, _30192_, _30123_);
  nor (_30194_, _30193_, _05788_);
  nor (_30195_, _30194_, _16625_);
  not (_30196_, _30195_);
  nor (_30197_, _30196_, _30191_);
  nor (_30198_, _30197_, _30126_);
  or (_30200_, _30198_, _42672_);
  or (_30201_, _42668_, \oc8051_golden_model_1.PCON [0]);
  and (_30202_, _30201_, _43998_);
  and (_43519_, _30202_, _30200_);
  nor (_30203_, _04685_, \oc8051_golden_model_1.PCON [1]);
  not (_30204_, _30203_);
  and (_30205_, _11695_, _04685_);
  nor (_30206_, _30205_, _02838_);
  and (_30207_, _30206_, _30204_);
  and (_30208_, _04685_, _02551_);
  nor (_30210_, _30208_, _30203_);
  and (_30211_, _30210_, _03075_);
  nor (_30212_, _10462_, _04000_);
  or (_30213_, _30212_, _30203_);
  nor (_30214_, _30213_, _03336_);
  and (_30215_, _30210_, _03813_);
  not (_30216_, \oc8051_golden_model_1.PCON [1]);
  nor (_30217_, _03813_, _30216_);
  or (_30218_, _30217_, _30215_);
  and (_30219_, _30218_, _03810_);
  and (_30221_, _11606_, _04685_);
  nor (_30222_, _30221_, _30203_);
  and (_30223_, _30222_, _02974_);
  or (_30224_, _30223_, _30219_);
  and (_30225_, _30224_, _03336_);
  nor (_30226_, _30225_, _30214_);
  nor (_30227_, _30226_, _03075_);
  or (_30228_, _30227_, _06770_);
  nor (_30229_, _30228_, _30211_);
  and (_30230_, _30213_, _06770_);
  or (_30232_, _30230_, _02853_);
  nor (_30233_, _30232_, _30229_);
  or (_30234_, _10462_, _06151_);
  nor (_30235_, _30203_, _05540_);
  and (_30236_, _30235_, _30234_);
  or (_30237_, _30236_, _30233_);
  and (_30238_, _30237_, _02838_);
  nor (_30239_, _30238_, _30207_);
  nor (_30240_, _30239_, _02802_);
  and (_30241_, _04685_, _03698_);
  not (_30242_, _30241_);
  nor (_30243_, _30203_, _02803_);
  and (_30244_, _30243_, _30242_);
  nor (_30245_, _30244_, _30240_);
  nor (_30246_, _30245_, _02980_);
  nor (_30247_, _11710_, _10462_);
  nor (_30248_, _30247_, _03887_);
  and (_30249_, _30248_, _30204_);
  nor (_30250_, _30249_, _30246_);
  nor (_30251_, _30250_, _03127_);
  nor (_30254_, _11715_, _10462_);
  nor (_30255_, _30254_, _03128_);
  and (_30256_, _30255_, _30204_);
  nor (_30257_, _30256_, _30251_);
  nor (_30258_, _30257_, _02970_);
  nor (_30259_, _11709_, _10462_);
  nor (_30260_, _30259_, _03883_);
  and (_30261_, _30260_, _30204_);
  nor (_30262_, _30261_, _30258_);
  nor (_30263_, _30262_, _03135_);
  nor (_30265_, _04685_, _30216_);
  nor (_30266_, _30265_, _13722_);
  nor (_30267_, _30266_, _03137_);
  and (_30268_, _30267_, _30210_);
  nor (_30269_, _30268_, _30263_);
  or (_30270_, _30269_, _17961_);
  and (_30271_, _30208_, _05178_);
  or (_30272_, _30271_, _05788_);
  or (_30273_, _30272_, _30203_);
  and (_30274_, _30273_, _03906_);
  and (_30276_, _30241_, _05178_);
  or (_30277_, _30203_, _05783_);
  or (_30278_, _30277_, _30276_);
  and (_30279_, _30278_, _30274_);
  and (_30280_, _30279_, _30270_);
  nor (_30281_, _30222_, _03906_);
  nor (_30282_, _30281_, _30280_);
  and (_30283_, _30282_, _02890_);
  nor (_30284_, _30221_, _30265_);
  nor (_30285_, _30284_, _02890_);
  or (_30287_, _30285_, _30283_);
  or (_30288_, _30287_, _42672_);
  or (_30289_, _42668_, \oc8051_golden_model_1.PCON [1]);
  and (_30290_, _30289_, _43998_);
  and (_43520_, _30290_, _30288_);
  not (_30291_, \oc8051_golden_model_1.PCON [2]);
  nor (_30292_, _04685_, _30291_);
  nor (_30293_, _30292_, _05130_);
  not (_30294_, _30293_);
  and (_30295_, _04685_, _05701_);
  nor (_30297_, _30295_, _30292_);
  nor (_30298_, _30297_, _03883_);
  and (_30299_, _30298_, _30294_);
  and (_30300_, _04685_, _04435_);
  nor (_30301_, _30300_, _30292_);
  and (_30302_, _30301_, _06770_);
  nor (_30303_, _11801_, _10462_);
  nor (_30304_, _30303_, _30292_);
  nor (_30305_, _30304_, _03810_);
  nor (_30306_, _03813_, _30291_);
  and (_30308_, _04685_, \oc8051_golden_model_1.ACC [2]);
  nor (_30309_, _30308_, _30292_);
  nor (_30310_, _30309_, _03814_);
  nor (_30311_, _30310_, _30306_);
  nor (_30312_, _30311_, _02974_);
  or (_30313_, _30312_, _30305_);
  and (_30314_, _30313_, _03336_);
  nor (_30315_, _30301_, _03336_);
  or (_30316_, _30315_, _30314_);
  and (_30317_, _30316_, _03084_);
  nor (_30319_, _30309_, _03084_);
  nor (_30320_, _30319_, _06770_);
  not (_30321_, _30320_);
  nor (_30322_, _30321_, _30317_);
  nor (_30323_, _30322_, _30302_);
  nor (_30324_, _30323_, _02853_);
  and (_30325_, _04685_, _06155_);
  nor (_30326_, _30292_, _05540_);
  not (_30327_, _30326_);
  nor (_30328_, _30327_, _30325_);
  nor (_30330_, _30328_, _30324_);
  and (_30331_, _30330_, _02838_);
  nor (_30332_, _11906_, _10462_);
  nor (_30333_, _30332_, _30292_);
  nor (_30334_, _30333_, _02838_);
  or (_30335_, _30334_, _30331_);
  and (_30336_, _30335_, _02803_);
  nor (_30337_, _30297_, _02803_);
  or (_30338_, _30337_, _30336_);
  and (_30339_, _30338_, _03887_);
  and (_30341_, _11921_, _04685_);
  nor (_30342_, _30341_, _30292_);
  nor (_30343_, _30342_, _03887_);
  or (_30344_, _30343_, _30339_);
  and (_30345_, _30344_, _03128_);
  and (_30346_, _11927_, _04685_);
  nor (_30347_, _30346_, _30292_);
  nor (_30348_, _30347_, _03128_);
  or (_30349_, _30348_, _30345_);
  and (_30350_, _30349_, _03883_);
  nor (_30352_, _30350_, _30299_);
  nor (_30353_, _30352_, _03135_);
  nor (_30354_, _30309_, _03137_);
  and (_30355_, _30354_, _30294_);
  or (_30356_, _30355_, _30353_);
  and (_30357_, _30356_, _05783_);
  nor (_30358_, _11919_, _10462_);
  nor (_30359_, _30358_, _30292_);
  nor (_30360_, _30359_, _05783_);
  or (_30361_, _30360_, _30357_);
  and (_30363_, _30361_, _05788_);
  nor (_30364_, _11926_, _10462_);
  nor (_30365_, _30364_, _30292_);
  nor (_30366_, _30365_, _05788_);
  or (_30367_, _30366_, _03163_);
  nor (_30368_, _30367_, _30363_);
  and (_30369_, _30304_, _03163_);
  or (_30370_, _30369_, _02888_);
  nor (_30371_, _30370_, _30368_);
  and (_30372_, _11985_, _04685_);
  nor (_30374_, _30372_, _30292_);
  nor (_30375_, _30374_, _02890_);
  or (_30376_, _30375_, _30371_);
  or (_30377_, _30376_, _42672_);
  or (_30378_, _42668_, \oc8051_golden_model_1.PCON [2]);
  and (_30379_, _30378_, _43998_);
  and (_43522_, _30379_, _30377_);
  not (_30380_, \oc8051_golden_model_1.PCON [3]);
  nor (_30381_, _04685_, _30380_);
  and (_30382_, _12133_, _04685_);
  nor (_30384_, _30382_, _30381_);
  nor (_30385_, _30384_, _03128_);
  and (_30386_, _04685_, \oc8051_golden_model_1.ACC [3]);
  nor (_30387_, _30386_, _30381_);
  nor (_30388_, _30387_, _03084_);
  nor (_30389_, _30387_, _03814_);
  nor (_30390_, _03813_, _30380_);
  or (_30391_, _30390_, _30389_);
  and (_30392_, _30391_, _03810_);
  nor (_30393_, _12017_, _10462_);
  nor (_30395_, _30393_, _30381_);
  nor (_30396_, _30395_, _03810_);
  or (_30397_, _30396_, _30392_);
  and (_30398_, _30397_, _03336_);
  and (_30399_, _04685_, _04241_);
  nor (_30400_, _30399_, _30381_);
  nor (_30401_, _30400_, _03336_);
  nor (_30402_, _30401_, _30398_);
  nor (_30403_, _30402_, _03075_);
  or (_30404_, _30403_, _06770_);
  nor (_30406_, _30404_, _30388_);
  and (_30407_, _30400_, _06770_);
  or (_30408_, _30407_, _02853_);
  nor (_30409_, _30408_, _30406_);
  and (_30410_, _04685_, _06154_);
  or (_30411_, _30410_, _30381_);
  and (_30412_, _30411_, _02853_);
  or (_30413_, _30412_, _02579_);
  or (_30414_, _30413_, _30409_);
  nor (_30415_, _12112_, _10462_);
  or (_30417_, _30381_, _02838_);
  or (_30418_, _30417_, _30415_);
  and (_30419_, _30418_, _02803_);
  and (_30420_, _30419_, _30414_);
  and (_30421_, _04685_, _05658_);
  nor (_30422_, _30421_, _30381_);
  nor (_30423_, _30422_, _02803_);
  or (_30424_, _30423_, _30420_);
  and (_30425_, _30424_, _03887_);
  and (_30426_, _12127_, _04685_);
  nor (_30428_, _30426_, _30381_);
  nor (_30429_, _30428_, _03887_);
  or (_30430_, _30429_, _30425_);
  and (_30431_, _30430_, _03128_);
  nor (_30432_, _30431_, _30385_);
  nor (_30433_, _30432_, _02970_);
  nor (_30434_, _30381_, _05079_);
  not (_30435_, _30434_);
  nor (_30436_, _30422_, _03883_);
  and (_30437_, _30436_, _30435_);
  nor (_30439_, _30437_, _30433_);
  nor (_30440_, _30439_, _03135_);
  nor (_30441_, _30387_, _03137_);
  and (_30442_, _30441_, _30435_);
  or (_30443_, _30442_, _30440_);
  and (_30444_, _30443_, _05783_);
  nor (_30445_, _12125_, _10462_);
  nor (_30446_, _30445_, _30381_);
  nor (_30447_, _30446_, _05783_);
  or (_30448_, _30447_, _30444_);
  and (_30450_, _30448_, _05788_);
  nor (_30451_, _12132_, _10462_);
  nor (_30452_, _30451_, _30381_);
  nor (_30453_, _30452_, _05788_);
  or (_30454_, _30453_, _03163_);
  nor (_30455_, _30454_, _30450_);
  and (_30456_, _30395_, _03163_);
  or (_30457_, _30456_, _02888_);
  nor (_30458_, _30457_, _30455_);
  and (_30459_, _12183_, _04685_);
  nor (_30461_, _30459_, _30381_);
  nor (_30462_, _30461_, _02890_);
  or (_30463_, _30462_, _30458_);
  or (_30464_, _30463_, _42672_);
  or (_30465_, _42668_, \oc8051_golden_model_1.PCON [3]);
  and (_30466_, _30465_, _43998_);
  and (_43523_, _30466_, _30464_);
  not (_30467_, \oc8051_golden_model_1.PCON [4]);
  nor (_30468_, _04685_, _30467_);
  and (_30469_, _12207_, _04685_);
  nor (_30471_, _30469_, _30468_);
  nor (_30472_, _30471_, _03128_);
  and (_30473_, _04685_, _04982_);
  nor (_30474_, _30473_, _30468_);
  and (_30475_, _30474_, _06770_);
  and (_30476_, _04685_, \oc8051_golden_model_1.ACC [4]);
  nor (_30477_, _30476_, _30468_);
  nor (_30478_, _30477_, _03084_);
  nor (_30479_, _30477_, _03814_);
  nor (_30480_, _03813_, _30467_);
  or (_30482_, _30480_, _30479_);
  and (_30483_, _30482_, _03810_);
  nor (_30484_, _12217_, _10462_);
  nor (_30485_, _30484_, _30468_);
  nor (_30486_, _30485_, _03810_);
  or (_30487_, _30486_, _30483_);
  and (_30488_, _30487_, _03336_);
  nor (_30489_, _30474_, _03336_);
  nor (_30490_, _30489_, _30488_);
  nor (_30491_, _30490_, _03075_);
  or (_30493_, _30491_, _06770_);
  nor (_30494_, _30493_, _30478_);
  nor (_30495_, _30494_, _30475_);
  nor (_30496_, _30495_, _02853_);
  and (_30497_, _04685_, _06159_);
  nor (_30498_, _30468_, _05540_);
  not (_30499_, _30498_);
  nor (_30500_, _30499_, _30497_);
  or (_30501_, _30500_, _02579_);
  nor (_30502_, _30501_, _30496_);
  nor (_30504_, _12321_, _10462_);
  nor (_30505_, _30504_, _30468_);
  nor (_30506_, _30505_, _02838_);
  or (_30507_, _30506_, _02802_);
  or (_30508_, _30507_, _30502_);
  and (_30509_, _05666_, _04685_);
  nor (_30510_, _30509_, _30468_);
  nand (_30511_, _30510_, _02802_);
  and (_30512_, _30511_, _30508_);
  and (_30513_, _30512_, _03887_);
  and (_30515_, _12211_, _04685_);
  nor (_30516_, _30515_, _30468_);
  nor (_30517_, _30516_, _03887_);
  or (_30518_, _30517_, _30513_);
  and (_30519_, _30518_, _03128_);
  nor (_30520_, _30519_, _30472_);
  nor (_30521_, _30520_, _02970_);
  nor (_30522_, _30468_, _05031_);
  not (_30523_, _30522_);
  nor (_30524_, _30510_, _03883_);
  and (_30526_, _30524_, _30523_);
  nor (_30527_, _30526_, _30521_);
  nor (_30528_, _30527_, _03135_);
  nor (_30529_, _30477_, _03137_);
  and (_30530_, _30529_, _30523_);
  or (_30531_, _30530_, _30528_);
  and (_30532_, _30531_, _05783_);
  nor (_30533_, _12209_, _10462_);
  nor (_30534_, _30533_, _30468_);
  nor (_30535_, _30534_, _05783_);
  or (_30537_, _30535_, _30532_);
  and (_30538_, _30537_, _05788_);
  nor (_30539_, _12206_, _10462_);
  nor (_30540_, _30539_, _30468_);
  nor (_30541_, _30540_, _05788_);
  or (_30542_, _30541_, _03163_);
  nor (_30543_, _30542_, _30538_);
  and (_30544_, _30485_, _03163_);
  or (_30545_, _30544_, _02888_);
  nor (_30546_, _30545_, _30543_);
  and (_30548_, _12389_, _04685_);
  nor (_30549_, _30548_, _30468_);
  nor (_30550_, _30549_, _02890_);
  or (_30551_, _30550_, _30546_);
  or (_30552_, _30551_, _42672_);
  or (_30553_, _42668_, \oc8051_golden_model_1.PCON [4]);
  and (_30554_, _30553_, _43998_);
  and (_43524_, _30554_, _30552_);
  not (_30555_, \oc8051_golden_model_1.PCON [5]);
  nor (_30556_, _04685_, _30555_);
  and (_30558_, _12411_, _04685_);
  nor (_30559_, _30558_, _30556_);
  nor (_30560_, _30559_, _03128_);
  and (_30561_, _04685_, \oc8051_golden_model_1.ACC [5]);
  nor (_30562_, _30561_, _30556_);
  nor (_30563_, _30562_, _03084_);
  nor (_30564_, _30562_, _03814_);
  nor (_30565_, _03813_, _30555_);
  or (_30566_, _30565_, _30564_);
  and (_30567_, _30566_, _03810_);
  nor (_30568_, _12407_, _10462_);
  nor (_30569_, _30568_, _30556_);
  nor (_30570_, _30569_, _03810_);
  or (_30571_, _30570_, _30567_);
  and (_30572_, _30571_, _03336_);
  and (_30573_, _04685_, _04877_);
  nor (_30574_, _30573_, _30556_);
  nor (_30575_, _30574_, _03336_);
  nor (_30576_, _30575_, _30572_);
  nor (_30577_, _30576_, _03075_);
  or (_30580_, _30577_, _06770_);
  nor (_30581_, _30580_, _30563_);
  and (_30582_, _30574_, _06770_);
  nor (_30583_, _30582_, _30581_);
  nor (_30584_, _30583_, _02853_);
  and (_30585_, _04685_, _06158_);
  nor (_30586_, _30556_, _05540_);
  not (_30587_, _30586_);
  nor (_30588_, _30587_, _30585_);
  or (_30589_, _30588_, _02579_);
  nor (_30591_, _30589_, _30584_);
  nor (_30592_, _12527_, _10462_);
  nor (_30593_, _30592_, _30556_);
  nor (_30594_, _30593_, _02838_);
  or (_30595_, _30594_, _02802_);
  or (_30596_, _30595_, _30591_);
  and (_30597_, _05614_, _04685_);
  nor (_30598_, _30597_, _30556_);
  nand (_30599_, _30598_, _02802_);
  and (_30600_, _30599_, _30596_);
  and (_30602_, _30600_, _03887_);
  and (_30603_, _12415_, _04685_);
  nor (_30604_, _30603_, _30556_);
  nor (_30605_, _30604_, _03887_);
  or (_30606_, _30605_, _30602_);
  and (_30607_, _30606_, _03128_);
  nor (_30608_, _30607_, _30560_);
  nor (_30609_, _30608_, _02970_);
  nor (_30610_, _30556_, _04924_);
  not (_30611_, _30610_);
  nor (_30613_, _30598_, _03883_);
  and (_30614_, _30613_, _30611_);
  nor (_30615_, _30614_, _30609_);
  nor (_30616_, _30615_, _03135_);
  nor (_30617_, _30562_, _03137_);
  and (_30618_, _30617_, _30611_);
  or (_30619_, _30618_, _30616_);
  and (_30620_, _30619_, _05783_);
  nor (_30621_, _12413_, _10462_);
  nor (_30622_, _30621_, _30556_);
  nor (_30624_, _30622_, _05783_);
  or (_30625_, _30624_, _30620_);
  and (_30626_, _30625_, _05788_);
  nor (_30627_, _12410_, _10462_);
  nor (_30628_, _30627_, _30556_);
  nor (_30629_, _30628_, _05788_);
  or (_30630_, _30629_, _03163_);
  nor (_30631_, _30630_, _30626_);
  and (_30632_, _30569_, _03163_);
  or (_30633_, _30632_, _02888_);
  nor (_30635_, _30633_, _30631_);
  and (_30636_, _12589_, _04685_);
  nor (_30637_, _30636_, _30556_);
  nor (_30638_, _30637_, _02890_);
  or (_30639_, _30638_, _30635_);
  or (_30640_, _30639_, _42672_);
  or (_30641_, _42668_, \oc8051_golden_model_1.PCON [5]);
  and (_30642_, _30641_, _43998_);
  and (_43525_, _30642_, _30640_);
  not (_30643_, \oc8051_golden_model_1.PCON [6]);
  nor (_30645_, _04685_, _30643_);
  and (_30646_, _12613_, _04685_);
  nor (_30647_, _30646_, _30645_);
  nor (_30648_, _30647_, _03128_);
  and (_30649_, _04685_, _04770_);
  nor (_30650_, _30649_, _30645_);
  and (_30651_, _30650_, _06770_);
  and (_30652_, _04685_, \oc8051_golden_model_1.ACC [6]);
  nor (_30653_, _30652_, _30645_);
  nor (_30654_, _30653_, _03814_);
  nor (_30656_, _03813_, _30643_);
  or (_30657_, _30656_, _30654_);
  and (_30658_, _30657_, _03810_);
  nor (_30659_, _12603_, _10462_);
  nor (_30660_, _30659_, _30645_);
  nor (_30661_, _30660_, _03810_);
  or (_30662_, _30661_, _30658_);
  and (_30663_, _30662_, _03336_);
  nor (_30664_, _30650_, _03336_);
  nor (_30665_, _30664_, _30663_);
  nor (_30667_, _30665_, _03075_);
  nor (_30668_, _30653_, _03084_);
  nor (_30669_, _30668_, _06770_);
  not (_30670_, _30669_);
  nor (_30671_, _30670_, _30667_);
  nor (_30672_, _30671_, _30651_);
  nor (_30673_, _30672_, _02853_);
  and (_30674_, _04685_, _05849_);
  nor (_30675_, _30645_, _05540_);
  not (_30676_, _30675_);
  nor (_30678_, _30676_, _30674_);
  or (_30679_, _30678_, _02579_);
  nor (_30680_, _30679_, _30673_);
  nor (_30681_, _12722_, _10462_);
  nor (_30682_, _30681_, _30645_);
  nor (_30683_, _30682_, _02838_);
  or (_30684_, _30683_, _02802_);
  or (_30685_, _30684_, _30680_);
  and (_30686_, _12729_, _04685_);
  nor (_30687_, _30686_, _30645_);
  nand (_30689_, _30687_, _02802_);
  and (_30690_, _30689_, _30685_);
  and (_30691_, _30690_, _03887_);
  and (_30692_, _12739_, _04685_);
  nor (_30693_, _30692_, _30645_);
  nor (_30694_, _30693_, _03887_);
  or (_30695_, _30694_, _30691_);
  and (_30696_, _30695_, _03128_);
  nor (_30697_, _30696_, _30648_);
  nor (_30698_, _30697_, _02970_);
  nor (_30700_, _30645_, _04819_);
  not (_30701_, _30700_);
  nor (_30702_, _30687_, _03883_);
  and (_30703_, _30702_, _30701_);
  nor (_30704_, _30703_, _30698_);
  nor (_30705_, _30704_, _03135_);
  nor (_30706_, _30653_, _03137_);
  and (_30707_, _30706_, _30701_);
  or (_30708_, _30707_, _30705_);
  and (_30709_, _30708_, _05783_);
  nor (_30711_, _12737_, _10462_);
  nor (_30712_, _30711_, _30645_);
  nor (_30713_, _30712_, _05783_);
  or (_30714_, _30713_, _30709_);
  and (_30715_, _30714_, _05788_);
  nor (_30716_, _12612_, _10462_);
  nor (_30717_, _30716_, _30645_);
  nor (_30718_, _30717_, _05788_);
  or (_30719_, _30718_, _03163_);
  nor (_30720_, _30719_, _30715_);
  and (_30722_, _30660_, _03163_);
  or (_30723_, _30722_, _02888_);
  nor (_30724_, _30723_, _30720_);
  and (_30725_, _12794_, _04685_);
  nor (_30726_, _30725_, _30645_);
  nor (_30727_, _30726_, _02890_);
  or (_30728_, _30727_, _30724_);
  or (_30729_, _30728_, _42672_);
  or (_30730_, _42668_, \oc8051_golden_model_1.PCON [6]);
  and (_30731_, _30730_, _43998_);
  and (_43526_, _30731_, _30729_);
  not (_30733_, \oc8051_golden_model_1.SBUF [0]);
  nor (_30734_, _04700_, _30733_);
  and (_30735_, _05226_, _04700_);
  nor (_30736_, _30735_, _30734_);
  and (_30737_, _30736_, _16625_);
  and (_30738_, _04700_, _05672_);
  nor (_30739_, _30738_, _30734_);
  or (_30740_, _30739_, _03883_);
  nor (_30741_, _30740_, _30735_);
  and (_30742_, _04700_, \oc8051_golden_model_1.ACC [0]);
  nor (_30743_, _30742_, _30734_);
  nor (_30744_, _30743_, _03084_);
  nor (_30745_, _30743_, _03814_);
  nor (_30746_, _03813_, _30733_);
  or (_30747_, _30746_, _30745_);
  and (_30748_, _30747_, _03810_);
  nor (_30749_, _30736_, _03810_);
  or (_30750_, _30749_, _30748_);
  and (_30751_, _30750_, _03336_);
  and (_30753_, _04700_, _03808_);
  nor (_30754_, _30753_, _30734_);
  nor (_30755_, _30754_, _03336_);
  nor (_30756_, _30755_, _30751_);
  nor (_30757_, _30756_, _03075_);
  or (_30758_, _30757_, _06770_);
  nor (_30759_, _30758_, _30744_);
  and (_30760_, _30754_, _06770_);
  nor (_30761_, _30760_, _30759_);
  nor (_30762_, _30761_, _02853_);
  and (_30764_, _04700_, _06152_);
  nor (_30765_, _30734_, _05540_);
  not (_30766_, _30765_);
  nor (_30767_, _30766_, _30764_);
  nor (_30768_, _30767_, _30762_);
  and (_30769_, _30768_, _02838_);
  nor (_30770_, _11505_, _10543_);
  nor (_30771_, _30770_, _30734_);
  nor (_30772_, _30771_, _02838_);
  or (_30773_, _30772_, _30769_);
  and (_30775_, _30773_, _02803_);
  nor (_30776_, _30739_, _02803_);
  or (_30777_, _30776_, _30775_);
  and (_30778_, _30777_, _03887_);
  and (_30779_, _11399_, _04700_);
  nor (_30780_, _30779_, _30734_);
  nor (_30781_, _30780_, _03887_);
  or (_30782_, _30781_, _30778_);
  and (_30783_, _30782_, _03128_);
  and (_30784_, _11522_, _04700_);
  nor (_30786_, _30784_, _30734_);
  nor (_30787_, _30786_, _03128_);
  or (_30788_, _30787_, _30783_);
  and (_30789_, _30788_, _03883_);
  nor (_30790_, _30789_, _30741_);
  nor (_30791_, _30790_, _03135_);
  nor (_30792_, _30734_, _09409_);
  or (_30793_, _30792_, _03137_);
  nor (_30794_, _30793_, _30743_);
  or (_30795_, _30794_, _30791_);
  and (_30797_, _30795_, _05783_);
  nor (_30798_, _11396_, _10543_);
  nor (_30799_, _30798_, _30734_);
  nor (_30800_, _30799_, _05783_);
  or (_30801_, _30800_, _30797_);
  and (_30802_, _30801_, _05788_);
  nor (_30803_, _11520_, _10543_);
  nor (_30804_, _30803_, _30734_);
  nor (_30805_, _30804_, _05788_);
  nor (_30806_, _30805_, _16625_);
  not (_30808_, _30806_);
  nor (_30809_, _30808_, _30802_);
  nor (_30810_, _30809_, _30737_);
  or (_30811_, _30810_, _42672_);
  or (_30812_, _42668_, \oc8051_golden_model_1.SBUF [0]);
  and (_30813_, _30812_, _43998_);
  and (_43528_, _30813_, _30811_);
  nor (_30814_, _04700_, \oc8051_golden_model_1.SBUF [1]);
  not (_30815_, _30814_);
  nor (_30816_, _11715_, _10543_);
  nor (_30818_, _30816_, _03128_);
  and (_30819_, _30818_, _30815_);
  and (_30820_, _04700_, _03698_);
  not (_30821_, _30820_);
  nor (_30822_, _30814_, _02803_);
  and (_30823_, _30822_, _30821_);
  and (_30824_, _11695_, _04700_);
  nor (_30825_, _30824_, _02838_);
  and (_30826_, _30825_, _30815_);
  and (_30827_, _04700_, _06151_);
  not (_30829_, \oc8051_golden_model_1.SBUF [1]);
  nor (_30830_, _04700_, _30829_);
  nor (_30831_, _30830_, _05540_);
  not (_30832_, _30831_);
  nor (_30833_, _30832_, _30827_);
  not (_30834_, _30833_);
  and (_30835_, _04700_, _04000_);
  or (_30836_, _30830_, _30142_);
  nor (_30837_, _30836_, _30835_);
  and (_30838_, _04700_, _02551_);
  nor (_30840_, _30838_, _30814_);
  and (_30841_, _30840_, _03075_);
  nor (_30842_, _30841_, _06770_);
  and (_30843_, _11606_, _04700_);
  nor (_30844_, _30843_, _30814_);
  and (_30845_, _30844_, _02974_);
  and (_30846_, _30840_, _03813_);
  nor (_30847_, _03813_, _30829_);
  nor (_30848_, _30847_, _30846_);
  nor (_30849_, _30848_, _02974_);
  or (_30851_, _30849_, _03069_);
  nor (_30852_, _30851_, _30845_);
  or (_30853_, _30852_, _03075_);
  and (_30854_, _30853_, _30842_);
  nor (_30855_, _30854_, _30837_);
  nor (_30856_, _30855_, _02853_);
  nor (_30857_, _30856_, _02579_);
  and (_30858_, _30857_, _30834_);
  nor (_30859_, _30858_, _30826_);
  nor (_30860_, _30859_, _02802_);
  nor (_30862_, _30860_, _30823_);
  nor (_30863_, _30862_, _02980_);
  nor (_30864_, _11710_, _10543_);
  nor (_30865_, _30864_, _03887_);
  and (_30866_, _30865_, _30815_);
  nor (_30867_, _30866_, _30863_);
  nor (_30868_, _30867_, _03127_);
  nor (_30869_, _30868_, _30819_);
  nor (_30870_, _30869_, _02970_);
  nor (_30871_, _11709_, _10543_);
  nor (_30873_, _30871_, _03883_);
  and (_30874_, _30873_, _30815_);
  nor (_30875_, _30874_, _30870_);
  nor (_30876_, _30875_, _03135_);
  nor (_30877_, _30830_, _13722_);
  nor (_30878_, _30877_, _03137_);
  and (_30879_, _30878_, _30840_);
  nor (_30880_, _30879_, _30876_);
  or (_30881_, _30880_, _17961_);
  and (_30882_, _11714_, _04700_);
  or (_30884_, _30882_, _05788_);
  or (_30885_, _30884_, _30814_);
  and (_30886_, _30885_, _03906_);
  and (_30887_, _30820_, _05178_);
  or (_30888_, _30814_, _05783_);
  or (_30889_, _30888_, _30887_);
  and (_30890_, _30889_, _30886_);
  and (_30891_, _30890_, _30881_);
  nor (_30892_, _30844_, _03906_);
  nor (_30893_, _30892_, _30891_);
  nor (_30895_, _30893_, _02888_);
  nor (_30896_, _30843_, _30830_);
  and (_30897_, _30896_, _02888_);
  nor (_30898_, _30897_, _30895_);
  or (_30899_, _30898_, _42672_);
  or (_30900_, _42668_, \oc8051_golden_model_1.SBUF [1]);
  and (_30901_, _30900_, _43998_);
  and (_43529_, _30901_, _30899_);
  not (_30902_, \oc8051_golden_model_1.SBUF [2]);
  nor (_30903_, _04700_, _30902_);
  and (_30905_, _04700_, _06155_);
  nor (_30906_, _30905_, _30903_);
  or (_30907_, _30906_, _05540_);
  and (_30908_, _04700_, \oc8051_golden_model_1.ACC [2]);
  nor (_30909_, _30908_, _30903_);
  nor (_30910_, _30909_, _03814_);
  nor (_30911_, _03813_, _30902_);
  or (_30912_, _30911_, _30910_);
  and (_30913_, _30912_, _03810_);
  nor (_30914_, _11801_, _10543_);
  nor (_30916_, _30914_, _30903_);
  nor (_30917_, _30916_, _03810_);
  or (_30918_, _30917_, _30913_);
  and (_30919_, _30918_, _03336_);
  and (_30920_, _04700_, _04435_);
  nor (_30921_, _30920_, _30903_);
  nor (_30922_, _30921_, _03336_);
  nor (_30923_, _30922_, _30919_);
  nor (_30924_, _30923_, _03075_);
  nor (_30925_, _30909_, _03084_);
  nor (_30927_, _30925_, _06770_);
  not (_30928_, _30927_);
  nor (_30929_, _30928_, _30924_);
  and (_30930_, _30921_, _06770_);
  or (_30931_, _30930_, _02853_);
  or (_30932_, _30931_, _30929_);
  and (_30933_, _30932_, _02838_);
  and (_30934_, _30933_, _30907_);
  nor (_30935_, _11906_, _10543_);
  or (_30936_, _30903_, _02838_);
  or (_30938_, _30936_, _30935_);
  and (_30939_, _30938_, _02803_);
  not (_30940_, _30939_);
  nor (_30941_, _30940_, _30934_);
  and (_30942_, _04700_, _05701_);
  nor (_30943_, _30942_, _30903_);
  nor (_30944_, _30943_, _02803_);
  or (_30945_, _30944_, _30941_);
  and (_30946_, _30945_, _03887_);
  and (_30947_, _11921_, _04700_);
  nor (_30949_, _30947_, _30903_);
  nor (_30950_, _30949_, _03887_);
  or (_30951_, _30950_, _30946_);
  and (_30952_, _30951_, _03128_);
  and (_30953_, _11927_, _04700_);
  nor (_30954_, _30953_, _30903_);
  nor (_30955_, _30954_, _03128_);
  or (_30956_, _30955_, _30952_);
  and (_30957_, _30956_, _03883_);
  nor (_30958_, _30903_, _05130_);
  or (_30960_, _30943_, _03883_);
  nor (_30961_, _30960_, _30958_);
  nor (_30962_, _30961_, _30957_);
  nor (_30963_, _30962_, _03135_);
  or (_30964_, _30958_, _03137_);
  nor (_30965_, _30964_, _30909_);
  or (_30966_, _30965_, _30963_);
  and (_30967_, _30966_, _05783_);
  nor (_30968_, _11919_, _10543_);
  nor (_30969_, _30968_, _30903_);
  nor (_30971_, _30969_, _05783_);
  or (_30972_, _30971_, _30967_);
  and (_30973_, _30972_, _05788_);
  nor (_30974_, _11926_, _10543_);
  nor (_30975_, _30974_, _30903_);
  nor (_30976_, _30975_, _05788_);
  or (_30977_, _30976_, _03163_);
  nor (_30978_, _30977_, _30973_);
  and (_30979_, _30916_, _03163_);
  or (_30980_, _30979_, _02888_);
  nor (_30982_, _30980_, _30978_);
  and (_30983_, _11985_, _04700_);
  nor (_30984_, _30983_, _30903_);
  nor (_30985_, _30984_, _02890_);
  or (_30986_, _30985_, _30982_);
  or (_30987_, _30986_, _42672_);
  or (_30988_, _42668_, \oc8051_golden_model_1.SBUF [2]);
  and (_30989_, _30988_, _43998_);
  and (_43530_, _30989_, _30987_);
  not (_30990_, \oc8051_golden_model_1.SBUF [3]);
  nor (_30992_, _04700_, _30990_);
  and (_30993_, _12133_, _04700_);
  nor (_30994_, _30993_, _30992_);
  nor (_30995_, _30994_, _03128_);
  and (_30996_, _04700_, \oc8051_golden_model_1.ACC [3]);
  nor (_30997_, _30996_, _30992_);
  nor (_30998_, _30997_, _03084_);
  nor (_30999_, _30997_, _03814_);
  nor (_31000_, _03813_, _30990_);
  or (_31001_, _31000_, _30999_);
  and (_31003_, _31001_, _03810_);
  nor (_31004_, _12017_, _10543_);
  nor (_31005_, _31004_, _30992_);
  nor (_31006_, _31005_, _03810_);
  or (_31007_, _31006_, _31003_);
  and (_31008_, _31007_, _03336_);
  and (_31009_, _04700_, _04241_);
  nor (_31010_, _31009_, _30992_);
  nor (_31011_, _31010_, _03336_);
  nor (_31012_, _31011_, _31008_);
  nor (_31014_, _31012_, _03075_);
  or (_31015_, _31014_, _06770_);
  nor (_31016_, _31015_, _30998_);
  and (_31017_, _31010_, _06770_);
  or (_31018_, _31017_, _02853_);
  nor (_31019_, _31018_, _31016_);
  and (_31020_, _04700_, _06154_);
  or (_31021_, _31020_, _30992_);
  and (_31022_, _31021_, _02853_);
  or (_31023_, _31022_, _02579_);
  or (_31025_, _31023_, _31019_);
  nor (_31026_, _12112_, _10543_);
  or (_31027_, _30992_, _02838_);
  or (_31028_, _31027_, _31026_);
  and (_31029_, _31028_, _02803_);
  and (_31030_, _31029_, _31025_);
  and (_31031_, _04700_, _05658_);
  nor (_31032_, _31031_, _30992_);
  nor (_31033_, _31032_, _02803_);
  or (_31034_, _31033_, _31030_);
  and (_31036_, _31034_, _03887_);
  and (_31037_, _12127_, _04700_);
  nor (_31038_, _31037_, _30992_);
  nor (_31039_, _31038_, _03887_);
  or (_31040_, _31039_, _31036_);
  and (_31041_, _31040_, _03128_);
  nor (_31042_, _31041_, _30995_);
  nor (_31043_, _31042_, _02970_);
  nor (_31044_, _30992_, _05079_);
  not (_31045_, _31044_);
  nor (_31046_, _31032_, _03883_);
  and (_31047_, _31046_, _31045_);
  nor (_31048_, _31047_, _31043_);
  nor (_31049_, _31048_, _03135_);
  nor (_31050_, _30997_, _03137_);
  and (_31051_, _31050_, _31045_);
  nor (_31052_, _31051_, _02965_);
  not (_31053_, _31052_);
  nor (_31054_, _31053_, _31049_);
  nor (_31055_, _12125_, _10543_);
  or (_31058_, _30992_, _05783_);
  nor (_31059_, _31058_, _31055_);
  or (_31060_, _31059_, _03123_);
  nor (_31061_, _31060_, _31054_);
  nor (_31062_, _12132_, _10543_);
  nor (_31063_, _31062_, _30992_);
  nor (_31064_, _31063_, _05788_);
  or (_31065_, _31064_, _03163_);
  nor (_31066_, _31065_, _31061_);
  and (_31067_, _31005_, _03163_);
  or (_31069_, _31067_, _02888_);
  nor (_31070_, _31069_, _31066_);
  and (_31071_, _12183_, _04700_);
  nor (_31072_, _31071_, _30992_);
  nor (_31073_, _31072_, _02890_);
  or (_31074_, _31073_, _31070_);
  or (_31075_, _31074_, _42672_);
  or (_31076_, _42668_, \oc8051_golden_model_1.SBUF [3]);
  and (_31077_, _31076_, _43998_);
  and (_43531_, _31077_, _31075_);
  not (_31079_, \oc8051_golden_model_1.SBUF [4]);
  nor (_31080_, _04700_, _31079_);
  and (_31081_, _12207_, _04700_);
  nor (_31082_, _31081_, _31080_);
  nor (_31083_, _31082_, _03128_);
  and (_31084_, _04700_, _04982_);
  nor (_31085_, _31084_, _31080_);
  and (_31086_, _31085_, _06770_);
  and (_31087_, _04700_, \oc8051_golden_model_1.ACC [4]);
  nor (_31088_, _31087_, _31080_);
  nor (_31090_, _31088_, _03084_);
  nor (_31091_, _31088_, _03814_);
  nor (_31092_, _03813_, _31079_);
  or (_31093_, _31092_, _31091_);
  and (_31094_, _31093_, _03810_);
  nor (_31095_, _12217_, _10543_);
  nor (_31096_, _31095_, _31080_);
  nor (_31097_, _31096_, _03810_);
  or (_31098_, _31097_, _31094_);
  and (_31099_, _31098_, _03336_);
  nor (_31101_, _31085_, _03336_);
  nor (_31102_, _31101_, _31099_);
  nor (_31103_, _31102_, _03075_);
  or (_31104_, _31103_, _06770_);
  nor (_31105_, _31104_, _31090_);
  nor (_31106_, _31105_, _31086_);
  nor (_31107_, _31106_, _02853_);
  and (_31108_, _04700_, _06159_);
  nor (_31109_, _31080_, _05540_);
  not (_31110_, _31109_);
  nor (_31112_, _31110_, _31108_);
  or (_31113_, _31112_, _02579_);
  nor (_31114_, _31113_, _31107_);
  nor (_31115_, _12321_, _10543_);
  nor (_31116_, _31115_, _31080_);
  nor (_31117_, _31116_, _02838_);
  or (_31118_, _31117_, _02802_);
  or (_31119_, _31118_, _31114_);
  and (_31120_, _05666_, _04700_);
  nor (_31121_, _31120_, _31080_);
  nand (_31123_, _31121_, _02802_);
  and (_31124_, _31123_, _31119_);
  and (_31125_, _31124_, _03887_);
  and (_31126_, _12211_, _04700_);
  nor (_31127_, _31126_, _31080_);
  nor (_31128_, _31127_, _03887_);
  or (_31129_, _31128_, _31125_);
  and (_31130_, _31129_, _03128_);
  nor (_31131_, _31130_, _31083_);
  nor (_31132_, _31131_, _02970_);
  nor (_31134_, _31080_, _05031_);
  not (_31135_, _31134_);
  nor (_31136_, _31121_, _03883_);
  and (_31137_, _31136_, _31135_);
  nor (_31138_, _31137_, _31132_);
  nor (_31139_, _31138_, _03135_);
  nor (_31140_, _31088_, _03137_);
  and (_31141_, _31140_, _31135_);
  or (_31142_, _31141_, _31139_);
  and (_31143_, _31142_, _05783_);
  nor (_31145_, _12209_, _10543_);
  nor (_31146_, _31145_, _31080_);
  nor (_31147_, _31146_, _05783_);
  or (_31148_, _31147_, _31143_);
  and (_31149_, _31148_, _05788_);
  nor (_31150_, _12206_, _10543_);
  nor (_31151_, _31150_, _31080_);
  nor (_31152_, _31151_, _05788_);
  or (_31153_, _31152_, _03163_);
  nor (_31154_, _31153_, _31149_);
  and (_31156_, _31096_, _03163_);
  or (_31157_, _31156_, _02888_);
  nor (_31158_, _31157_, _31154_);
  and (_31159_, _12389_, _04700_);
  nor (_31160_, _31159_, _31080_);
  nor (_31161_, _31160_, _02890_);
  or (_31162_, _31161_, _31158_);
  or (_31163_, _31162_, _42672_);
  or (_31164_, _42668_, \oc8051_golden_model_1.SBUF [4]);
  and (_31165_, _31164_, _43998_);
  and (_43532_, _31165_, _31163_);
  not (_31167_, \oc8051_golden_model_1.SBUF [5]);
  nor (_31168_, _04700_, _31167_);
  and (_31169_, _12411_, _04700_);
  nor (_31170_, _31169_, _31168_);
  nor (_31171_, _31170_, _03128_);
  and (_31172_, _04700_, _04877_);
  nor (_31173_, _31172_, _31168_);
  and (_31174_, _31173_, _06770_);
  nor (_31175_, _12407_, _10543_);
  nor (_31177_, _31175_, _31168_);
  and (_31178_, _31177_, _02974_);
  and (_31179_, _04700_, \oc8051_golden_model_1.ACC [5]);
  nor (_31180_, _31179_, _31168_);
  or (_31181_, _31180_, _03814_);
  or (_31182_, _03813_, _31167_);
  and (_31183_, _31182_, _03810_);
  and (_31184_, _31183_, _31181_);
  or (_31185_, _31184_, _03069_);
  nor (_31186_, _31185_, _31178_);
  nor (_31188_, _31173_, _03336_);
  nor (_31189_, _31188_, _31186_);
  nor (_31190_, _31189_, _03075_);
  nor (_31191_, _31180_, _03084_);
  nor (_31192_, _31191_, _06770_);
  not (_31193_, _31192_);
  nor (_31194_, _31193_, _31190_);
  nor (_31195_, _31194_, _31174_);
  nor (_31196_, _31195_, _02853_);
  and (_31197_, _04700_, _06158_);
  nor (_31199_, _31168_, _05540_);
  not (_31200_, _31199_);
  nor (_31201_, _31200_, _31197_);
  or (_31202_, _31201_, _02579_);
  nor (_31203_, _31202_, _31196_);
  nor (_31204_, _12527_, _10543_);
  nor (_31205_, _31204_, _31168_);
  nor (_31206_, _31205_, _02838_);
  or (_31207_, _31206_, _02802_);
  or (_31208_, _31207_, _31203_);
  and (_31210_, _05614_, _04700_);
  nor (_31211_, _31210_, _31168_);
  nand (_31212_, _31211_, _02802_);
  and (_31213_, _31212_, _31208_);
  and (_31214_, _31213_, _03887_);
  and (_31215_, _12415_, _04700_);
  nor (_31216_, _31215_, _31168_);
  nor (_31217_, _31216_, _03887_);
  or (_31218_, _31217_, _31214_);
  and (_31219_, _31218_, _03128_);
  nor (_31221_, _31219_, _31171_);
  nor (_31222_, _31221_, _02970_);
  nor (_31223_, _31168_, _04924_);
  not (_31224_, _31223_);
  nor (_31225_, _31211_, _03883_);
  and (_31226_, _31225_, _31224_);
  nor (_31227_, _31226_, _31222_);
  nor (_31228_, _31227_, _03135_);
  nor (_31229_, _31180_, _03137_);
  and (_31230_, _31229_, _31224_);
  or (_31232_, _31230_, _31228_);
  and (_31233_, _31232_, _05783_);
  nor (_31234_, _12413_, _10543_);
  nor (_31235_, _31234_, _31168_);
  nor (_31236_, _31235_, _05783_);
  or (_31237_, _31236_, _31233_);
  and (_31238_, _31237_, _05788_);
  nor (_31239_, _12410_, _10543_);
  nor (_31240_, _31239_, _31168_);
  nor (_31241_, _31240_, _05788_);
  or (_31243_, _31241_, _03163_);
  nor (_31244_, _31243_, _31238_);
  and (_31245_, _31177_, _03163_);
  or (_31246_, _31245_, _02888_);
  nor (_31247_, _31246_, _31244_);
  and (_31248_, _12589_, _04700_);
  nor (_31249_, _31248_, _31168_);
  nor (_31250_, _31249_, _02890_);
  or (_31251_, _31250_, _31247_);
  or (_31252_, _31251_, _42672_);
  or (_31254_, _42668_, \oc8051_golden_model_1.SBUF [5]);
  and (_31255_, _31254_, _43998_);
  and (_43533_, _31255_, _31252_);
  not (_31256_, \oc8051_golden_model_1.SBUF [6]);
  nor (_31257_, _04700_, _31256_);
  and (_31258_, _12613_, _04700_);
  nor (_31259_, _31258_, _31257_);
  nor (_31260_, _31259_, _03128_);
  and (_31261_, _04700_, _04770_);
  nor (_31262_, _31261_, _31257_);
  and (_31264_, _31262_, _06770_);
  and (_31265_, _04700_, \oc8051_golden_model_1.ACC [6]);
  nor (_31266_, _31265_, _31257_);
  nor (_31267_, _31266_, _03814_);
  nor (_31268_, _03813_, _31256_);
  or (_31269_, _31268_, _31267_);
  and (_31270_, _31269_, _03810_);
  nor (_31271_, _12603_, _10543_);
  nor (_31272_, _31271_, _31257_);
  nor (_31273_, _31272_, _03810_);
  or (_31274_, _31273_, _31270_);
  and (_31275_, _31274_, _03336_);
  nor (_31276_, _31262_, _03336_);
  nor (_31277_, _31276_, _31275_);
  nor (_31278_, _31277_, _03075_);
  nor (_31279_, _31266_, _03084_);
  nor (_31280_, _31279_, _06770_);
  not (_31281_, _31280_);
  nor (_31282_, _31281_, _31278_);
  nor (_31283_, _31282_, _31264_);
  nor (_31286_, _31283_, _02853_);
  and (_31287_, _04700_, _05849_);
  nor (_31288_, _31257_, _05540_);
  not (_31289_, _31288_);
  nor (_31290_, _31289_, _31287_);
  or (_31291_, _31290_, _02579_);
  nor (_31292_, _31291_, _31286_);
  nor (_31293_, _12722_, _10543_);
  nor (_31294_, _31293_, _31257_);
  nor (_31295_, _31294_, _02838_);
  or (_31297_, _31295_, _02802_);
  or (_31298_, _31297_, _31292_);
  and (_31299_, _12729_, _04700_);
  nor (_31300_, _31299_, _31257_);
  nand (_31301_, _31300_, _02802_);
  and (_31302_, _31301_, _31298_);
  and (_31303_, _31302_, _03887_);
  and (_31304_, _12739_, _04700_);
  nor (_31305_, _31304_, _31257_);
  nor (_31306_, _31305_, _03887_);
  or (_31308_, _31306_, _31303_);
  and (_31309_, _31308_, _03128_);
  nor (_31310_, _31309_, _31260_);
  nor (_31311_, _31310_, _02970_);
  nor (_31312_, _31257_, _04819_);
  not (_31313_, _31312_);
  nor (_31314_, _31300_, _03883_);
  and (_31315_, _31314_, _31313_);
  nor (_31316_, _31315_, _31311_);
  nor (_31317_, _31316_, _03135_);
  nor (_31319_, _31266_, _03137_);
  and (_31320_, _31319_, _31313_);
  or (_31321_, _31320_, _31317_);
  and (_31322_, _31321_, _05783_);
  nor (_31323_, _12737_, _10543_);
  nor (_31324_, _31323_, _31257_);
  nor (_31325_, _31324_, _05783_);
  or (_31326_, _31325_, _31322_);
  and (_31327_, _31326_, _05788_);
  nor (_31328_, _12612_, _10543_);
  nor (_31330_, _31328_, _31257_);
  nor (_31331_, _31330_, _05788_);
  or (_31332_, _31331_, _03163_);
  nor (_31333_, _31332_, _31327_);
  and (_31334_, _31272_, _03163_);
  or (_31335_, _31334_, _02888_);
  nor (_31336_, _31335_, _31333_);
  and (_31337_, _12794_, _04700_);
  nor (_31338_, _31337_, _31257_);
  nor (_31339_, _31338_, _02890_);
  or (_31341_, _31339_, _31336_);
  or (_31342_, _31341_, _42672_);
  or (_31343_, _42668_, \oc8051_golden_model_1.SBUF [6]);
  and (_31344_, _31343_, _43998_);
  and (_43534_, _31344_, _31342_);
  not (_31345_, \oc8051_golden_model_1.SCON [0]);
  nor (_31346_, _04666_, _31345_);
  and (_31347_, _11522_, _04666_);
  nor (_31348_, _31347_, _31346_);
  nor (_31349_, _31348_, _03128_);
  and (_31351_, _04666_, _03808_);
  nor (_31352_, _31351_, _31346_);
  and (_31353_, _31352_, _06770_);
  and (_31354_, _04666_, \oc8051_golden_model_1.ACC [0]);
  nor (_31355_, _31354_, _31346_);
  nor (_31356_, _31355_, _03814_);
  nor (_31357_, _03813_, _31345_);
  or (_31358_, _31357_, _31356_);
  and (_31359_, _31358_, _03810_);
  and (_31360_, _05226_, _04666_);
  nor (_31362_, _31360_, _31346_);
  nor (_31363_, _31362_, _03810_);
  or (_31364_, _31363_, _31359_);
  and (_31365_, _31364_, _02881_);
  nor (_31366_, _05338_, _31345_);
  and (_31367_, _11417_, _05338_);
  nor (_31368_, _31367_, _31366_);
  nor (_31369_, _31368_, _02881_);
  nor (_31370_, _31369_, _31365_);
  nor (_31371_, _31370_, _03069_);
  nor (_31373_, _31352_, _03336_);
  or (_31374_, _31373_, _31371_);
  and (_31375_, _31374_, _03084_);
  nor (_31376_, _31355_, _03084_);
  or (_31377_, _31376_, _31375_);
  and (_31378_, _31377_, _02877_);
  and (_31379_, _31346_, _02876_);
  or (_31380_, _31379_, _31378_);
  and (_31381_, _31380_, _02870_);
  nor (_31382_, _31362_, _02870_);
  or (_31384_, _31382_, _31381_);
  and (_31385_, _31384_, _02864_);
  nor (_31386_, _11448_, _10633_);
  nor (_31387_, _31386_, _31366_);
  nor (_31388_, _31387_, _02864_);
  or (_31389_, _31388_, _06770_);
  nor (_31390_, _31389_, _31385_);
  nor (_31391_, _31390_, _31353_);
  nor (_31392_, _31391_, _02853_);
  and (_31393_, _04666_, _06152_);
  nor (_31395_, _31346_, _05540_);
  not (_31396_, _31395_);
  nor (_31397_, _31396_, _31393_);
  or (_31398_, _31397_, _02579_);
  nor (_31399_, _31398_, _31392_);
  nor (_31400_, _11505_, _10649_);
  nor (_31401_, _31400_, _31346_);
  nor (_31402_, _31401_, _02838_);
  or (_31403_, _31402_, _02802_);
  or (_31404_, _31403_, _31399_);
  and (_31406_, _04666_, _05672_);
  nor (_31407_, _31406_, _31346_);
  nand (_31408_, _31407_, _02802_);
  and (_31409_, _31408_, _31404_);
  and (_31410_, _31409_, _03887_);
  and (_31411_, _11399_, _04666_);
  nor (_31412_, _31411_, _31346_);
  nor (_31413_, _31412_, _03887_);
  or (_31414_, _31413_, _31410_);
  and (_31415_, _31414_, _03128_);
  nor (_31417_, _31415_, _31349_);
  nor (_31418_, _31417_, _02970_);
  or (_31419_, _31407_, _03883_);
  nor (_31420_, _31419_, _31360_);
  nor (_31421_, _31420_, _31418_);
  nor (_31422_, _31421_, _03135_);
  nor (_31423_, _31346_, _09409_);
  or (_31424_, _31423_, _03137_);
  nor (_31425_, _31424_, _31355_);
  or (_31426_, _31425_, _31422_);
  and (_31428_, _31426_, _05783_);
  nor (_31429_, _11396_, _10649_);
  nor (_31430_, _31429_, _31346_);
  nor (_31431_, _31430_, _05783_);
  or (_31432_, _31431_, _31428_);
  and (_31433_, _31432_, _05788_);
  nor (_31434_, _11520_, _10649_);
  nor (_31435_, _31434_, _31346_);
  nor (_31436_, _31435_, _05788_);
  or (_31437_, _31436_, _31433_);
  and (_31439_, _31437_, _03906_);
  nor (_31440_, _31362_, _03906_);
  or (_31441_, _31440_, _31439_);
  and (_31442_, _31441_, _02498_);
  and (_31443_, _31346_, _02497_);
  or (_31444_, _31443_, _31442_);
  and (_31445_, _31444_, _02890_);
  nor (_31446_, _31362_, _02890_);
  or (_31447_, _31446_, _31445_);
  or (_31448_, _31447_, _42672_);
  or (_31450_, _42668_, \oc8051_golden_model_1.SCON [0]);
  and (_31451_, _31450_, _43998_);
  and (_43536_, _31451_, _31448_);
  and (_31452_, _04666_, _03698_);
  not (_31453_, _31452_);
  nor (_31454_, _04666_, \oc8051_golden_model_1.SCON [1]);
  nor (_31455_, _31454_, _02803_);
  and (_31456_, _31455_, _31453_);
  not (_31457_, \oc8051_golden_model_1.SCON [1]);
  nor (_31458_, _04666_, _31457_);
  and (_31460_, _04666_, _06151_);
  or (_31461_, _31460_, _31458_);
  and (_31462_, _31461_, _02853_);
  and (_31463_, _04666_, _02551_);
  nor (_31464_, _31463_, _31454_);
  and (_31465_, _31464_, _03813_);
  nor (_31466_, _03813_, _31457_);
  or (_31467_, _31466_, _31465_);
  and (_31468_, _31467_, _03810_);
  and (_31469_, _11606_, _04666_);
  nor (_31471_, _31469_, _31454_);
  and (_31472_, _31471_, _02974_);
  or (_31473_, _31472_, _31468_);
  and (_31474_, _31473_, _02881_);
  nor (_31475_, _05338_, _31457_);
  and (_31476_, _11592_, _05338_);
  nor (_31477_, _31476_, _31475_);
  nor (_31478_, _31477_, _02881_);
  or (_31479_, _31478_, _31474_);
  and (_31480_, _31479_, _03336_);
  and (_31482_, _04666_, _04000_);
  nor (_31483_, _31482_, _31458_);
  nor (_31484_, _31483_, _03336_);
  or (_31485_, _31484_, _31480_);
  and (_31486_, _31485_, _03084_);
  and (_31487_, _31464_, _03075_);
  or (_31488_, _31487_, _31486_);
  and (_31489_, _31488_, _02877_);
  and (_31490_, _11595_, _05338_);
  nor (_31491_, _31490_, _31475_);
  nor (_31493_, _31491_, _02877_);
  or (_31494_, _31493_, _02869_);
  or (_31495_, _31494_, _31489_);
  and (_31496_, _31476_, _11591_);
  or (_31497_, _31475_, _02870_);
  or (_31498_, _31497_, _31496_);
  and (_31499_, _31498_, _31495_);
  and (_31500_, _31499_, _02864_);
  nor (_31501_, _11638_, _10633_);
  nor (_31502_, _31475_, _31501_);
  nor (_31504_, _31502_, _02864_);
  or (_31505_, _31504_, _06770_);
  nor (_31506_, _31505_, _31500_);
  and (_31507_, _31483_, _06770_);
  or (_31508_, _31507_, _02853_);
  nor (_31509_, _31508_, _31506_);
  or (_31510_, _31509_, _31462_);
  and (_31511_, _31510_, _02838_);
  nor (_31512_, _11695_, _10649_);
  nor (_31513_, _31512_, _31458_);
  nor (_31515_, _31513_, _02838_);
  nor (_31516_, _31515_, _31511_);
  nor (_31517_, _31516_, _02802_);
  nor (_31518_, _31517_, _31456_);
  nor (_31519_, _31518_, _02980_);
  nor (_31520_, _11710_, _10649_);
  or (_31521_, _31520_, _03887_);
  nor (_31522_, _31521_, _31454_);
  nor (_31523_, _31522_, _31519_);
  nor (_31524_, _31523_, _03127_);
  and (_31526_, _11715_, _04666_);
  or (_31527_, _31526_, _31458_);
  and (_31528_, _31527_, _03127_);
  nor (_31529_, _31528_, _31524_);
  nor (_31530_, _31529_, _02970_);
  nor (_31531_, _11709_, _10649_);
  or (_31532_, _31531_, _03883_);
  nor (_31533_, _31532_, _31454_);
  nor (_31534_, _31533_, _31530_);
  nor (_31535_, _31534_, _03135_);
  nor (_31537_, _31458_, _13722_);
  nor (_31538_, _31537_, _03137_);
  and (_31539_, _31538_, _31464_);
  nor (_31540_, _31539_, _31535_);
  or (_31541_, _31540_, _17961_);
  nor (_31542_, _11708_, _10649_);
  or (_31543_, _31542_, _31458_);
  and (_31544_, _31543_, _02965_);
  not (_31545_, _31544_);
  and (_31546_, _11714_, _04666_);
  or (_31547_, _31546_, _05788_);
  or (_31548_, _31547_, _31454_);
  and (_31549_, _31548_, _03906_);
  and (_31550_, _31549_, _31545_);
  and (_31551_, _31550_, _31541_);
  nor (_31552_, _31471_, _03906_);
  or (_31553_, _31552_, _02497_);
  nor (_31554_, _31553_, _31551_);
  nor (_31555_, _31491_, _02498_);
  or (_31556_, _31555_, _02888_);
  nor (_31558_, _31556_, _31554_);
  nor (_31559_, _31469_, _31458_);
  and (_31560_, _31559_, _02888_);
  nor (_31561_, _31560_, _31558_);
  or (_31562_, _31561_, _42672_);
  or (_31563_, _42668_, \oc8051_golden_model_1.SCON [1]);
  and (_31564_, _31563_, _43998_);
  and (_43537_, _31564_, _31562_);
  not (_31565_, \oc8051_golden_model_1.SCON [2]);
  nor (_31566_, _04666_, _31565_);
  and (_31568_, _11927_, _04666_);
  nor (_31569_, _31568_, _31566_);
  nor (_31570_, _31569_, _03128_);
  and (_31571_, _04666_, _04435_);
  nor (_31572_, _31571_, _31566_);
  and (_31573_, _31572_, _06770_);
  and (_31574_, _04666_, \oc8051_golden_model_1.ACC [2]);
  nor (_31575_, _31574_, _31566_);
  nor (_31576_, _31575_, _03814_);
  nor (_31577_, _03813_, _31565_);
  or (_31579_, _31577_, _31576_);
  and (_31580_, _31579_, _03810_);
  nor (_31581_, _11801_, _10649_);
  nor (_31582_, _31581_, _31566_);
  nor (_31583_, _31582_, _03810_);
  or (_31584_, _31583_, _31580_);
  and (_31585_, _31584_, _02881_);
  nor (_31586_, _05338_, _31565_);
  and (_31587_, _11815_, _05338_);
  nor (_31588_, _31587_, _31586_);
  nor (_31590_, _31588_, _02881_);
  or (_31591_, _31590_, _31585_);
  and (_31592_, _31591_, _03336_);
  nor (_31593_, _31572_, _03336_);
  or (_31594_, _31593_, _31592_);
  and (_31595_, _31594_, _03084_);
  nor (_31596_, _31575_, _03084_);
  or (_31597_, _31596_, _31595_);
  and (_31598_, _31597_, _02877_);
  and (_31599_, _11797_, _05338_);
  nor (_31601_, _31599_, _31586_);
  nor (_31602_, _31601_, _02877_);
  or (_31603_, _31602_, _02869_);
  or (_31604_, _31603_, _31598_);
  and (_31605_, _31587_, _11830_);
  or (_31606_, _31586_, _02870_);
  or (_31607_, _31606_, _31605_);
  and (_31608_, _31607_, _02864_);
  and (_31609_, _31608_, _31604_);
  nor (_31610_, _11848_, _10633_);
  nor (_31612_, _31610_, _31586_);
  nor (_31613_, _31612_, _02864_);
  nor (_31614_, _31613_, _06770_);
  not (_31615_, _31614_);
  nor (_31616_, _31615_, _31609_);
  nor (_31617_, _31616_, _31573_);
  nor (_31618_, _31617_, _02853_);
  and (_31619_, _04666_, _06155_);
  nor (_31620_, _31566_, _05540_);
  not (_31621_, _31620_);
  nor (_31623_, _31621_, _31619_);
  or (_31624_, _31623_, _02579_);
  nor (_31625_, _31624_, _31618_);
  nor (_31626_, _11906_, _10649_);
  nor (_31627_, _31626_, _31566_);
  nor (_31628_, _31627_, _02838_);
  or (_31629_, _31628_, _02802_);
  or (_31630_, _31629_, _31625_);
  and (_31631_, _04666_, _05701_);
  nor (_31632_, _31631_, _31566_);
  nand (_31634_, _31632_, _02802_);
  and (_31635_, _31634_, _31630_);
  and (_31636_, _31635_, _03887_);
  and (_31637_, _11921_, _04666_);
  nor (_31638_, _31637_, _31566_);
  nor (_31639_, _31638_, _03887_);
  or (_31640_, _31639_, _31636_);
  and (_31641_, _31640_, _03128_);
  nor (_31642_, _31641_, _31570_);
  nor (_31643_, _31642_, _02970_);
  nor (_31645_, _31566_, _05130_);
  not (_31646_, _31645_);
  nor (_31647_, _31632_, _03883_);
  and (_31648_, _31647_, _31646_);
  nor (_31649_, _31648_, _31643_);
  nor (_31650_, _31649_, _03135_);
  nor (_31651_, _31575_, _03137_);
  and (_31652_, _31651_, _31646_);
  nor (_31653_, _31652_, _02965_);
  not (_31654_, _31653_);
  nor (_31656_, _31654_, _31650_);
  nor (_31657_, _11919_, _10649_);
  or (_31658_, _31566_, _05783_);
  nor (_31659_, _31658_, _31657_);
  or (_31660_, _31659_, _03123_);
  nor (_31661_, _31660_, _31656_);
  nor (_31662_, _11926_, _10649_);
  nor (_31663_, _31662_, _31566_);
  nor (_31664_, _31663_, _05788_);
  or (_31665_, _31664_, _31661_);
  and (_31667_, _31665_, _03906_);
  nor (_31668_, _31582_, _03906_);
  or (_31669_, _31668_, _31667_);
  and (_31670_, _31669_, _02498_);
  nor (_31671_, _31601_, _02498_);
  or (_31672_, _31671_, _31670_);
  and (_31673_, _31672_, _02890_);
  and (_31674_, _11985_, _04666_);
  nor (_31675_, _31674_, _31566_);
  nor (_31676_, _31675_, _02890_);
  or (_31678_, _31676_, _31673_);
  or (_31679_, _31678_, _42672_);
  or (_31680_, _42668_, \oc8051_golden_model_1.SCON [2]);
  and (_31681_, _31680_, _43998_);
  and (_43538_, _31681_, _31679_);
  not (_31682_, \oc8051_golden_model_1.SCON [3]);
  nor (_31683_, _04666_, _31682_);
  and (_31684_, _12133_, _04666_);
  nor (_31685_, _31684_, _31683_);
  nor (_31686_, _31685_, _03128_);
  and (_31688_, _04666_, _04241_);
  nor (_31689_, _31688_, _31683_);
  and (_31690_, _31689_, _06770_);
  and (_31691_, _04666_, \oc8051_golden_model_1.ACC [3]);
  nor (_31692_, _31691_, _31683_);
  nor (_31693_, _31692_, _03814_);
  nor (_31694_, _03813_, _31682_);
  or (_31695_, _31694_, _31693_);
  and (_31696_, _31695_, _03810_);
  nor (_31697_, _12017_, _10649_);
  nor (_31699_, _31697_, _31683_);
  nor (_31700_, _31699_, _03810_);
  or (_31701_, _31700_, _31696_);
  and (_31702_, _31701_, _02881_);
  nor (_31703_, _05338_, _31682_);
  and (_31704_, _12021_, _05338_);
  nor (_31705_, _31704_, _31703_);
  nor (_31706_, _31705_, _02881_);
  or (_31707_, _31706_, _03069_);
  or (_31708_, _31707_, _31702_);
  nand (_31710_, _31689_, _03069_);
  and (_31711_, _31710_, _31708_);
  and (_31712_, _31711_, _03084_);
  nor (_31713_, _31692_, _03084_);
  or (_31714_, _31713_, _31712_);
  and (_31715_, _31714_, _02877_);
  and (_31716_, _12005_, _05338_);
  nor (_31717_, _31716_, _31703_);
  nor (_31718_, _31717_, _02877_);
  or (_31719_, _31718_, _02869_);
  or (_31721_, _31719_, _31715_);
  nor (_31722_, _31703_, _12036_);
  nor (_31723_, _31722_, _31705_);
  or (_31724_, _31723_, _02870_);
  and (_31725_, _31724_, _02864_);
  and (_31726_, _31725_, _31721_);
  nor (_31727_, _12054_, _10633_);
  nor (_31728_, _31727_, _31703_);
  nor (_31729_, _31728_, _02864_);
  nor (_31730_, _31729_, _06770_);
  not (_31732_, _31730_);
  nor (_31733_, _31732_, _31726_);
  nor (_31734_, _31733_, _31690_);
  nor (_31735_, _31734_, _02853_);
  and (_31736_, _04666_, _06154_);
  nor (_31737_, _31683_, _05540_);
  not (_31738_, _31737_);
  nor (_31739_, _31738_, _31736_);
  or (_31740_, _31739_, _02579_);
  nor (_31741_, _31740_, _31735_);
  nor (_31743_, _12112_, _10649_);
  nor (_31744_, _31743_, _31683_);
  nor (_31745_, _31744_, _02838_);
  or (_31746_, _31745_, _02802_);
  or (_31747_, _31746_, _31741_);
  and (_31748_, _04666_, _05658_);
  nor (_31749_, _31748_, _31683_);
  nand (_31750_, _31749_, _02802_);
  and (_31751_, _31750_, _31747_);
  and (_31752_, _31751_, _03887_);
  and (_31754_, _12127_, _04666_);
  nor (_31755_, _31754_, _31683_);
  nor (_31756_, _31755_, _03887_);
  or (_31757_, _31756_, _31752_);
  and (_31758_, _31757_, _03128_);
  nor (_31759_, _31758_, _31686_);
  nor (_31760_, _31759_, _02970_);
  nor (_31761_, _31683_, _05079_);
  not (_31762_, _31761_);
  nor (_31763_, _31749_, _03883_);
  and (_31765_, _31763_, _31762_);
  nor (_31766_, _31765_, _31760_);
  nor (_31767_, _31766_, _03135_);
  nor (_31768_, _31692_, _03137_);
  and (_31769_, _31768_, _31762_);
  or (_31770_, _31769_, _31767_);
  and (_31771_, _31770_, _05783_);
  nor (_31772_, _12125_, _10649_);
  nor (_31773_, _31772_, _31683_);
  nor (_31774_, _31773_, _05783_);
  or (_31776_, _31774_, _31771_);
  and (_31777_, _31776_, _05788_);
  nor (_31778_, _12132_, _10649_);
  nor (_31779_, _31778_, _31683_);
  nor (_31780_, _31779_, _05788_);
  or (_31781_, _31780_, _31777_);
  and (_31782_, _31781_, _03906_);
  nor (_31783_, _31699_, _03906_);
  or (_31784_, _31783_, _31782_);
  and (_31785_, _31784_, _02498_);
  nor (_31787_, _31717_, _02498_);
  or (_31788_, _31787_, _31785_);
  and (_31789_, _31788_, _02890_);
  and (_31790_, _12183_, _04666_);
  nor (_31791_, _31790_, _31683_);
  nor (_31792_, _31791_, _02890_);
  or (_31793_, _31792_, _31789_);
  or (_31794_, _31793_, _42672_);
  or (_31795_, _42668_, \oc8051_golden_model_1.SCON [3]);
  and (_31796_, _31795_, _43998_);
  and (_43539_, _31796_, _31794_);
  not (_31798_, \oc8051_golden_model_1.SCON [4]);
  nor (_31799_, _04666_, _31798_);
  and (_31800_, _12207_, _04666_);
  nor (_31801_, _31800_, _31799_);
  nor (_31802_, _31801_, _03128_);
  and (_31803_, _04666_, _04982_);
  nor (_31804_, _31803_, _31799_);
  and (_31805_, _31804_, _06770_);
  nor (_31806_, _05338_, _31798_);
  and (_31808_, _12213_, _05338_);
  nor (_31809_, _31808_, _31806_);
  nor (_31810_, _31809_, _02877_);
  and (_31811_, _04666_, \oc8051_golden_model_1.ACC [4]);
  nor (_31812_, _31811_, _31799_);
  nor (_31813_, _31812_, _03814_);
  nor (_31814_, _03813_, _31798_);
  or (_31815_, _31814_, _31813_);
  and (_31816_, _31815_, _03810_);
  nor (_31817_, _12217_, _10649_);
  nor (_31819_, _31817_, _31799_);
  nor (_31820_, _31819_, _03810_);
  or (_31821_, _31820_, _31816_);
  and (_31822_, _31821_, _02881_);
  and (_31823_, _12231_, _05338_);
  nor (_31824_, _31823_, _31806_);
  nor (_31825_, _31824_, _02881_);
  or (_31826_, _31825_, _03069_);
  or (_31827_, _31826_, _31822_);
  nand (_31828_, _31804_, _03069_);
  and (_31830_, _31828_, _31827_);
  and (_31831_, _31830_, _03084_);
  nor (_31832_, _31812_, _03084_);
  or (_31833_, _31832_, _31831_);
  and (_31834_, _31833_, _02877_);
  nor (_31835_, _31834_, _31810_);
  nor (_31836_, _31835_, _02869_);
  and (_31837_, _12247_, _05338_);
  nor (_31838_, _31837_, _31806_);
  nor (_31839_, _31838_, _02870_);
  nor (_31841_, _31839_, _31836_);
  nor (_31842_, _31841_, _02863_);
  nor (_31843_, _12264_, _10633_);
  nor (_31844_, _31843_, _31806_);
  nor (_31845_, _31844_, _02864_);
  nor (_31846_, _31845_, _06770_);
  not (_31847_, _31846_);
  nor (_31848_, _31847_, _31842_);
  nor (_31849_, _31848_, _31805_);
  nor (_31850_, _31849_, _02853_);
  and (_31851_, _04666_, _06159_);
  nor (_31852_, _31799_, _05540_);
  not (_31853_, _31852_);
  nor (_31854_, _31853_, _31851_);
  nor (_31855_, _31854_, _02579_);
  not (_31856_, _31855_);
  nor (_31857_, _31856_, _31850_);
  nor (_31858_, _12321_, _10649_);
  nor (_31859_, _31858_, _31799_);
  nor (_31860_, _31859_, _02838_);
  or (_31863_, _31860_, _02802_);
  or (_31864_, _31863_, _31857_);
  and (_31865_, _05666_, _04666_);
  nor (_31866_, _31865_, _31799_);
  nand (_31867_, _31866_, _02802_);
  and (_31868_, _31867_, _31864_);
  and (_31869_, _31868_, _03887_);
  and (_31870_, _12211_, _04666_);
  nor (_31871_, _31870_, _31799_);
  nor (_31872_, _31871_, _03887_);
  or (_31874_, _31872_, _31869_);
  and (_31875_, _31874_, _03128_);
  nor (_31876_, _31875_, _31802_);
  nor (_31877_, _31876_, _02970_);
  nor (_31878_, _31799_, _05031_);
  not (_31879_, _31878_);
  nor (_31880_, _31866_, _03883_);
  and (_31881_, _31880_, _31879_);
  nor (_31882_, _31881_, _31877_);
  nor (_31883_, _31882_, _03135_);
  nor (_31885_, _31812_, _03137_);
  and (_31886_, _31885_, _31879_);
  or (_31887_, _31886_, _31883_);
  and (_31888_, _31887_, _05783_);
  nor (_31889_, _12209_, _10649_);
  nor (_31890_, _31889_, _31799_);
  nor (_31891_, _31890_, _05783_);
  or (_31892_, _31891_, _31888_);
  and (_31893_, _31892_, _05788_);
  nor (_31894_, _12206_, _10649_);
  nor (_31896_, _31894_, _31799_);
  nor (_31897_, _31896_, _05788_);
  or (_31898_, _31897_, _31893_);
  and (_31899_, _31898_, _03906_);
  nor (_31900_, _31819_, _03906_);
  or (_31901_, _31900_, _31899_);
  and (_31902_, _31901_, _02498_);
  nor (_31903_, _31809_, _02498_);
  or (_31904_, _31903_, _31902_);
  and (_31905_, _31904_, _02890_);
  and (_31907_, _12389_, _04666_);
  nor (_31908_, _31907_, _31799_);
  nor (_31909_, _31908_, _02890_);
  or (_31910_, _31909_, _31905_);
  or (_31911_, _31910_, _42672_);
  or (_31912_, _42668_, \oc8051_golden_model_1.SCON [4]);
  and (_31913_, _31912_, _43998_);
  and (_43540_, _31913_, _31911_);
  not (_31914_, \oc8051_golden_model_1.SCON [5]);
  nor (_31915_, _04666_, _31914_);
  and (_31917_, _12411_, _04666_);
  nor (_31918_, _31917_, _31915_);
  nor (_31919_, _31918_, _03128_);
  and (_31920_, _04666_, _06158_);
  or (_31921_, _31920_, _31915_);
  and (_31922_, _31921_, _02853_);
  nor (_31923_, _12407_, _10649_);
  nor (_31924_, _31923_, _31915_);
  and (_31925_, _31924_, _02974_);
  and (_31926_, _04666_, \oc8051_golden_model_1.ACC [5]);
  nor (_31928_, _31926_, _31915_);
  or (_31929_, _31928_, _03814_);
  or (_31930_, _03813_, _31914_);
  and (_31931_, _31930_, _03810_);
  and (_31932_, _31931_, _31929_);
  or (_31933_, _31932_, _02880_);
  nor (_31934_, _31933_, _31925_);
  nor (_31935_, _05338_, _31914_);
  and (_31936_, _12435_, _05338_);
  nor (_31937_, _31936_, _31935_);
  nor (_31939_, _31937_, _02881_);
  or (_31940_, _31939_, _03069_);
  or (_31941_, _31940_, _31934_);
  and (_31942_, _04666_, _04877_);
  nor (_31943_, _31942_, _31915_);
  nand (_31944_, _31943_, _03069_);
  and (_31945_, _31944_, _31941_);
  and (_31946_, _31945_, _03084_);
  nor (_31947_, _31928_, _03084_);
  or (_31948_, _31947_, _31946_);
  and (_31950_, _31948_, _02877_);
  and (_31951_, _12417_, _05338_);
  nor (_31952_, _31951_, _31935_);
  nor (_31953_, _31952_, _02877_);
  or (_31954_, _31953_, _02869_);
  or (_31955_, _31954_, _31950_);
  nor (_31956_, _31935_, _12450_);
  nor (_31957_, _31956_, _31937_);
  or (_31958_, _31957_, _02870_);
  and (_31959_, _31958_, _02864_);
  and (_31961_, _31959_, _31955_);
  nor (_31962_, _12468_, _10633_);
  nor (_31963_, _31962_, _31935_);
  nor (_31964_, _31963_, _02864_);
  nor (_31965_, _31964_, _06770_);
  not (_31966_, _31965_);
  nor (_31967_, _31966_, _31961_);
  and (_31968_, _31943_, _06770_);
  or (_31969_, _31968_, _02853_);
  nor (_31970_, _31969_, _31967_);
  or (_31972_, _31970_, _31922_);
  and (_31973_, _31972_, _02838_);
  nor (_31974_, _12527_, _10649_);
  nor (_31975_, _31974_, _31915_);
  nor (_31976_, _31975_, _02838_);
  or (_31977_, _31976_, _02802_);
  or (_31978_, _31977_, _31973_);
  and (_31979_, _05614_, _04666_);
  nor (_31980_, _31979_, _31915_);
  nand (_31981_, _31980_, _02802_);
  and (_31983_, _31981_, _31978_);
  and (_31984_, _31983_, _03887_);
  and (_31985_, _12415_, _04666_);
  nor (_31986_, _31985_, _31915_);
  nor (_31987_, _31986_, _03887_);
  or (_31988_, _31987_, _31984_);
  and (_31989_, _31988_, _03128_);
  nor (_31990_, _31989_, _31919_);
  nor (_31991_, _31990_, _02970_);
  nor (_31992_, _31915_, _04924_);
  not (_31994_, _31992_);
  nor (_31995_, _31980_, _03883_);
  and (_31996_, _31995_, _31994_);
  nor (_31997_, _31996_, _31991_);
  nor (_31998_, _31997_, _03135_);
  nor (_31999_, _31928_, _03137_);
  and (_32000_, _31999_, _31994_);
  or (_32001_, _32000_, _31998_);
  and (_32002_, _32001_, _05783_);
  nor (_32003_, _12413_, _10649_);
  nor (_32005_, _32003_, _31915_);
  nor (_32006_, _32005_, _05783_);
  or (_32007_, _32006_, _32002_);
  and (_32008_, _32007_, _05788_);
  nor (_32009_, _12410_, _10649_);
  nor (_32010_, _32009_, _31915_);
  nor (_32011_, _32010_, _05788_);
  or (_32012_, _32011_, _32008_);
  and (_32013_, _32012_, _03906_);
  nor (_32014_, _31924_, _03906_);
  or (_32016_, _32014_, _32013_);
  and (_32017_, _32016_, _02498_);
  nor (_32018_, _31952_, _02498_);
  or (_32019_, _32018_, _32017_);
  and (_32020_, _32019_, _02890_);
  and (_32021_, _12589_, _04666_);
  nor (_32022_, _32021_, _31915_);
  nor (_32023_, _32022_, _02890_);
  or (_32024_, _32023_, _32020_);
  or (_32025_, _32024_, _42672_);
  or (_32027_, _42668_, \oc8051_golden_model_1.SCON [5]);
  and (_32028_, _32027_, _43998_);
  and (_43541_, _32028_, _32025_);
  not (_32029_, \oc8051_golden_model_1.SCON [6]);
  nor (_32030_, _04666_, _32029_);
  and (_32031_, _12613_, _04666_);
  nor (_32032_, _32031_, _32030_);
  nor (_32033_, _32032_, _03128_);
  and (_32034_, _04666_, _05849_);
  or (_32035_, _32034_, _32030_);
  and (_32037_, _32035_, _02853_);
  and (_32038_, _04666_, \oc8051_golden_model_1.ACC [6]);
  nor (_32039_, _32038_, _32030_);
  nor (_32040_, _32039_, _03814_);
  nor (_32041_, _03813_, _32029_);
  or (_32042_, _32041_, _32040_);
  and (_32043_, _32042_, _03810_);
  nor (_32044_, _12603_, _10649_);
  nor (_32045_, _32044_, _32030_);
  nor (_32046_, _32045_, _03810_);
  or (_32048_, _32046_, _32043_);
  and (_32049_, _32048_, _02881_);
  nor (_32050_, _05338_, _32029_);
  and (_32051_, _12618_, _05338_);
  nor (_32052_, _32051_, _32050_);
  nor (_32053_, _32052_, _02881_);
  or (_32054_, _32053_, _03069_);
  or (_32055_, _32054_, _32049_);
  and (_32056_, _04666_, _04770_);
  nor (_32057_, _32056_, _32030_);
  nand (_32059_, _32057_, _03069_);
  and (_32060_, _32059_, _32055_);
  and (_32061_, _32060_, _03084_);
  nor (_32062_, _32039_, _03084_);
  or (_32063_, _32062_, _32061_);
  and (_32064_, _32063_, _02877_);
  and (_32065_, _12616_, _05338_);
  nor (_32066_, _32065_, _32050_);
  nor (_32067_, _32066_, _02877_);
  or (_32068_, _32067_, _32064_);
  and (_32070_, _32068_, _02870_);
  nor (_32071_, _32050_, _12646_);
  nor (_32072_, _32071_, _32052_);
  and (_32073_, _32072_, _02869_);
  or (_32074_, _32073_, _32070_);
  and (_32075_, _32074_, _02864_);
  nor (_32076_, _12664_, _10633_);
  nor (_32077_, _32076_, _32050_);
  nor (_32078_, _32077_, _02864_);
  nor (_32079_, _32078_, _06770_);
  not (_32081_, _32079_);
  nor (_32082_, _32081_, _32075_);
  and (_32083_, _32057_, _06770_);
  or (_32084_, _32083_, _02853_);
  nor (_32085_, _32084_, _32082_);
  or (_32086_, _32085_, _32037_);
  and (_32087_, _32086_, _02838_);
  nor (_32088_, _12722_, _10649_);
  nor (_32089_, _32088_, _32030_);
  nor (_32090_, _32089_, _02838_);
  or (_32092_, _32090_, _02802_);
  or (_32093_, _32092_, _32087_);
  and (_32094_, _12729_, _04666_);
  nor (_32095_, _32094_, _32030_);
  nand (_32096_, _32095_, _02802_);
  and (_32097_, _32096_, _32093_);
  and (_32098_, _32097_, _03887_);
  and (_32099_, _12739_, _04666_);
  nor (_32100_, _32099_, _32030_);
  nor (_32101_, _32100_, _03887_);
  or (_32103_, _32101_, _32098_);
  and (_32104_, _32103_, _03128_);
  nor (_32105_, _32104_, _32033_);
  nor (_32106_, _32105_, _02970_);
  nor (_32107_, _32030_, _04819_);
  not (_32108_, _32107_);
  nor (_32109_, _32095_, _03883_);
  and (_32110_, _32109_, _32108_);
  nor (_32111_, _32110_, _32106_);
  nor (_32112_, _32111_, _03135_);
  nor (_32114_, _32039_, _03137_);
  and (_32115_, _32114_, _32108_);
  or (_32116_, _32115_, _32112_);
  and (_32117_, _32116_, _05783_);
  nor (_32118_, _12737_, _10649_);
  nor (_32119_, _32118_, _32030_);
  nor (_32120_, _32119_, _05783_);
  or (_32121_, _32120_, _32117_);
  and (_32122_, _32121_, _05788_);
  nor (_32123_, _12612_, _10649_);
  nor (_32125_, _32123_, _32030_);
  nor (_32126_, _32125_, _05788_);
  or (_32127_, _32126_, _32122_);
  and (_32128_, _32127_, _03906_);
  nor (_32129_, _32045_, _03906_);
  or (_32130_, _32129_, _32128_);
  and (_32131_, _32130_, _02498_);
  nor (_32132_, _32066_, _02498_);
  or (_32133_, _32132_, _32131_);
  and (_32134_, _32133_, _02890_);
  and (_32136_, _12794_, _04666_);
  nor (_32137_, _32136_, _32030_);
  nor (_32138_, _32137_, _02890_);
  or (_32139_, _32138_, _32134_);
  or (_32140_, _32139_, _42672_);
  or (_32141_, _42668_, \oc8051_golden_model_1.SCON [6]);
  and (_32142_, _32141_, _43998_);
  and (_43542_, _32142_, _32140_);
  nor (_32143_, _04617_, _02866_);
  and (_32144_, _05226_, _04617_);
  nor (_32146_, _32144_, _32143_);
  and (_32147_, _32146_, _16625_);
  and (_32148_, _04617_, \oc8051_golden_model_1.ACC [0]);
  nor (_32149_, _32148_, _32143_);
  nor (_32150_, _32149_, _03814_);
  nor (_32151_, _03813_, _02866_);
  or (_32152_, _32151_, _32150_);
  and (_32153_, _32152_, _03810_);
  nor (_32154_, _32146_, _03810_);
  or (_32155_, _32154_, _32153_);
  and (_32157_, _32155_, _03336_);
  or (_32158_, _32157_, _03395_);
  and (_32159_, _32158_, _03084_);
  nor (_32160_, _32149_, _03084_);
  or (_32161_, _32160_, _32159_);
  and (_32162_, _32161_, _03941_);
  nor (_32163_, _03851_, _06770_);
  not (_32164_, _32163_);
  nor (_32165_, _32164_, _32162_);
  and (_32166_, _04617_, _03808_);
  or (_32168_, _32143_, _05535_);
  nor (_32169_, _32168_, _32166_);
  nor (_32170_, _32169_, _32165_);
  nor (_32171_, _32170_, _02853_);
  and (_32172_, _04617_, _06152_);
  nor (_32173_, _32143_, _05540_);
  not (_32174_, _32173_);
  nor (_32175_, _32174_, _32172_);
  nor (_32176_, _32175_, _32171_);
  and (_32177_, _32176_, _02838_);
  nor (_32179_, _11505_, _10777_);
  nor (_32180_, _32179_, _32143_);
  nor (_32181_, _32180_, _02838_);
  or (_32182_, _32181_, _32177_);
  and (_32183_, _32182_, _02803_);
  and (_32184_, _04617_, _05672_);
  nor (_32185_, _32184_, _32143_);
  nor (_32186_, _32185_, _02803_);
  or (_32187_, _32186_, _32183_);
  and (_32188_, _32187_, _03887_);
  and (_32190_, _11399_, _04617_);
  nor (_32191_, _32190_, _32143_);
  nor (_32192_, _32191_, _03887_);
  or (_32193_, _32192_, _32188_);
  and (_32194_, _32193_, _03128_);
  and (_32195_, _11522_, _04617_);
  nor (_32196_, _32195_, _32143_);
  nor (_32197_, _32196_, _03128_);
  or (_32198_, _32197_, _32194_);
  and (_32199_, _32198_, _03883_);
  or (_32201_, _32185_, _03883_);
  nor (_32202_, _32201_, _32144_);
  nor (_32203_, _32202_, _32199_);
  nor (_32204_, _32203_, _03135_);
  and (_32205_, _11521_, _04617_);
  or (_32206_, _32205_, _32143_);
  and (_32207_, _32206_, _03135_);
  or (_32208_, _32207_, _32204_);
  and (_32209_, _32208_, _05783_);
  nor (_32210_, _11396_, _10777_);
  nor (_32212_, _32210_, _32143_);
  nor (_32213_, _32212_, _05783_);
  or (_32214_, _32213_, _32209_);
  and (_32215_, _32214_, _05788_);
  nor (_32216_, _11520_, _10777_);
  nor (_32217_, _32216_, _32143_);
  nor (_32218_, _32217_, _05788_);
  nor (_32219_, _32218_, _16625_);
  not (_32220_, _32219_);
  nor (_32221_, _32220_, _32215_);
  nor (_32223_, _32221_, _32147_);
  and (_32224_, _32223_, _42668_);
  nor (_32225_, \oc8051_golden_model_1.SP [0], rst);
  nor (_32226_, _32225_, _00000_);
  or (_43544_, _32226_, _32224_);
  nor (_32227_, _04617_, _03700_);
  and (_32228_, _11606_, _04617_);
  nor (_32229_, _32228_, _32227_);
  nor (_32230_, _32229_, _02890_);
  not (_32231_, _29014_);
  nor (_32233_, _04617_, \oc8051_golden_model_1.SP [1]);
  not (_32234_, _32233_);
  nor (_32235_, _11715_, _10777_);
  nor (_32236_, _32235_, _03128_);
  and (_32237_, _32236_, _32234_);
  and (_32238_, _02514_, _03700_);
  nor (_32239_, _11695_, _10777_);
  or (_32240_, _32239_, _32227_);
  and (_32241_, _32240_, _02579_);
  and (_32242_, _04617_, _02551_);
  nor (_32244_, _32242_, _32233_);
  nor (_32245_, _32244_, _03814_);
  nor (_32246_, _09434_, \oc8051_golden_model_1.SP [1]);
  and (_32247_, _02611_, \oc8051_golden_model_1.SP [1]);
  nor (_32248_, _32247_, _32246_);
  nor (_32249_, _32248_, _32245_);
  and (_32250_, _32249_, _03810_);
  nor (_32251_, _32233_, _32228_);
  and (_32252_, _32251_, _02974_);
  or (_32253_, _32252_, _32250_);
  and (_32255_, _32253_, _02609_);
  nor (_32256_, _02609_, \oc8051_golden_model_1.SP [1]);
  or (_32257_, _32256_, _03069_);
  or (_32258_, _32257_, _32255_);
  nand (_32259_, _03069_, _03939_);
  and (_32260_, _32259_, _32258_);
  and (_32261_, _32260_, _03084_);
  and (_32262_, _32244_, _03075_);
  or (_32263_, _32262_, _32261_);
  and (_32264_, _32263_, _03941_);
  nor (_32266_, _10750_, _03940_);
  not (_32267_, _32266_);
  nor (_32268_, _32267_, _32264_);
  nand (_32269_, _10750_, \oc8051_golden_model_1.SP [1]);
  and (_32270_, _32269_, _05535_);
  not (_32271_, _32270_);
  nor (_32272_, _32271_, _32268_);
  or (_32273_, _10777_, _04000_);
  nor (_32274_, _32233_, _05535_);
  and (_32275_, _32274_, _32273_);
  nor (_32277_, _32275_, _02853_);
  not (_32278_, _32277_);
  nor (_32279_, _32278_, _32272_);
  and (_32280_, _04617_, _06151_);
  nor (_32281_, _32227_, _05540_);
  not (_32282_, _32281_);
  nor (_32283_, _32282_, _32280_);
  nor (_32284_, _32283_, _02579_);
  not (_32285_, _32284_);
  nor (_32286_, _32285_, _32279_);
  nor (_32288_, _32286_, _32241_);
  nor (_32289_, _32288_, _02802_);
  and (_32290_, _04617_, _03698_);
  not (_32291_, _32290_);
  nor (_32292_, _32233_, _02803_);
  and (_32293_, _32292_, _32291_);
  or (_32294_, _32293_, _32289_);
  and (_32295_, _32294_, _04093_);
  or (_32296_, _32295_, _32238_);
  and (_32297_, _32296_, _03887_);
  nor (_32299_, _11710_, _10777_);
  nor (_32300_, _32299_, _03887_);
  and (_32301_, _32300_, _32234_);
  nor (_32302_, _32301_, _32297_);
  nor (_32303_, _32302_, _03127_);
  nor (_32304_, _32303_, _32237_);
  nor (_32305_, _32304_, _02970_);
  nor (_32306_, _11709_, _10777_);
  nor (_32307_, _32306_, _03883_);
  and (_32308_, _32307_, _32234_);
  nor (_32310_, _32308_, _32305_);
  nor (_32311_, _32310_, _09689_);
  nor (_32312_, _02532_, \oc8051_golden_model_1.SP [1]);
  nor (_32313_, _32227_, _13722_);
  nor (_32314_, _32313_, _03137_);
  and (_32315_, _32314_, _32244_);
  nor (_32316_, _32315_, _32312_);
  not (_32317_, _32316_);
  nor (_32318_, _32317_, _32311_);
  or (_32319_, _32318_, _17961_);
  and (_32321_, _32290_, _05178_);
  nor (_32322_, _32321_, _05783_);
  and (_32323_, _32322_, _32234_);
  nand (_32324_, _32242_, _05178_);
  nor (_32325_, _32233_, _05788_);
  and (_32326_, _32325_, _32324_);
  nor (_32327_, _32326_, _32323_);
  and (_32328_, _32327_, _32319_);
  nor (_32329_, _32328_, _32231_);
  nor (_32330_, _29014_, \oc8051_golden_model_1.SP [1]);
  nor (_32332_, _32330_, _02892_);
  not (_32333_, _32332_);
  nor (_32334_, _32333_, _32329_);
  and (_32335_, _02892_, \oc8051_golden_model_1.SP [1]);
  nor (_32336_, _32335_, _03163_);
  not (_32337_, _32336_);
  nor (_32338_, _32337_, _32334_);
  and (_32339_, _32251_, _03163_);
  nor (_32340_, _32339_, _04337_);
  not (_32341_, _32340_);
  nor (_32343_, _32341_, _32338_);
  nor (_32344_, _03915_, _03700_);
  nor (_32345_, _32344_, _02888_);
  not (_32346_, _32345_);
  nor (_32347_, _32346_, _32343_);
  nor (_32348_, _32347_, _32230_);
  nor (_32349_, _32348_, _42672_);
  nor (_32350_, \oc8051_golden_model_1.SP [1], rst);
  nor (_32351_, _32350_, _00000_);
  or (_43545_, _32351_, _32349_);
  nor (_32353_, _13156_, _02529_);
  nor (_32354_, _13156_, _02532_);
  nor (_32355_, _32354_, _02965_);
  nor (_32356_, _04617_, _03335_);
  and (_32357_, _11927_, _04617_);
  nor (_32358_, _32357_, _32356_);
  nor (_32359_, _32358_, _03128_);
  and (_32360_, _13156_, _02514_);
  and (_32361_, _04617_, _04435_);
  or (_32362_, _32356_, _05535_);
  nor (_32363_, _32362_, _32361_);
  nor (_32364_, _13156_, _02614_);
  nor (_32365_, _11801_, _10777_);
  nor (_32366_, _32365_, _32356_);
  and (_32367_, _32366_, _02974_);
  and (_32368_, _04617_, \oc8051_golden_model_1.ACC [2]);
  nor (_32369_, _32368_, _32356_);
  or (_32370_, _32369_, _03814_);
  nand (_32371_, _09434_, \oc8051_golden_model_1.SP [2]);
  nor (_32372_, _13156_, _02611_);
  nor (_32374_, _32372_, _02974_);
  and (_32375_, _32374_, _32371_);
  and (_32376_, _32375_, _32370_);
  or (_32377_, _32376_, _04252_);
  nor (_32378_, _32377_, _32367_);
  nor (_32379_, _13156_, _02609_);
  nor (_32380_, _32379_, _32378_);
  nor (_32381_, _32380_, _03069_);
  nor (_32382_, _05393_, _03336_);
  or (_32383_, _32382_, _32381_);
  and (_32385_, _32383_, _03084_);
  nor (_32386_, _32369_, _03084_);
  or (_32387_, _32386_, _32385_);
  and (_32388_, _32387_, _03941_);
  or (_32389_, _32388_, _04365_);
  and (_32390_, _32389_, _02614_);
  or (_32391_, _32390_, _32364_);
  and (_32392_, _32391_, _04251_);
  and (_32393_, _04539_, _02581_);
  nor (_32394_, _32393_, _06770_);
  not (_32396_, _32394_);
  nor (_32397_, _32396_, _32392_);
  nor (_32398_, _32397_, _32363_);
  nor (_32399_, _32398_, _02853_);
  and (_32400_, _04617_, _06155_);
  nor (_32401_, _32356_, _05540_);
  not (_32402_, _32401_);
  nor (_32403_, _32402_, _32400_);
  or (_32404_, _32403_, _02579_);
  nor (_32405_, _32404_, _32399_);
  nor (_32407_, _11906_, _10777_);
  nor (_32408_, _32407_, _32356_);
  nor (_32409_, _32408_, _02838_);
  or (_32410_, _32409_, _02802_);
  or (_32411_, _32410_, _32405_);
  and (_32412_, _04617_, _05701_);
  nor (_32413_, _32412_, _32356_);
  nand (_32414_, _32413_, _02802_);
  and (_32415_, _32414_, _32411_);
  nor (_32416_, _32415_, _02514_);
  nor (_32418_, _32416_, _32360_);
  and (_32419_, _32418_, _03887_);
  and (_32420_, _11921_, _04617_);
  nor (_32421_, _32420_, _32356_);
  nor (_32422_, _32421_, _03887_);
  or (_32423_, _32422_, _32419_);
  and (_32424_, _32423_, _03128_);
  nor (_32425_, _32424_, _32359_);
  nor (_32426_, _32425_, _02970_);
  nor (_32427_, _32356_, _05130_);
  not (_32429_, _32427_);
  nor (_32430_, _32413_, _03883_);
  and (_32431_, _32430_, _32429_);
  nor (_32432_, _32431_, _32426_);
  nor (_32433_, _32432_, _09689_);
  nor (_32434_, _32369_, _03137_);
  and (_32435_, _32434_, _32429_);
  nor (_32436_, _32435_, _32433_);
  and (_32437_, _32436_, _32355_);
  nor (_32438_, _11919_, _10777_);
  nor (_32440_, _32438_, _32356_);
  and (_32441_, _32440_, _02965_);
  nor (_32442_, _32441_, _32437_);
  and (_32443_, _32442_, _05788_);
  nor (_32444_, _11926_, _10777_);
  nor (_32445_, _32444_, _32356_);
  nor (_32446_, _32445_, _05788_);
  or (_32447_, _32446_, _32443_);
  and (_32448_, _32447_, _09726_);
  and (_32449_, _13156_, _03145_);
  or (_32451_, _32449_, _32448_);
  and (_32452_, _32451_, _02529_);
  or (_32453_, _32452_, _32353_);
  and (_32454_, _32453_, _02893_);
  and (_32455_, _13156_, _02892_);
  or (_32456_, _32455_, _03163_);
  nor (_32457_, _32456_, _32454_);
  and (_32458_, _32366_, _03163_);
  nor (_32459_, _32458_, _04337_);
  not (_32460_, _32459_);
  nor (_32462_, _32460_, _32457_);
  nor (_32463_, _13156_, _03915_);
  nor (_32464_, _32463_, _02888_);
  not (_32465_, _32464_);
  nor (_32466_, _32465_, _32462_);
  and (_32467_, _11985_, _04617_);
  nor (_32468_, _32467_, _32356_);
  and (_32469_, _32468_, _02888_);
  nor (_32470_, _32469_, _32466_);
  and (_32471_, _32470_, _42668_);
  nor (_32473_, \oc8051_golden_model_1.SP [2], rst);
  nor (_32474_, _32473_, _00000_);
  or (_43546_, _32474_, _32471_);
  nor (_32475_, _04542_, _03915_);
  nor (_32476_, _04617_, _03068_);
  and (_32477_, _12133_, _04617_);
  nor (_32478_, _32477_, _32476_);
  nor (_32479_, _32478_, _03128_);
  and (_32480_, _12976_, _02514_);
  nor (_32481_, _12017_, _10777_);
  nor (_32482_, _32481_, _32476_);
  and (_32483_, _32482_, _02974_);
  and (_32484_, _04617_, \oc8051_golden_model_1.ACC [3]);
  nor (_32485_, _32484_, _32476_);
  or (_32486_, _32485_, _03814_);
  nand (_32487_, _09434_, \oc8051_golden_model_1.SP [3]);
  nor (_32488_, _12976_, _02611_);
  nor (_32489_, _32488_, _02974_);
  and (_32490_, _32489_, _32487_);
  and (_32491_, _32490_, _32486_);
  nor (_32494_, _32491_, _04252_);
  not (_32495_, _32494_);
  nor (_32496_, _32495_, _32483_);
  nor (_32497_, _12976_, _02609_);
  or (_32498_, _32497_, _03069_);
  nor (_32499_, _32498_, _32496_);
  and (_32500_, _05382_, _03069_);
  nor (_32501_, _32500_, _32499_);
  and (_32502_, _32501_, _03084_);
  nor (_32503_, _32485_, _03084_);
  or (_32505_, _32503_, _32502_);
  and (_32506_, _32505_, _03941_);
  nor (_32507_, _04289_, _10750_);
  not (_32508_, _32507_);
  nor (_32509_, _32508_, _32506_);
  nand (_32510_, _12976_, _10750_);
  and (_32511_, _32510_, _05535_);
  not (_32512_, _32511_);
  nor (_32513_, _32512_, _32509_);
  and (_32514_, _04617_, _04241_);
  nor (_32516_, _32514_, _32476_);
  nor (_32517_, _32516_, _05535_);
  nor (_32518_, _32517_, _02853_);
  not (_32519_, _32518_);
  nor (_32520_, _32519_, _32513_);
  and (_32521_, _04617_, _06154_);
  nor (_32522_, _32476_, _05540_);
  not (_32523_, _32522_);
  nor (_32524_, _32523_, _32521_);
  or (_32525_, _32524_, _02579_);
  nor (_32527_, _32525_, _32520_);
  nor (_32528_, _12112_, _10777_);
  nor (_32529_, _32528_, _32476_);
  nor (_32530_, _32529_, _02838_);
  or (_32531_, _32530_, _02802_);
  or (_32532_, _32531_, _32527_);
  and (_32533_, _04617_, _05658_);
  nor (_32534_, _32533_, _32476_);
  nand (_32535_, _32534_, _02802_);
  and (_32536_, _32535_, _32532_);
  nor (_32538_, _32536_, _02514_);
  nor (_32539_, _32538_, _32480_);
  and (_32540_, _32539_, _03887_);
  and (_32541_, _12127_, _04617_);
  nor (_32542_, _32541_, _32476_);
  nor (_32543_, _32542_, _03887_);
  or (_32544_, _32543_, _32540_);
  and (_32545_, _32544_, _03128_);
  nor (_32546_, _32545_, _32479_);
  nor (_32547_, _32546_, _02970_);
  nor (_32549_, _32476_, _05079_);
  not (_32550_, _32549_);
  nor (_32551_, _32534_, _03883_);
  and (_32552_, _32551_, _32550_);
  nor (_32553_, _32552_, _32547_);
  nor (_32554_, _32553_, _09689_);
  nor (_32555_, _12976_, _02532_);
  or (_32556_, _32549_, _03137_);
  nor (_32557_, _32556_, _32485_);
  nor (_32558_, _32557_, _32555_);
  and (_32560_, _32558_, _05783_);
  not (_32561_, _32560_);
  nor (_32562_, _32561_, _32554_);
  nor (_32563_, _12125_, _10777_);
  or (_32564_, _32476_, _05783_);
  nor (_32565_, _32564_, _32563_);
  nor (_32566_, _32565_, _32562_);
  and (_32567_, _32566_, _05788_);
  nor (_32568_, _12132_, _10777_);
  nor (_32569_, _32568_, _32476_);
  nor (_32571_, _32569_, _05788_);
  or (_32572_, _32571_, _32567_);
  and (_32573_, _32572_, _09726_);
  nor (_32574_, _05379_, _03068_);
  nor (_32575_, _32574_, _05380_);
  and (_32576_, _32575_, _02529_);
  nor (_32577_, _32576_, _29014_);
  nor (_32578_, _32577_, _32573_);
  nor (_32579_, _04542_, _02529_);
  nor (_32580_, _32579_, _32578_);
  and (_32582_, _32580_, _02893_);
  nor (_32583_, _32575_, _02893_);
  or (_32584_, _32583_, _32582_);
  and (_32585_, _32584_, _03906_);
  nor (_32586_, _32482_, _03906_);
  nor (_32587_, _32586_, _04337_);
  not (_32588_, _32587_);
  nor (_32589_, _32588_, _32585_);
  nor (_32590_, _32589_, _32475_);
  and (_32591_, _32590_, _02890_);
  and (_32593_, _12183_, _04617_);
  nor (_32594_, _32593_, _32476_);
  nor (_32595_, _32594_, _02890_);
  or (_32596_, _32595_, _32591_);
  or (_32597_, _32596_, _42672_);
  or (_32598_, _42668_, \oc8051_golden_model_1.SP [3]);
  and (_32599_, _32598_, _43998_);
  and (_43547_, _32599_, _32597_);
  nor (_32600_, _04247_, \oc8051_golden_model_1.SP [4]);
  nor (_32601_, _32600_, _10701_);
  nor (_32603_, _32601_, _03915_);
  nor (_32604_, _04617_, _10734_);
  and (_32605_, _12207_, _04617_);
  nor (_32606_, _32605_, _32604_);
  nor (_32607_, _32606_, _03128_);
  nor (_32608_, _12217_, _10777_);
  nor (_32609_, _32608_, _32604_);
  and (_32610_, _32609_, _02974_);
  and (_32611_, _04617_, \oc8051_golden_model_1.ACC [4]);
  nor (_32612_, _32611_, _32604_);
  or (_32614_, _32612_, _03814_);
  nand (_32615_, _09434_, \oc8051_golden_model_1.SP [4]);
  not (_32616_, _32601_);
  nor (_32617_, _32616_, _02611_);
  nor (_32618_, _32617_, _02974_);
  and (_32619_, _32618_, _32615_);
  and (_32620_, _32619_, _32614_);
  nor (_32621_, _32620_, _04252_);
  not (_32622_, _32621_);
  nor (_32623_, _32622_, _32610_);
  nor (_32625_, _32616_, _02609_);
  or (_32626_, _32625_, _03069_);
  nor (_32627_, _32626_, _32623_);
  and (_32628_, _10735_, _02866_);
  nor (_32629_, _05381_, _10734_);
  nor (_32630_, _32629_, _32628_);
  and (_32631_, _32630_, _03069_);
  nor (_32632_, _32631_, _32627_);
  and (_32633_, _32632_, _03084_);
  nor (_32634_, _32612_, _03084_);
  or (_32636_, _32634_, _32633_);
  and (_32637_, _32636_, _03941_);
  nor (_32638_, _04248_, _10734_);
  and (_32639_, _04248_, _10734_);
  nor (_32640_, _32639_, _32638_);
  and (_32641_, _32640_, _02875_);
  nor (_32642_, _32641_, _10750_);
  not (_32643_, _32642_);
  nor (_32644_, _32643_, _32637_);
  nand (_32645_, _32616_, _10750_);
  and (_32647_, _32645_, _05535_);
  not (_32648_, _32647_);
  nor (_32649_, _32648_, _32644_);
  and (_32650_, _04617_, _04982_);
  nor (_32651_, _32650_, _32604_);
  nor (_32652_, _32651_, _05535_);
  nor (_32653_, _32652_, _02853_);
  not (_32654_, _32653_);
  nor (_32655_, _32654_, _32649_);
  and (_32656_, _04617_, _06159_);
  nor (_32658_, _32604_, _05540_);
  not (_32659_, _32658_);
  nor (_32660_, _32659_, _32656_);
  or (_32661_, _32660_, _02579_);
  nor (_32662_, _32661_, _32655_);
  nor (_32663_, _12321_, _10777_);
  nor (_32664_, _32663_, _32604_);
  nor (_32665_, _32664_, _02838_);
  or (_32666_, _32665_, _02802_);
  or (_32667_, _32666_, _32662_);
  and (_32669_, _05666_, _04617_);
  nor (_32670_, _32669_, _32604_);
  nand (_32671_, _32670_, _02802_);
  and (_32672_, _32671_, _32667_);
  nor (_32673_, _32672_, _02514_);
  and (_32674_, _32616_, _02514_);
  nor (_32675_, _32674_, _32673_);
  and (_32676_, _32675_, _03887_);
  and (_32677_, _12211_, _04617_);
  nor (_32678_, _32677_, _32604_);
  nor (_32680_, _32678_, _03887_);
  or (_32681_, _32680_, _32676_);
  and (_32682_, _32681_, _03128_);
  nor (_32683_, _32682_, _32607_);
  nor (_32684_, _32683_, _02970_);
  nor (_32685_, _32604_, _05031_);
  not (_32686_, _32685_);
  nor (_32687_, _32670_, _03883_);
  and (_32688_, _32687_, _32686_);
  nor (_32689_, _32688_, _32684_);
  nor (_32691_, _32689_, _09689_);
  nor (_32692_, _32612_, _03137_);
  and (_32693_, _32692_, _32686_);
  nor (_32694_, _32616_, _02532_);
  nor (_32695_, _32694_, _32693_);
  and (_32696_, _32695_, _05783_);
  not (_32697_, _32696_);
  nor (_32698_, _32697_, _32691_);
  nor (_32699_, _12209_, _10777_);
  or (_32700_, _32604_, _05783_);
  nor (_32702_, _32700_, _32699_);
  nor (_32703_, _32702_, _32698_);
  and (_32704_, _32703_, _05788_);
  nor (_32705_, _12206_, _10777_);
  nor (_32706_, _32705_, _32604_);
  nor (_32707_, _32706_, _05788_);
  or (_32708_, _32707_, _32704_);
  and (_32709_, _32708_, _09726_);
  nor (_32710_, _05380_, _10734_);
  nor (_32711_, _32710_, _10735_);
  and (_32713_, _32711_, _02529_);
  nor (_32714_, _32713_, _29014_);
  nor (_32715_, _32714_, _32709_);
  nor (_32716_, _32601_, _02529_);
  nor (_32717_, _32716_, _32715_);
  and (_32718_, _32717_, _02893_);
  nor (_32719_, _32711_, _02893_);
  or (_32720_, _32719_, _32718_);
  and (_32721_, _32720_, _03906_);
  nor (_32722_, _32609_, _03906_);
  nor (_32724_, _32722_, _04337_);
  not (_32725_, _32724_);
  nor (_32726_, _32725_, _32721_);
  nor (_32727_, _32726_, _32603_);
  and (_32728_, _32727_, _02890_);
  and (_32729_, _12389_, _04617_);
  nor (_32730_, _32729_, _32604_);
  nor (_32731_, _32730_, _02890_);
  or (_32732_, _32731_, _32728_);
  or (_32733_, _32732_, _42672_);
  or (_32735_, _42668_, \oc8051_golden_model_1.SP [4]);
  and (_32736_, _32735_, _43998_);
  and (_43548_, _32736_, _32733_);
  nor (_32737_, _10701_, \oc8051_golden_model_1.SP [5]);
  nor (_32738_, _32737_, _10702_);
  nor (_32739_, _32738_, _03915_);
  nor (_32740_, _04617_, _10733_);
  and (_32741_, _12411_, _04617_);
  nor (_32742_, _32741_, _32740_);
  nor (_32743_, _32742_, _03128_);
  nor (_32745_, _12407_, _10777_);
  nor (_32746_, _32745_, _32740_);
  and (_32747_, _32746_, _02974_);
  and (_32748_, _04617_, \oc8051_golden_model_1.ACC [5]);
  nor (_32749_, _32748_, _32740_);
  or (_32750_, _32749_, _03814_);
  nand (_32751_, _09434_, \oc8051_golden_model_1.SP [5]);
  not (_32752_, _32738_);
  nor (_32753_, _32752_, _02611_);
  nor (_32754_, _32753_, _02974_);
  and (_32756_, _32754_, _32751_);
  and (_32757_, _32756_, _32750_);
  nor (_32758_, _32757_, _04252_);
  not (_32759_, _32758_);
  nor (_32760_, _32759_, _32747_);
  nor (_32761_, _32752_, _02609_);
  or (_32762_, _32761_, _32760_);
  and (_32763_, _32762_, _03336_);
  and (_32764_, _10736_, _02866_);
  nor (_32765_, _32628_, _10733_);
  nor (_32767_, _32765_, _32764_);
  nor (_32768_, _32767_, _03336_);
  or (_32769_, _32768_, _32763_);
  and (_32770_, _32769_, _03084_);
  nor (_32771_, _32749_, _03084_);
  or (_32772_, _32771_, _32770_);
  and (_32773_, _32772_, _03941_);
  and (_32774_, _10702_, \oc8051_golden_model_1.SP [0]);
  nor (_32775_, _32638_, \oc8051_golden_model_1.SP [5]);
  nor (_32776_, _32775_, _32774_);
  and (_32778_, _32776_, _02875_);
  nor (_32779_, _32778_, _10750_);
  not (_32780_, _32779_);
  nor (_32781_, _32780_, _32773_);
  nand (_32782_, _32752_, _10750_);
  and (_32783_, _32782_, _05535_);
  not (_32784_, _32783_);
  nor (_32785_, _32784_, _32781_);
  and (_32786_, _04617_, _04877_);
  nor (_32787_, _32786_, _32740_);
  nor (_32788_, _32787_, _05535_);
  nor (_32789_, _32788_, _02853_);
  not (_32790_, _32789_);
  nor (_32791_, _32790_, _32785_);
  and (_32792_, _04617_, _06158_);
  nor (_32793_, _32740_, _05540_);
  not (_32794_, _32793_);
  nor (_32795_, _32794_, _32792_);
  or (_32796_, _32795_, _02579_);
  nor (_32797_, _32796_, _32791_);
  nor (_32800_, _12527_, _10777_);
  nor (_32801_, _32800_, _32740_);
  nor (_32802_, _32801_, _02838_);
  or (_32803_, _32802_, _02802_);
  or (_32804_, _32803_, _32797_);
  and (_32805_, _05614_, _04617_);
  nor (_32806_, _32805_, _32740_);
  nand (_32807_, _32806_, _02802_);
  and (_32808_, _32807_, _32804_);
  nor (_32809_, _32808_, _02514_);
  and (_32811_, _32752_, _02514_);
  nor (_32812_, _32811_, _32809_);
  and (_32813_, _32812_, _03887_);
  and (_32814_, _12415_, _04617_);
  nor (_32815_, _32814_, _32740_);
  nor (_32816_, _32815_, _03887_);
  or (_32817_, _32816_, _32813_);
  and (_32818_, _32817_, _03128_);
  nor (_32819_, _32818_, _32743_);
  nor (_32820_, _32819_, _02970_);
  nor (_32822_, _32740_, _04924_);
  not (_32823_, _32822_);
  nor (_32824_, _32806_, _03883_);
  and (_32825_, _32824_, _32823_);
  nor (_32826_, _32825_, _32820_);
  nor (_32827_, _32826_, _09689_);
  nor (_32828_, _32749_, _03137_);
  and (_32829_, _32828_, _32823_);
  nor (_32830_, _32752_, _02532_);
  nor (_32831_, _32830_, _32829_);
  and (_32833_, _32831_, _05783_);
  not (_32834_, _32833_);
  nor (_32835_, _32834_, _32827_);
  nor (_32836_, _12413_, _10777_);
  or (_32837_, _32740_, _05783_);
  nor (_32838_, _32837_, _32836_);
  nor (_32839_, _32838_, _32835_);
  and (_32840_, _32839_, _05788_);
  nor (_32841_, _12410_, _10777_);
  nor (_32842_, _32841_, _32740_);
  nor (_32844_, _32842_, _05788_);
  or (_32845_, _32844_, _32840_);
  and (_32846_, _32845_, _09726_);
  nor (_32847_, _10735_, _10733_);
  nor (_32848_, _32847_, _10736_);
  and (_32849_, _32848_, _02529_);
  nor (_32850_, _32849_, _29014_);
  nor (_32851_, _32850_, _32846_);
  nor (_32852_, _32738_, _02529_);
  nor (_32853_, _32852_, _32851_);
  and (_32855_, _32853_, _02893_);
  nor (_32856_, _32848_, _02893_);
  or (_32857_, _32856_, _32855_);
  and (_32858_, _32857_, _03906_);
  nor (_32859_, _32746_, _03906_);
  nor (_32860_, _32859_, _04337_);
  not (_32861_, _32860_);
  nor (_32862_, _32861_, _32858_);
  nor (_32863_, _32862_, _32739_);
  nor (_32864_, _32863_, _02888_);
  and (_32866_, _12589_, _04617_);
  nor (_32867_, _32866_, _32740_);
  and (_32868_, _32867_, _02888_);
  nor (_32869_, _32868_, _32864_);
  or (_32870_, _32869_, _42672_);
  or (_32871_, _42668_, \oc8051_golden_model_1.SP [5]);
  and (_32872_, _32871_, _43998_);
  and (_43549_, _32872_, _32870_);
  nor (_32873_, _04617_, _10732_);
  and (_32874_, _12613_, _04617_);
  nor (_32876_, _32874_, _32873_);
  nor (_32877_, _32876_, _03128_);
  and (_32878_, _04617_, _05849_);
  or (_32879_, _32878_, _32873_);
  and (_32880_, _32879_, _02853_);
  nor (_32881_, _12603_, _10777_);
  nor (_32882_, _32881_, _32873_);
  and (_32883_, _32882_, _02974_);
  and (_32884_, _04617_, \oc8051_golden_model_1.ACC [6]);
  nor (_32885_, _32884_, _32873_);
  or (_32887_, _32885_, _03814_);
  nand (_32888_, _09434_, \oc8051_golden_model_1.SP [6]);
  nor (_32889_, _10702_, \oc8051_golden_model_1.SP [6]);
  nor (_32890_, _32889_, _10703_);
  not (_32891_, _32890_);
  nor (_32892_, _32891_, _02611_);
  nor (_32893_, _32892_, _02974_);
  and (_32894_, _32893_, _32888_);
  and (_32895_, _32894_, _32887_);
  nor (_32896_, _32895_, _04252_);
  not (_32898_, _32896_);
  nor (_32899_, _32898_, _32883_);
  nor (_32900_, _32891_, _02609_);
  or (_32901_, _32900_, _03069_);
  nor (_32902_, _32901_, _32899_);
  nor (_32903_, _32764_, _10732_);
  nor (_32904_, _32903_, _10739_);
  and (_32905_, _32904_, _03069_);
  nor (_32906_, _32905_, _32902_);
  and (_32907_, _32906_, _03084_);
  nor (_32909_, _32885_, _03084_);
  or (_32910_, _32909_, _32907_);
  and (_32911_, _32910_, _03941_);
  nor (_32912_, _32774_, \oc8051_golden_model_1.SP [6]);
  nor (_32913_, _32912_, _10751_);
  and (_32914_, _32913_, _02875_);
  nor (_32915_, _32914_, _32911_);
  nor (_32916_, _32915_, _10750_);
  nand (_32917_, _32890_, _10750_);
  and (_32918_, _32917_, _05535_);
  not (_32920_, _32918_);
  nor (_32921_, _32920_, _32916_);
  and (_32922_, _04617_, _04770_);
  or (_32923_, _32873_, _05535_);
  nor (_32924_, _32923_, _32922_);
  or (_32925_, _32924_, _02853_);
  nor (_32926_, _32925_, _32921_);
  or (_32927_, _32926_, _32880_);
  and (_32928_, _32927_, _02838_);
  nor (_32929_, _12722_, _10777_);
  nor (_32931_, _32929_, _32873_);
  nor (_32932_, _32931_, _02838_);
  or (_32933_, _32932_, _02802_);
  or (_32934_, _32933_, _32928_);
  and (_32935_, _12729_, _04617_);
  nor (_32936_, _32935_, _32873_);
  nand (_32937_, _32936_, _02802_);
  and (_32938_, _32937_, _32934_);
  nor (_32939_, _32938_, _02514_);
  and (_32940_, _32891_, _02514_);
  nor (_32942_, _32940_, _32939_);
  and (_32943_, _32942_, _03887_);
  and (_32944_, _12739_, _04617_);
  nor (_32945_, _32944_, _32873_);
  nor (_32946_, _32945_, _03887_);
  or (_32947_, _32946_, _32943_);
  and (_32948_, _32947_, _03128_);
  nor (_32949_, _32948_, _32877_);
  nor (_32950_, _32949_, _02970_);
  nor (_32951_, _32873_, _04819_);
  not (_32953_, _32951_);
  nor (_32954_, _32936_, _03883_);
  and (_32955_, _32954_, _32953_);
  nor (_32956_, _32955_, _32950_);
  nor (_32957_, _32956_, _09689_);
  nor (_32958_, _32885_, _03137_);
  and (_32959_, _32958_, _32953_);
  nor (_32960_, _32891_, _02532_);
  nor (_32961_, _32960_, _32959_);
  and (_32962_, _32961_, _05783_);
  not (_32964_, _32962_);
  nor (_32965_, _32964_, _32957_);
  nor (_32966_, _12737_, _10777_);
  nor (_32967_, _32966_, _32873_);
  and (_32968_, _32967_, _02965_);
  nor (_32969_, _32968_, _32965_);
  and (_32970_, _32969_, _05788_);
  nor (_32971_, _12612_, _10777_);
  nor (_32972_, _32971_, _32873_);
  nor (_32973_, _32972_, _05788_);
  or (_32975_, _32973_, _32970_);
  and (_32976_, _32975_, _09726_);
  nor (_32977_, _10736_, _10732_);
  nor (_32978_, _32977_, _10738_);
  not (_32979_, _32978_);
  and (_32980_, _32979_, _03145_);
  or (_32981_, _32980_, _03898_);
  nor (_32982_, _32981_, _32976_);
  nor (_32983_, _32890_, _02529_);
  or (_32984_, _32983_, _02892_);
  nor (_32986_, _32984_, _32982_);
  and (_32987_, _32979_, _02892_);
  or (_32988_, _32987_, _03163_);
  nor (_32989_, _32988_, _32986_);
  and (_32990_, _32882_, _03163_);
  nor (_32991_, _32990_, _04337_);
  not (_32992_, _32991_);
  nor (_32993_, _32992_, _32989_);
  nor (_32994_, _32891_, _03915_);
  nor (_32995_, _32994_, _02888_);
  not (_32997_, _32995_);
  nor (_32998_, _32997_, _32993_);
  and (_32999_, _12794_, _04617_);
  or (_33000_, _32873_, _02890_);
  nor (_33001_, _33000_, _32999_);
  nor (_33002_, _33001_, _32998_);
  or (_33003_, _33002_, _42672_);
  or (_33004_, _42668_, \oc8051_golden_model_1.SP [6]);
  and (_33005_, _33004_, _43998_);
  and (_43550_, _33005_, _33003_);
  not (_33007_, \oc8051_golden_model_1.TCON [0]);
  nor (_33008_, _04622_, _33007_);
  and (_33009_, _11522_, _04622_);
  nor (_33010_, _33009_, _33008_);
  nor (_33011_, _33010_, _03128_);
  and (_33012_, _04622_, _03808_);
  nor (_33013_, _33012_, _33008_);
  and (_33014_, _33013_, _06770_);
  and (_33015_, _04622_, \oc8051_golden_model_1.ACC [0]);
  nor (_33016_, _33015_, _33008_);
  nor (_33018_, _33016_, _03814_);
  nor (_33019_, _03813_, _33007_);
  or (_33020_, _33019_, _33018_);
  and (_33021_, _33020_, _03810_);
  and (_33022_, _05226_, _04622_);
  nor (_33023_, _33022_, _33008_);
  nor (_33024_, _33023_, _03810_);
  or (_33025_, _33024_, _33021_);
  and (_33026_, _33025_, _02881_);
  nor (_33027_, _05320_, _33007_);
  and (_33029_, _11417_, _05320_);
  nor (_33030_, _33029_, _33027_);
  nor (_33031_, _33030_, _02881_);
  nor (_33032_, _33031_, _33026_);
  nor (_33033_, _33032_, _03069_);
  nor (_33034_, _33013_, _03336_);
  or (_33035_, _33034_, _33033_);
  and (_33036_, _33035_, _03084_);
  nor (_33037_, _33016_, _03084_);
  or (_33038_, _33037_, _33036_);
  and (_33040_, _33038_, _02877_);
  and (_33041_, _33008_, _02876_);
  or (_33042_, _33041_, _33040_);
  and (_33043_, _33042_, _02870_);
  nor (_33044_, _33023_, _02870_);
  or (_33045_, _33044_, _33043_);
  and (_33046_, _33045_, _02864_);
  nor (_33047_, _11448_, _10889_);
  nor (_33048_, _33047_, _33027_);
  nor (_33049_, _33048_, _02864_);
  or (_33051_, _33049_, _06770_);
  nor (_33052_, _33051_, _33046_);
  nor (_33053_, _33052_, _33014_);
  nor (_33054_, _33053_, _02853_);
  and (_33055_, _04622_, _06152_);
  nor (_33056_, _33008_, _05540_);
  not (_33057_, _33056_);
  nor (_33058_, _33057_, _33055_);
  or (_33059_, _33058_, _02579_);
  nor (_33060_, _33059_, _33054_);
  nor (_33062_, _11505_, _10905_);
  nor (_33063_, _33062_, _33008_);
  nor (_33064_, _33063_, _02838_);
  or (_33065_, _33064_, _02802_);
  or (_33066_, _33065_, _33060_);
  and (_33067_, _04622_, _05672_);
  nor (_33068_, _33067_, _33008_);
  nand (_33069_, _33068_, _02802_);
  and (_33070_, _33069_, _33066_);
  and (_33071_, _33070_, _03887_);
  and (_33073_, _11399_, _04622_);
  nor (_33074_, _33073_, _33008_);
  nor (_33075_, _33074_, _03887_);
  or (_33076_, _33075_, _33071_);
  and (_33077_, _33076_, _03128_);
  nor (_33078_, _33077_, _33011_);
  nor (_33079_, _33078_, _02970_);
  nor (_33080_, _33068_, _03883_);
  not (_33081_, _33080_);
  nor (_33082_, _33081_, _33022_);
  nor (_33084_, _33082_, _33079_);
  nor (_33085_, _33084_, _03135_);
  nor (_33086_, _33008_, _09409_);
  or (_33087_, _33086_, _03137_);
  nor (_33088_, _33087_, _33016_);
  or (_33089_, _33088_, _33085_);
  and (_33090_, _33089_, _05783_);
  nor (_33091_, _11396_, _10905_);
  nor (_33092_, _33091_, _33008_);
  nor (_33093_, _33092_, _05783_);
  or (_33095_, _33093_, _33090_);
  and (_33096_, _33095_, _05788_);
  nor (_33097_, _11520_, _10905_);
  nor (_33098_, _33097_, _33008_);
  nor (_33099_, _33098_, _05788_);
  or (_33100_, _33099_, _33096_);
  and (_33101_, _33100_, _03906_);
  nor (_33102_, _33023_, _03906_);
  or (_33103_, _33102_, _33101_);
  and (_33104_, _33103_, _02498_);
  and (_33106_, _33008_, _02497_);
  or (_33107_, _33106_, _33104_);
  and (_33108_, _33107_, _02890_);
  nor (_33109_, _33023_, _02890_);
  or (_33110_, _33109_, _33108_);
  or (_33111_, _33110_, _42672_);
  or (_33112_, _42668_, \oc8051_golden_model_1.TCON [0]);
  and (_33113_, _33112_, _43998_);
  and (_43552_, _33113_, _33111_);
  nand (_33114_, _04622_, _03698_);
  or (_33116_, _04622_, \oc8051_golden_model_1.TCON [1]);
  and (_33117_, _33116_, _02802_);
  and (_33118_, _33117_, _33114_);
  nand (_33119_, _11695_, _04622_);
  and (_33120_, _33116_, _02579_);
  and (_33121_, _33120_, _33119_);
  not (_33122_, \oc8051_golden_model_1.TCON [1]);
  nor (_33123_, _04622_, _33122_);
  and (_33124_, _04622_, _04000_);
  or (_33125_, _33124_, _33123_);
  or (_33127_, _33125_, _03336_);
  and (_33128_, _11606_, _04622_);
  not (_33129_, _33128_);
  and (_33130_, _33129_, _33116_);
  or (_33131_, _33130_, _03810_);
  nand (_33132_, _04622_, _02551_);
  and (_33133_, _33132_, _33116_);
  and (_33134_, _33133_, _03813_);
  nor (_33135_, _03813_, _33122_);
  or (_33136_, _33135_, _02974_);
  or (_33137_, _33136_, _33134_);
  and (_33138_, _33137_, _02881_);
  and (_33139_, _33138_, _33131_);
  nor (_33140_, _05320_, _33122_);
  and (_33141_, _11592_, _05320_);
  or (_33142_, _33141_, _33140_);
  and (_33143_, _33142_, _02880_);
  or (_33144_, _33143_, _03069_);
  or (_33145_, _33144_, _33139_);
  and (_33146_, _33145_, _33127_);
  or (_33148_, _33146_, _03075_);
  or (_33149_, _33133_, _03084_);
  and (_33150_, _33149_, _02877_);
  and (_33151_, _33150_, _33148_);
  and (_33152_, _11595_, _05320_);
  or (_33153_, _33152_, _33140_);
  and (_33154_, _33153_, _02876_);
  or (_33155_, _33154_, _02869_);
  or (_33156_, _33155_, _33151_);
  and (_33157_, _33141_, _11591_);
  or (_33159_, _33140_, _02870_);
  or (_33160_, _33159_, _33157_);
  and (_33161_, _33160_, _33156_);
  and (_33162_, _33161_, _02864_);
  nor (_33163_, _11638_, _10889_);
  or (_33164_, _33140_, _33163_);
  and (_33165_, _33164_, _02863_);
  or (_33166_, _33165_, _06770_);
  or (_33167_, _33166_, _33162_);
  or (_33168_, _33125_, _05535_);
  and (_33170_, _33168_, _33167_);
  or (_33171_, _33170_, _02853_);
  and (_33172_, _04622_, _06151_);
  or (_33173_, _33123_, _05540_);
  or (_33174_, _33173_, _33172_);
  and (_33175_, _33174_, _02838_);
  and (_33176_, _33175_, _33171_);
  or (_33177_, _33176_, _33121_);
  and (_33178_, _33177_, _02803_);
  or (_33179_, _33178_, _33118_);
  and (_33181_, _33179_, _03887_);
  or (_33182_, _11710_, _10905_);
  and (_33183_, _33116_, _02980_);
  and (_33184_, _33183_, _33182_);
  or (_33185_, _33184_, _33181_);
  and (_33186_, _33185_, _03128_);
  or (_33187_, _11715_, _10905_);
  and (_33188_, _33116_, _03127_);
  and (_33189_, _33188_, _33187_);
  or (_33190_, _33189_, _33186_);
  and (_33192_, _33190_, _03883_);
  or (_33193_, _11709_, _10905_);
  and (_33194_, _33116_, _02970_);
  and (_33195_, _33194_, _33193_);
  or (_33196_, _33195_, _33192_);
  and (_33197_, _33196_, _03137_);
  or (_33198_, _33123_, _13722_);
  and (_33199_, _33133_, _03135_);
  and (_33200_, _33199_, _33198_);
  or (_33201_, _33200_, _33197_);
  and (_33203_, _33201_, _03124_);
  or (_33204_, _33132_, _13722_);
  and (_33205_, _33116_, _03123_);
  and (_33206_, _33205_, _33204_);
  or (_33207_, _33206_, _03163_);
  or (_33208_, _33114_, _13722_);
  and (_33209_, _33116_, _02965_);
  and (_33210_, _33209_, _33208_);
  or (_33211_, _33210_, _33207_);
  or (_33212_, _33211_, _33203_);
  or (_33214_, _33130_, _03906_);
  and (_33215_, _33214_, _02498_);
  and (_33216_, _33215_, _33212_);
  and (_33217_, _33153_, _02497_);
  or (_33218_, _33217_, _02888_);
  or (_33219_, _33218_, _33216_);
  or (_33220_, _33128_, _33123_);
  or (_33221_, _33220_, _02890_);
  and (_33222_, _33221_, _33219_);
  or (_33223_, _33222_, _42672_);
  or (_33225_, _42668_, \oc8051_golden_model_1.TCON [1]);
  and (_33226_, _33225_, _43998_);
  and (_43553_, _33226_, _33223_);
  not (_33227_, \oc8051_golden_model_1.TCON [2]);
  nor (_33228_, _04622_, _33227_);
  and (_33229_, _11927_, _04622_);
  nor (_33230_, _33229_, _33228_);
  nor (_33231_, _33230_, _03128_);
  and (_33232_, _04622_, _04435_);
  nor (_33233_, _33232_, _33228_);
  and (_33235_, _33233_, _06770_);
  and (_33236_, _04622_, \oc8051_golden_model_1.ACC [2]);
  nor (_33237_, _33236_, _33228_);
  nor (_33238_, _33237_, _03814_);
  nor (_33239_, _03813_, _33227_);
  or (_33240_, _33239_, _33238_);
  and (_33241_, _33240_, _03810_);
  nor (_33242_, _11801_, _10905_);
  nor (_33243_, _33242_, _33228_);
  nor (_33244_, _33243_, _03810_);
  or (_33246_, _33244_, _33241_);
  and (_33247_, _33246_, _02881_);
  nor (_33248_, _05320_, _33227_);
  and (_33249_, _11815_, _05320_);
  nor (_33250_, _33249_, _33248_);
  nor (_33251_, _33250_, _02881_);
  or (_33252_, _33251_, _33247_);
  and (_33253_, _33252_, _03336_);
  nor (_33254_, _33233_, _03336_);
  or (_33255_, _33254_, _33253_);
  and (_33257_, _33255_, _03084_);
  nor (_33258_, _33237_, _03084_);
  or (_33259_, _33258_, _33257_);
  and (_33260_, _33259_, _02877_);
  and (_33261_, _11797_, _05320_);
  nor (_33262_, _33261_, _33248_);
  nor (_33263_, _33262_, _02877_);
  or (_33264_, _33263_, _02869_);
  or (_33265_, _33264_, _33260_);
  and (_33266_, _33249_, _11830_);
  or (_33268_, _33248_, _02870_);
  or (_33269_, _33268_, _33266_);
  and (_33270_, _33269_, _02864_);
  and (_33271_, _33270_, _33265_);
  nor (_33272_, _11848_, _10889_);
  nor (_33273_, _33272_, _33248_);
  nor (_33274_, _33273_, _02864_);
  nor (_33275_, _33274_, _06770_);
  not (_33276_, _33275_);
  nor (_33277_, _33276_, _33271_);
  nor (_33279_, _33277_, _33235_);
  nor (_33280_, _33279_, _02853_);
  and (_33281_, _04622_, _06155_);
  nor (_33282_, _33228_, _05540_);
  not (_33283_, _33282_);
  nor (_33284_, _33283_, _33281_);
  or (_33285_, _33284_, _02579_);
  nor (_33286_, _33285_, _33280_);
  nor (_33287_, _11906_, _10905_);
  nor (_33288_, _33287_, _33228_);
  nor (_33290_, _33288_, _02838_);
  or (_33291_, _33290_, _02802_);
  or (_33292_, _33291_, _33286_);
  and (_33293_, _04622_, _05701_);
  nor (_33294_, _33293_, _33228_);
  nand (_33295_, _33294_, _02802_);
  and (_33296_, _33295_, _33292_);
  and (_33297_, _33296_, _03887_);
  and (_33298_, _11921_, _04622_);
  nor (_33299_, _33298_, _33228_);
  nor (_33301_, _33299_, _03887_);
  or (_33302_, _33301_, _33297_);
  and (_33303_, _33302_, _03128_);
  nor (_33304_, _33303_, _33231_);
  nor (_33305_, _33304_, _02970_);
  nor (_33306_, _33228_, _05130_);
  not (_33307_, _33306_);
  nor (_33308_, _33294_, _03883_);
  and (_33309_, _33308_, _33307_);
  nor (_33310_, _33309_, _33305_);
  nor (_33312_, _33310_, _03135_);
  nor (_33313_, _33237_, _03137_);
  and (_33314_, _33313_, _33307_);
  nor (_33315_, _33314_, _02965_);
  not (_33316_, _33315_);
  nor (_33317_, _33316_, _33312_);
  nor (_33318_, _11919_, _10905_);
  or (_33319_, _33228_, _05783_);
  nor (_33320_, _33319_, _33318_);
  or (_33321_, _33320_, _03123_);
  nor (_33323_, _33321_, _33317_);
  nor (_33324_, _11926_, _10905_);
  nor (_33325_, _33324_, _33228_);
  nor (_33326_, _33325_, _05788_);
  or (_33327_, _33326_, _33323_);
  and (_33328_, _33327_, _03906_);
  nor (_33329_, _33243_, _03906_);
  or (_33330_, _33329_, _33328_);
  and (_33331_, _33330_, _02498_);
  nor (_33332_, _33262_, _02498_);
  or (_33334_, _33332_, _33331_);
  and (_33335_, _33334_, _02890_);
  and (_33336_, _11985_, _04622_);
  nor (_33337_, _33336_, _33228_);
  nor (_33338_, _33337_, _02890_);
  or (_33339_, _33338_, _33335_);
  or (_33340_, _33339_, _42672_);
  or (_33341_, _42668_, \oc8051_golden_model_1.TCON [2]);
  and (_33342_, _33341_, _43998_);
  and (_43554_, _33342_, _33340_);
  not (_33344_, \oc8051_golden_model_1.TCON [3]);
  nor (_33345_, _04622_, _33344_);
  and (_33346_, _12133_, _04622_);
  nor (_33347_, _33346_, _33345_);
  nor (_33348_, _33347_, _03128_);
  and (_33349_, _04622_, _04241_);
  nor (_33350_, _33349_, _33345_);
  and (_33351_, _33350_, _06770_);
  and (_33352_, _04622_, \oc8051_golden_model_1.ACC [3]);
  nor (_33353_, _33352_, _33345_);
  nor (_33355_, _33353_, _03814_);
  nor (_33356_, _03813_, _33344_);
  or (_33357_, _33356_, _33355_);
  and (_33358_, _33357_, _03810_);
  nor (_33359_, _12017_, _10905_);
  nor (_33360_, _33359_, _33345_);
  nor (_33361_, _33360_, _03810_);
  or (_33362_, _33361_, _33358_);
  and (_33363_, _33362_, _02881_);
  nor (_33364_, _05320_, _33344_);
  and (_33366_, _12021_, _05320_);
  nor (_33367_, _33366_, _33364_);
  nor (_33368_, _33367_, _02881_);
  or (_33369_, _33368_, _03069_);
  or (_33370_, _33369_, _33363_);
  nand (_33371_, _33350_, _03069_);
  and (_33372_, _33371_, _33370_);
  and (_33373_, _33372_, _03084_);
  nor (_33374_, _33353_, _03084_);
  or (_33375_, _33374_, _33373_);
  and (_33377_, _33375_, _02877_);
  and (_33378_, _12005_, _05320_);
  nor (_33379_, _33378_, _33364_);
  nor (_33380_, _33379_, _02877_);
  or (_33381_, _33380_, _02869_);
  or (_33382_, _33381_, _33377_);
  nor (_33383_, _33364_, _12036_);
  nor (_33384_, _33383_, _33367_);
  or (_33385_, _33384_, _02870_);
  and (_33386_, _33385_, _02864_);
  and (_33388_, _33386_, _33382_);
  nor (_33389_, _12054_, _10889_);
  nor (_33390_, _33389_, _33364_);
  nor (_33391_, _33390_, _02864_);
  nor (_33392_, _33391_, _06770_);
  not (_33393_, _33392_);
  nor (_33394_, _33393_, _33388_);
  nor (_33395_, _33394_, _33351_);
  nor (_33396_, _33395_, _02853_);
  and (_33397_, _04622_, _06154_);
  nor (_33399_, _33345_, _05540_);
  not (_33400_, _33399_);
  nor (_33401_, _33400_, _33397_);
  or (_33402_, _33401_, _02579_);
  nor (_33403_, _33402_, _33396_);
  nor (_33404_, _12112_, _10905_);
  nor (_33405_, _33404_, _33345_);
  nor (_33406_, _33405_, _02838_);
  or (_33407_, _33406_, _02802_);
  or (_33408_, _33407_, _33403_);
  and (_33410_, _04622_, _05658_);
  nor (_33411_, _33410_, _33345_);
  nand (_33412_, _33411_, _02802_);
  and (_33413_, _33412_, _33408_);
  and (_33414_, _33413_, _03887_);
  and (_33415_, _12127_, _04622_);
  nor (_33416_, _33415_, _33345_);
  nor (_33417_, _33416_, _03887_);
  or (_33418_, _33417_, _33414_);
  and (_33419_, _33418_, _03128_);
  nor (_33421_, _33419_, _33348_);
  nor (_33422_, _33421_, _02970_);
  nor (_33423_, _33345_, _05079_);
  not (_33424_, _33423_);
  nor (_33425_, _33411_, _03883_);
  and (_33426_, _33425_, _33424_);
  nor (_33427_, _33426_, _33422_);
  nor (_33428_, _33427_, _03135_);
  nor (_33429_, _33353_, _03137_);
  and (_33430_, _33429_, _33424_);
  or (_33432_, _33430_, _33428_);
  and (_33433_, _33432_, _05783_);
  nor (_33434_, _12125_, _10905_);
  nor (_33435_, _33434_, _33345_);
  nor (_33436_, _33435_, _05783_);
  or (_33437_, _33436_, _33433_);
  and (_33438_, _33437_, _05788_);
  nor (_33439_, _12132_, _10905_);
  nor (_33440_, _33439_, _33345_);
  nor (_33441_, _33440_, _05788_);
  or (_33443_, _33441_, _33438_);
  and (_33444_, _33443_, _03906_);
  nor (_33445_, _33360_, _03906_);
  or (_33446_, _33445_, _33444_);
  and (_33447_, _33446_, _02498_);
  nor (_33448_, _33379_, _02498_);
  or (_33449_, _33448_, _33447_);
  and (_33450_, _33449_, _02890_);
  and (_33451_, _12183_, _04622_);
  nor (_33452_, _33451_, _33345_);
  nor (_33454_, _33452_, _02890_);
  or (_33455_, _33454_, _33450_);
  or (_33456_, _33455_, _42672_);
  or (_33457_, _42668_, \oc8051_golden_model_1.TCON [3]);
  and (_33458_, _33457_, _43998_);
  and (_43555_, _33458_, _33456_);
  not (_33459_, \oc8051_golden_model_1.TCON [4]);
  nor (_33460_, _04622_, _33459_);
  and (_33461_, _12207_, _04622_);
  nor (_33462_, _33461_, _33460_);
  nor (_33464_, _33462_, _03128_);
  and (_33465_, _04622_, _04982_);
  nor (_33466_, _33465_, _33460_);
  and (_33467_, _33466_, _06770_);
  nor (_33468_, _05320_, _33459_);
  and (_33469_, _12213_, _05320_);
  nor (_33470_, _33469_, _33468_);
  nor (_33471_, _33470_, _02877_);
  and (_33472_, _04622_, \oc8051_golden_model_1.ACC [4]);
  nor (_33473_, _33472_, _33460_);
  nor (_33475_, _33473_, _03814_);
  nor (_33476_, _03813_, _33459_);
  or (_33477_, _33476_, _33475_);
  and (_33478_, _33477_, _03810_);
  nor (_33479_, _12217_, _10905_);
  nor (_33480_, _33479_, _33460_);
  nor (_33481_, _33480_, _03810_);
  or (_33482_, _33481_, _33478_);
  and (_33483_, _33482_, _02881_);
  and (_33484_, _12231_, _05320_);
  nor (_33486_, _33484_, _33468_);
  nor (_33487_, _33486_, _02881_);
  or (_33488_, _33487_, _03069_);
  or (_33489_, _33488_, _33483_);
  nand (_33490_, _33466_, _03069_);
  and (_33491_, _33490_, _33489_);
  and (_33492_, _33491_, _03084_);
  nor (_33493_, _33473_, _03084_);
  or (_33494_, _33493_, _33492_);
  and (_33495_, _33494_, _02877_);
  nor (_33497_, _33495_, _33471_);
  nor (_33498_, _33497_, _02869_);
  and (_33499_, _12247_, _05320_);
  nor (_33500_, _33499_, _33468_);
  nor (_33501_, _33500_, _02870_);
  nor (_33502_, _33501_, _33498_);
  nor (_33503_, _33502_, _02863_);
  nor (_33504_, _12264_, _10889_);
  nor (_33505_, _33504_, _33468_);
  nor (_33506_, _33505_, _02864_);
  nor (_33507_, _33506_, _06770_);
  not (_33508_, _33507_);
  nor (_33509_, _33508_, _33503_);
  nor (_33510_, _33509_, _33467_);
  nor (_33511_, _33510_, _02853_);
  and (_33512_, _04622_, _06159_);
  nor (_33513_, _33460_, _05540_);
  not (_33514_, _33513_);
  nor (_33515_, _33514_, _33512_);
  nor (_33516_, _33515_, _02579_);
  not (_33519_, _33516_);
  nor (_33520_, _33519_, _33511_);
  nor (_33521_, _12321_, _10905_);
  nor (_33522_, _33521_, _33460_);
  nor (_33523_, _33522_, _02838_);
  or (_33524_, _33523_, _02802_);
  or (_33525_, _33524_, _33520_);
  and (_33526_, _05666_, _04622_);
  nor (_33527_, _33526_, _33460_);
  nand (_33528_, _33527_, _02802_);
  and (_33530_, _33528_, _33525_);
  and (_33531_, _33530_, _03887_);
  and (_33532_, _12211_, _04622_);
  nor (_33533_, _33532_, _33460_);
  nor (_33534_, _33533_, _03887_);
  or (_33535_, _33534_, _33531_);
  and (_33536_, _33535_, _03128_);
  nor (_33537_, _33536_, _33464_);
  nor (_33538_, _33537_, _02970_);
  nor (_33539_, _33460_, _05031_);
  not (_33541_, _33539_);
  nor (_33542_, _33527_, _03883_);
  and (_33543_, _33542_, _33541_);
  nor (_33544_, _33543_, _33538_);
  nor (_33545_, _33544_, _03135_);
  nor (_33546_, _33473_, _03137_);
  and (_33547_, _33546_, _33541_);
  nor (_33548_, _33547_, _02965_);
  not (_33549_, _33548_);
  nor (_33550_, _33549_, _33545_);
  nor (_33552_, _12209_, _10905_);
  or (_33553_, _33460_, _05783_);
  nor (_33554_, _33553_, _33552_);
  or (_33555_, _33554_, _03123_);
  nor (_33556_, _33555_, _33550_);
  nor (_33557_, _12206_, _10905_);
  nor (_33558_, _33557_, _33460_);
  nor (_33559_, _33558_, _05788_);
  or (_33560_, _33559_, _33556_);
  and (_33561_, _33560_, _03906_);
  nor (_33563_, _33480_, _03906_);
  or (_33564_, _33563_, _33561_);
  and (_33565_, _33564_, _02498_);
  nor (_33566_, _33470_, _02498_);
  or (_33567_, _33566_, _33565_);
  and (_33568_, _33567_, _02890_);
  and (_33569_, _12389_, _04622_);
  nor (_33570_, _33569_, _33460_);
  nor (_33571_, _33570_, _02890_);
  or (_33572_, _33571_, _33568_);
  or (_33574_, _33572_, _42672_);
  or (_33575_, _42668_, \oc8051_golden_model_1.TCON [4]);
  and (_33576_, _33575_, _43998_);
  and (_43556_, _33576_, _33574_);
  not (_33577_, \oc8051_golden_model_1.TCON [5]);
  nor (_33578_, _04622_, _33577_);
  and (_33579_, _12411_, _04622_);
  nor (_33580_, _33579_, _33578_);
  nor (_33581_, _33580_, _03128_);
  and (_33582_, _04622_, _06158_);
  or (_33584_, _33582_, _33578_);
  and (_33585_, _33584_, _02853_);
  nor (_33586_, _12407_, _10905_);
  nor (_33587_, _33586_, _33578_);
  and (_33588_, _33587_, _02974_);
  and (_33589_, _04622_, \oc8051_golden_model_1.ACC [5]);
  nor (_33590_, _33589_, _33578_);
  or (_33591_, _33590_, _03814_);
  or (_33592_, _03813_, _33577_);
  and (_33593_, _33592_, _03810_);
  and (_33595_, _33593_, _33591_);
  or (_33596_, _33595_, _02880_);
  nor (_33597_, _33596_, _33588_);
  nor (_33598_, _05320_, _33577_);
  and (_33599_, _12435_, _05320_);
  nor (_33600_, _33599_, _33598_);
  nor (_33601_, _33600_, _02881_);
  or (_33602_, _33601_, _03069_);
  or (_33603_, _33602_, _33597_);
  and (_33604_, _04622_, _04877_);
  nor (_33606_, _33604_, _33578_);
  nand (_33607_, _33606_, _03069_);
  and (_33608_, _33607_, _33603_);
  and (_33609_, _33608_, _03084_);
  nor (_33610_, _33590_, _03084_);
  or (_33611_, _33610_, _33609_);
  and (_33612_, _33611_, _02877_);
  and (_33613_, _12417_, _05320_);
  nor (_33614_, _33613_, _33598_);
  nor (_33615_, _33614_, _02877_);
  or (_33617_, _33615_, _33612_);
  and (_33618_, _33617_, _02870_);
  nor (_33619_, _33598_, _12450_);
  nor (_33620_, _33619_, _33600_);
  and (_33621_, _33620_, _02869_);
  or (_33622_, _33621_, _33618_);
  and (_33623_, _33622_, _02864_);
  nor (_33624_, _12468_, _10889_);
  nor (_33625_, _33624_, _33598_);
  nor (_33626_, _33625_, _02864_);
  nor (_33628_, _33626_, _06770_);
  not (_33629_, _33628_);
  nor (_33630_, _33629_, _33623_);
  and (_33631_, _33606_, _06770_);
  or (_33632_, _33631_, _02853_);
  nor (_33633_, _33632_, _33630_);
  or (_33634_, _33633_, _33585_);
  and (_33635_, _33634_, _02838_);
  nor (_33636_, _12527_, _10905_);
  nor (_33637_, _33636_, _33578_);
  nor (_33639_, _33637_, _02838_);
  or (_33640_, _33639_, _02802_);
  or (_33641_, _33640_, _33635_);
  and (_33642_, _05614_, _04622_);
  nor (_33643_, _33642_, _33578_);
  nand (_33644_, _33643_, _02802_);
  and (_33645_, _33644_, _33641_);
  and (_33646_, _33645_, _03887_);
  and (_33647_, _12415_, _04622_);
  nor (_33648_, _33647_, _33578_);
  nor (_33650_, _33648_, _03887_);
  or (_33651_, _33650_, _33646_);
  and (_33652_, _33651_, _03128_);
  nor (_33653_, _33652_, _33581_);
  nor (_33654_, _33653_, _02970_);
  nor (_33655_, _33578_, _04924_);
  not (_33656_, _33655_);
  nor (_33657_, _33643_, _03883_);
  and (_33658_, _33657_, _33656_);
  nor (_33659_, _33658_, _33654_);
  nor (_33661_, _33659_, _03135_);
  nor (_33662_, _33590_, _03137_);
  and (_33663_, _33662_, _33656_);
  or (_33664_, _33663_, _33661_);
  and (_33665_, _33664_, _05783_);
  nor (_33666_, _12413_, _10905_);
  nor (_33667_, _33666_, _33578_);
  nor (_33668_, _33667_, _05783_);
  or (_33669_, _33668_, _33665_);
  and (_33670_, _33669_, _05788_);
  nor (_33672_, _12410_, _10905_);
  nor (_33673_, _33672_, _33578_);
  nor (_33674_, _33673_, _05788_);
  or (_33675_, _33674_, _33670_);
  and (_33676_, _33675_, _03906_);
  nor (_33677_, _33587_, _03906_);
  or (_33678_, _33677_, _33676_);
  and (_33679_, _33678_, _02498_);
  nor (_33680_, _33614_, _02498_);
  nor (_33681_, _33680_, _02888_);
  not (_33683_, _33681_);
  nor (_33684_, _33683_, _33679_);
  and (_33685_, _12589_, _04622_);
  or (_33686_, _33578_, _02890_);
  nor (_33687_, _33686_, _33685_);
  nor (_33688_, _33687_, _33684_);
  or (_33689_, _33688_, _42672_);
  or (_33690_, _42668_, \oc8051_golden_model_1.TCON [5]);
  and (_33691_, _33690_, _43998_);
  and (_43557_, _33691_, _33689_);
  not (_33693_, \oc8051_golden_model_1.TCON [6]);
  nor (_33694_, _04622_, _33693_);
  and (_33695_, _12613_, _04622_);
  nor (_33696_, _33695_, _33694_);
  nor (_33697_, _33696_, _03128_);
  and (_33698_, _04622_, _05849_);
  or (_33699_, _33698_, _33694_);
  and (_33700_, _33699_, _02853_);
  and (_33701_, _04622_, \oc8051_golden_model_1.ACC [6]);
  nor (_33702_, _33701_, _33694_);
  nor (_33704_, _33702_, _03814_);
  nor (_33705_, _03813_, _33693_);
  or (_33706_, _33705_, _33704_);
  and (_33707_, _33706_, _03810_);
  nor (_33708_, _12603_, _10905_);
  nor (_33709_, _33708_, _33694_);
  nor (_33710_, _33709_, _03810_);
  or (_33711_, _33710_, _33707_);
  and (_33712_, _33711_, _02881_);
  nor (_33713_, _05320_, _33693_);
  and (_33715_, _12618_, _05320_);
  nor (_33716_, _33715_, _33713_);
  nor (_33717_, _33716_, _02881_);
  or (_33718_, _33717_, _03069_);
  or (_33719_, _33718_, _33712_);
  and (_33720_, _04622_, _04770_);
  nor (_33721_, _33720_, _33694_);
  nand (_33722_, _33721_, _03069_);
  and (_33723_, _33722_, _33719_);
  and (_33724_, _33723_, _03084_);
  nor (_33726_, _33702_, _03084_);
  or (_33727_, _33726_, _33724_);
  and (_33728_, _33727_, _02877_);
  and (_33729_, _12616_, _05320_);
  nor (_33730_, _33729_, _33713_);
  nor (_33731_, _33730_, _02877_);
  or (_33732_, _33731_, _33728_);
  and (_33733_, _33732_, _02870_);
  nor (_33734_, _33713_, _12646_);
  nor (_33735_, _33734_, _33716_);
  and (_33737_, _33735_, _02869_);
  or (_33738_, _33737_, _33733_);
  and (_33739_, _33738_, _02864_);
  nor (_33740_, _12664_, _10889_);
  nor (_33741_, _33740_, _33713_);
  nor (_33742_, _33741_, _02864_);
  nor (_33743_, _33742_, _06770_);
  not (_33744_, _33743_);
  nor (_33745_, _33744_, _33739_);
  and (_33746_, _33721_, _06770_);
  or (_33748_, _33746_, _02853_);
  nor (_33749_, _33748_, _33745_);
  or (_33750_, _33749_, _33700_);
  and (_33751_, _33750_, _02838_);
  nor (_33752_, _12722_, _10905_);
  nor (_33753_, _33752_, _33694_);
  nor (_33754_, _33753_, _02838_);
  or (_33755_, _33754_, _02802_);
  or (_33756_, _33755_, _33751_);
  and (_33757_, _12729_, _04622_);
  nor (_33759_, _33757_, _33694_);
  nand (_33760_, _33759_, _02802_);
  and (_33761_, _33760_, _33756_);
  and (_33762_, _33761_, _03887_);
  and (_33763_, _12739_, _04622_);
  nor (_33764_, _33763_, _33694_);
  nor (_33765_, _33764_, _03887_);
  or (_33766_, _33765_, _33762_);
  and (_33767_, _33766_, _03128_);
  nor (_33768_, _33767_, _33697_);
  nor (_33770_, _33768_, _02970_);
  nor (_33771_, _33694_, _04819_);
  not (_33772_, _33771_);
  nor (_33773_, _33759_, _03883_);
  and (_33774_, _33773_, _33772_);
  nor (_33775_, _33774_, _33770_);
  nor (_33776_, _33775_, _03135_);
  nor (_33777_, _33702_, _03137_);
  and (_33778_, _33777_, _33772_);
  or (_33779_, _33778_, _33776_);
  and (_33781_, _33779_, _05783_);
  nor (_33782_, _12737_, _10905_);
  nor (_33783_, _33782_, _33694_);
  nor (_33784_, _33783_, _05783_);
  or (_33785_, _33784_, _33781_);
  and (_33786_, _33785_, _05788_);
  nor (_33787_, _12612_, _10905_);
  nor (_33788_, _33787_, _33694_);
  nor (_33789_, _33788_, _05788_);
  or (_33790_, _33789_, _33786_);
  and (_33792_, _33790_, _03906_);
  nor (_33793_, _33709_, _03906_);
  or (_33794_, _33793_, _33792_);
  and (_33795_, _33794_, _02498_);
  nor (_33796_, _33730_, _02498_);
  or (_33797_, _33796_, _33795_);
  and (_33798_, _33797_, _02890_);
  and (_33799_, _12794_, _04622_);
  nor (_33800_, _33799_, _33694_);
  nor (_33801_, _33800_, _02890_);
  or (_33803_, _33801_, _33798_);
  or (_33804_, _33803_, _42672_);
  or (_33805_, _42668_, \oc8051_golden_model_1.TCON [6]);
  and (_33806_, _33805_, _43998_);
  and (_43559_, _33806_, _33804_);
  not (_33807_, \oc8051_golden_model_1.TH0 [0]);
  nor (_33808_, _04679_, _33807_);
  and (_33809_, _05226_, _04679_);
  nor (_33810_, _33809_, _33808_);
  and (_33811_, _33810_, _16625_);
  and (_33813_, _04679_, \oc8051_golden_model_1.ACC [0]);
  nor (_33814_, _33813_, _33808_);
  nor (_33815_, _33814_, _03084_);
  nor (_33816_, _33814_, _03814_);
  nor (_33817_, _03813_, _33807_);
  or (_33818_, _33817_, _33816_);
  and (_33819_, _33818_, _03810_);
  nor (_33820_, _33810_, _03810_);
  or (_33821_, _33820_, _33819_);
  and (_33822_, _33821_, _03336_);
  and (_33824_, _04679_, _03808_);
  nor (_33825_, _33824_, _33808_);
  nor (_33826_, _33825_, _03336_);
  nor (_33827_, _33826_, _33822_);
  nor (_33828_, _33827_, _03075_);
  or (_33829_, _33828_, _06770_);
  nor (_33830_, _33829_, _33815_);
  and (_33831_, _33825_, _06770_);
  nor (_33832_, _33831_, _33830_);
  nor (_33833_, _33832_, _02853_);
  and (_33835_, _04679_, _06152_);
  nor (_33836_, _33808_, _05540_);
  not (_33837_, _33836_);
  nor (_33838_, _33837_, _33835_);
  nor (_33839_, _33838_, _33833_);
  and (_33840_, _33839_, _02838_);
  nor (_33841_, _11505_, _10989_);
  nor (_33842_, _33841_, _33808_);
  nor (_33843_, _33842_, _02838_);
  or (_33844_, _33843_, _33840_);
  and (_33846_, _33844_, _02803_);
  and (_33847_, _04679_, _05672_);
  nor (_33848_, _33847_, _33808_);
  nor (_33849_, _33848_, _02803_);
  or (_33850_, _33849_, _33846_);
  and (_33851_, _33850_, _03887_);
  and (_33852_, _11399_, _04679_);
  nor (_33853_, _33852_, _33808_);
  nor (_33854_, _33853_, _03887_);
  or (_33855_, _33854_, _33851_);
  and (_33857_, _33855_, _03128_);
  and (_33858_, _11522_, _04679_);
  nor (_33859_, _33858_, _33808_);
  nor (_33860_, _33859_, _03128_);
  or (_33861_, _33860_, _33857_);
  and (_33862_, _33861_, _03883_);
  or (_33863_, _33848_, _03883_);
  nor (_33864_, _33863_, _33809_);
  nor (_33865_, _33864_, _33862_);
  nor (_33866_, _33865_, _03135_);
  nor (_33868_, _33808_, _09409_);
  or (_33869_, _33868_, _03137_);
  nor (_33870_, _33869_, _33814_);
  or (_33871_, _33870_, _33866_);
  and (_33872_, _33871_, _05783_);
  nor (_33873_, _11396_, _10989_);
  nor (_33874_, _33873_, _33808_);
  nor (_33875_, _33874_, _05783_);
  or (_33876_, _33875_, _33872_);
  and (_33877_, _33876_, _05788_);
  nor (_33879_, _11520_, _10989_);
  nor (_33880_, _33879_, _33808_);
  nor (_33881_, _33880_, _05788_);
  nor (_33882_, _33881_, _16625_);
  not (_33883_, _33882_);
  nor (_33884_, _33883_, _33877_);
  nor (_33885_, _33884_, _33811_);
  or (_33886_, _33885_, _42672_);
  or (_33887_, _42668_, \oc8051_golden_model_1.TH0 [0]);
  and (_33888_, _33887_, _43998_);
  and (_43560_, _33888_, _33886_);
  not (_33890_, \oc8051_golden_model_1.TH0 [1]);
  nor (_33891_, _04679_, _33890_);
  and (_33892_, _11715_, _04679_);
  or (_33893_, _33892_, _33891_);
  and (_33894_, _33893_, _03127_);
  and (_33895_, _04679_, _03698_);
  not (_33896_, _33895_);
  nor (_33897_, _04679_, \oc8051_golden_model_1.TH0 [1]);
  nor (_33898_, _33897_, _02803_);
  and (_33900_, _33898_, _33896_);
  and (_33901_, _04679_, _06151_);
  nor (_33902_, _33891_, _05540_);
  not (_33903_, _33902_);
  nor (_33904_, _33903_, _33901_);
  not (_33905_, _33904_);
  and (_33906_, _04679_, _04000_);
  or (_33907_, _33891_, _30142_);
  nor (_33908_, _33907_, _33906_);
  and (_33909_, _04679_, _02551_);
  nor (_33911_, _33909_, _33897_);
  and (_33912_, _33911_, _03075_);
  nor (_33913_, _33912_, _06770_);
  and (_33914_, _11606_, _04679_);
  nor (_33915_, _33914_, _33897_);
  and (_33916_, _33915_, _02974_);
  and (_33917_, _33911_, _03813_);
  nor (_33918_, _03813_, _33890_);
  nor (_33919_, _33918_, _33917_);
  nor (_33920_, _33919_, _02974_);
  or (_33922_, _33920_, _03069_);
  nor (_33923_, _33922_, _33916_);
  or (_33924_, _33923_, _03075_);
  and (_33925_, _33924_, _33913_);
  nor (_33926_, _33925_, _33908_);
  nor (_33927_, _33926_, _02853_);
  nor (_33928_, _33927_, _02579_);
  and (_33929_, _33928_, _33905_);
  and (_33930_, _11695_, _04679_);
  or (_33931_, _33930_, _02838_);
  nor (_33933_, _33931_, _33897_);
  nor (_33934_, _33933_, _33929_);
  nor (_33935_, _33934_, _02802_);
  nor (_33936_, _33935_, _33900_);
  nor (_33937_, _33936_, _02980_);
  nor (_33938_, _11710_, _10989_);
  or (_33939_, _33938_, _03887_);
  nor (_33940_, _33939_, _33897_);
  nor (_33941_, _33940_, _33937_);
  nor (_33942_, _33941_, _03127_);
  nor (_33944_, _33942_, _33894_);
  nor (_33945_, _33944_, _02970_);
  and (_33946_, _11709_, _04679_);
  or (_33947_, _33946_, _33891_);
  and (_33948_, _33947_, _02970_);
  nor (_33949_, _33948_, _33945_);
  nor (_33950_, _33949_, _03135_);
  nor (_33951_, _33891_, _13722_);
  nor (_33952_, _33951_, _03137_);
  and (_33953_, _33952_, _33911_);
  nor (_33955_, _33953_, _33950_);
  or (_33956_, _33955_, _17961_);
  nor (_33957_, _11708_, _10989_);
  or (_33958_, _33957_, _33891_);
  and (_33959_, _33958_, _02965_);
  not (_33960_, _33959_);
  and (_33961_, _11714_, _04679_);
  or (_33962_, _33961_, _05788_);
  or (_33963_, _33962_, _33897_);
  and (_33964_, _33963_, _03906_);
  and (_33966_, _33964_, _33960_);
  and (_33967_, _33966_, _33956_);
  nor (_33968_, _33915_, _03906_);
  nor (_33969_, _33968_, _33967_);
  and (_33970_, _33969_, _02890_);
  nor (_33971_, _33914_, _33891_);
  nor (_33972_, _33971_, _02890_);
  or (_33973_, _33972_, _33970_);
  or (_33974_, _33973_, _42672_);
  or (_33975_, _42668_, \oc8051_golden_model_1.TH0 [1]);
  and (_33977_, _33975_, _43998_);
  and (_43561_, _33977_, _33974_);
  not (_33978_, \oc8051_golden_model_1.TH0 [2]);
  nor (_33979_, _04679_, _33978_);
  and (_33980_, _11927_, _04679_);
  nor (_33981_, _33980_, _33979_);
  nor (_33982_, _33981_, _03128_);
  and (_33983_, _04679_, \oc8051_golden_model_1.ACC [2]);
  nor (_33984_, _33983_, _33979_);
  nor (_33985_, _33984_, _03084_);
  nor (_33987_, _33984_, _03814_);
  nor (_33988_, _03813_, _33978_);
  or (_33989_, _33988_, _33987_);
  and (_33990_, _33989_, _03810_);
  nor (_33991_, _11801_, _10989_);
  nor (_33992_, _33991_, _33979_);
  nor (_33993_, _33992_, _03810_);
  or (_33994_, _33993_, _33990_);
  and (_33995_, _33994_, _03336_);
  and (_33996_, _04679_, _04435_);
  nor (_33998_, _33996_, _33979_);
  nor (_33999_, _33998_, _03336_);
  nor (_34000_, _33999_, _33995_);
  nor (_34001_, _34000_, _03075_);
  or (_34002_, _34001_, _06770_);
  nor (_34003_, _34002_, _33985_);
  and (_34004_, _33998_, _06770_);
  nor (_34005_, _34004_, _34003_);
  nor (_34006_, _34005_, _02853_);
  and (_34007_, _04679_, _06155_);
  nor (_34009_, _33979_, _05540_);
  not (_34010_, _34009_);
  nor (_34011_, _34010_, _34007_);
  or (_34012_, _34011_, _02579_);
  nor (_34013_, _34012_, _34006_);
  nor (_34014_, _11906_, _10989_);
  nor (_34015_, _34014_, _33979_);
  nor (_34016_, _34015_, _02838_);
  or (_34017_, _34016_, _02802_);
  or (_34018_, _34017_, _34013_);
  and (_34020_, _04679_, _05701_);
  nor (_34021_, _34020_, _33979_);
  nand (_34022_, _34021_, _02802_);
  and (_34023_, _34022_, _34018_);
  and (_34024_, _34023_, _03887_);
  and (_34025_, _11921_, _04679_);
  nor (_34026_, _34025_, _33979_);
  nor (_34027_, _34026_, _03887_);
  or (_34028_, _34027_, _34024_);
  and (_34029_, _34028_, _03128_);
  nor (_34030_, _34029_, _33982_);
  nor (_34031_, _34030_, _02970_);
  nor (_34032_, _33979_, _05130_);
  not (_34033_, _34032_);
  nor (_34034_, _34021_, _03883_);
  and (_34035_, _34034_, _34033_);
  nor (_34036_, _34035_, _34031_);
  nor (_34037_, _34036_, _03135_);
  nor (_34038_, _33984_, _03137_);
  and (_34039_, _34038_, _34033_);
  or (_34042_, _34039_, _34037_);
  and (_34043_, _34042_, _05783_);
  nor (_34044_, _11919_, _10989_);
  nor (_34045_, _34044_, _33979_);
  nor (_34046_, _34045_, _05783_);
  or (_34047_, _34046_, _34043_);
  and (_34048_, _34047_, _05788_);
  nor (_34049_, _11926_, _10989_);
  nor (_34050_, _34049_, _33979_);
  nor (_34051_, _34050_, _05788_);
  or (_34053_, _34051_, _03163_);
  nor (_34054_, _34053_, _34048_);
  and (_34055_, _33992_, _03163_);
  or (_34056_, _34055_, _02888_);
  nor (_34057_, _34056_, _34054_);
  and (_34058_, _11985_, _04679_);
  nor (_34059_, _34058_, _33979_);
  nor (_34060_, _34059_, _02890_);
  or (_34061_, _34060_, _34057_);
  or (_34062_, _34061_, _42672_);
  or (_34064_, _42668_, \oc8051_golden_model_1.TH0 [2]);
  and (_34065_, _34064_, _43998_);
  and (_43562_, _34065_, _34062_);
  not (_34066_, \oc8051_golden_model_1.TH0 [3]);
  nor (_34067_, _04679_, _34066_);
  and (_34068_, _12133_, _04679_);
  nor (_34069_, _34068_, _34067_);
  nor (_34070_, _34069_, _03128_);
  and (_34071_, _04679_, \oc8051_golden_model_1.ACC [3]);
  nor (_34072_, _34071_, _34067_);
  nor (_34074_, _34072_, _03814_);
  nor (_34075_, _03813_, _34066_);
  or (_34076_, _34075_, _34074_);
  and (_34077_, _34076_, _03810_);
  nor (_34078_, _12017_, _10989_);
  nor (_34079_, _34078_, _34067_);
  nor (_34080_, _34079_, _03810_);
  or (_34081_, _34080_, _34077_);
  and (_34082_, _34081_, _03336_);
  and (_34083_, _04679_, _04241_);
  nor (_34085_, _34083_, _34067_);
  nor (_34086_, _34085_, _03336_);
  nor (_34087_, _34086_, _34082_);
  nor (_34088_, _34087_, _03075_);
  nor (_34089_, _34072_, _03084_);
  nor (_34090_, _34089_, _06770_);
  not (_34091_, _34090_);
  nor (_34092_, _34091_, _34088_);
  and (_34093_, _34085_, _06770_);
  or (_34094_, _34093_, _02853_);
  nor (_34096_, _34094_, _34092_);
  and (_34097_, _04679_, _06154_);
  or (_34098_, _34097_, _34067_);
  and (_34099_, _34098_, _02853_);
  or (_34100_, _34099_, _02579_);
  or (_34101_, _34100_, _34096_);
  nor (_34102_, _12112_, _10989_);
  or (_34103_, _34067_, _02838_);
  or (_34104_, _34103_, _34102_);
  and (_34105_, _34104_, _02803_);
  and (_34107_, _34105_, _34101_);
  and (_34108_, _04679_, _05658_);
  nor (_34109_, _34108_, _34067_);
  nor (_34110_, _34109_, _02803_);
  or (_34111_, _34110_, _34107_);
  and (_34112_, _34111_, _03887_);
  and (_34113_, _12127_, _04679_);
  nor (_34114_, _34113_, _34067_);
  nor (_34115_, _34114_, _03887_);
  or (_34116_, _34115_, _34112_);
  and (_34118_, _34116_, _03128_);
  nor (_34119_, _34118_, _34070_);
  nor (_34120_, _34119_, _02970_);
  nor (_34121_, _34067_, _05079_);
  not (_34122_, _34121_);
  nor (_34123_, _34109_, _03883_);
  and (_34124_, _34123_, _34122_);
  nor (_34125_, _34124_, _34120_);
  nor (_34126_, _34125_, _03135_);
  nor (_34127_, _34072_, _03137_);
  and (_34129_, _34127_, _34122_);
  or (_34130_, _34129_, _34126_);
  and (_34131_, _34130_, _05783_);
  nor (_34132_, _12125_, _10989_);
  nor (_34133_, _34132_, _34067_);
  nor (_34134_, _34133_, _05783_);
  or (_34135_, _34134_, _34131_);
  and (_34136_, _34135_, _05788_);
  nor (_34137_, _12132_, _10989_);
  nor (_34138_, _34137_, _34067_);
  nor (_34140_, _34138_, _05788_);
  or (_34141_, _34140_, _03163_);
  nor (_34142_, _34141_, _34136_);
  and (_34143_, _34079_, _03163_);
  or (_34144_, _34143_, _02888_);
  nor (_34145_, _34144_, _34142_);
  and (_34146_, _12183_, _04679_);
  nor (_34147_, _34146_, _34067_);
  nor (_34148_, _34147_, _02890_);
  or (_34149_, _34148_, _34145_);
  or (_34151_, _34149_, _42672_);
  or (_34152_, _42668_, \oc8051_golden_model_1.TH0 [3]);
  and (_34153_, _34152_, _43998_);
  and (_43563_, _34153_, _34151_);
  not (_34154_, \oc8051_golden_model_1.TH0 [4]);
  nor (_34155_, _04679_, _34154_);
  and (_34156_, _12207_, _04679_);
  nor (_34157_, _34156_, _34155_);
  nor (_34158_, _34157_, _03128_);
  and (_34159_, _04679_, _04982_);
  nor (_34161_, _34159_, _34155_);
  and (_34162_, _34161_, _06770_);
  and (_34163_, _04679_, \oc8051_golden_model_1.ACC [4]);
  nor (_34164_, _34163_, _34155_);
  nor (_34165_, _34164_, _03814_);
  nor (_34166_, _03813_, _34154_);
  or (_34167_, _34166_, _34165_);
  and (_34168_, _34167_, _03810_);
  nor (_34169_, _12217_, _10989_);
  nor (_34170_, _34169_, _34155_);
  nor (_34172_, _34170_, _03810_);
  or (_34173_, _34172_, _34168_);
  and (_34174_, _34173_, _03336_);
  nor (_34175_, _34161_, _03336_);
  nor (_34176_, _34175_, _34174_);
  nor (_34177_, _34176_, _03075_);
  nor (_34178_, _34164_, _03084_);
  nor (_34179_, _34178_, _06770_);
  not (_34180_, _34179_);
  nor (_34181_, _34180_, _34177_);
  nor (_34183_, _34181_, _34162_);
  nor (_34184_, _34183_, _02853_);
  and (_34185_, _04679_, _06159_);
  nor (_34186_, _34155_, _05540_);
  not (_34187_, _34186_);
  nor (_34188_, _34187_, _34185_);
  or (_34189_, _34188_, _02579_);
  nor (_34190_, _34189_, _34184_);
  nor (_34191_, _12321_, _10989_);
  nor (_34192_, _34191_, _34155_);
  nor (_34194_, _34192_, _02838_);
  or (_34195_, _34194_, _02802_);
  or (_34196_, _34195_, _34190_);
  and (_34197_, _05666_, _04679_);
  nor (_34198_, _34197_, _34155_);
  nand (_34199_, _34198_, _02802_);
  and (_34200_, _34199_, _34196_);
  and (_34201_, _34200_, _03887_);
  and (_34202_, _12211_, _04679_);
  nor (_34203_, _34202_, _34155_);
  nor (_34205_, _34203_, _03887_);
  or (_34206_, _34205_, _34201_);
  and (_34207_, _34206_, _03128_);
  nor (_34208_, _34207_, _34158_);
  nor (_34209_, _34208_, _02970_);
  nor (_34210_, _34155_, _05031_);
  not (_34211_, _34210_);
  nor (_34212_, _34198_, _03883_);
  and (_34213_, _34212_, _34211_);
  nor (_34214_, _34213_, _34209_);
  nor (_34216_, _34214_, _03135_);
  nor (_34217_, _34164_, _03137_);
  and (_34218_, _34217_, _34211_);
  or (_34219_, _34218_, _34216_);
  and (_34220_, _34219_, _05783_);
  nor (_34221_, _12209_, _10989_);
  nor (_34222_, _34221_, _34155_);
  nor (_34223_, _34222_, _05783_);
  or (_34224_, _34223_, _34220_);
  and (_34225_, _34224_, _05788_);
  nor (_34227_, _12206_, _10989_);
  nor (_34228_, _34227_, _34155_);
  nor (_34229_, _34228_, _05788_);
  or (_34230_, _34229_, _03163_);
  nor (_34231_, _34230_, _34225_);
  and (_34232_, _34170_, _03163_);
  or (_34233_, _34232_, _02888_);
  nor (_34234_, _34233_, _34231_);
  and (_34235_, _12389_, _04679_);
  nor (_34236_, _34235_, _34155_);
  nor (_34238_, _34236_, _02890_);
  or (_34239_, _34238_, _34234_);
  or (_34240_, _34239_, _42672_);
  or (_34241_, _42668_, \oc8051_golden_model_1.TH0 [4]);
  and (_34242_, _34241_, _43998_);
  and (_43564_, _34242_, _34240_);
  not (_34243_, \oc8051_golden_model_1.TH0 [5]);
  nor (_34244_, _04679_, _34243_);
  and (_34245_, _12411_, _04679_);
  nor (_34246_, _34245_, _34244_);
  nor (_34248_, _34246_, _03128_);
  and (_34249_, _04679_, _04877_);
  nor (_34250_, _34249_, _34244_);
  and (_34251_, _34250_, _06770_);
  nor (_34252_, _12407_, _10989_);
  nor (_34253_, _34252_, _34244_);
  and (_34254_, _34253_, _02974_);
  and (_34255_, _04679_, \oc8051_golden_model_1.ACC [5]);
  nor (_34256_, _34255_, _34244_);
  or (_34257_, _34256_, _03814_);
  or (_34259_, _03813_, _34243_);
  and (_34260_, _34259_, _03810_);
  and (_34261_, _34260_, _34257_);
  or (_34262_, _34261_, _03069_);
  nor (_34263_, _34262_, _34254_);
  nor (_34264_, _34250_, _03336_);
  nor (_34265_, _34264_, _34263_);
  nor (_34266_, _34265_, _03075_);
  nor (_34267_, _34256_, _03084_);
  nor (_34268_, _34267_, _06770_);
  not (_34270_, _34268_);
  nor (_34271_, _34270_, _34266_);
  nor (_34272_, _34271_, _34251_);
  nor (_34273_, _34272_, _02853_);
  and (_34274_, _04679_, _06158_);
  nor (_34275_, _34244_, _05540_);
  not (_34276_, _34275_);
  nor (_34277_, _34276_, _34274_);
  or (_34278_, _34277_, _02579_);
  nor (_34279_, _34278_, _34273_);
  nor (_34281_, _12527_, _10989_);
  nor (_34282_, _34281_, _34244_);
  nor (_34283_, _34282_, _02838_);
  or (_34284_, _34283_, _02802_);
  or (_34285_, _34284_, _34279_);
  and (_34286_, _05614_, _04679_);
  nor (_34287_, _34286_, _34244_);
  nand (_34288_, _34287_, _02802_);
  and (_34289_, _34288_, _34285_);
  and (_34290_, _34289_, _03887_);
  and (_34292_, _12415_, _04679_);
  nor (_34293_, _34292_, _34244_);
  nor (_34294_, _34293_, _03887_);
  or (_34295_, _34294_, _34290_);
  and (_34296_, _34295_, _03128_);
  nor (_34297_, _34296_, _34248_);
  nor (_34298_, _34297_, _02970_);
  nor (_34299_, _34244_, _04924_);
  not (_34300_, _34299_);
  nor (_34301_, _34287_, _03883_);
  and (_34302_, _34301_, _34300_);
  nor (_34303_, _34302_, _34298_);
  nor (_34304_, _34303_, _03135_);
  nor (_34305_, _34256_, _03137_);
  and (_34306_, _34305_, _34300_);
  nor (_34307_, _34306_, _02965_);
  not (_34308_, _34307_);
  nor (_34309_, _34308_, _34304_);
  nor (_34310_, _12413_, _10989_);
  or (_34311_, _34244_, _05783_);
  nor (_34314_, _34311_, _34310_);
  or (_34315_, _34314_, _03123_);
  nor (_34316_, _34315_, _34309_);
  nor (_34317_, _12410_, _10989_);
  nor (_34318_, _34317_, _34244_);
  nor (_34319_, _34318_, _05788_);
  or (_34320_, _34319_, _03163_);
  nor (_34321_, _34320_, _34316_);
  and (_34322_, _34253_, _03163_);
  or (_34323_, _34322_, _02888_);
  nor (_34325_, _34323_, _34321_);
  and (_34326_, _12589_, _04679_);
  nor (_34327_, _34326_, _34244_);
  nor (_34328_, _34327_, _02890_);
  or (_34329_, _34328_, _34325_);
  or (_34330_, _34329_, _42672_);
  or (_34331_, _42668_, \oc8051_golden_model_1.TH0 [5]);
  and (_34332_, _34331_, _43998_);
  and (_43565_, _34332_, _34330_);
  not (_34333_, \oc8051_golden_model_1.TH0 [6]);
  nor (_34335_, _04679_, _34333_);
  and (_34336_, _12613_, _04679_);
  nor (_34337_, _34336_, _34335_);
  nor (_34338_, _34337_, _03128_);
  and (_34339_, _04679_, \oc8051_golden_model_1.ACC [6]);
  nor (_34340_, _34339_, _34335_);
  nor (_34341_, _34340_, _03084_);
  nor (_34342_, _34340_, _03814_);
  nor (_34343_, _03813_, _34333_);
  or (_34344_, _34343_, _34342_);
  and (_34346_, _34344_, _03810_);
  nor (_34347_, _12603_, _10989_);
  nor (_34348_, _34347_, _34335_);
  nor (_34349_, _34348_, _03810_);
  or (_34350_, _34349_, _34346_);
  and (_34351_, _34350_, _03336_);
  and (_34352_, _04679_, _04770_);
  nor (_34353_, _34352_, _34335_);
  nor (_34354_, _34353_, _03336_);
  nor (_34355_, _34354_, _34351_);
  nor (_34357_, _34355_, _03075_);
  or (_34358_, _34357_, _06770_);
  nor (_34359_, _34358_, _34341_);
  and (_34360_, _34353_, _06770_);
  nor (_34361_, _34360_, _34359_);
  nor (_34362_, _34361_, _02853_);
  and (_34363_, _04679_, _05849_);
  nor (_34364_, _34335_, _05540_);
  not (_34365_, _34364_);
  nor (_34366_, _34365_, _34363_);
  or (_34368_, _34366_, _02579_);
  nor (_34369_, _34368_, _34362_);
  nor (_34370_, _12722_, _10989_);
  nor (_34371_, _34370_, _34335_);
  nor (_34372_, _34371_, _02838_);
  or (_34373_, _34372_, _02802_);
  or (_34374_, _34373_, _34369_);
  and (_34375_, _12729_, _04679_);
  nor (_34376_, _34375_, _34335_);
  nand (_34377_, _34376_, _02802_);
  and (_34379_, _34377_, _34374_);
  and (_34380_, _34379_, _03887_);
  and (_34381_, _12739_, _04679_);
  nor (_34382_, _34381_, _34335_);
  nor (_34383_, _34382_, _03887_);
  or (_34384_, _34383_, _34380_);
  and (_34385_, _34384_, _03128_);
  nor (_34386_, _34385_, _34338_);
  nor (_34387_, _34386_, _02970_);
  nor (_34388_, _34335_, _04819_);
  not (_34390_, _34388_);
  nor (_34391_, _34376_, _03883_);
  and (_34392_, _34391_, _34390_);
  nor (_34393_, _34392_, _34387_);
  nor (_34394_, _34393_, _03135_);
  nor (_34395_, _34340_, _03137_);
  and (_34396_, _34395_, _34390_);
  or (_34397_, _34396_, _34394_);
  and (_34398_, _34397_, _05783_);
  nor (_34399_, _12737_, _10989_);
  nor (_34401_, _34399_, _34335_);
  nor (_34402_, _34401_, _05783_);
  or (_34403_, _34402_, _34398_);
  and (_34404_, _34403_, _05788_);
  nor (_34405_, _12612_, _10989_);
  nor (_34406_, _34405_, _34335_);
  nor (_34407_, _34406_, _05788_);
  or (_34408_, _34407_, _03163_);
  nor (_34409_, _34408_, _34404_);
  and (_34410_, _34348_, _03163_);
  or (_34412_, _34410_, _02888_);
  nor (_34413_, _34412_, _34409_);
  and (_34414_, _12794_, _04679_);
  nor (_34415_, _34414_, _34335_);
  nor (_34416_, _34415_, _02890_);
  or (_34417_, _34416_, _34413_);
  or (_34418_, _34417_, _42672_);
  or (_34419_, _42668_, \oc8051_golden_model_1.TH0 [6]);
  and (_34420_, _34419_, _43998_);
  and (_43566_, _34420_, _34418_);
  not (_34422_, \oc8051_golden_model_1.TH1 [0]);
  nor (_34423_, _04660_, _34422_);
  and (_34424_, _05226_, _04660_);
  nor (_34425_, _34424_, _34423_);
  and (_34426_, _34425_, _16625_);
  and (_34427_, _04660_, _05672_);
  nor (_34428_, _34427_, _34423_);
  or (_34429_, _34428_, _03883_);
  nor (_34430_, _34429_, _34424_);
  and (_34431_, _04660_, \oc8051_golden_model_1.ACC [0]);
  nor (_34433_, _34431_, _34423_);
  nor (_34434_, _34433_, _03084_);
  nor (_34435_, _34433_, _03814_);
  nor (_34436_, _03813_, _34422_);
  or (_34437_, _34436_, _34435_);
  and (_34438_, _34437_, _03810_);
  nor (_34439_, _34425_, _03810_);
  or (_34440_, _34439_, _34438_);
  and (_34441_, _34440_, _03336_);
  and (_34442_, _04660_, _03808_);
  nor (_34444_, _34442_, _34423_);
  nor (_34445_, _34444_, _03336_);
  nor (_34446_, _34445_, _34441_);
  nor (_34447_, _34446_, _03075_);
  or (_34448_, _34447_, _06770_);
  nor (_34449_, _34448_, _34434_);
  and (_34450_, _34444_, _06770_);
  nor (_34451_, _34450_, _34449_);
  nor (_34452_, _34451_, _02853_);
  and (_34453_, _04660_, _06152_);
  nor (_34455_, _34423_, _05540_);
  not (_34456_, _34455_);
  nor (_34457_, _34456_, _34453_);
  nor (_34458_, _34457_, _34452_);
  and (_34459_, _34458_, _02838_);
  nor (_34460_, _11505_, _11071_);
  nor (_34461_, _34460_, _34423_);
  nor (_34462_, _34461_, _02838_);
  or (_34463_, _34462_, _34459_);
  and (_34464_, _34463_, _02803_);
  nor (_34466_, _34428_, _02803_);
  or (_34467_, _34466_, _34464_);
  and (_34468_, _34467_, _03887_);
  and (_34469_, _11399_, _04660_);
  nor (_34470_, _34469_, _34423_);
  nor (_34471_, _34470_, _03887_);
  or (_34472_, _34471_, _34468_);
  and (_34473_, _34472_, _03128_);
  and (_34474_, _11522_, _04660_);
  nor (_34475_, _34474_, _34423_);
  nor (_34477_, _34475_, _03128_);
  or (_34478_, _34477_, _34473_);
  and (_34479_, _34478_, _03883_);
  nor (_34480_, _34479_, _34430_);
  nor (_34481_, _34480_, _03135_);
  nor (_34482_, _34423_, _09409_);
  or (_34483_, _34482_, _03137_);
  nor (_34484_, _34483_, _34433_);
  or (_34485_, _34484_, _34481_);
  and (_34486_, _34485_, _05783_);
  nor (_34488_, _11396_, _11071_);
  nor (_34489_, _34488_, _34423_);
  nor (_34490_, _34489_, _05783_);
  or (_34491_, _34490_, _34486_);
  and (_34492_, _34491_, _05788_);
  nor (_34493_, _11520_, _11071_);
  nor (_34494_, _34493_, _34423_);
  nor (_34495_, _34494_, _05788_);
  nor (_34496_, _34495_, _16625_);
  not (_34497_, _34496_);
  nor (_34499_, _34497_, _34492_);
  nor (_34500_, _34499_, _34426_);
  or (_34501_, _34500_, _42672_);
  or (_34502_, _42668_, \oc8051_golden_model_1.TH1 [0]);
  and (_34503_, _34502_, _43998_);
  and (_43568_, _34503_, _34501_);
  nor (_34504_, _04660_, \oc8051_golden_model_1.TH1 [1]);
  nor (_34505_, _11071_, _04000_);
  or (_34506_, _34505_, _34504_);
  nor (_34507_, _34506_, _03336_);
  and (_34509_, _04660_, _02551_);
  nor (_34510_, _34509_, _34504_);
  and (_34511_, _34510_, _03813_);
  not (_34512_, \oc8051_golden_model_1.TH1 [1]);
  nor (_34513_, _03813_, _34512_);
  or (_34514_, _34513_, _34511_);
  and (_34515_, _34514_, _03810_);
  and (_34516_, _11606_, _04660_);
  nor (_34517_, _34516_, _34504_);
  and (_34518_, _34517_, _02974_);
  or (_34520_, _34518_, _34515_);
  and (_34521_, _34520_, _03336_);
  nor (_34522_, _34521_, _34507_);
  nor (_34523_, _34522_, _03075_);
  and (_34524_, _34510_, _03075_);
  nor (_34525_, _34524_, _06770_);
  not (_34526_, _34525_);
  nor (_34527_, _34526_, _34523_);
  and (_34528_, _34506_, _06770_);
  or (_34529_, _34528_, _02853_);
  nor (_34531_, _34529_, _34527_);
  or (_34532_, _11071_, _06151_);
  nor (_34533_, _34504_, _05540_);
  and (_34534_, _34533_, _34532_);
  or (_34535_, _34534_, _34531_);
  and (_34536_, _34535_, _02838_);
  and (_34537_, _11695_, _04660_);
  or (_34538_, _34537_, _02838_);
  nor (_34539_, _34538_, _34504_);
  nor (_34540_, _34539_, _34536_);
  nor (_34542_, _34540_, _02802_);
  and (_34543_, _04660_, _03698_);
  not (_34544_, _34543_);
  nor (_34545_, _34504_, _02803_);
  and (_34546_, _34545_, _34544_);
  nor (_34547_, _34546_, _34542_);
  nor (_34548_, _34547_, _02980_);
  nor (_34549_, _11710_, _11071_);
  or (_34550_, _34549_, _03887_);
  nor (_34551_, _34550_, _34504_);
  nor (_34553_, _34551_, _34548_);
  nor (_34554_, _34553_, _03127_);
  nor (_34555_, _04660_, _34512_);
  and (_34556_, _11715_, _04660_);
  or (_34557_, _34556_, _34555_);
  and (_34558_, _34557_, _03127_);
  nor (_34559_, _34558_, _34554_);
  nor (_34560_, _34559_, _02970_);
  and (_34561_, _11709_, _04660_);
  or (_34562_, _34561_, _34555_);
  and (_34564_, _34562_, _02970_);
  nor (_34565_, _34564_, _34560_);
  nor (_34566_, _34565_, _03135_);
  nor (_34567_, _34555_, _13722_);
  nor (_34568_, _34567_, _03137_);
  and (_34569_, _34568_, _34510_);
  nor (_34570_, _34569_, _34566_);
  or (_34571_, _34570_, _17961_);
  nor (_34572_, _11708_, _11071_);
  or (_34573_, _34572_, _34555_);
  and (_34575_, _34573_, _02965_);
  not (_34576_, _34575_);
  and (_34577_, _11714_, _04660_);
  or (_34578_, _34577_, _05788_);
  or (_34579_, _34578_, _34504_);
  and (_34580_, _34579_, _03906_);
  and (_34581_, _34580_, _34576_);
  and (_34582_, _34581_, _34571_);
  nor (_34583_, _34517_, _03906_);
  nor (_34584_, _34583_, _34582_);
  and (_34586_, _34584_, _02890_);
  nor (_34587_, _34516_, _34555_);
  nor (_34588_, _34587_, _02890_);
  or (_34589_, _34588_, _34586_);
  or (_34590_, _34589_, _42672_);
  or (_34591_, _42668_, \oc8051_golden_model_1.TH1 [1]);
  and (_34592_, _34591_, _43998_);
  and (_43569_, _34592_, _34590_);
  not (_34593_, \oc8051_golden_model_1.TH1 [2]);
  nor (_34594_, _04660_, _34593_);
  and (_34596_, _11927_, _04660_);
  nor (_34597_, _34596_, _34594_);
  nor (_34598_, _34597_, _03128_);
  and (_34599_, _04660_, _04435_);
  nor (_34600_, _34599_, _34594_);
  and (_34601_, _34600_, _06770_);
  and (_34602_, _04660_, \oc8051_golden_model_1.ACC [2]);
  nor (_34603_, _34602_, _34594_);
  nor (_34604_, _34603_, _03084_);
  nor (_34605_, _34603_, _03814_);
  nor (_34607_, _03813_, _34593_);
  or (_34608_, _34607_, _34605_);
  and (_34609_, _34608_, _03810_);
  nor (_34610_, _11801_, _11071_);
  nor (_34611_, _34610_, _34594_);
  nor (_34612_, _34611_, _03810_);
  or (_34613_, _34612_, _34609_);
  and (_34614_, _34613_, _03336_);
  nor (_34615_, _34600_, _03336_);
  nor (_34616_, _34615_, _34614_);
  nor (_34618_, _34616_, _03075_);
  or (_34619_, _34618_, _06770_);
  nor (_34620_, _34619_, _34604_);
  nor (_34621_, _34620_, _34601_);
  nor (_34622_, _34621_, _02853_);
  and (_34623_, _04660_, _06155_);
  nor (_34624_, _34594_, _05540_);
  not (_34625_, _34624_);
  nor (_34626_, _34625_, _34623_);
  or (_34627_, _34626_, _02579_);
  nor (_34629_, _34627_, _34622_);
  nor (_34630_, _11906_, _11071_);
  nor (_34631_, _34630_, _34594_);
  nor (_34632_, _34631_, _02838_);
  or (_34633_, _34632_, _02802_);
  or (_34634_, _34633_, _34629_);
  and (_34635_, _04660_, _05701_);
  nor (_34636_, _34635_, _34594_);
  nand (_34637_, _34636_, _02802_);
  and (_34638_, _34637_, _34634_);
  and (_34640_, _34638_, _03887_);
  and (_34641_, _11921_, _04660_);
  nor (_34642_, _34641_, _34594_);
  nor (_34643_, _34642_, _03887_);
  or (_34644_, _34643_, _34640_);
  and (_34645_, _34644_, _03128_);
  nor (_34646_, _34645_, _34598_);
  nor (_34647_, _34646_, _02970_);
  nor (_34648_, _34594_, _05130_);
  not (_34649_, _34648_);
  nor (_34651_, _34636_, _03883_);
  and (_34652_, _34651_, _34649_);
  nor (_34653_, _34652_, _34647_);
  nor (_34654_, _34653_, _03135_);
  nor (_34655_, _34603_, _03137_);
  and (_34656_, _34655_, _34649_);
  or (_34657_, _34656_, _34654_);
  and (_34658_, _34657_, _05783_);
  nor (_34659_, _11919_, _11071_);
  nor (_34660_, _34659_, _34594_);
  nor (_34662_, _34660_, _05783_);
  or (_34663_, _34662_, _34658_);
  and (_34664_, _34663_, _05788_);
  nor (_34665_, _11926_, _11071_);
  nor (_34666_, _34665_, _34594_);
  nor (_34667_, _34666_, _05788_);
  or (_34668_, _34667_, _03163_);
  nor (_34669_, _34668_, _34664_);
  and (_34670_, _34611_, _03163_);
  or (_34671_, _34670_, _02888_);
  nor (_34673_, _34671_, _34669_);
  and (_34674_, _11985_, _04660_);
  nor (_34675_, _34674_, _34594_);
  nor (_34676_, _34675_, _02890_);
  or (_34677_, _34676_, _34673_);
  or (_34678_, _34677_, _42672_);
  or (_34679_, _42668_, \oc8051_golden_model_1.TH1 [2]);
  and (_34680_, _34679_, _43998_);
  and (_43570_, _34680_, _34678_);
  not (_34681_, \oc8051_golden_model_1.TH1 [3]);
  nor (_34683_, _04660_, _34681_);
  and (_34684_, _12133_, _04660_);
  nor (_34685_, _34684_, _34683_);
  nor (_34686_, _34685_, _03128_);
  and (_34687_, _04660_, \oc8051_golden_model_1.ACC [3]);
  nor (_34688_, _34687_, _34683_);
  nor (_34689_, _34688_, _03814_);
  nor (_34690_, _03813_, _34681_);
  or (_34691_, _34690_, _34689_);
  and (_34692_, _34691_, _03810_);
  nor (_34694_, _12017_, _11071_);
  nor (_34695_, _34694_, _34683_);
  nor (_34696_, _34695_, _03810_);
  or (_34697_, _34696_, _34692_);
  and (_34698_, _34697_, _03336_);
  and (_34699_, _04660_, _04241_);
  nor (_34700_, _34699_, _34683_);
  nor (_34701_, _34700_, _03336_);
  nor (_34702_, _34701_, _34698_);
  nor (_34703_, _34702_, _03075_);
  nor (_34705_, _34688_, _03084_);
  nor (_34706_, _34705_, _06770_);
  not (_34707_, _34706_);
  nor (_34708_, _34707_, _34703_);
  and (_34709_, _34700_, _06770_);
  or (_34710_, _34709_, _02853_);
  nor (_34711_, _34710_, _34708_);
  and (_34712_, _04660_, _06154_);
  or (_34713_, _34712_, _34683_);
  and (_34714_, _34713_, _02853_);
  or (_34716_, _34714_, _02579_);
  or (_34717_, _34716_, _34711_);
  nor (_34718_, _12112_, _11071_);
  or (_34719_, _34683_, _02838_);
  or (_34720_, _34719_, _34718_);
  and (_34721_, _34720_, _02803_);
  and (_34722_, _34721_, _34717_);
  and (_34723_, _04660_, _05658_);
  nor (_34724_, _34723_, _34683_);
  nor (_34725_, _34724_, _02803_);
  or (_34727_, _34725_, _34722_);
  and (_34728_, _34727_, _03887_);
  and (_34729_, _12127_, _04660_);
  nor (_34730_, _34729_, _34683_);
  nor (_34731_, _34730_, _03887_);
  or (_34732_, _34731_, _34728_);
  and (_34733_, _34732_, _03128_);
  nor (_34734_, _34733_, _34686_);
  nor (_34735_, _34734_, _02970_);
  nor (_34736_, _34683_, _05079_);
  not (_34738_, _34736_);
  nor (_34739_, _34724_, _03883_);
  and (_34740_, _34739_, _34738_);
  nor (_34741_, _34740_, _34735_);
  nor (_34742_, _34741_, _03135_);
  nor (_34743_, _34688_, _03137_);
  and (_34744_, _34743_, _34738_);
  or (_34745_, _34744_, _34742_);
  and (_34746_, _34745_, _05783_);
  nor (_34747_, _12125_, _11071_);
  nor (_34749_, _34747_, _34683_);
  nor (_34750_, _34749_, _05783_);
  or (_34751_, _34750_, _34746_);
  and (_34752_, _34751_, _05788_);
  nor (_34753_, _12132_, _11071_);
  nor (_34754_, _34753_, _34683_);
  nor (_34755_, _34754_, _05788_);
  or (_34756_, _34755_, _03163_);
  nor (_34757_, _34756_, _34752_);
  and (_34758_, _34695_, _03163_);
  or (_34760_, _34758_, _02888_);
  nor (_34761_, _34760_, _34757_);
  and (_34762_, _12183_, _04660_);
  nor (_34763_, _34762_, _34683_);
  nor (_34764_, _34763_, _02890_);
  or (_34765_, _34764_, _34761_);
  or (_34766_, _34765_, _42672_);
  or (_34767_, _42668_, \oc8051_golden_model_1.TH1 [3]);
  and (_34768_, _34767_, _43998_);
  and (_43571_, _34768_, _34766_);
  not (_34770_, \oc8051_golden_model_1.TH1 [4]);
  nor (_34771_, _04660_, _34770_);
  nor (_34772_, _34771_, _05031_);
  not (_34773_, _34772_);
  and (_34774_, _05666_, _04660_);
  nor (_34775_, _34774_, _34771_);
  nor (_34776_, _34775_, _03883_);
  and (_34777_, _34776_, _34773_);
  and (_34778_, _12207_, _04660_);
  nor (_34779_, _34778_, _34771_);
  nor (_34781_, _34779_, _03128_);
  and (_34782_, _04660_, _04982_);
  nor (_34783_, _34782_, _34771_);
  and (_34784_, _34783_, _06770_);
  and (_34785_, _04660_, \oc8051_golden_model_1.ACC [4]);
  nor (_34786_, _34785_, _34771_);
  nor (_34787_, _34786_, _03084_);
  nor (_34788_, _34786_, _03814_);
  nor (_34789_, _03813_, _34770_);
  or (_34790_, _34789_, _34788_);
  and (_34792_, _34790_, _03810_);
  nor (_34793_, _12217_, _11071_);
  nor (_34794_, _34793_, _34771_);
  nor (_34795_, _34794_, _03810_);
  or (_34796_, _34795_, _34792_);
  and (_34797_, _34796_, _03336_);
  nor (_34798_, _34783_, _03336_);
  nor (_34799_, _34798_, _34797_);
  nor (_34800_, _34799_, _03075_);
  or (_34801_, _34800_, _06770_);
  nor (_34803_, _34801_, _34787_);
  nor (_34804_, _34803_, _34784_);
  nor (_34805_, _34804_, _02853_);
  and (_34806_, _04660_, _06159_);
  nor (_34807_, _34771_, _05540_);
  not (_34808_, _34807_);
  nor (_34809_, _34808_, _34806_);
  or (_34810_, _34809_, _02579_);
  nor (_34811_, _34810_, _34805_);
  nor (_34812_, _12321_, _11071_);
  nor (_34814_, _34812_, _34771_);
  nor (_34815_, _34814_, _02838_);
  or (_34816_, _34815_, _02802_);
  or (_34817_, _34816_, _34811_);
  nand (_34818_, _34775_, _02802_);
  and (_34819_, _34818_, _34817_);
  and (_34820_, _34819_, _03887_);
  and (_34821_, _12211_, _04660_);
  nor (_34822_, _34821_, _34771_);
  nor (_34823_, _34822_, _03887_);
  or (_34825_, _34823_, _34820_);
  and (_34826_, _34825_, _03128_);
  nor (_34827_, _34826_, _34781_);
  nor (_34828_, _34827_, _02970_);
  nor (_34829_, _34828_, _34777_);
  nor (_34830_, _34829_, _03135_);
  nor (_34831_, _34786_, _03137_);
  and (_34832_, _34831_, _34773_);
  nor (_34833_, _34832_, _02965_);
  not (_34834_, _34833_);
  nor (_34836_, _34834_, _34830_);
  nor (_34837_, _12209_, _11071_);
  or (_34838_, _34771_, _05783_);
  nor (_34839_, _34838_, _34837_);
  or (_34840_, _34839_, _03123_);
  nor (_34841_, _34840_, _34836_);
  nor (_34842_, _12206_, _11071_);
  nor (_34843_, _34842_, _34771_);
  nor (_34844_, _34843_, _05788_);
  or (_34845_, _34844_, _03163_);
  nor (_34847_, _34845_, _34841_);
  and (_34848_, _34794_, _03163_);
  or (_34849_, _34848_, _02888_);
  nor (_34850_, _34849_, _34847_);
  and (_34851_, _12389_, _04660_);
  nor (_34852_, _34851_, _34771_);
  nor (_34853_, _34852_, _02890_);
  or (_34854_, _34853_, _34850_);
  or (_34855_, _34854_, _42672_);
  or (_34856_, _42668_, \oc8051_golden_model_1.TH1 [4]);
  and (_34858_, _34856_, _43998_);
  and (_43572_, _34858_, _34855_);
  not (_34859_, \oc8051_golden_model_1.TH1 [5]);
  nor (_34860_, _04660_, _34859_);
  and (_34861_, _12411_, _04660_);
  nor (_34862_, _34861_, _34860_);
  nor (_34863_, _34862_, _03128_);
  and (_34864_, _04660_, _04877_);
  nor (_34865_, _34864_, _34860_);
  and (_34866_, _34865_, _06770_);
  nor (_34868_, _12407_, _11071_);
  nor (_34869_, _34868_, _34860_);
  and (_34870_, _34869_, _02974_);
  and (_34871_, _04660_, \oc8051_golden_model_1.ACC [5]);
  nor (_34872_, _34871_, _34860_);
  or (_34873_, _34872_, _03814_);
  or (_34874_, _03813_, _34859_);
  and (_34875_, _34874_, _03810_);
  and (_34876_, _34875_, _34873_);
  or (_34877_, _34876_, _03069_);
  nor (_34879_, _34877_, _34870_);
  nor (_34880_, _34865_, _03336_);
  nor (_34881_, _34880_, _34879_);
  nor (_34882_, _34881_, _03075_);
  nor (_34883_, _34872_, _03084_);
  nor (_34884_, _34883_, _06770_);
  not (_34885_, _34884_);
  nor (_34886_, _34885_, _34882_);
  nor (_34887_, _34886_, _34866_);
  nor (_34888_, _34887_, _02853_);
  and (_34890_, _04660_, _06158_);
  nor (_34891_, _34860_, _05540_);
  not (_34892_, _34891_);
  nor (_34893_, _34892_, _34890_);
  or (_34894_, _34893_, _02579_);
  nor (_34895_, _34894_, _34888_);
  nor (_34896_, _12527_, _11071_);
  nor (_34897_, _34896_, _34860_);
  nor (_34898_, _34897_, _02838_);
  or (_34899_, _34898_, _02802_);
  or (_34901_, _34899_, _34895_);
  and (_34902_, _05614_, _04660_);
  nor (_34903_, _34902_, _34860_);
  nand (_34904_, _34903_, _02802_);
  and (_34905_, _34904_, _34901_);
  and (_34906_, _34905_, _03887_);
  and (_34907_, _12415_, _04660_);
  nor (_34908_, _34907_, _34860_);
  nor (_34909_, _34908_, _03887_);
  or (_34910_, _34909_, _34906_);
  and (_34912_, _34910_, _03128_);
  nor (_34913_, _34912_, _34863_);
  nor (_34914_, _34913_, _02970_);
  nor (_34915_, _34860_, _04924_);
  not (_34916_, _34915_);
  nor (_34917_, _34903_, _03883_);
  and (_34918_, _34917_, _34916_);
  nor (_34919_, _34918_, _34914_);
  nor (_34920_, _34919_, _03135_);
  nor (_34921_, _34872_, _03137_);
  and (_34922_, _34921_, _34916_);
  nor (_34923_, _34922_, _02965_);
  not (_34924_, _34923_);
  nor (_34925_, _34924_, _34920_);
  nor (_34926_, _12413_, _11071_);
  or (_34927_, _34860_, _05783_);
  nor (_34928_, _34927_, _34926_);
  or (_34929_, _34928_, _03123_);
  nor (_34930_, _34929_, _34925_);
  nor (_34931_, _12410_, _11071_);
  nor (_34934_, _34931_, _34860_);
  nor (_34935_, _34934_, _05788_);
  or (_34936_, _34935_, _03163_);
  nor (_34937_, _34936_, _34930_);
  and (_34938_, _34869_, _03163_);
  or (_34939_, _34938_, _02888_);
  nor (_34940_, _34939_, _34937_);
  and (_34941_, _12589_, _04660_);
  nor (_34942_, _34941_, _34860_);
  nor (_34943_, _34942_, _02890_);
  or (_34945_, _34943_, _34940_);
  or (_34946_, _34945_, _42672_);
  or (_34947_, _42668_, \oc8051_golden_model_1.TH1 [5]);
  and (_34948_, _34947_, _43998_);
  and (_43573_, _34948_, _34946_);
  not (_34949_, \oc8051_golden_model_1.TH1 [6]);
  nor (_34950_, _04660_, _34949_);
  and (_34951_, _12613_, _04660_);
  nor (_34952_, _34951_, _34950_);
  nor (_34953_, _34952_, _03128_);
  and (_34955_, _04660_, \oc8051_golden_model_1.ACC [6]);
  nor (_34956_, _34955_, _34950_);
  nor (_34957_, _34956_, _03084_);
  nor (_34958_, _34956_, _03814_);
  nor (_34959_, _03813_, _34949_);
  or (_34960_, _34959_, _34958_);
  and (_34961_, _34960_, _03810_);
  nor (_34962_, _12603_, _11071_);
  nor (_34963_, _34962_, _34950_);
  nor (_34964_, _34963_, _03810_);
  or (_34966_, _34964_, _34961_);
  and (_34967_, _34966_, _03336_);
  and (_34968_, _04660_, _04770_);
  nor (_34969_, _34968_, _34950_);
  nor (_34970_, _34969_, _03336_);
  nor (_34971_, _34970_, _34967_);
  nor (_34972_, _34971_, _03075_);
  or (_34973_, _34972_, _06770_);
  nor (_34974_, _34973_, _34957_);
  and (_34975_, _34969_, _06770_);
  nor (_34977_, _34975_, _34974_);
  nor (_34978_, _34977_, _02853_);
  and (_34979_, _04660_, _05849_);
  nor (_34980_, _34950_, _05540_);
  not (_34981_, _34980_);
  nor (_34982_, _34981_, _34979_);
  or (_34983_, _34982_, _02579_);
  nor (_34984_, _34983_, _34978_);
  nor (_34985_, _12722_, _11071_);
  nor (_34986_, _34985_, _34950_);
  nor (_34988_, _34986_, _02838_);
  or (_34989_, _34988_, _02802_);
  or (_34990_, _34989_, _34984_);
  and (_34991_, _12729_, _04660_);
  nor (_34992_, _34991_, _34950_);
  nand (_34993_, _34992_, _02802_);
  and (_34994_, _34993_, _34990_);
  and (_34995_, _34994_, _03887_);
  and (_34996_, _12739_, _04660_);
  nor (_34997_, _34996_, _34950_);
  nor (_34999_, _34997_, _03887_);
  or (_35000_, _34999_, _34995_);
  and (_35001_, _35000_, _03128_);
  nor (_35002_, _35001_, _34953_);
  nor (_35003_, _35002_, _02970_);
  nor (_35004_, _34950_, _04819_);
  not (_35005_, _35004_);
  nor (_35006_, _34992_, _03883_);
  and (_35007_, _35006_, _35005_);
  nor (_35008_, _35007_, _35003_);
  nor (_35010_, _35008_, _03135_);
  nor (_35011_, _34956_, _03137_);
  and (_35012_, _35011_, _35005_);
  or (_35013_, _35012_, _35010_);
  and (_35014_, _35013_, _05783_);
  nor (_35015_, _12737_, _11071_);
  nor (_35016_, _35015_, _34950_);
  nor (_35017_, _35016_, _05783_);
  or (_35018_, _35017_, _35014_);
  and (_35019_, _35018_, _05788_);
  nor (_35021_, _12612_, _11071_);
  nor (_35022_, _35021_, _34950_);
  nor (_35023_, _35022_, _05788_);
  or (_35024_, _35023_, _03163_);
  nor (_35025_, _35024_, _35019_);
  and (_35026_, _34963_, _03163_);
  or (_35027_, _35026_, _02888_);
  nor (_35028_, _35027_, _35025_);
  and (_35029_, _12794_, _04660_);
  nor (_35030_, _35029_, _34950_);
  nor (_35032_, _35030_, _02890_);
  or (_35033_, _35032_, _35028_);
  or (_35034_, _35033_, _42672_);
  or (_35035_, _42668_, \oc8051_golden_model_1.TH1 [6]);
  and (_35036_, _35035_, _43998_);
  and (_43574_, _35036_, _35034_);
  not (_35037_, \oc8051_golden_model_1.TL0 [0]);
  nor (_35038_, _04676_, _35037_);
  and (_35039_, _05226_, _04676_);
  nor (_35040_, _35039_, _35038_);
  and (_35042_, _35040_, _16625_);
  and (_35043_, _04676_, \oc8051_golden_model_1.ACC [0]);
  nor (_35044_, _35043_, _35038_);
  nor (_35045_, _35044_, _03084_);
  nor (_35046_, _35044_, _03814_);
  nor (_35047_, _03813_, _35037_);
  or (_35048_, _35047_, _35046_);
  and (_35049_, _35048_, _03810_);
  nor (_35050_, _35040_, _03810_);
  or (_35051_, _35050_, _35049_);
  and (_35053_, _35051_, _03336_);
  and (_35054_, _04676_, _03808_);
  nor (_35055_, _35054_, _35038_);
  nor (_35056_, _35055_, _03336_);
  nor (_35057_, _35056_, _35053_);
  nor (_35058_, _35057_, _03075_);
  or (_35059_, _35058_, _06770_);
  nor (_35060_, _35059_, _35045_);
  and (_35061_, _35055_, _06770_);
  nor (_35062_, _35061_, _35060_);
  nor (_35064_, _35062_, _02853_);
  and (_35065_, _04676_, _06152_);
  nor (_35066_, _35038_, _05540_);
  not (_35067_, _35066_);
  nor (_35068_, _35067_, _35065_);
  nor (_35069_, _35068_, _35064_);
  and (_35070_, _35069_, _02838_);
  nor (_35071_, _11505_, _11152_);
  nor (_35072_, _35071_, _35038_);
  nor (_35073_, _35072_, _02838_);
  or (_35075_, _35073_, _35070_);
  and (_35076_, _35075_, _02803_);
  and (_35077_, _04676_, _05672_);
  nor (_35078_, _35077_, _35038_);
  nor (_35079_, _35078_, _02803_);
  or (_35080_, _35079_, _35076_);
  and (_35081_, _35080_, _03887_);
  and (_35082_, _11399_, _04676_);
  nor (_35083_, _35082_, _35038_);
  nor (_35084_, _35083_, _03887_);
  or (_35086_, _35084_, _35081_);
  and (_35087_, _35086_, _03128_);
  and (_35088_, _11522_, _04676_);
  nor (_35089_, _35088_, _35038_);
  nor (_35090_, _35089_, _03128_);
  or (_35091_, _35090_, _35087_);
  and (_35092_, _35091_, _03883_);
  or (_35093_, _35078_, _03883_);
  nor (_35094_, _35093_, _35039_);
  nor (_35095_, _35094_, _35092_);
  nor (_35097_, _35095_, _03135_);
  nor (_35098_, _35038_, _09409_);
  or (_35099_, _35098_, _03137_);
  nor (_35100_, _35099_, _35044_);
  or (_35101_, _35100_, _35097_);
  and (_35102_, _35101_, _05783_);
  nor (_35103_, _11396_, _11152_);
  nor (_35104_, _35103_, _35038_);
  nor (_35105_, _35104_, _05783_);
  or (_35106_, _35105_, _35102_);
  and (_35108_, _35106_, _05788_);
  nor (_35109_, _11520_, _11152_);
  nor (_35110_, _35109_, _35038_);
  nor (_35111_, _35110_, _05788_);
  nor (_35112_, _35111_, _16625_);
  not (_35113_, _35112_);
  nor (_35114_, _35113_, _35108_);
  nor (_35115_, _35114_, _35042_);
  or (_35116_, _35115_, _42672_);
  or (_35117_, _42668_, \oc8051_golden_model_1.TL0 [0]);
  and (_35119_, _35117_, _43998_);
  and (_43576_, _35119_, _35116_);
  nor (_35120_, _04676_, \oc8051_golden_model_1.TL0 [1]);
  nor (_35121_, _11152_, _04000_);
  or (_35122_, _35121_, _35120_);
  nor (_35123_, _35122_, _03336_);
  and (_35124_, _04676_, _02551_);
  nor (_35125_, _35124_, _35120_);
  and (_35126_, _35125_, _03813_);
  not (_35127_, \oc8051_golden_model_1.TL0 [1]);
  nor (_35129_, _03813_, _35127_);
  or (_35130_, _35129_, _35126_);
  and (_35131_, _35130_, _03810_);
  and (_35132_, _11606_, _04676_);
  nor (_35133_, _35132_, _35120_);
  and (_35134_, _35133_, _02974_);
  or (_35135_, _35134_, _35131_);
  and (_35136_, _35135_, _03336_);
  nor (_35137_, _35136_, _35123_);
  nor (_35138_, _35137_, _03075_);
  and (_35140_, _35125_, _03075_);
  nor (_35141_, _35140_, _06770_);
  not (_35142_, _35141_);
  nor (_35143_, _35142_, _35138_);
  and (_35144_, _35122_, _06770_);
  or (_35145_, _35144_, _02853_);
  nor (_35146_, _35145_, _35143_);
  or (_35147_, _11152_, _06151_);
  nor (_35148_, _35120_, _05540_);
  and (_35149_, _35148_, _35147_);
  or (_35151_, _35149_, _35146_);
  and (_35152_, _35151_, _02838_);
  not (_35153_, _35120_);
  and (_35154_, _11695_, _04676_);
  nor (_35155_, _35154_, _02838_);
  and (_35156_, _35155_, _35153_);
  nor (_35157_, _35156_, _35152_);
  nor (_35158_, _35157_, _02802_);
  and (_35159_, _04676_, _03698_);
  not (_35160_, _35159_);
  nor (_35162_, _35120_, _02803_);
  and (_35163_, _35162_, _35160_);
  nor (_35164_, _35163_, _35158_);
  nor (_35165_, _35164_, _02980_);
  nor (_35166_, _11710_, _11152_);
  nor (_35167_, _35166_, _03887_);
  and (_35168_, _35167_, _35153_);
  nor (_35169_, _35168_, _35165_);
  nor (_35170_, _35169_, _03127_);
  nor (_35171_, _11715_, _11152_);
  nor (_35173_, _35171_, _03128_);
  and (_35174_, _35173_, _35153_);
  nor (_35175_, _35174_, _35170_);
  nor (_35176_, _35175_, _02970_);
  nor (_35177_, _11709_, _11152_);
  nor (_35178_, _35177_, _03883_);
  and (_35179_, _35178_, _35153_);
  nor (_35180_, _35179_, _35176_);
  nor (_35181_, _35180_, _03135_);
  nor (_35182_, _04676_, _35127_);
  nor (_35184_, _35182_, _13722_);
  nor (_35185_, _35184_, _03137_);
  and (_35186_, _35185_, _35125_);
  nor (_35187_, _35186_, _35181_);
  or (_35188_, _35187_, _17961_);
  and (_35189_, _35124_, _05178_);
  or (_35190_, _35189_, _05788_);
  or (_35191_, _35190_, _35120_);
  and (_35192_, _35191_, _03906_);
  and (_35193_, _35159_, _05178_);
  or (_35195_, _35120_, _05783_);
  or (_35196_, _35195_, _35193_);
  and (_35197_, _35196_, _35192_);
  and (_35198_, _35197_, _35188_);
  nor (_35199_, _35133_, _03906_);
  nor (_35200_, _35199_, _35198_);
  nor (_35201_, _35200_, _02888_);
  nor (_35202_, _35132_, _35182_);
  and (_35203_, _35202_, _02888_);
  nor (_35204_, _35203_, _35201_);
  or (_35206_, _35204_, _42672_);
  or (_35207_, _42668_, \oc8051_golden_model_1.TL0 [1]);
  and (_35208_, _35207_, _43998_);
  and (_43577_, _35208_, _35206_);
  not (_35209_, \oc8051_golden_model_1.TL0 [2]);
  nor (_35210_, _04676_, _35209_);
  nor (_35211_, _35210_, _05130_);
  not (_35212_, _35211_);
  and (_35213_, _04676_, _05701_);
  nor (_35214_, _35213_, _35210_);
  nor (_35216_, _35214_, _03883_);
  and (_35217_, _35216_, _35212_);
  and (_35218_, _11927_, _04676_);
  nor (_35219_, _35218_, _35210_);
  nor (_35220_, _35219_, _03128_);
  and (_35221_, _04676_, \oc8051_golden_model_1.ACC [2]);
  nor (_35222_, _35221_, _35210_);
  nor (_35223_, _35222_, _03084_);
  nor (_35224_, _35222_, _03814_);
  nor (_35225_, _03813_, _35209_);
  or (_35227_, _35225_, _35224_);
  and (_35228_, _35227_, _03810_);
  nor (_35229_, _11801_, _11152_);
  nor (_35230_, _35229_, _35210_);
  nor (_35231_, _35230_, _03810_);
  or (_35232_, _35231_, _35228_);
  and (_35233_, _35232_, _03336_);
  and (_35234_, _04676_, _04435_);
  nor (_35235_, _35234_, _35210_);
  nor (_35236_, _35235_, _03336_);
  nor (_35238_, _35236_, _35233_);
  nor (_35239_, _35238_, _03075_);
  or (_35240_, _35239_, _06770_);
  nor (_35241_, _35240_, _35223_);
  and (_35242_, _35235_, _06770_);
  nor (_35243_, _35242_, _35241_);
  nor (_35244_, _35243_, _02853_);
  and (_35245_, _04676_, _06155_);
  nor (_35246_, _35210_, _05540_);
  not (_35247_, _35246_);
  nor (_35249_, _35247_, _35245_);
  or (_35250_, _35249_, _02579_);
  nor (_35251_, _35250_, _35244_);
  nor (_35252_, _11906_, _11152_);
  nor (_35253_, _35252_, _35210_);
  nor (_35254_, _35253_, _02838_);
  or (_35255_, _35254_, _02802_);
  or (_35256_, _35255_, _35251_);
  nand (_35257_, _35214_, _02802_);
  and (_35258_, _35257_, _35256_);
  and (_35260_, _35258_, _03887_);
  and (_35261_, _11921_, _04676_);
  nor (_35262_, _35261_, _35210_);
  nor (_35263_, _35262_, _03887_);
  or (_35264_, _35263_, _35260_);
  and (_35265_, _35264_, _03128_);
  nor (_35266_, _35265_, _35220_);
  nor (_35267_, _35266_, _02970_);
  nor (_35268_, _35267_, _35217_);
  nor (_35269_, _35268_, _03135_);
  nor (_35271_, _35222_, _03137_);
  and (_35272_, _35271_, _35212_);
  or (_35273_, _35272_, _35269_);
  and (_35274_, _35273_, _05783_);
  nor (_35275_, _11919_, _11152_);
  nor (_35276_, _35275_, _35210_);
  nor (_35277_, _35276_, _05783_);
  or (_35278_, _35277_, _35274_);
  and (_35279_, _35278_, _05788_);
  nor (_35280_, _11926_, _11152_);
  nor (_35282_, _35280_, _35210_);
  nor (_35283_, _35282_, _05788_);
  or (_35284_, _35283_, _03163_);
  nor (_35285_, _35284_, _35279_);
  and (_35286_, _35230_, _03163_);
  or (_35287_, _35286_, _02888_);
  nor (_35288_, _35287_, _35285_);
  and (_35289_, _11985_, _04676_);
  nor (_35290_, _35289_, _35210_);
  nor (_35291_, _35290_, _02890_);
  or (_35293_, _35291_, _35288_);
  or (_35294_, _35293_, _42672_);
  or (_35295_, _42668_, \oc8051_golden_model_1.TL0 [2]);
  and (_35296_, _35295_, _43998_);
  and (_43578_, _35296_, _35294_);
  not (_35297_, \oc8051_golden_model_1.TL0 [3]);
  nor (_35298_, _04676_, _35297_);
  and (_35299_, _12133_, _04676_);
  nor (_35300_, _35299_, _35298_);
  nor (_35301_, _35300_, _03128_);
  and (_35303_, _04676_, \oc8051_golden_model_1.ACC [3]);
  nor (_35304_, _35303_, _35298_);
  nor (_35305_, _35304_, _03814_);
  nor (_35306_, _03813_, _35297_);
  or (_35307_, _35306_, _35305_);
  and (_35308_, _35307_, _03810_);
  nor (_35309_, _12017_, _11152_);
  nor (_35310_, _35309_, _35298_);
  nor (_35311_, _35310_, _03810_);
  or (_35312_, _35311_, _35308_);
  and (_35314_, _35312_, _03336_);
  and (_35315_, _04676_, _04241_);
  nor (_35316_, _35315_, _35298_);
  nor (_35317_, _35316_, _03336_);
  nor (_35318_, _35317_, _35314_);
  nor (_35319_, _35318_, _03075_);
  nor (_35320_, _35304_, _03084_);
  nor (_35321_, _35320_, _06770_);
  not (_35322_, _35321_);
  nor (_35323_, _35322_, _35319_);
  and (_35325_, _35316_, _06770_);
  or (_35326_, _35325_, _02853_);
  nor (_35327_, _35326_, _35323_);
  and (_35328_, _04676_, _06154_);
  or (_35329_, _35328_, _35298_);
  and (_35330_, _35329_, _02853_);
  or (_35331_, _35330_, _02579_);
  or (_35332_, _35331_, _35327_);
  nor (_35333_, _12112_, _11152_);
  or (_35334_, _35298_, _02838_);
  or (_35336_, _35334_, _35333_);
  and (_35337_, _35336_, _02803_);
  and (_35338_, _35337_, _35332_);
  and (_35339_, _04676_, _05658_);
  nor (_35340_, _35339_, _35298_);
  nor (_35341_, _35340_, _02803_);
  or (_35342_, _35341_, _35338_);
  and (_35343_, _35342_, _03887_);
  and (_35344_, _12127_, _04676_);
  nor (_35345_, _35344_, _35298_);
  nor (_35347_, _35345_, _03887_);
  or (_35348_, _35347_, _35343_);
  and (_35349_, _35348_, _03128_);
  nor (_35350_, _35349_, _35301_);
  nor (_35351_, _35350_, _02970_);
  nor (_35352_, _35298_, _05079_);
  not (_35353_, _35352_);
  nor (_35354_, _35340_, _03883_);
  and (_35355_, _35354_, _35353_);
  nor (_35356_, _35355_, _35351_);
  nor (_35358_, _35356_, _03135_);
  nor (_35359_, _35304_, _03137_);
  and (_35360_, _35359_, _35353_);
  or (_35361_, _35360_, _35358_);
  and (_35362_, _35361_, _05783_);
  nor (_35363_, _12125_, _11152_);
  nor (_35364_, _35363_, _35298_);
  nor (_35365_, _35364_, _05783_);
  or (_35366_, _35365_, _35362_);
  and (_35367_, _35366_, _05788_);
  nor (_35369_, _12132_, _11152_);
  nor (_35370_, _35369_, _35298_);
  nor (_35371_, _35370_, _05788_);
  or (_35372_, _35371_, _03163_);
  nor (_35373_, _35372_, _35367_);
  and (_35374_, _35310_, _03163_);
  or (_35375_, _35374_, _02888_);
  nor (_35376_, _35375_, _35373_);
  and (_35377_, _12183_, _04676_);
  nor (_35378_, _35377_, _35298_);
  nor (_35380_, _35378_, _02890_);
  or (_35381_, _35380_, _35376_);
  or (_35382_, _35381_, _42672_);
  or (_35383_, _42668_, \oc8051_golden_model_1.TL0 [3]);
  and (_35384_, _35383_, _43998_);
  and (_43579_, _35384_, _35382_);
  not (_35385_, \oc8051_golden_model_1.TL0 [4]);
  nor (_35386_, _04676_, _35385_);
  nor (_35387_, _35386_, _05031_);
  not (_35388_, _35387_);
  and (_35390_, _05666_, _04676_);
  nor (_35391_, _35390_, _35386_);
  nor (_35392_, _35391_, _03883_);
  and (_35393_, _35392_, _35388_);
  and (_35394_, _12207_, _04676_);
  nor (_35395_, _35394_, _35386_);
  nor (_35396_, _35395_, _03128_);
  and (_35397_, _04676_, \oc8051_golden_model_1.ACC [4]);
  nor (_35398_, _35397_, _35386_);
  nor (_35399_, _35398_, _03084_);
  nor (_35401_, _35398_, _03814_);
  nor (_35402_, _03813_, _35385_);
  or (_35403_, _35402_, _35401_);
  and (_35404_, _35403_, _03810_);
  nor (_35405_, _12217_, _11152_);
  nor (_35406_, _35405_, _35386_);
  nor (_35407_, _35406_, _03810_);
  or (_35408_, _35407_, _35404_);
  and (_35409_, _35408_, _03336_);
  and (_35410_, _04676_, _04982_);
  nor (_35412_, _35410_, _35386_);
  nor (_35413_, _35412_, _03336_);
  nor (_35414_, _35413_, _35409_);
  nor (_35415_, _35414_, _03075_);
  or (_35416_, _35415_, _06770_);
  nor (_35417_, _35416_, _35399_);
  and (_35418_, _35412_, _06770_);
  nor (_35419_, _35418_, _35417_);
  nor (_35420_, _35419_, _02853_);
  and (_35421_, _04676_, _06159_);
  nor (_35423_, _35386_, _05540_);
  not (_35424_, _35423_);
  nor (_35425_, _35424_, _35421_);
  or (_35426_, _35425_, _02579_);
  nor (_35427_, _35426_, _35420_);
  nor (_35428_, _12321_, _11152_);
  nor (_35429_, _35428_, _35386_);
  nor (_35430_, _35429_, _02838_);
  or (_35431_, _35430_, _02802_);
  or (_35432_, _35431_, _35427_);
  nand (_35434_, _35391_, _02802_);
  and (_35435_, _35434_, _35432_);
  and (_35436_, _35435_, _03887_);
  and (_35437_, _12211_, _04676_);
  nor (_35438_, _35437_, _35386_);
  nor (_35439_, _35438_, _03887_);
  or (_35440_, _35439_, _35436_);
  and (_35441_, _35440_, _03128_);
  nor (_35442_, _35441_, _35396_);
  nor (_35443_, _35442_, _02970_);
  nor (_35445_, _35443_, _35393_);
  nor (_35446_, _35445_, _03135_);
  nor (_35447_, _35398_, _03137_);
  and (_35448_, _35447_, _35388_);
  or (_35449_, _35448_, _35446_);
  and (_35450_, _35449_, _05783_);
  nor (_35451_, _12209_, _11152_);
  nor (_35452_, _35451_, _35386_);
  nor (_35453_, _35452_, _05783_);
  or (_35454_, _35453_, _35450_);
  and (_35456_, _35454_, _05788_);
  nor (_35457_, _12206_, _11152_);
  nor (_35458_, _35457_, _35386_);
  nor (_35459_, _35458_, _05788_);
  or (_35460_, _35459_, _03163_);
  nor (_35461_, _35460_, _35456_);
  and (_35462_, _35406_, _03163_);
  or (_35463_, _35462_, _02888_);
  nor (_35464_, _35463_, _35461_);
  and (_35465_, _12389_, _04676_);
  nor (_35467_, _35465_, _35386_);
  nor (_35468_, _35467_, _02890_);
  or (_35469_, _35468_, _35464_);
  or (_35470_, _35469_, _42672_);
  or (_35471_, _42668_, \oc8051_golden_model_1.TL0 [4]);
  and (_35472_, _35471_, _43998_);
  and (_43581_, _35472_, _35470_);
  not (_35473_, \oc8051_golden_model_1.TL0 [5]);
  nor (_35474_, _04676_, _35473_);
  and (_35475_, _12411_, _04676_);
  nor (_35477_, _35475_, _35474_);
  nor (_35478_, _35477_, _03128_);
  and (_35479_, _04676_, \oc8051_golden_model_1.ACC [5]);
  nor (_35480_, _35479_, _35474_);
  nor (_35481_, _35480_, _03084_);
  nor (_35482_, _12407_, _11152_);
  nor (_35483_, _35482_, _35474_);
  and (_35484_, _35483_, _02974_);
  or (_35485_, _35480_, _03814_);
  or (_35486_, _03813_, _35473_);
  and (_35488_, _35486_, _03810_);
  and (_35489_, _35488_, _35485_);
  or (_35490_, _35489_, _03069_);
  nor (_35491_, _35490_, _35484_);
  and (_35492_, _04676_, _04877_);
  nor (_35493_, _35492_, _35474_);
  nor (_35494_, _35493_, _03336_);
  nor (_35495_, _35494_, _35491_);
  nor (_35496_, _35495_, _03075_);
  or (_35497_, _35496_, _06770_);
  nor (_35499_, _35497_, _35481_);
  and (_35500_, _35493_, _06770_);
  nor (_35501_, _35500_, _35499_);
  nor (_35502_, _35501_, _02853_);
  and (_35503_, _04676_, _06158_);
  nor (_35504_, _35474_, _05540_);
  not (_35505_, _35504_);
  nor (_35506_, _35505_, _35503_);
  or (_35507_, _35506_, _02579_);
  nor (_35508_, _35507_, _35502_);
  nor (_35510_, _12527_, _11152_);
  nor (_35511_, _35510_, _35474_);
  nor (_35512_, _35511_, _02838_);
  or (_35513_, _35512_, _02802_);
  or (_35514_, _35513_, _35508_);
  and (_35515_, _05614_, _04676_);
  nor (_35516_, _35515_, _35474_);
  nand (_35517_, _35516_, _02802_);
  and (_35518_, _35517_, _35514_);
  and (_35519_, _35518_, _03887_);
  and (_35521_, _12415_, _04676_);
  nor (_35522_, _35521_, _35474_);
  nor (_35523_, _35522_, _03887_);
  or (_35524_, _35523_, _35519_);
  and (_35525_, _35524_, _03128_);
  nor (_35526_, _35525_, _35478_);
  nor (_35527_, _35526_, _02970_);
  nor (_35528_, _35474_, _04924_);
  not (_35529_, _35528_);
  nor (_35530_, _35516_, _03883_);
  and (_35532_, _35530_, _35529_);
  nor (_35533_, _35532_, _35527_);
  nor (_35534_, _35533_, _03135_);
  nor (_35535_, _35480_, _03137_);
  and (_35536_, _35535_, _35529_);
  or (_35537_, _35536_, _35534_);
  and (_35538_, _35537_, _05783_);
  nor (_35539_, _12413_, _11152_);
  nor (_35540_, _35539_, _35474_);
  nor (_35541_, _35540_, _05783_);
  or (_35543_, _35541_, _35538_);
  and (_35544_, _35543_, _05788_);
  nor (_35545_, _12410_, _11152_);
  nor (_35546_, _35545_, _35474_);
  nor (_35547_, _35546_, _05788_);
  or (_35548_, _35547_, _03163_);
  nor (_35549_, _35548_, _35544_);
  and (_35550_, _35483_, _03163_);
  or (_35551_, _35550_, _02888_);
  nor (_35552_, _35551_, _35549_);
  and (_35554_, _12589_, _04676_);
  nor (_35555_, _35554_, _35474_);
  nor (_35556_, _35555_, _02890_);
  or (_35557_, _35556_, _35552_);
  or (_35558_, _35557_, _42672_);
  or (_35559_, _42668_, \oc8051_golden_model_1.TL0 [5]);
  and (_35560_, _35559_, _43998_);
  and (_43582_, _35560_, _35558_);
  not (_35561_, \oc8051_golden_model_1.TL0 [6]);
  nor (_35562_, _04676_, _35561_);
  and (_35564_, _12613_, _04676_);
  nor (_35565_, _35564_, _35562_);
  nor (_35566_, _35565_, _03128_);
  and (_35567_, _04676_, \oc8051_golden_model_1.ACC [6]);
  nor (_35568_, _35567_, _35562_);
  nor (_35569_, _35568_, _03084_);
  nor (_35570_, _35568_, _03814_);
  nor (_35571_, _03813_, _35561_);
  or (_35572_, _35571_, _35570_);
  and (_35573_, _35572_, _03810_);
  nor (_35575_, _12603_, _11152_);
  nor (_35576_, _35575_, _35562_);
  nor (_35577_, _35576_, _03810_);
  or (_35578_, _35577_, _35573_);
  and (_35579_, _35578_, _03336_);
  and (_35580_, _04676_, _04770_);
  nor (_35581_, _35580_, _35562_);
  nor (_35582_, _35581_, _03336_);
  nor (_35583_, _35582_, _35579_);
  nor (_35584_, _35583_, _03075_);
  or (_35586_, _35584_, _06770_);
  nor (_35587_, _35586_, _35569_);
  and (_35588_, _35581_, _06770_);
  nor (_35589_, _35588_, _35587_);
  nor (_35590_, _35589_, _02853_);
  and (_35591_, _04676_, _05849_);
  nor (_35592_, _35562_, _05540_);
  not (_35593_, _35592_);
  nor (_35594_, _35593_, _35591_);
  or (_35595_, _35594_, _02579_);
  nor (_35597_, _35595_, _35590_);
  nor (_35598_, _12722_, _11152_);
  nor (_35599_, _35598_, _35562_);
  nor (_35600_, _35599_, _02838_);
  or (_35601_, _35600_, _02802_);
  or (_35602_, _35601_, _35597_);
  and (_35603_, _12729_, _04676_);
  nor (_35604_, _35603_, _35562_);
  nand (_35605_, _35604_, _02802_);
  and (_35606_, _35605_, _35602_);
  and (_35608_, _35606_, _03887_);
  and (_35609_, _12739_, _04676_);
  nor (_35610_, _35609_, _35562_);
  nor (_35611_, _35610_, _03887_);
  or (_35612_, _35611_, _35608_);
  and (_35613_, _35612_, _03128_);
  nor (_35614_, _35613_, _35566_);
  nor (_35615_, _35614_, _02970_);
  nor (_35616_, _35562_, _04819_);
  not (_35617_, _35616_);
  nor (_35619_, _35604_, _03883_);
  and (_35620_, _35619_, _35617_);
  nor (_35621_, _35620_, _35615_);
  nor (_35622_, _35621_, _03135_);
  nor (_35623_, _35568_, _03137_);
  and (_35624_, _35623_, _35617_);
  or (_35625_, _35624_, _35622_);
  and (_35626_, _35625_, _05783_);
  nor (_35627_, _12737_, _11152_);
  nor (_35628_, _35627_, _35562_);
  nor (_35630_, _35628_, _05783_);
  or (_35631_, _35630_, _35626_);
  and (_35632_, _35631_, _05788_);
  nor (_35633_, _12612_, _11152_);
  nor (_35634_, _35633_, _35562_);
  nor (_35635_, _35634_, _05788_);
  or (_35636_, _35635_, _03163_);
  nor (_35637_, _35636_, _35632_);
  and (_35638_, _35576_, _03163_);
  or (_35639_, _35638_, _02888_);
  nor (_35642_, _35639_, _35637_);
  and (_35643_, _12794_, _04676_);
  nor (_35644_, _35643_, _35562_);
  nor (_35645_, _35644_, _02890_);
  or (_35646_, _35645_, _35642_);
  or (_35647_, _35646_, _42672_);
  or (_35648_, _42668_, \oc8051_golden_model_1.TL0 [6]);
  and (_35649_, _35648_, _43998_);
  and (_43583_, _35649_, _35647_);
  not (_35650_, \oc8051_golden_model_1.TL1 [0]);
  nor (_35652_, _04656_, _35650_);
  and (_35653_, _05226_, _04656_);
  nor (_35654_, _35653_, _35652_);
  and (_35655_, _35654_, _16625_);
  and (_35656_, _04656_, _03808_);
  nor (_35657_, _35656_, _35652_);
  and (_35658_, _35657_, _06770_);
  and (_35659_, _04656_, \oc8051_golden_model_1.ACC [0]);
  nor (_35660_, _35659_, _35652_);
  nor (_35661_, _35660_, _03814_);
  nor (_35664_, _03813_, _35650_);
  or (_35665_, _35664_, _35661_);
  and (_35666_, _35665_, _03810_);
  nor (_35667_, _35654_, _03810_);
  or (_35668_, _35667_, _35666_);
  and (_35669_, _35668_, _03336_);
  nor (_35670_, _35657_, _03336_);
  nor (_35671_, _35670_, _35669_);
  nor (_35672_, _35671_, _03075_);
  nor (_35673_, _35660_, _03084_);
  nor (_35675_, _35673_, _06770_);
  not (_35676_, _35675_);
  nor (_35677_, _35676_, _35672_);
  nor (_35678_, _35677_, _35658_);
  nor (_35679_, _35678_, _02853_);
  and (_35680_, _04656_, _06152_);
  nor (_35681_, _35652_, _05540_);
  not (_35682_, _35681_);
  nor (_35683_, _35682_, _35680_);
  nor (_35684_, _35683_, _35679_);
  and (_35687_, _35684_, _02838_);
  nor (_35688_, _11505_, _11233_);
  nor (_35689_, _35688_, _35652_);
  nor (_35690_, _35689_, _02838_);
  or (_35691_, _35690_, _35687_);
  and (_35692_, _35691_, _02803_);
  and (_35693_, _04656_, _05672_);
  nor (_35694_, _35693_, _35652_);
  nor (_35695_, _35694_, _02803_);
  or (_35696_, _35695_, _35692_);
  and (_35698_, _35696_, _03887_);
  and (_35699_, _11399_, _04656_);
  nor (_35700_, _35699_, _35652_);
  nor (_35701_, _35700_, _03887_);
  or (_35702_, _35701_, _35698_);
  and (_35703_, _35702_, _03128_);
  and (_35704_, _11522_, _04656_);
  nor (_35705_, _35704_, _35652_);
  nor (_35706_, _35705_, _03128_);
  or (_35707_, _35706_, _35703_);
  and (_35710_, _35707_, _03883_);
  or (_35711_, _35694_, _03883_);
  nor (_35712_, _35711_, _35653_);
  nor (_35713_, _35712_, _35710_);
  nor (_35714_, _35713_, _03135_);
  nor (_35715_, _35652_, _09409_);
  or (_35716_, _35715_, _03137_);
  nor (_35717_, _35716_, _35660_);
  or (_35718_, _35717_, _35714_);
  and (_35719_, _35718_, _05783_);
  nor (_35721_, _11396_, _11233_);
  nor (_35722_, _35721_, _35652_);
  nor (_35723_, _35722_, _05783_);
  or (_35724_, _35723_, _35719_);
  and (_35725_, _35724_, _05788_);
  nor (_35726_, _11520_, _11233_);
  nor (_35727_, _35726_, _35652_);
  nor (_35728_, _35727_, _05788_);
  nor (_35729_, _35728_, _16625_);
  not (_35730_, _35729_);
  nor (_35732_, _35730_, _35725_);
  nor (_35733_, _35732_, _35655_);
  or (_35734_, _35733_, _42672_);
  or (_35735_, _42668_, \oc8051_golden_model_1.TL1 [0]);
  and (_35736_, _35735_, _43998_);
  and (_43584_, _35736_, _35734_);
  nor (_35737_, _04656_, \oc8051_golden_model_1.TL1 [1]);
  and (_35738_, _04656_, _02551_);
  nor (_35739_, _35738_, _35737_);
  and (_35740_, _35739_, _03075_);
  nor (_35742_, _11233_, _04000_);
  or (_35743_, _35742_, _35737_);
  nor (_35744_, _35743_, _03336_);
  and (_35745_, _35739_, _03813_);
  not (_35746_, \oc8051_golden_model_1.TL1 [1]);
  nor (_35747_, _03813_, _35746_);
  or (_35748_, _35747_, _35745_);
  and (_35749_, _35748_, _03810_);
  and (_35750_, _11606_, _04656_);
  nor (_35751_, _35750_, _35737_);
  and (_35753_, _35751_, _02974_);
  or (_35754_, _35753_, _35749_);
  and (_35755_, _35754_, _03336_);
  nor (_35756_, _35755_, _35744_);
  nor (_35757_, _35756_, _03075_);
  or (_35758_, _35757_, _06770_);
  nor (_35759_, _35758_, _35740_);
  and (_35760_, _35743_, _06770_);
  or (_35761_, _35760_, _02853_);
  nor (_35762_, _35761_, _35759_);
  or (_35764_, _11233_, _06151_);
  nor (_35765_, _35737_, _05540_);
  and (_35766_, _35765_, _35764_);
  or (_35767_, _35766_, _35762_);
  and (_35768_, _35767_, _02838_);
  not (_35769_, _35737_);
  and (_35770_, _11695_, _04656_);
  nor (_35771_, _35770_, _02838_);
  and (_35772_, _35771_, _35769_);
  nor (_35773_, _35772_, _35768_);
  nor (_35775_, _35773_, _02802_);
  and (_35776_, _04656_, _03698_);
  not (_35777_, _35776_);
  nor (_35778_, _35737_, _02803_);
  and (_35779_, _35778_, _35777_);
  nor (_35780_, _35779_, _35775_);
  nor (_35781_, _35780_, _02980_);
  nor (_35782_, _11710_, _11233_);
  nor (_35783_, _35782_, _03887_);
  and (_35784_, _35783_, _35769_);
  nor (_35786_, _35784_, _35781_);
  nor (_35787_, _35786_, _03127_);
  nor (_35788_, _11715_, _11233_);
  nor (_35789_, _35788_, _03128_);
  and (_35790_, _35789_, _35769_);
  nor (_35791_, _35790_, _35787_);
  nor (_35792_, _35791_, _02970_);
  nor (_35793_, _11709_, _11233_);
  nor (_35794_, _35793_, _03883_);
  and (_35795_, _35794_, _35769_);
  nor (_35797_, _35795_, _35792_);
  nor (_35798_, _35797_, _03135_);
  nor (_35799_, _04656_, _35746_);
  nor (_35800_, _35799_, _13722_);
  nor (_35801_, _35800_, _03137_);
  and (_35802_, _35801_, _35739_);
  nor (_35803_, _35802_, _35798_);
  or (_35804_, _35803_, _17961_);
  and (_35805_, _11714_, _04656_);
  or (_35806_, _35805_, _05788_);
  or (_35808_, _35806_, _35737_);
  and (_35809_, _35808_, _03906_);
  and (_35810_, _35776_, _05178_);
  or (_35811_, _35737_, _05783_);
  or (_35812_, _35811_, _35810_);
  and (_35813_, _35812_, _35809_);
  and (_35814_, _35813_, _35804_);
  nor (_35815_, _35751_, _03906_);
  nor (_35816_, _35815_, _35814_);
  and (_35817_, _35816_, _02890_);
  nor (_35819_, _35750_, _35799_);
  nor (_35820_, _35819_, _02890_);
  or (_35821_, _35820_, _35817_);
  or (_35822_, _35821_, _42672_);
  or (_35823_, _42668_, \oc8051_golden_model_1.TL1 [1]);
  and (_35824_, _35823_, _43998_);
  and (_43585_, _35824_, _35822_);
  not (_35825_, \oc8051_golden_model_1.TL1 [2]);
  nor (_35826_, _04656_, _35825_);
  nor (_35827_, _35826_, _05130_);
  not (_35829_, _35827_);
  and (_35830_, _04656_, _05701_);
  nor (_35831_, _35830_, _35826_);
  nor (_35832_, _35831_, _03883_);
  and (_35833_, _35832_, _35829_);
  and (_35834_, _04656_, _04435_);
  nor (_35835_, _35834_, _35826_);
  and (_35836_, _35835_, _06770_);
  nor (_35837_, _11801_, _11233_);
  nor (_35838_, _35837_, _35826_);
  nor (_35840_, _35838_, _03810_);
  nor (_35841_, _03813_, _35825_);
  and (_35842_, _04656_, \oc8051_golden_model_1.ACC [2]);
  nor (_35843_, _35842_, _35826_);
  nor (_35844_, _35843_, _03814_);
  nor (_35845_, _35844_, _35841_);
  nor (_35846_, _35845_, _02974_);
  or (_35847_, _35846_, _35840_);
  and (_35848_, _35847_, _03336_);
  nor (_35849_, _35835_, _03336_);
  or (_35851_, _35849_, _35848_);
  and (_35852_, _35851_, _03084_);
  nor (_35853_, _35843_, _03084_);
  nor (_35854_, _35853_, _06770_);
  not (_35855_, _35854_);
  nor (_35856_, _35855_, _35852_);
  nor (_35857_, _35856_, _35836_);
  nor (_35858_, _35857_, _02853_);
  and (_35859_, _04656_, _06155_);
  nor (_35860_, _35826_, _05540_);
  not (_35862_, _35860_);
  nor (_35863_, _35862_, _35859_);
  nor (_35864_, _35863_, _35858_);
  and (_35865_, _35864_, _02838_);
  nor (_35866_, _11906_, _11233_);
  nor (_35867_, _35866_, _35826_);
  nor (_35868_, _35867_, _02838_);
  or (_35869_, _35868_, _35865_);
  and (_35870_, _35869_, _02803_);
  nor (_35871_, _35831_, _02803_);
  or (_35873_, _35871_, _35870_);
  and (_35874_, _35873_, _03887_);
  and (_35875_, _11921_, _04656_);
  nor (_35876_, _35875_, _35826_);
  nor (_35877_, _35876_, _03887_);
  or (_35878_, _35877_, _35874_);
  and (_35879_, _35878_, _03128_);
  and (_35880_, _11927_, _04656_);
  nor (_35881_, _35880_, _35826_);
  nor (_35882_, _35881_, _03128_);
  or (_35884_, _35882_, _35879_);
  and (_35885_, _35884_, _03883_);
  nor (_35886_, _35885_, _35833_);
  nor (_35887_, _35886_, _03135_);
  nor (_35888_, _35843_, _03137_);
  and (_35889_, _35888_, _35829_);
  or (_35890_, _35889_, _35887_);
  and (_35891_, _35890_, _05783_);
  nor (_35892_, _11919_, _11233_);
  nor (_35893_, _35892_, _35826_);
  nor (_35895_, _35893_, _05783_);
  or (_35896_, _35895_, _35891_);
  and (_35897_, _35896_, _05788_);
  nor (_35898_, _11926_, _11233_);
  nor (_35899_, _35898_, _35826_);
  nor (_35900_, _35899_, _05788_);
  or (_35901_, _35900_, _03163_);
  nor (_35902_, _35901_, _35897_);
  and (_35903_, _35838_, _03163_);
  or (_35904_, _35903_, _02888_);
  nor (_35906_, _35904_, _35902_);
  and (_35907_, _11985_, _04656_);
  nor (_35908_, _35907_, _35826_);
  nor (_35909_, _35908_, _02890_);
  or (_35910_, _35909_, _35906_);
  or (_35911_, _35910_, _42672_);
  or (_35912_, _42668_, \oc8051_golden_model_1.TL1 [2]);
  and (_35913_, _35912_, _43998_);
  and (_43586_, _35913_, _35911_);
  not (_35914_, \oc8051_golden_model_1.TL1 [3]);
  nor (_35916_, _04656_, _35914_);
  and (_35917_, _12133_, _04656_);
  nor (_35918_, _35917_, _35916_);
  nor (_35919_, _35918_, _03128_);
  and (_35920_, _04656_, _04241_);
  nor (_35921_, _35920_, _35916_);
  and (_35922_, _35921_, _06770_);
  and (_35923_, _04656_, \oc8051_golden_model_1.ACC [3]);
  nor (_35924_, _35923_, _35916_);
  nor (_35925_, _35924_, _03084_);
  nor (_35927_, _35924_, _03814_);
  nor (_35928_, _03813_, _35914_);
  or (_35929_, _35928_, _35927_);
  and (_35930_, _35929_, _03810_);
  nor (_35931_, _12017_, _11233_);
  nor (_35932_, _35931_, _35916_);
  nor (_35933_, _35932_, _03810_);
  or (_35934_, _35933_, _35930_);
  and (_35935_, _35934_, _03336_);
  nor (_35936_, _35921_, _03336_);
  nor (_35938_, _35936_, _35935_);
  nor (_35939_, _35938_, _03075_);
  or (_35940_, _35939_, _06770_);
  nor (_35941_, _35940_, _35925_);
  or (_35942_, _35941_, _02853_);
  nor (_35943_, _35942_, _35922_);
  and (_35944_, _04656_, _06154_);
  nor (_35945_, _35944_, _35916_);
  nor (_35946_, _35945_, _05540_);
  nor (_35947_, _35946_, _02579_);
  not (_35949_, _35947_);
  nor (_35950_, _35949_, _35943_);
  nor (_35951_, _12112_, _11233_);
  or (_35952_, _35916_, _02838_);
  nor (_35953_, _35952_, _35951_);
  or (_35954_, _35953_, _02802_);
  nor (_35955_, _35954_, _35950_);
  and (_35956_, _04656_, _05658_);
  nor (_35957_, _35956_, _35916_);
  nor (_35958_, _35957_, _02803_);
  or (_35960_, _35958_, _35955_);
  and (_35961_, _35960_, _03887_);
  and (_35962_, _12127_, _04656_);
  nor (_35963_, _35962_, _35916_);
  nor (_35964_, _35963_, _03887_);
  or (_35965_, _35964_, _35961_);
  and (_35966_, _35965_, _03128_);
  nor (_35967_, _35966_, _35919_);
  nor (_35968_, _35967_, _02970_);
  nor (_35969_, _35916_, _05079_);
  not (_35971_, _35969_);
  nor (_35972_, _35957_, _03883_);
  and (_35973_, _35972_, _35971_);
  nor (_35974_, _35973_, _35968_);
  nor (_35975_, _35974_, _03135_);
  nor (_35976_, _35924_, _03137_);
  and (_35977_, _35976_, _35971_);
  or (_35978_, _35977_, _35975_);
  and (_35979_, _35978_, _05783_);
  nor (_35980_, _12125_, _11233_);
  nor (_35982_, _35980_, _35916_);
  nor (_35983_, _35982_, _05783_);
  or (_35984_, _35983_, _35979_);
  and (_35985_, _35984_, _05788_);
  nor (_35986_, _12132_, _11233_);
  nor (_35987_, _35986_, _35916_);
  nor (_35988_, _35987_, _05788_);
  or (_35989_, _35988_, _03163_);
  nor (_35990_, _35989_, _35985_);
  and (_35991_, _35932_, _03163_);
  or (_35993_, _35991_, _02888_);
  nor (_35994_, _35993_, _35990_);
  and (_35995_, _12183_, _04656_);
  nor (_35996_, _35995_, _35916_);
  nor (_35997_, _35996_, _02890_);
  or (_35998_, _35997_, _35994_);
  or (_35999_, _35998_, _42672_);
  or (_36000_, _42668_, \oc8051_golden_model_1.TL1 [3]);
  and (_36001_, _36000_, _43998_);
  and (_43587_, _36001_, _35999_);
  not (_36003_, \oc8051_golden_model_1.TL1 [4]);
  nor (_36004_, _04656_, _36003_);
  nor (_36005_, _36004_, _05031_);
  not (_36006_, _36005_);
  and (_36007_, _05666_, _04656_);
  nor (_36008_, _36007_, _36004_);
  nor (_36009_, _36008_, _03883_);
  and (_36010_, _36009_, _36006_);
  and (_36011_, _12207_, _04656_);
  nor (_36012_, _36011_, _36004_);
  nor (_36014_, _36012_, _03128_);
  and (_36015_, _04656_, \oc8051_golden_model_1.ACC [4]);
  nor (_36016_, _36015_, _36004_);
  nor (_36017_, _36016_, _03084_);
  nor (_36018_, _36016_, _03814_);
  nor (_36019_, _03813_, _36003_);
  or (_36020_, _36019_, _36018_);
  and (_36021_, _36020_, _03810_);
  nor (_36022_, _12217_, _11233_);
  nor (_36023_, _36022_, _36004_);
  nor (_36025_, _36023_, _03810_);
  or (_36026_, _36025_, _36021_);
  and (_36027_, _36026_, _03336_);
  and (_36028_, _04656_, _04982_);
  nor (_36029_, _36028_, _36004_);
  nor (_36030_, _36029_, _03336_);
  nor (_36031_, _36030_, _36027_);
  nor (_36032_, _36031_, _03075_);
  or (_36033_, _36032_, _06770_);
  nor (_36034_, _36033_, _36017_);
  and (_36036_, _36029_, _06770_);
  nor (_36037_, _36036_, _36034_);
  nor (_36038_, _36037_, _02853_);
  and (_36039_, _04656_, _06159_);
  nor (_36040_, _36004_, _05540_);
  not (_36041_, _36040_);
  nor (_36042_, _36041_, _36039_);
  or (_36043_, _36042_, _02579_);
  nor (_36044_, _36043_, _36038_);
  nor (_36045_, _12321_, _11233_);
  nor (_36047_, _36045_, _36004_);
  nor (_36048_, _36047_, _02838_);
  or (_36049_, _36048_, _02802_);
  or (_36050_, _36049_, _36044_);
  nand (_36051_, _36008_, _02802_);
  and (_36052_, _36051_, _36050_);
  and (_36053_, _36052_, _03887_);
  and (_36054_, _12211_, _04656_);
  nor (_36055_, _36054_, _36004_);
  nor (_36056_, _36055_, _03887_);
  or (_36058_, _36056_, _36053_);
  and (_36059_, _36058_, _03128_);
  nor (_36060_, _36059_, _36014_);
  nor (_36061_, _36060_, _02970_);
  nor (_36062_, _36061_, _36010_);
  nor (_36063_, _36062_, _03135_);
  nor (_36064_, _36016_, _03137_);
  and (_36065_, _36064_, _36006_);
  nor (_36066_, _36065_, _02965_);
  not (_36067_, _36066_);
  nor (_36069_, _36067_, _36063_);
  nor (_36070_, _12209_, _11233_);
  or (_36071_, _36004_, _05783_);
  nor (_36072_, _36071_, _36070_);
  or (_36073_, _36072_, _03123_);
  nor (_36074_, _36073_, _36069_);
  nor (_36075_, _12206_, _11233_);
  nor (_36076_, _36075_, _36004_);
  nor (_36077_, _36076_, _05788_);
  or (_36078_, _36077_, _03163_);
  nor (_36080_, _36078_, _36074_);
  and (_36081_, _36023_, _03163_);
  or (_36082_, _36081_, _02888_);
  nor (_36083_, _36082_, _36080_);
  and (_36084_, _12389_, _04656_);
  nor (_36085_, _36084_, _36004_);
  nor (_36086_, _36085_, _02890_);
  or (_36087_, _36086_, _36083_);
  or (_36088_, _36087_, _42672_);
  or (_36089_, _42668_, \oc8051_golden_model_1.TL1 [4]);
  and (_36091_, _36089_, _43998_);
  and (_43588_, _36091_, _36088_);
  not (_36092_, \oc8051_golden_model_1.TL1 [5]);
  nor (_36093_, _04656_, _36092_);
  and (_36094_, _12411_, _04656_);
  nor (_36095_, _36094_, _36093_);
  nor (_36096_, _36095_, _03128_);
  and (_36097_, _04656_, _04877_);
  nor (_36098_, _36097_, _36093_);
  and (_36099_, _36098_, _06770_);
  and (_36101_, _04656_, \oc8051_golden_model_1.ACC [5]);
  nor (_36102_, _36101_, _36093_);
  nor (_36103_, _36102_, _03084_);
  nor (_36104_, _12407_, _11233_);
  nor (_36105_, _36104_, _36093_);
  and (_36106_, _36105_, _02974_);
  or (_36107_, _36102_, _03814_);
  or (_36108_, _03813_, _36092_);
  and (_36109_, _36108_, _03810_);
  and (_36110_, _36109_, _36107_);
  or (_36112_, _36110_, _03069_);
  nor (_36113_, _36112_, _36106_);
  nor (_36114_, _36098_, _03336_);
  nor (_36115_, _36114_, _36113_);
  nor (_36116_, _36115_, _03075_);
  or (_36117_, _36116_, _06770_);
  nor (_36118_, _36117_, _36103_);
  nor (_36119_, _36118_, _36099_);
  nor (_36120_, _36119_, _02853_);
  and (_36121_, _04656_, _06158_);
  nor (_36123_, _36093_, _05540_);
  not (_36124_, _36123_);
  nor (_36125_, _36124_, _36121_);
  or (_36126_, _36125_, _02579_);
  nor (_36127_, _36126_, _36120_);
  nor (_36128_, _12527_, _11233_);
  nor (_36129_, _36128_, _36093_);
  nor (_36130_, _36129_, _02838_);
  or (_36131_, _36130_, _02802_);
  or (_36132_, _36131_, _36127_);
  and (_36134_, _05614_, _04656_);
  nor (_36135_, _36134_, _36093_);
  nand (_36136_, _36135_, _02802_);
  and (_36137_, _36136_, _36132_);
  and (_36138_, _36137_, _03887_);
  and (_36139_, _12415_, _04656_);
  nor (_36140_, _36139_, _36093_);
  nor (_36141_, _36140_, _03887_);
  or (_36142_, _36141_, _36138_);
  and (_36143_, _36142_, _03128_);
  nor (_36145_, _36143_, _36096_);
  nor (_36146_, _36145_, _02970_);
  nor (_36147_, _36093_, _04924_);
  not (_36148_, _36147_);
  nor (_36149_, _36135_, _03883_);
  and (_36150_, _36149_, _36148_);
  nor (_36151_, _36150_, _36146_);
  nor (_36152_, _36151_, _03135_);
  nor (_36153_, _36102_, _03137_);
  and (_36154_, _36153_, _36148_);
  or (_36156_, _36154_, _36152_);
  and (_36157_, _36156_, _05783_);
  nor (_36158_, _12413_, _11233_);
  nor (_36159_, _36158_, _36093_);
  nor (_36160_, _36159_, _05783_);
  or (_36161_, _36160_, _36157_);
  and (_36162_, _36161_, _05788_);
  nor (_36163_, _12410_, _11233_);
  nor (_36164_, _36163_, _36093_);
  nor (_36165_, _36164_, _05788_);
  or (_36167_, _36165_, _03163_);
  nor (_36168_, _36167_, _36162_);
  and (_36169_, _36105_, _03163_);
  or (_36170_, _36169_, _02888_);
  nor (_36171_, _36170_, _36168_);
  and (_36172_, _12589_, _04656_);
  nor (_36173_, _36172_, _36093_);
  nor (_36174_, _36173_, _02890_);
  or (_36175_, _36174_, _36171_);
  or (_36176_, _36175_, _42672_);
  or (_36178_, _42668_, \oc8051_golden_model_1.TL1 [5]);
  and (_36179_, _36178_, _43998_);
  and (_43589_, _36179_, _36176_);
  not (_36180_, \oc8051_golden_model_1.TL1 [6]);
  nor (_36181_, _04656_, _36180_);
  and (_36182_, _04656_, \oc8051_golden_model_1.ACC [6]);
  nor (_36183_, _36182_, _36181_);
  nor (_36184_, _36183_, _03814_);
  nor (_36185_, _03813_, _36180_);
  or (_36186_, _36185_, _36184_);
  and (_36188_, _36186_, _03810_);
  nor (_36189_, _12603_, _11233_);
  nor (_36190_, _36189_, _36181_);
  nor (_36191_, _36190_, _03810_);
  or (_36192_, _36191_, _36188_);
  and (_36193_, _36192_, _03336_);
  and (_36194_, _04656_, _04770_);
  nor (_36195_, _36194_, _36181_);
  nor (_36196_, _36195_, _03336_);
  nor (_36197_, _36196_, _36193_);
  nor (_36199_, _36197_, _03075_);
  nor (_36200_, _36183_, _03084_);
  nor (_36201_, _36200_, _06770_);
  not (_36202_, _36201_);
  nor (_36203_, _36202_, _36199_);
  or (_36204_, _36195_, _02853_);
  and (_36205_, _36204_, _09582_);
  or (_36206_, _36205_, _36203_);
  and (_36207_, _04656_, _05849_);
  nor (_36208_, _36207_, _36181_);
  or (_36210_, _36208_, _05540_);
  and (_36211_, _36210_, _02838_);
  and (_36212_, _36211_, _36206_);
  nor (_36213_, _12722_, _11233_);
  or (_36214_, _36181_, _02838_);
  nor (_36215_, _36214_, _36213_);
  or (_36216_, _36215_, _02802_);
  nor (_36217_, _36216_, _36212_);
  and (_36218_, _12729_, _04656_);
  nor (_36219_, _36218_, _36181_);
  nor (_36221_, _36219_, _02803_);
  or (_36222_, _36221_, _02980_);
  nor (_36223_, _36222_, _36217_);
  and (_36224_, _12739_, _04656_);
  nor (_36225_, _36224_, _36181_);
  and (_36226_, _36225_, _02980_);
  nor (_36227_, _36226_, _36223_);
  and (_36228_, _36227_, _03128_);
  and (_36229_, _12613_, _04656_);
  nor (_36230_, _36229_, _36181_);
  nor (_36232_, _36230_, _03128_);
  or (_36233_, _36232_, _36228_);
  and (_36234_, _36233_, _03883_);
  nor (_36235_, _36181_, _04819_);
  not (_36236_, _36235_);
  nor (_36237_, _36219_, _03883_);
  and (_36238_, _36237_, _36236_);
  nor (_36239_, _36238_, _36234_);
  nor (_36240_, _36239_, _03135_);
  nor (_36241_, _36183_, _03137_);
  and (_36243_, _36241_, _36236_);
  nor (_36244_, _36243_, _02965_);
  not (_36245_, _36244_);
  nor (_36246_, _36245_, _36240_);
  nor (_36247_, _12737_, _11233_);
  or (_36248_, _36181_, _05783_);
  nor (_36249_, _36248_, _36247_);
  or (_36250_, _36249_, _03123_);
  nor (_36251_, _36250_, _36246_);
  nor (_36252_, _12612_, _11233_);
  nor (_36254_, _36252_, _36181_);
  nor (_36255_, _36254_, _05788_);
  or (_36256_, _36255_, _03163_);
  nor (_36257_, _36256_, _36251_);
  and (_36258_, _36190_, _03163_);
  or (_36259_, _36258_, _02888_);
  nor (_36260_, _36259_, _36257_);
  and (_36261_, _12794_, _04656_);
  nor (_36262_, _36261_, _36181_);
  nor (_36263_, _36262_, _02890_);
  or (_36265_, _36263_, _36260_);
  or (_36266_, _36265_, _42672_);
  or (_36267_, _42668_, \oc8051_golden_model_1.TL1 [6]);
  and (_36268_, _36267_, _43998_);
  and (_43590_, _36268_, _36266_);
  not (_36269_, \oc8051_golden_model_1.TMOD [0]);
  nor (_36270_, _04664_, _36269_);
  and (_36271_, _05226_, _04664_);
  nor (_36272_, _36271_, _36270_);
  and (_36273_, _36272_, _16625_);
  and (_36275_, _04664_, _05672_);
  nor (_36276_, _36275_, _36270_);
  or (_36277_, _36276_, _03883_);
  nor (_36278_, _36277_, _36271_);
  and (_36279_, _04664_, \oc8051_golden_model_1.ACC [0]);
  nor (_36280_, _36279_, _36270_);
  nor (_36281_, _36280_, _03084_);
  nor (_36282_, _36281_, _06770_);
  nor (_36283_, _36272_, _03810_);
  nor (_36284_, _03813_, _36269_);
  nor (_36286_, _36280_, _03814_);
  nor (_36287_, _36286_, _36284_);
  nor (_36288_, _36287_, _02974_);
  or (_36289_, _36288_, _03069_);
  nor (_36290_, _36289_, _36283_);
  or (_36291_, _36290_, _03075_);
  and (_36292_, _36291_, _36282_);
  and (_36293_, _04664_, _03808_);
  or (_36294_, _36270_, _30142_);
  nor (_36295_, _36294_, _36293_);
  nor (_36297_, _36295_, _36292_);
  nor (_36298_, _36297_, _02853_);
  and (_36299_, _04664_, _06152_);
  nor (_36300_, _36270_, _05540_);
  not (_36301_, _36300_);
  nor (_36302_, _36301_, _36299_);
  nor (_36303_, _36302_, _36298_);
  and (_36304_, _36303_, _02838_);
  nor (_36305_, _11505_, _11315_);
  nor (_36306_, _36305_, _36270_);
  nor (_36308_, _36306_, _02838_);
  or (_36309_, _36308_, _36304_);
  and (_36310_, _36309_, _02803_);
  nor (_36311_, _36276_, _02803_);
  or (_36312_, _36311_, _36310_);
  and (_36313_, _36312_, _03887_);
  and (_36314_, _11399_, _04664_);
  nor (_36315_, _36314_, _36270_);
  nor (_36316_, _36315_, _03887_);
  or (_36317_, _36316_, _36313_);
  and (_36319_, _36317_, _03128_);
  and (_36320_, _11522_, _04664_);
  nor (_36321_, _36320_, _36270_);
  nor (_36322_, _36321_, _03128_);
  or (_36323_, _36322_, _36319_);
  and (_36324_, _36323_, _03883_);
  nor (_36325_, _36324_, _36278_);
  nor (_36326_, _36325_, _03135_);
  nor (_36327_, _36270_, _09409_);
  or (_36328_, _36327_, _03137_);
  nor (_36330_, _36328_, _36280_);
  or (_36331_, _36330_, _36326_);
  and (_36332_, _36331_, _05783_);
  nor (_36333_, _11396_, _11315_);
  nor (_36334_, _36333_, _36270_);
  nor (_36335_, _36334_, _05783_);
  or (_36336_, _36335_, _36332_);
  and (_36337_, _36336_, _05788_);
  nor (_36338_, _11520_, _11315_);
  nor (_36339_, _36338_, _36270_);
  nor (_36341_, _36339_, _05788_);
  nor (_36342_, _36341_, _16625_);
  not (_36343_, _36342_);
  nor (_36344_, _36343_, _36337_);
  nor (_36345_, _36344_, _36273_);
  or (_36346_, _36345_, _42672_);
  or (_36347_, _42668_, \oc8051_golden_model_1.TMOD [0]);
  and (_36348_, _36347_, _43998_);
  and (_43592_, _36348_, _36346_);
  nor (_36349_, _04664_, \oc8051_golden_model_1.TMOD [1]);
  not (_36351_, _36349_);
  and (_36352_, _11695_, _04664_);
  nor (_36353_, _36352_, _02838_);
  and (_36354_, _36353_, _36351_);
  and (_36355_, _04664_, _02551_);
  nor (_36356_, _36355_, _36349_);
  and (_36357_, _36356_, _03075_);
  nor (_36358_, _11315_, _04000_);
  or (_36359_, _36358_, _36349_);
  nor (_36360_, _36359_, _03336_);
  and (_36362_, _36356_, _03813_);
  not (_36363_, \oc8051_golden_model_1.TMOD [1]);
  nor (_36364_, _03813_, _36363_);
  or (_36365_, _36364_, _36362_);
  and (_36366_, _36365_, _03810_);
  and (_36367_, _11606_, _04664_);
  nor (_36368_, _36367_, _36349_);
  and (_36369_, _36368_, _02974_);
  or (_36370_, _36369_, _36366_);
  and (_36371_, _36370_, _03336_);
  nor (_36373_, _36371_, _36360_);
  nor (_36374_, _36373_, _03075_);
  or (_36375_, _36374_, _06770_);
  nor (_36376_, _36375_, _36357_);
  and (_36377_, _36359_, _06770_);
  or (_36378_, _36377_, _02853_);
  nor (_36379_, _36378_, _36376_);
  or (_36380_, _11315_, _06151_);
  nor (_36381_, _36349_, _05540_);
  and (_36382_, _36381_, _36380_);
  or (_36384_, _36382_, _36379_);
  and (_36385_, _36384_, _02838_);
  nor (_36386_, _36385_, _36354_);
  nor (_36387_, _36386_, _02802_);
  and (_36388_, _04664_, _03698_);
  not (_36389_, _36388_);
  nor (_36390_, _36349_, _02803_);
  and (_36391_, _36390_, _36389_);
  nor (_36392_, _36391_, _36387_);
  nor (_36393_, _36392_, _02980_);
  nor (_36395_, _11710_, _11315_);
  nor (_36396_, _36395_, _03887_);
  and (_36397_, _36396_, _36351_);
  nor (_36398_, _36397_, _36393_);
  nor (_36399_, _36398_, _03127_);
  nor (_36400_, _11715_, _11315_);
  nor (_36401_, _36400_, _03128_);
  and (_36402_, _36401_, _36351_);
  nor (_36403_, _36402_, _36399_);
  nor (_36404_, _36403_, _02970_);
  nor (_36406_, _11709_, _11315_);
  nor (_36407_, _36406_, _03883_);
  and (_36408_, _36407_, _36351_);
  nor (_36409_, _36408_, _36404_);
  nor (_36410_, _36409_, _03135_);
  nor (_36411_, _04664_, _36363_);
  nor (_36412_, _36411_, _13722_);
  nor (_36413_, _36412_, _03137_);
  and (_36414_, _36413_, _36356_);
  nor (_36415_, _36414_, _36410_);
  or (_36417_, _36415_, _17961_);
  and (_36418_, _11714_, _04664_);
  or (_36419_, _36418_, _05788_);
  or (_36420_, _36419_, _36349_);
  and (_36421_, _36420_, _03906_);
  and (_36422_, _36388_, _05178_);
  or (_36423_, _36349_, _05783_);
  or (_36424_, _36423_, _36422_);
  and (_36425_, _36424_, _36421_);
  and (_36426_, _36425_, _36417_);
  nor (_36428_, _36368_, _03906_);
  nor (_36429_, _36428_, _36426_);
  and (_36430_, _36429_, _02890_);
  nor (_36431_, _36367_, _36411_);
  nor (_36432_, _36431_, _02890_);
  or (_36433_, _36432_, _36430_);
  or (_36434_, _36433_, _42672_);
  or (_36435_, _42668_, \oc8051_golden_model_1.TMOD [1]);
  and (_36436_, _36435_, _43998_);
  and (_43593_, _36436_, _36434_);
  not (_36438_, \oc8051_golden_model_1.TMOD [2]);
  nor (_36439_, _04664_, _36438_);
  nor (_36440_, _36439_, _05130_);
  not (_36441_, _36440_);
  and (_36442_, _04664_, _05701_);
  nor (_36443_, _36442_, _36439_);
  nor (_36444_, _36443_, _03883_);
  and (_36445_, _36444_, _36441_);
  and (_36446_, _04664_, _04435_);
  nor (_36447_, _36446_, _36439_);
  and (_36449_, _36447_, _06770_);
  nor (_36450_, _11801_, _11315_);
  nor (_36451_, _36450_, _36439_);
  nor (_36452_, _36451_, _03810_);
  nor (_36453_, _03813_, _36438_);
  and (_36454_, _04664_, \oc8051_golden_model_1.ACC [2]);
  nor (_36455_, _36454_, _36439_);
  nor (_36456_, _36455_, _03814_);
  nor (_36457_, _36456_, _36453_);
  nor (_36458_, _36457_, _02974_);
  or (_36460_, _36458_, _36452_);
  and (_36461_, _36460_, _03336_);
  nor (_36462_, _36447_, _03336_);
  or (_36463_, _36462_, _36461_);
  and (_36464_, _36463_, _03084_);
  nor (_36465_, _36455_, _03084_);
  nor (_36466_, _36465_, _06770_);
  not (_36467_, _36466_);
  nor (_36468_, _36467_, _36464_);
  nor (_36469_, _36468_, _36449_);
  nor (_36471_, _36469_, _02853_);
  and (_36472_, _04664_, _06155_);
  nor (_36473_, _36439_, _05540_);
  not (_36474_, _36473_);
  nor (_36475_, _36474_, _36472_);
  nor (_36476_, _36475_, _36471_);
  and (_36477_, _36476_, _02838_);
  nor (_36478_, _11906_, _11315_);
  nor (_36479_, _36478_, _36439_);
  nor (_36480_, _36479_, _02838_);
  or (_36482_, _36480_, _36477_);
  and (_36483_, _36482_, _02803_);
  nor (_36484_, _36443_, _02803_);
  or (_36485_, _36484_, _36483_);
  and (_36486_, _36485_, _03887_);
  and (_36487_, _11921_, _04664_);
  nor (_36488_, _36487_, _36439_);
  nor (_36489_, _36488_, _03887_);
  or (_36490_, _36489_, _36486_);
  and (_36491_, _36490_, _03128_);
  and (_36493_, _11927_, _04664_);
  nor (_36494_, _36493_, _36439_);
  nor (_36495_, _36494_, _03128_);
  or (_36496_, _36495_, _36491_);
  and (_36497_, _36496_, _03883_);
  nor (_36498_, _36497_, _36445_);
  nor (_36499_, _36498_, _03135_);
  nor (_36500_, _36455_, _03137_);
  and (_36501_, _36500_, _36441_);
  or (_36502_, _36501_, _36499_);
  and (_36504_, _36502_, _05783_);
  nor (_36505_, _11919_, _11315_);
  nor (_36506_, _36505_, _36439_);
  nor (_36507_, _36506_, _05783_);
  or (_36508_, _36507_, _36504_);
  and (_36509_, _36508_, _05788_);
  nor (_36510_, _11926_, _11315_);
  nor (_36511_, _36510_, _36439_);
  nor (_36512_, _36511_, _05788_);
  or (_36513_, _36512_, _03163_);
  nor (_36515_, _36513_, _36509_);
  and (_36516_, _36451_, _03163_);
  or (_36517_, _36516_, _02888_);
  nor (_36518_, _36517_, _36515_);
  and (_36519_, _11985_, _04664_);
  nor (_36520_, _36519_, _36439_);
  nor (_36521_, _36520_, _02890_);
  or (_36522_, _36521_, _36518_);
  or (_36523_, _36522_, _42672_);
  or (_36524_, _42668_, \oc8051_golden_model_1.TMOD [2]);
  and (_36526_, _36524_, _43998_);
  and (_43594_, _36526_, _36523_);
  not (_36527_, \oc8051_golden_model_1.TMOD [3]);
  nor (_36528_, _04664_, _36527_);
  nor (_36529_, _36528_, _05079_);
  not (_36530_, _36529_);
  and (_36531_, _04664_, _05658_);
  nor (_36532_, _36531_, _36528_);
  nor (_36533_, _36532_, _03883_);
  and (_36534_, _36533_, _36530_);
  and (_36536_, _12133_, _04664_);
  nor (_36537_, _36536_, _36528_);
  nor (_36538_, _36537_, _03128_);
  and (_36539_, _04664_, \oc8051_golden_model_1.ACC [3]);
  nor (_36540_, _36539_, _36528_);
  nor (_36541_, _36540_, _03084_);
  nor (_36542_, _36540_, _03814_);
  nor (_36543_, _03813_, _36527_);
  or (_36544_, _36543_, _36542_);
  and (_36545_, _36544_, _03810_);
  nor (_36547_, _12017_, _11315_);
  nor (_36548_, _36547_, _36528_);
  nor (_36549_, _36548_, _03810_);
  or (_36550_, _36549_, _36545_);
  and (_36551_, _36550_, _03336_);
  and (_36552_, _04664_, _04241_);
  nor (_36553_, _36552_, _36528_);
  nor (_36554_, _36553_, _03336_);
  nor (_36555_, _36554_, _36551_);
  nor (_36556_, _36555_, _03075_);
  or (_36558_, _36556_, _06770_);
  nor (_36559_, _36558_, _36541_);
  and (_36560_, _36553_, _06770_);
  or (_36561_, _36560_, _02853_);
  nor (_36562_, _36561_, _36559_);
  and (_36563_, _04664_, _06154_);
  or (_36564_, _36563_, _36528_);
  and (_36565_, _36564_, _02853_);
  or (_36566_, _36565_, _02579_);
  or (_36567_, _36566_, _36562_);
  nor (_36569_, _12112_, _11315_);
  or (_36570_, _36528_, _02838_);
  or (_36571_, _36570_, _36569_);
  and (_36572_, _36571_, _02803_);
  and (_36573_, _36572_, _36567_);
  nor (_36574_, _36532_, _02803_);
  or (_36575_, _36574_, _36573_);
  and (_36576_, _36575_, _03887_);
  and (_36577_, _12127_, _04664_);
  nor (_36578_, _36577_, _36528_);
  nor (_36580_, _36578_, _03887_);
  or (_36581_, _36580_, _36576_);
  and (_36582_, _36581_, _03128_);
  nor (_36583_, _36582_, _36538_);
  nor (_36584_, _36583_, _02970_);
  nor (_36585_, _36584_, _36534_);
  nor (_36586_, _36585_, _03135_);
  nor (_36587_, _36540_, _03137_);
  and (_36588_, _36587_, _36530_);
  or (_36589_, _36588_, _36586_);
  and (_36591_, _36589_, _05783_);
  nor (_36592_, _12125_, _11315_);
  nor (_36593_, _36592_, _36528_);
  nor (_36594_, _36593_, _05783_);
  or (_36595_, _36594_, _36591_);
  and (_36596_, _36595_, _05788_);
  nor (_36597_, _12132_, _11315_);
  nor (_36598_, _36597_, _36528_);
  nor (_36599_, _36598_, _05788_);
  or (_36600_, _36599_, _03163_);
  nor (_36602_, _36600_, _36596_);
  and (_36603_, _36548_, _03163_);
  or (_36604_, _36603_, _02888_);
  nor (_36605_, _36604_, _36602_);
  and (_36606_, _12183_, _04664_);
  nor (_36607_, _36606_, _36528_);
  nor (_36608_, _36607_, _02890_);
  or (_36609_, _36608_, _36605_);
  or (_36610_, _36609_, _42672_);
  or (_36611_, _42668_, \oc8051_golden_model_1.TMOD [3]);
  and (_36613_, _36611_, _43998_);
  and (_43595_, _36613_, _36610_);
  not (_36614_, \oc8051_golden_model_1.TMOD [4]);
  nor (_36615_, _04664_, _36614_);
  nor (_36616_, _36615_, _05031_);
  not (_36617_, _36616_);
  and (_36618_, _05666_, _04664_);
  nor (_36619_, _36618_, _36615_);
  nor (_36620_, _36619_, _03883_);
  and (_36621_, _36620_, _36617_);
  and (_36623_, _04664_, _06159_);
  nor (_36624_, _36623_, _36615_);
  nor (_36625_, _36624_, _05540_);
  and (_36626_, _04664_, \oc8051_golden_model_1.ACC [4]);
  nor (_36627_, _36626_, _36615_);
  nor (_36628_, _36627_, _03814_);
  nor (_36629_, _03813_, _36614_);
  or (_36630_, _36629_, _36628_);
  and (_36631_, _36630_, _03810_);
  nor (_36632_, _12217_, _11315_);
  nor (_36634_, _36632_, _36615_);
  nor (_36635_, _36634_, _03810_);
  or (_36636_, _36635_, _36631_);
  and (_36637_, _36636_, _03336_);
  and (_36638_, _04664_, _04982_);
  nor (_36639_, _36638_, _36615_);
  nor (_36640_, _36639_, _03336_);
  nor (_36641_, _36640_, _36637_);
  nor (_36642_, _36641_, _03075_);
  nor (_36643_, _36627_, _03084_);
  nor (_36645_, _36643_, _06770_);
  not (_36646_, _36645_);
  nor (_36647_, _36646_, _36642_);
  nor (_36648_, _36639_, _02853_);
  nor (_36649_, _36648_, _02857_);
  nor (_36650_, _36649_, _36647_);
  or (_36651_, _36650_, _36625_);
  and (_36652_, _36651_, _02838_);
  nor (_36653_, _12321_, _11315_);
  nor (_36654_, _36653_, _36615_);
  nor (_36656_, _36654_, _02838_);
  or (_36657_, _36656_, _36652_);
  and (_36658_, _36657_, _02803_);
  nor (_36659_, _36619_, _02803_);
  or (_36660_, _36659_, _36658_);
  and (_36661_, _36660_, _03887_);
  and (_36662_, _12211_, _04664_);
  nor (_36663_, _36662_, _36615_);
  nor (_36664_, _36663_, _03887_);
  or (_36665_, _36664_, _36661_);
  and (_36667_, _36665_, _03128_);
  and (_36668_, _12207_, _04664_);
  nor (_36669_, _36668_, _36615_);
  nor (_36670_, _36669_, _03128_);
  or (_36671_, _36670_, _36667_);
  and (_36672_, _36671_, _03883_);
  nor (_36673_, _36672_, _36621_);
  nor (_36674_, _36673_, _03135_);
  nor (_36675_, _36627_, _03137_);
  and (_36676_, _36675_, _36617_);
  or (_36678_, _36676_, _36674_);
  and (_36679_, _36678_, _05783_);
  nor (_36680_, _12209_, _11315_);
  nor (_36681_, _36680_, _36615_);
  nor (_36682_, _36681_, _05783_);
  or (_36683_, _36682_, _36679_);
  and (_36684_, _36683_, _05788_);
  nor (_36685_, _12206_, _11315_);
  nor (_36686_, _36685_, _36615_);
  nor (_36687_, _36686_, _05788_);
  or (_36689_, _36687_, _03163_);
  nor (_36690_, _36689_, _36684_);
  and (_36691_, _36634_, _03163_);
  or (_36692_, _36691_, _02888_);
  nor (_36693_, _36692_, _36690_);
  and (_36694_, _12389_, _04664_);
  nor (_36695_, _36694_, _36615_);
  nor (_36696_, _36695_, _02890_);
  or (_36697_, _36696_, _36693_);
  or (_36698_, _36697_, _42672_);
  or (_36700_, _42668_, \oc8051_golden_model_1.TMOD [4]);
  and (_36701_, _36700_, _43998_);
  and (_43596_, _36701_, _36698_);
  not (_36702_, \oc8051_golden_model_1.TMOD [5]);
  nor (_36703_, _04664_, _36702_);
  and (_36704_, _12411_, _04664_);
  nor (_36705_, _36704_, _36703_);
  nor (_36706_, _36705_, _03128_);
  and (_36707_, _04664_, _04877_);
  nor (_36708_, _36707_, _36703_);
  and (_36710_, _36708_, _06770_);
  and (_36711_, _04664_, \oc8051_golden_model_1.ACC [5]);
  nor (_36712_, _36711_, _36703_);
  nor (_36713_, _36712_, _03084_);
  nor (_36714_, _12407_, _11315_);
  nor (_36715_, _36714_, _36703_);
  and (_36716_, _36715_, _02974_);
  or (_36717_, _36712_, _03814_);
  or (_36718_, _03813_, _36702_);
  and (_36719_, _36718_, _03810_);
  and (_36721_, _36719_, _36717_);
  or (_36722_, _36721_, _03069_);
  nor (_36723_, _36722_, _36716_);
  nor (_36724_, _36708_, _03336_);
  nor (_36725_, _36724_, _36723_);
  nor (_36726_, _36725_, _03075_);
  or (_36727_, _36726_, _06770_);
  nor (_36728_, _36727_, _36713_);
  or (_36729_, _36728_, _02853_);
  or (_36730_, _36729_, _36710_);
  and (_36732_, _04664_, _06158_);
  nor (_36733_, _36732_, _36703_);
  or (_36734_, _36733_, _05540_);
  and (_36735_, _36734_, _02838_);
  and (_36736_, _36735_, _36730_);
  nor (_36737_, _12527_, _11315_);
  or (_36738_, _36703_, _02838_);
  nor (_36739_, _36738_, _36737_);
  or (_36740_, _36739_, _02802_);
  nor (_36741_, _36740_, _36736_);
  and (_36743_, _05614_, _04664_);
  nor (_36744_, _36743_, _36703_);
  nor (_36745_, _36744_, _02803_);
  or (_36746_, _36745_, _36741_);
  and (_36747_, _36746_, _03887_);
  and (_36748_, _12415_, _04664_);
  nor (_36749_, _36748_, _36703_);
  nor (_36750_, _36749_, _03887_);
  or (_36751_, _36750_, _36747_);
  and (_36752_, _36751_, _03128_);
  nor (_36754_, _36752_, _36706_);
  nor (_36755_, _36754_, _02970_);
  nor (_36756_, _36703_, _04924_);
  not (_36757_, _36756_);
  nor (_36758_, _36744_, _03883_);
  and (_36759_, _36758_, _36757_);
  nor (_36760_, _36759_, _36755_);
  nor (_36761_, _36760_, _03135_);
  nor (_36762_, _36712_, _03137_);
  and (_36763_, _36762_, _36757_);
  or (_36765_, _36763_, _36761_);
  and (_36766_, _36765_, _05783_);
  nor (_36767_, _12413_, _11315_);
  nor (_36768_, _36767_, _36703_);
  nor (_36769_, _36768_, _05783_);
  or (_36770_, _36769_, _36766_);
  and (_36771_, _36770_, _05788_);
  nor (_36772_, _12410_, _11315_);
  nor (_36773_, _36772_, _36703_);
  nor (_36774_, _36773_, _05788_);
  or (_36776_, _36774_, _03163_);
  nor (_36777_, _36776_, _36771_);
  and (_36778_, _36715_, _03163_);
  or (_36779_, _36778_, _02888_);
  nor (_36780_, _36779_, _36777_);
  and (_36781_, _12589_, _04664_);
  nor (_36782_, _36781_, _36703_);
  nor (_36783_, _36782_, _02890_);
  or (_36784_, _36783_, _36780_);
  or (_36785_, _36784_, _42672_);
  or (_36787_, _42668_, \oc8051_golden_model_1.TMOD [5]);
  and (_36788_, _36787_, _43998_);
  and (_43597_, _36788_, _36785_);
  not (_36789_, \oc8051_golden_model_1.TMOD [6]);
  nor (_36790_, _04664_, _36789_);
  and (_36791_, _12613_, _04664_);
  nor (_36792_, _36791_, _36790_);
  nor (_36793_, _36792_, _03128_);
  and (_36794_, _04664_, _04770_);
  nor (_36795_, _36794_, _36790_);
  and (_36797_, _36795_, _06770_);
  and (_36798_, _04664_, \oc8051_golden_model_1.ACC [6]);
  nor (_36799_, _36798_, _36790_);
  nor (_36800_, _36799_, _03814_);
  nor (_36801_, _03813_, _36789_);
  or (_36802_, _36801_, _36800_);
  and (_36803_, _36802_, _03810_);
  nor (_36804_, _12603_, _11315_);
  nor (_36805_, _36804_, _36790_);
  nor (_36806_, _36805_, _03810_);
  or (_36808_, _36806_, _36803_);
  and (_36809_, _36808_, _03336_);
  nor (_36810_, _36795_, _03336_);
  nor (_36811_, _36810_, _36809_);
  nor (_36812_, _36811_, _03075_);
  nor (_36813_, _36799_, _03084_);
  nor (_36814_, _36813_, _06770_);
  not (_36815_, _36814_);
  nor (_36816_, _36815_, _36812_);
  nor (_36817_, _36816_, _36797_);
  nor (_36819_, _36817_, _02853_);
  and (_36820_, _04664_, _05849_);
  nor (_36821_, _36790_, _05540_);
  not (_36822_, _36821_);
  nor (_36823_, _36822_, _36820_);
  or (_36824_, _36823_, _02579_);
  nor (_36825_, _36824_, _36819_);
  nor (_36826_, _12722_, _11315_);
  nor (_36827_, _36826_, _36790_);
  nor (_36828_, _36827_, _02838_);
  or (_36830_, _36828_, _02802_);
  or (_36831_, _36830_, _36825_);
  and (_36832_, _12729_, _04664_);
  nor (_36833_, _36832_, _36790_);
  nand (_36834_, _36833_, _02802_);
  and (_36835_, _36834_, _36831_);
  and (_36836_, _36835_, _03887_);
  and (_36837_, _12739_, _04664_);
  nor (_36838_, _36837_, _36790_);
  nor (_36839_, _36838_, _03887_);
  or (_36841_, _36839_, _36836_);
  and (_36842_, _36841_, _03128_);
  nor (_36843_, _36842_, _36793_);
  nor (_36844_, _36843_, _02970_);
  nor (_36845_, _36790_, _04819_);
  not (_36846_, _36845_);
  nor (_36847_, _36833_, _03883_);
  and (_36848_, _36847_, _36846_);
  nor (_36849_, _36848_, _36844_);
  nor (_36850_, _36849_, _03135_);
  nor (_36852_, _36799_, _03137_);
  and (_36853_, _36852_, _36846_);
  or (_36854_, _36853_, _36850_);
  and (_36855_, _36854_, _05783_);
  nor (_36856_, _12737_, _11315_);
  nor (_36857_, _36856_, _36790_);
  nor (_36858_, _36857_, _05783_);
  or (_36859_, _36858_, _36855_);
  and (_36860_, _36859_, _05788_);
  nor (_36861_, _12612_, _11315_);
  nor (_36863_, _36861_, _36790_);
  nor (_36864_, _36863_, _05788_);
  or (_36865_, _36864_, _03163_);
  nor (_36866_, _36865_, _36860_);
  and (_36867_, _36805_, _03163_);
  or (_36868_, _36867_, _02888_);
  nor (_36869_, _36868_, _36866_);
  and (_36870_, _12794_, _04664_);
  nor (_36871_, _36870_, _36790_);
  nor (_36872_, _36871_, _02890_);
  or (_36874_, _36872_, _36869_);
  or (_36875_, _36874_, _42672_);
  or (_36876_, _42668_, \oc8051_golden_model_1.TMOD [6]);
  and (_36877_, _36876_, _43998_);
  and (_43599_, _36877_, _36875_);
  and (_36878_, _42672_, \oc8051_golden_model_1.P0INREG [0]);
  or (_36879_, _36878_, _00628_);
  and (_43600_, _36879_, _43998_);
  and (_36880_, _42672_, \oc8051_golden_model_1.P0INREG [1]);
  or (_36881_, _36880_, _00643_);
  and (_43601_, _36881_, _43998_);
  and (_36883_, _42672_, \oc8051_golden_model_1.P0INREG [2]);
  or (_36884_, _36883_, _00636_);
  and (_43603_, _36884_, _43998_);
  and (_36885_, _42672_, \oc8051_golden_model_1.P0INREG [3]);
  or (_36886_, _36885_, _00650_);
  and (_43604_, _36886_, _43998_);
  and (_36887_, _42672_, \oc8051_golden_model_1.P0INREG [4]);
  or (_36888_, _36887_, _00663_);
  and (_43605_, _36888_, _43998_);
  and (_36890_, _42672_, \oc8051_golden_model_1.P0INREG [5]);
  or (_36891_, _36890_, _00678_);
  and (_43606_, _36891_, _43998_);
  and (_36892_, _42672_, \oc8051_golden_model_1.P0INREG [6]);
  or (_36893_, _36892_, _00671_);
  and (_43607_, _36893_, _43998_);
  and (_36894_, _42672_, \oc8051_golden_model_1.P1INREG [0]);
  or (_36895_, _36894_, _00595_);
  and (_43608_, _36895_, _43998_);
  and (_36896_, _42672_, \oc8051_golden_model_1.P1INREG [1]);
  or (_36898_, _36896_, _00585_);
  and (_43609_, _36898_, _43998_);
  and (_36899_, _42672_, \oc8051_golden_model_1.P1INREG [2]);
  or (_36900_, _36899_, _00604_);
  and (_43610_, _36900_, _43998_);
  and (_36901_, _42672_, \oc8051_golden_model_1.P1INREG [3]);
  or (_36902_, _36901_, _00614_);
  and (_43611_, _36902_, _43998_);
  and (_36903_, _42672_, \oc8051_golden_model_1.P1INREG [4]);
  or (_36904_, _36903_, _00555_);
  and (_43612_, _36904_, _43998_);
  and (_36906_, _42672_, \oc8051_golden_model_1.P1INREG [5]);
  or (_36907_, _36906_, _00545_);
  and (_43613_, _36907_, _43998_);
  and (_36908_, _42672_, \oc8051_golden_model_1.P1INREG [6]);
  or (_36909_, _36908_, _00565_);
  and (_43614_, _36909_, _43998_);
  and (_36910_, _42672_, \oc8051_golden_model_1.P2INREG [0]);
  or (_36911_, _36910_, _00720_);
  and (_43616_, _36911_, _43998_);
  and (_36913_, _42672_, \oc8051_golden_model_1.P2INREG [1]);
  or (_36914_, _36913_, _00713_);
  and (_43617_, _36914_, _43998_);
  and (_36915_, _42672_, \oc8051_golden_model_1.P2INREG [2]);
  or (_36916_, _36915_, _00698_);
  and (_43618_, _36916_, _43998_);
  and (_36917_, _42672_, \oc8051_golden_model_1.P2INREG [3]);
  or (_36918_, _36917_, _00706_);
  and (_43619_, _36918_, _43998_);
  and (_36919_, _42672_, \oc8051_golden_model_1.P2INREG [4]);
  or (_36921_, _36919_, _00741_);
  and (_43621_, _36921_, _43998_);
  and (_36922_, _42672_, \oc8051_golden_model_1.P2INREG [5]);
  or (_36923_, _36922_, _00748_);
  and (_43622_, _36923_, _43998_);
  and (_36924_, _42672_, \oc8051_golden_model_1.P2INREG [6]);
  or (_36925_, _36924_, _00733_);
  and (_43623_, _36925_, _43998_);
  and (_36926_, _42672_, \oc8051_golden_model_1.P3INREG [0]);
  or (_36927_, _36926_, _00521_);
  and (_43625_, _36927_, _43998_);
  and (_36929_, _42672_, \oc8051_golden_model_1.P3INREG [1]);
  or (_36930_, _36929_, _00493_);
  and (_43626_, _36930_, _43998_);
  and (_36931_, _42672_, \oc8051_golden_model_1.P3INREG [2]);
  or (_36932_, _36931_, _00513_);
  and (_43627_, _36932_, _43998_);
  and (_36933_, _42672_, \oc8051_golden_model_1.P3INREG [3]);
  or (_36934_, _36933_, _00504_);
  and (_43628_, _36934_, _43998_);
  and (_36936_, _42672_, \oc8051_golden_model_1.P3INREG [4]);
  or (_36937_, _36936_, _00466_);
  and (_43629_, _36937_, _43998_);
  and (_36938_, _42672_, \oc8051_golden_model_1.P3INREG [5]);
  or (_36939_, _36938_, _00455_);
  and (_43630_, _36939_, _43998_);
  and (_36940_, _42672_, \oc8051_golden_model_1.P3INREG [6]);
  or (_36941_, _36940_, _00473_);
  and (_43631_, _36941_, _43998_);
  and (_00005_[6], _00474_, _43998_);
  and (_00005_[5], _00456_, _43998_);
  and (_00005_[4], _00467_, _43998_);
  and (_00005_[3], _00505_, _43998_);
  and (_00005_[2], _00514_, _43998_);
  and (_00005_[1], _00494_, _43998_);
  and (_00005_[0], _00522_, _43998_);
  and (_00004_[6], _00734_, _43998_);
  and (_00004_[5], _00749_, _43998_);
  and (_00004_[4], _00742_, _43998_);
  and (_00004_[3], _00707_, _43998_);
  and (_00004_[2], _00699_, _43998_);
  and (_00004_[1], _00714_, _43998_);
  and (_00004_[0], _00721_, _43998_);
  and (_00003_[6], _00566_, _43998_);
  and (_00003_[5], _00546_, _43998_);
  and (_00003_[4], _00557_, _43998_);
  and (_00003_[3], _00615_, _43998_);
  and (_00003_[2], _00606_, _43998_);
  and (_00003_[1], _00586_, _43998_);
  and (_00003_[0], _00596_, _43998_);
  and (_00002_[6], _00672_, _43998_);
  and (_00002_[5], _00679_, _43998_);
  and (_00002_[4], _00664_, _43998_);
  and (_00002_[3], _00651_, _43998_);
  and (_00002_[2], _00637_, _43998_);
  and (_00002_[1], _00644_, _43998_);
  and (_00002_[0], _00629_, _43998_);
  nor (_36945_, _08606_, _08497_);
  nor (_36946_, _10952_, _10697_);
  and (_36947_, _36946_, _36945_);
  not (_36949_, _33688_);
  nand (_36950_, _36949_, _33222_);
  nor (_36951_, _36950_, _33803_);
  nor (_36952_, _31561_, _19452_);
  nor (_36953_, _32139_, _32024_);
  and (_36954_, _36953_, _36952_);
  nor (_36955_, _18652_, _18536_);
  nor (_36956_, _19337_, _18874_);
  and (_36957_, _36956_, _36955_);
  and (_36958_, _36957_, _36954_);
  and (_36960_, _36958_, _36951_);
  or (_36961_, _31910_, _19222_);
  nor (_36962_, _36961_, _33572_);
  nor (_36963_, _36265_, _36175_);
  nor (_36964_, _36874_, _36784_);
  and (_36965_, _36964_, _36963_);
  nor (_36966_, _35033_, _34945_);
  nor (_36967_, _35646_, _35557_);
  and (_36968_, _36967_, _36966_);
  and (_36969_, _36968_, _36965_);
  nor (_36971_, _18305_, _18189_);
  and (_36972_, _36971_, _36969_);
  nor (_36973_, _34677_, _34149_);
  nor (_36974_, _35293_, _34765_);
  and (_36975_, _36974_, _36973_);
  nor (_36976_, _35115_, _34500_);
  nor (_36977_, _36345_, _35733_);
  and (_36978_, _36977_, _36976_);
  or (_36979_, _09594_, _02301_);
  nor (_36980_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_36982_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_36983_, _36982_, _36980_);
  nor (_36984_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_36985_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_36986_, _36985_, _36984_);
  and (_36987_, _36986_, _36983_);
  nor (_36988_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_36989_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_36990_, _36989_, _36988_);
  nor (_36991_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_36993_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_36994_, _36993_, _36991_);
  and (_36995_, _36994_, _36990_);
  and (_36996_, _36995_, _36987_);
  nor (_36997_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_36998_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_36999_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_37000_, _36999_, _36998_);
  and (_37001_, _37000_, _36997_);
  nor (_37002_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37004_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_37005_, _37004_, _37002_);
  nor (_37006_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_37007_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_37008_, _37007_, _37006_);
  and (_37009_, _37008_, _37005_);
  and (_37010_, _37009_, _37001_);
  and (_37011_, _37010_, _36996_);
  nor (_37012_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37013_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_37015_, _37013_, _37012_);
  nor (_37016_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_37017_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_37018_, _37017_, _37016_);
  and (_37019_, _37018_, _37015_);
  nor (_37020_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  nor (_37021_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  and (_37022_, _37021_, _37020_);
  nor (_37023_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_37024_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_37026_, _37024_, _37023_);
  and (_37027_, _37026_, _37022_);
  and (_37028_, _37027_, _37019_);
  nor (_37029_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37030_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_37031_, _37030_, _37029_);
  nor (_37032_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  nor (_37033_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  and (_37034_, _37033_, _37032_);
  and (_37035_, _37034_, _37031_);
  nor (_37037_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_37038_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_37039_, _37038_, _37037_);
  nor (_37040_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_37041_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_37042_, _37041_, _37040_);
  and (_37043_, _37042_, _37039_);
  and (_37044_, _37043_, _37035_);
  and (_37045_, _37044_, _37028_);
  nor (_37046_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_37048_, _37046_, op0_cnst);
  nor (_37049_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_37050_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_37051_, _37050_, _37049_);
  nor (_37052_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_37053_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_37054_, _37053_, _37052_);
  and (_37055_, _37054_, _37051_);
  and (_37056_, _37055_, _37048_);
  nor (_37057_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37059_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_37060_, _37059_, _37057_);
  nor (_37061_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_37062_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_37063_, _37062_, _37061_);
  and (_37064_, _37063_, _37060_);
  and (_37065_, \oc8051_golden_model_1.TCON [1], _33007_);
  nor (_37066_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_37067_, _37066_, _37065_);
  nor (_37068_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_37070_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_37071_, _37070_, _37068_);
  and (_37072_, _37071_, _37067_);
  and (_37073_, _37072_, _37064_);
  and (_37074_, _37073_, _37056_);
  and (_37075_, _37074_, _37045_);
  and (_37076_, _37075_, _37011_);
  nand (_37077_, _37076_, _36979_);
  nor (_37078_, _37077_, _30198_);
  nor (_37079_, _33885_, _30810_);
  and (_37081_, _37079_, _37078_);
  nand (_37082_, _37081_, _36978_);
  nor (_37083_, _37082_, _30463_);
  nor (_37084_, _34061_, _31074_);
  and (_37085_, _37084_, _37083_);
  and (_37086_, _37085_, _36975_);
  or (_37087_, _35998_, _35381_);
  or (_37088_, _37087_, _36609_);
  nor (_37089_, _37088_, _30287_);
  and (_37090_, _37089_, _37086_);
  nor (_37092_, _30986_, _30376_);
  nor (_37093_, _36522_, _35910_);
  nand (_37094_, _37093_, _37092_);
  or (_37095_, _37094_, _30898_);
  or (_37096_, _37095_, _33973_);
  nor (_37097_, _37096_, _17957_);
  and (_37098_, _37097_, _37090_);
  nor (_37099_, _35204_, _34854_);
  nor (_37100_, _35821_, _35469_);
  and (_37101_, _37100_, _37099_);
  nor (_37103_, _31162_, _30551_);
  nor (_37104_, _34589_, _34239_);
  and (_37105_, _37104_, _37103_);
  and (_37106_, _37105_, _37101_);
  and (_37107_, _37106_, _37098_);
  nor (_37108_, _33110_, _31447_);
  nor (_37109_, _34417_, _34329_);
  and (_37110_, _37109_, _37108_);
  nor (_37111_, _30728_, _30639_);
  nor (_37112_, _31341_, _31251_);
  and (_37114_, _37112_, _37111_);
  and (_37115_, _37114_, _37110_);
  and (_37116_, _37115_, _37107_);
  and (_37117_, _37116_, _36972_);
  or (_37118_, _31793_, _19105_);
  or (_37119_, _37118_, _33455_);
  nor (_37120_, _37119_, _18072_);
  and (_37121_, _37120_, _37117_);
  not (_37122_, _18759_);
  nor (_37123_, _18990_, _37122_);
  nor (_37125_, _33339_, _31678_);
  and (_37126_, _37125_, _37123_);
  nor (_37127_, _11196_, _11115_);
  nor (_37128_, _11360_, _11277_);
  and (_37129_, _37128_, _37127_);
  or (_37130_, _36433_, _36087_);
  or (_37131_, _37130_, _36697_);
  nor (_37132_, _37131_, _10506_);
  nor (_37133_, _11034_, _10588_);
  and (_37134_, _37133_, _37132_);
  and (_37136_, _37134_, _37129_);
  nand (_37137_, _37136_, _37126_);
  nor (_37138_, _37137_, _18421_);
  and (_37139_, _37138_, _37121_);
  and (_37140_, _37139_, _36962_);
  and (_37141_, _37140_, _36960_);
  and (_37142_, _37141_, _36947_);
  and (_37143_, _37142_, _42668_);
  and (_37144_, _37143_, _43998_);
  and (_37145_, _32470_, _38470_);
  nor (_37147_, _32869_, _38488_);
  nor (_37148_, _32596_, _38476_);
  nor (_37149_, _32223_, _38401_);
  and (_37150_, _32223_, _38401_);
  or (_37151_, _37150_, _37149_);
  or (_37152_, _37151_, _37148_);
  or (_37153_, _37152_, _37147_);
  nor (_37154_, _32470_, _38470_);
  and (_37155_, _32869_, _38488_);
  or (_37156_, _32348_, _38464_);
  nand (_37158_, _32348_, _38464_);
  and (_37159_, _37158_, _37156_);
  or (_37160_, _37159_, _37155_);
  or (_37161_, _37160_, _37154_);
  or (_37162_, _37161_, _37153_);
  nor (_37163_, _33002_, _38494_);
  and (_37164_, _33002_, _38494_);
  or (_37165_, _37164_, _37163_);
  nor (_37166_, _10844_, _38306_);
  and (_37167_, _32596_, _38476_);
  or (_37169_, _37167_, _37166_);
  and (_37170_, _10844_, _38306_);
  nor (_37171_, _32732_, _38482_);
  and (_37172_, _32732_, _38482_);
  or (_37173_, _37172_, _37171_);
  or (_37174_, _37173_, _37170_);
  or (_37175_, _37174_, _37169_);
  or (_37176_, _37175_, _37165_);
  or (_37177_, _37176_, _37162_);
  or (_37178_, _37177_, _37145_);
  and (_00007_, _37178_, _37144_);
  and (_37180_, _10424_, _38910_);
  nor (_37181_, _10424_, _38910_);
  and (_37182_, _29591_, _38965_);
  nor (_37183_, _29591_, _38965_);
  or (_37184_, _30117_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_37185_, _30117_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_37186_, _37185_, _37184_);
  not (_37187_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_37188_, _29934_, _37187_);
  and (_37190_, _29334_, _38957_);
  nor (_37191_, _29934_, _37187_);
  or (_37192_, _37191_, _37190_);
  or (_37193_, _37192_, _37188_);
  and (_37194_, _29820_, _40152_);
  nor (_37195_, _29820_, _40152_);
  nor (_37196_, _29334_, _38957_);
  nor (_37197_, _29703_, _39001_);
  and (_37198_, _29703_, _39001_);
  or (_37199_, _37198_, _37197_);
  or (_37201_, _37199_, _37196_);
  or (_37202_, _37201_, _37195_);
  or (_37203_, _37202_, _37194_);
  or (_37204_, _37203_, _37193_);
  or (_37205_, _37204_, _37186_);
  or (_37206_, _37205_, _37183_);
  or (_37207_, _37206_, _37182_);
  or (_37208_, _37207_, _37181_);
  or (_37209_, _37208_, _37180_);
  and (_00006_, _37209_, _37144_);
  or (_00001_, _37142_, rst);
  and (_00005_[7], _00481_, _43998_);
  and (_00004_[7], _00756_, _43998_);
  and (_00003_[7], _00574_, _43998_);
  and (_00002_[7], _00686_, _43998_);
  or (_37211_, _03486_, _42560_);
  nand (_37212_, _03486_, _42560_);
  and (_37213_, _37212_, _37211_);
  not (_37214_, _42577_);
  nor (_37215_, _03698_, _37214_);
  and (_37217_, _03698_, _37214_);
  or (_37218_, _37217_, _37215_);
  or (_37219_, _37218_, _37213_);
  or (_37220_, _05613_, _42645_);
  nand (_37221_, _05613_, _42645_);
  and (_37222_, _37221_, _37220_);
  not (_37223_, _42628_);
  nor (_37224_, _05582_, _37223_);
  and (_37225_, _05582_, _37223_);
  or (_37226_, _37225_, _37224_);
  or (_37228_, _37226_, _37222_);
  or (_37229_, _37228_, _37219_);
  or (_37230_, _03297_, _42594_);
  nand (_37231_, _03297_, _42594_);
  and (_37232_, _37231_, _37230_);
  not (_37233_, _42611_);
  nor (_37234_, _03057_, _37233_);
  and (_37235_, _03057_, _37233_);
  or (_37236_, _37235_, _37234_);
  or (_37237_, _37236_, _37232_);
  or (_37239_, _05649_, _42662_);
  nand (_37240_, _05649_, _42662_);
  and (_37241_, _37240_, _37239_);
  nand (_37242_, _05311_, _42543_);
  or (_37243_, _05311_, _42543_);
  and (_37244_, _37243_, _37242_);
  or (_37245_, _37244_, _37241_);
  or (_37246_, _37245_, _37237_);
  or (_37247_, _37246_, _37229_);
  or (_37248_, _02992_, _42925_);
  nor (_37250_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_37251_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_37252_, _37251_, _37250_);
  or (_37253_, _37252_, _02987_);
  or (_37254_, _02462_, _35686_);
  nand (_37255_, _02462_, _35686_);
  and (_37256_, _37255_, _37254_);
  nor (_37257_, _02493_, _33802_);
  and (_37258_, _02493_, _33802_);
  or (_37259_, _37258_, _37257_);
  or (_37261_, _37259_, _37256_);
  or (_37262_, _02503_, _34313_);
  nand (_37263_, _02503_, _34313_);
  and (_37264_, _37263_, _37262_);
  or (_37265_, _02333_, _35052_);
  or (_37266_, _02502_, _43219_);
  and (_37267_, _37266_, _37265_);
  or (_37268_, _37267_, _37264_);
  or (_37269_, _37268_, _37261_);
  and (_37270_, _02429_, _33551_);
  nor (_37272_, _02429_, _33551_);
  or (_37273_, _37272_, _37270_);
  and (_37274_, _02398_, _34041_);
  nor (_37275_, _02398_, _34041_);
  or (_37276_, _37275_, _37274_);
  or (_37277_, _37276_, _37273_);
  nor (_37278_, _02506_, _34563_);
  and (_37279_, _02506_, _34563_);
  or (_37280_, _37279_, _37278_);
  not (_37281_, _02301_);
  and (_37283_, _37281_, _34802_);
  nor (_37284_, _37281_, _34802_);
  or (_37285_, _37284_, _37283_);
  or (_37286_, _37285_, _37280_);
  or (_37287_, _37286_, _37277_);
  or (_37288_, _37287_, _37269_);
  nor (_37289_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_37290_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_37291_, _37290_, _37289_);
  nor (_37292_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_37294_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_37295_, _37294_, _37292_);
  and (_37296_, _37295_, _37291_);
  or (_37297_, \oc8051_golden_model_1.PC [12], _38529_);
  or (_37298_, _26829_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_37299_, _37298_, _37297_);
  or (_37300_, \oc8051_golden_model_1.PC [13], _38504_);
  or (_37301_, _09090_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_37302_, _37301_, _37300_);
  and (_37303_, _37302_, _37299_);
  and (_37305_, _37303_, _37296_);
  and (_37306_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_37307_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_37308_, _37307_, _37306_);
  nor (_37309_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_37310_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_37311_, _37310_, _37309_);
  and (_37312_, _37311_, _37308_);
  and (_37313_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_37314_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_37316_, _37314_, _37313_);
  nor (_37317_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_37318_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_37319_, _37318_, _37317_);
  and (_37320_, _37319_, _37316_);
  and (_37321_, _37320_, _37312_);
  and (_37322_, _37321_, _37305_);
  or (_37323_, \oc8051_golden_model_1.PC [0], _42925_);
  or (_37324_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_37325_, _37324_, _37323_);
  nor (_37327_, _37325_, _37252_);
  or (_37328_, \oc8051_golden_model_1.PC [3], _42909_);
  or (_37329_, _02211_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_37330_, _37329_, _37328_);
  and (_37331_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_37332_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_37333_, _37332_, _37331_);
  and (_37334_, _37333_, _37330_);
  and (_37335_, _37334_, _37327_);
  or (_37336_, \oc8051_golden_model_1.PC [4], _42904_);
  or (_37338_, _24060_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_37339_, _37338_, _37336_);
  nand (_37340_, \oc8051_golden_model_1.PC [5], _42898_);
  or (_37341_, \oc8051_golden_model_1.PC [5], _42898_);
  and (_37342_, _37341_, _37340_);
  and (_37343_, _37342_, _37339_);
  or (_37344_, \oc8051_golden_model_1.PC [6], _42891_);
  or (_37345_, _24791_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_37346_, _37345_, _37344_);
  and (_37347_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_37348_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_37349_, _37348_, _37347_);
  and (_37350_, _37349_, _37346_);
  and (_37351_, _37350_, _37343_);
  and (_37352_, _37351_, _37335_);
  and (_37353_, _37352_, _37322_);
  and (_37354_, _37353_, _42668_);
  and (_37355_, _37354_, _37288_);
  and (_37356_, _37355_, _37253_);
  and (_37357_, _37356_, _37248_);
  and (_37359_, _37357_, _37247_);
  or (_37360_, _03665_, _40093_);
  nand (_37361_, _03665_, _40093_);
  and (_37362_, _37361_, _37360_);
  or (_37363_, _02837_, _39878_);
  nand (_37364_, _02837_, _39878_);
  and (_37365_, _37364_, _37363_);
  or (_37366_, _37365_, _37362_);
  not (_37367_, _40199_);
  nor (_37368_, _02927_, _37367_);
  and (_37370_, _02927_, _37367_);
  or (_37371_, _37370_, _37368_);
  and (_37372_, _02763_, _39938_);
  nor (_37373_, _02763_, _39938_);
  or (_37374_, _37373_, _37372_);
  or (_37375_, _37374_, _37371_);
  or (_37376_, _37375_, _37366_);
  or (_37377_, _02794_, _39972_);
  nand (_37378_, _02794_, _39972_);
  and (_37379_, _37378_, _37377_);
  or (_37381_, _03256_, _40021_);
  nand (_37382_, _03256_, _40021_);
  and (_37383_, _37382_, _37381_);
  or (_37384_, _37383_, _37379_);
  or (_37385_, _03211_, _40057_);
  nand (_37386_, _03211_, _40057_);
  and (_37387_, _37386_, _37385_);
  nand (_37388_, _03629_, _40147_);
  or (_37389_, _03629_, _40147_);
  and (_37390_, _37389_, _37388_);
  or (_37392_, _37390_, _37387_);
  or (_37393_, _37392_, _37384_);
  or (_37394_, _37393_, _37376_);
  and (_37395_, _42814_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_37396_, _37395_, _42962_);
  and (_37397_, _37396_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_37398_, _37397_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_37399_, _37398_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_37400_, _37398_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_37401_, _37400_, _37399_);
  and (_37403_, _25122_, \oc8051_golden_model_1.ACC [7]);
  nor (_37404_, _25122_, \oc8051_golden_model_1.ACC [7]);
  nor (_37405_, _37404_, _37403_);
  and (_37406_, _24767_, \oc8051_golden_model_1.ACC [6]);
  nor (_37407_, _24767_, \oc8051_golden_model_1.ACC [6]);
  nor (_37408_, _37407_, _37406_);
  and (_37409_, _24401_, \oc8051_golden_model_1.ACC [5]);
  nor (_37410_, _24401_, \oc8051_golden_model_1.ACC [5]);
  nor (_37411_, _37410_, _37409_);
  and (_37412_, _24036_, \oc8051_golden_model_1.ACC [4]);
  and (_37414_, _37412_, _37411_);
  nor (_37415_, _37414_, _37409_);
  nor (_37416_, _02569_, _02563_);
  nor (_37417_, _37416_, _02568_);
  not (_37418_, _37417_);
  nor (_37419_, _24036_, \oc8051_golden_model_1.ACC [4]);
  nor (_37420_, _37419_, _37412_);
  and (_37421_, _37420_, _37411_);
  nand (_37422_, _37421_, _37418_);
  nand (_37423_, _37422_, _37415_);
  and (_37425_, _37423_, _37408_);
  or (_37426_, _37425_, _37406_);
  and (_37427_, _37426_, _37405_);
  nor (_37428_, _37427_, _37403_);
  and (_37429_, _25830_, _25487_);
  and (_37430_, _26485_, _26161_);
  and (_37431_, _37430_, _37429_);
  not (_37432_, _37431_);
  nor (_37433_, _37432_, _37428_);
  and (_37434_, _37433_, _26794_);
  nor (_37436_, _37434_, _27111_);
  not (_37437_, _37436_);
  and (_37438_, _37434_, _27111_);
  nor (_37439_, _37438_, _02635_);
  and (_37440_, _37439_, _37437_);
  and (_37441_, _27262_, _02583_);
  not (_37442_, _02582_);
  and (_37443_, _27164_, _02624_);
  and (_37444_, _27173_, _02630_);
  nor (_37445_, _37444_, _37443_);
  and (_37447_, _37445_, _02605_);
  nor (_37448_, _37447_, _37442_);
  not (_37449_, _37448_);
  nor (_37450_, _37449_, _37441_);
  nor (_37451_, _09097_, _02582_);
  nor (_37452_, _37451_, _37450_);
  and (_37453_, _37452_, _02635_);
  nor (_37454_, _37453_, _37440_);
  nor (_37455_, _37454_, _02673_);
  nor (_37456_, _27164_, _02542_);
  or (_37458_, _37456_, _37455_);
  and (_37459_, _37458_, _37401_);
  nor (_37460_, _37458_, _37401_);
  or (_37461_, _37460_, _37459_);
  nor (_37462_, _37400_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_37463_, _37400_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_37464_, _37463_, _37462_);
  not (_37465_, _37464_);
  nor (_37466_, _27558_, _02605_);
  and (_37467_, _27415_, _02630_);
  and (_37469_, _12800_, _02624_);
  nor (_37470_, _37469_, _37467_);
  nor (_37471_, _37470_, _02583_);
  nor (_37472_, _37471_, _37442_);
  not (_37473_, _37472_);
  nor (_37474_, _37473_, _37466_);
  nor (_37475_, _12800_, _02582_);
  or (_37476_, _37475_, _02546_);
  nor (_37477_, _37476_, _37474_);
  and (_37478_, _37438_, _27414_);
  nor (_37480_, _37438_, _27414_);
  nor (_37481_, _37480_, _37478_);
  nor (_37482_, _37481_, _02635_);
  or (_37483_, _37482_, _02673_);
  nor (_37484_, _37483_, _37477_);
  nor (_37485_, _12800_, _02542_);
  or (_37486_, _37485_, _37484_);
  nand (_37487_, _37486_, _37465_);
  or (_37488_, _37486_, _37465_);
  and (_37489_, _37488_, _37487_);
  and (_37491_, _37489_, _37461_);
  and (_37492_, _37491_, _37394_);
  and (property_invalid_rom_pc, _37492_, _37359_);
  and (_37493_, _37142_, inst_finished_r);
  nor (_37494_, _38306_, \oc8051_golden_model_1.SP [7]);
  and (_37495_, _38306_, \oc8051_golden_model_1.SP [7]);
  or (_37496_, _37495_, _37494_);
  nor (_37497_, _38494_, \oc8051_golden_model_1.SP [6]);
  and (_37498_, _38494_, \oc8051_golden_model_1.SP [6]);
  or (_37499_, _37498_, _37497_);
  nor (_37501_, _38488_, \oc8051_golden_model_1.SP [5]);
  and (_37502_, _38488_, \oc8051_golden_model_1.SP [5]);
  or (_37503_, _37502_, _37501_);
  and (_37504_, _38476_, \oc8051_golden_model_1.SP [3]);
  nor (_37505_, _38476_, \oc8051_golden_model_1.SP [3]);
  or (_37506_, _37505_, _37504_);
  nor (_37507_, _38464_, \oc8051_golden_model_1.SP [1]);
  or (_37508_, _38401_, _02866_);
  nand (_37509_, _38401_, _02866_);
  and (_37510_, _37509_, _37508_);
  and (_37512_, _38464_, \oc8051_golden_model_1.SP [1]);
  or (_37513_, _37512_, _37510_);
  or (_37514_, _37513_, _37507_);
  and (_37515_, _38470_, \oc8051_golden_model_1.SP [2]);
  nor (_37516_, _38470_, \oc8051_golden_model_1.SP [2]);
  or (_37517_, _37516_, _37515_);
  or (_37518_, _37517_, _37514_);
  or (_37519_, _37518_, _37506_);
  nor (_37520_, _38482_, \oc8051_golden_model_1.SP [4]);
  and (_37521_, _38482_, \oc8051_golden_model_1.SP [4]);
  or (_37523_, _37521_, _37520_);
  or (_37524_, _37523_, _37519_);
  or (_37525_, _37524_, _37503_);
  or (_37526_, _37525_, _37499_);
  or (_37527_, _37526_, _37496_);
  and (_37528_, _37527_, property_invalid_sp_1_r);
  and (property_invalid_sp, _37528_, _37493_);
  nand (_37529_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_37530_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_37531_, _37530_, _37529_);
  and (_37533_, _29233_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_37534_, \oc8051_golden_model_1.PSW [1], _38957_);
  or (_37535_, _37534_, _37533_);
  or (_37536_, _37535_, _37531_);
  and (_37537_, _29707_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_37538_, \oc8051_golden_model_1.PSW [4], _40152_);
  or (_37539_, _37538_, _37537_);
  and (_37540_, _29595_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_37541_, \oc8051_golden_model_1.PSW [3], _39001_);
  or (_37542_, _37541_, _37540_);
  or (_37544_, _37542_, _37539_);
  or (_37545_, _37544_, _37536_);
  and (_37546_, _07293_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_37547_, \oc8051_golden_model_1.PSW [7], _38910_);
  or (_37548_, _37547_, _37546_);
  and (_37549_, _29824_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_37550_, \oc8051_golden_model_1.PSW [5], _37187_);
  or (_37551_, _37550_, _37549_);
  nand (_37552_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_37553_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_37555_, _37553_, _37552_);
  or (_37556_, _37555_, _37551_);
  or (_37557_, _37556_, _37548_);
  or (_37558_, _37557_, _37545_);
  and (_37559_, _37558_, property_invalid_psw_1_r);
  and (property_invalid_psw, _37559_, _37493_);
  nand (_37560_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_37561_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_37562_, _37561_, _37560_);
  and (_37563_, _22102_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_37565_, \oc8051_golden_model_1.P3 [2], _39739_);
  or (_37566_, _37565_, _37563_);
  or (_37567_, _37566_, _37562_);
  and (_37568_, \oc8051_golden_model_1.P3 [0], _39713_);
  and (_37569_, _21883_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_37570_, _37569_, _37568_);
  and (_37571_, _21989_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_37572_, \oc8051_golden_model_1.P3 [1], _39728_);
  or (_37573_, _37572_, _37571_);
  or (_37574_, _37573_, _37570_);
  or (_37576_, _37574_, _37567_);
  or (_37577_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_37578_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_37579_, _37578_, _37577_);
  or (_37580_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_37581_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_37582_, _37581_, _37580_);
  or (_37583_, _37582_, _37579_);
  and (_37584_, _08933_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_37585_, \oc8051_golden_model_1.P3 [7], _39400_);
  or (_37587_, _37585_, _37584_);
  nand (_37588_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_37589_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_37590_, _37589_, _37588_);
  or (_37591_, _37590_, _37587_);
  or (_37592_, _37591_, _37583_);
  or (_37593_, _37592_, _37576_);
  and (property_invalid_p3, _37593_, _37493_);
  nand (_37594_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_37595_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_37597_, _37595_, _37594_);
  and (_37598_, _21318_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_37599_, \oc8051_golden_model_1.P2 [2], _39640_);
  or (_37600_, _37599_, _37598_);
  or (_37601_, _37600_, _37597_);
  and (_37602_, \oc8051_golden_model_1.P2 [0], _39607_);
  and (_37603_, _21099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_37604_, _37603_, _37602_);
  and (_37605_, _21204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_37606_, \oc8051_golden_model_1.P2 [1], _39620_);
  or (_37608_, _37606_, _37605_);
  or (_37609_, _37608_, _37604_);
  or (_37610_, _37609_, _37601_);
  or (_37611_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_37612_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_37613_, _37612_, _37611_);
  or (_37614_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_37615_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_37616_, _37615_, _37614_);
  or (_37617_, _37616_, _37613_);
  and (_37619_, _08830_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_37620_, \oc8051_golden_model_1.P2 [7], _39392_);
  or (_37621_, _37620_, _37619_);
  nand (_37622_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_37623_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_37624_, _37623_, _37622_);
  or (_37625_, _37624_, _37621_);
  or (_37626_, _37625_, _37617_);
  or (_37627_, _37626_, _37610_);
  and (property_invalid_p2, _37627_, _37493_);
  nand (_37629_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_37630_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_37631_, _37630_, _37629_);
  and (_37632_, _20539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_37633_, \oc8051_golden_model_1.P1 [2], _39541_);
  or (_37634_, _37633_, _37632_);
  or (_37635_, _37634_, _37631_);
  and (_37636_, \oc8051_golden_model_1.P1 [0], _39514_);
  and (_37637_, _20320_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_37638_, _37637_, _37636_);
  and (_37640_, _20426_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_37641_, \oc8051_golden_model_1.P1 [1], _39527_);
  or (_37642_, _37641_, _37640_);
  or (_37643_, _37642_, _37638_);
  or (_37644_, _37643_, _37635_);
  or (_37645_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_37646_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_37647_, _37646_, _37645_);
  or (_37648_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_37649_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_37651_, _37649_, _37648_);
  or (_37652_, _37651_, _37647_);
  and (_37653_, _08727_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_37654_, \oc8051_golden_model_1.P1 [7], _39374_);
  or (_37655_, _37654_, _37653_);
  nand (_37656_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_37657_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_37658_, _37657_, _37656_);
  or (_37659_, _37658_, _37655_);
  or (_37660_, _37659_, _37652_);
  or (_37662_, _37660_, _37644_);
  and (property_invalid_p1, _37662_, _37493_);
  nand (_37663_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_37664_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_37665_, _37664_, _37663_);
  and (_37666_, _19696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_37667_, \oc8051_golden_model_1.P0 [2], _39451_);
  or (_37668_, _37667_, _37666_);
  or (_37669_, _37668_, _37665_);
  and (_37670_, \oc8051_golden_model_1.P0 [0], _39423_);
  and (_37672_, _19456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_37673_, _37672_, _37670_);
  and (_37674_, _19573_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_37675_, \oc8051_golden_model_1.P0 [1], _39435_);
  or (_37676_, _37675_, _37674_);
  or (_37677_, _37676_, _37673_);
  or (_37678_, _37677_, _37669_);
  or (_37679_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_37680_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_37681_, _37680_, _37679_);
  or (_37683_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_37684_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_37685_, _37684_, _37683_);
  or (_37686_, _37685_, _37681_);
  and (_37687_, _08610_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_37688_, \oc8051_golden_model_1.P0 [7], _39360_);
  or (_37689_, _37688_, _37687_);
  nand (_37690_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_37691_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_37692_, _37691_, _37690_);
  or (_37694_, _37692_, _37689_);
  or (_37695_, _37694_, _37686_);
  or (_37696_, _37695_, _37678_);
  and (property_invalid_p0, _37696_, _37493_);
  or (_37697_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_37698_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37699_, _37698_, _37697_);
  nand (_37700_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_37701_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37702_, _37701_, _37700_);
  or (_37704_, _37702_, _37699_);
  and (_37705_, _03353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_37706_, \oc8051_golden_model_1.IRAM[0] [0], _40311_);
  or (_37707_, _37706_, _37705_);
  and (_37708_, _03943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_37709_, \oc8051_golden_model_1.IRAM[0] [1], _40324_);
  or (_37710_, _37709_, _37708_);
  or (_37711_, _37710_, _37707_);
  or (_37712_, _37711_, _37704_);
  or (_37713_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_37715_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37716_, _37715_, _37713_);
  nand (_37717_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_37718_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_37719_, _37718_, _37717_);
  or (_37720_, _37719_, _37716_);
  or (_37721_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_37722_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_37723_, _37722_, _37721_);
  or (_37724_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_37726_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_37727_, _37726_, _37724_);
  or (_37728_, _37727_, _37723_);
  or (_37729_, _37728_, _37720_);
  or (_37730_, _37729_, _37712_);
  or (_37731_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_37732_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_37733_, _37732_, _37731_);
  or (_37734_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_37735_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_37737_, _37735_, _37734_);
  or (_37738_, _37737_, _37733_);
  or (_37739_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_37740_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_37741_, _37740_, _37739_);
  nand (_37742_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_37743_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_37744_, _37743_, _37742_);
  or (_37745_, _37744_, _37741_);
  or (_37746_, _37745_, _37738_);
  and (_37748_, _04927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_37749_, \oc8051_golden_model_1.IRAM[1] [4], _40396_);
  or (_37750_, _37749_, _37748_);
  and (_37751_, \oc8051_golden_model_1.IRAM[1] [5], _40400_);
  and (_37752_, _04822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_37753_, _37752_, _37751_);
  or (_37754_, _37753_, _37750_);
  or (_37755_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_37756_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_37757_, _37756_, _37755_);
  nand (_37759_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_37760_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_37761_, _37760_, _37759_);
  or (_37762_, _37761_, _37757_);
  or (_37763_, _37762_, _37754_);
  or (_37764_, _37763_, _37746_);
  or (_37765_, _37764_, _37730_);
  or (_37766_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_37767_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_37768_, _37767_, _37766_);
  or (_37770_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_37771_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37772_, _37771_, _37770_);
  or (_37773_, _37772_, _37768_);
  and (_37774_, \oc8051_golden_model_1.IRAM[2] [2], _40416_);
  and (_37775_, _04380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_37776_, _37775_, _37774_);
  nand (_37777_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_37778_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_37779_, _37778_, _37777_);
  or (_37781_, _37779_, _37776_);
  or (_37782_, _37781_, _37773_);
  and (_37783_, _04828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_37784_, \oc8051_golden_model_1.IRAM[2] [5], _40424_);
  or (_37785_, _37784_, _37783_);
  and (_37786_, _04933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_37787_, \oc8051_golden_model_1.IRAM[2] [4], _40421_);
  or (_37788_, _37787_, _37786_);
  or (_37789_, _37788_, _37785_);
  and (_37790_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_37792_, \oc8051_golden_model_1.IRAM[2] [7], _40430_);
  or (_37793_, _37792_, _37790_);
  nand (_37794_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_37795_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_37796_, _37795_, _37794_);
  or (_37797_, _37796_, _37793_);
  or (_37798_, _37797_, _37789_);
  or (_37799_, _37798_, _37782_);
  and (_37800_, \oc8051_golden_model_1.IRAM[3] [1], _40437_);
  and (_37801_, _03949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_37803_, _37801_, _37800_);
  and (_37804_, _03755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_37805_, \oc8051_golden_model_1.IRAM[3] [0], _40434_);
  or (_37806_, _37805_, _37804_);
  or (_37807_, _37806_, _37803_);
  and (_37808_, \oc8051_golden_model_1.IRAM[3] [2], _40440_);
  and (_37809_, _04377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_37810_, _37809_, _37808_);
  nand (_37811_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_37812_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_37814_, _37812_, _37811_);
  or (_37815_, _37814_, _37810_);
  or (_37816_, _37815_, _37807_);
  nand (_37817_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_37818_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_37819_, _37818_, _37817_);
  and (_37820_, _04556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_37821_, \oc8051_golden_model_1.IRAM[3] [7], _40227_);
  or (_37822_, _37821_, _37820_);
  or (_37823_, _37822_, _37819_);
  or (_37825_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_37826_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_37827_, _37826_, _37825_);
  or (_37828_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_37829_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_37830_, _37829_, _37828_);
  or (_37831_, _37830_, _37827_);
  or (_37832_, _37831_, _37823_);
  or (_37833_, _37832_, _37816_);
  or (_37834_, _37833_, _37799_);
  or (_37836_, _37834_, _37765_);
  and (_37837_, _03771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37838_, \oc8051_golden_model_1.IRAM[4] [0], _40457_);
  or (_37839_, _37838_, _37837_);
  and (_37840_, \oc8051_golden_model_1.IRAM[4] [1], _40460_);
  and (_37841_, _03963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_37842_, _37841_, _37840_);
  or (_37843_, _37842_, _37839_);
  or (_37844_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_37845_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_37847_, _37845_, _37844_);
  nand (_37848_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_37849_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_37850_, _37849_, _37848_);
  or (_37851_, _37850_, _37847_);
  or (_37852_, _37851_, _37843_);
  or (_37853_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_37854_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_37855_, _37854_, _37853_);
  or (_37856_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_37858_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_37859_, _37858_, _37856_);
  or (_37860_, _37859_, _37855_);
  or (_37861_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_37862_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_37863_, _37862_, _37861_);
  nand (_37864_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_37865_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_37866_, _37865_, _37864_);
  or (_37867_, _37866_, _37863_);
  or (_37869_, _37867_, _37860_);
  or (_37870_, _37869_, _37852_);
  or (_37871_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_37872_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_37873_, _37872_, _37871_);
  nand (_37874_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_37875_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_37876_, _37875_, _37874_);
  or (_37877_, _37876_, _37873_);
  or (_37878_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_37880_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37881_, _37880_, _37878_);
  or (_37882_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_37883_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_37884_, _37883_, _37882_);
  or (_37885_, _37884_, _37881_);
  or (_37886_, _37885_, _37877_);
  or (_37887_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_37888_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_37889_, _37888_, _37887_);
  nand (_37891_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_37892_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_37893_, _37892_, _37891_);
  or (_37894_, _37893_, _37889_);
  and (_37895_, _04948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_37896_, \oc8051_golden_model_1.IRAM[5] [4], _40515_);
  or (_37897_, _37896_, _37895_);
  and (_37898_, _04843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_37899_, \oc8051_golden_model_1.IRAM[5] [5], _40518_);
  or (_37900_, _37899_, _37898_);
  or (_37902_, _37900_, _37897_);
  or (_37903_, _37902_, _37894_);
  or (_37904_, _37903_, _37886_);
  or (_37905_, _37904_, _37870_);
  and (_37906_, \oc8051_golden_model_1.IRAM[6] [2], _40531_);
  and (_37907_, _04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_37908_, _37907_, _37906_);
  nand (_37909_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_37910_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37911_, _37910_, _37909_);
  or (_37913_, _37911_, _37908_);
  or (_37914_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_37915_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37916_, _37915_, _37914_);
  or (_37917_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_37918_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37919_, _37918_, _37917_);
  or (_37920_, _37919_, _37916_);
  or (_37921_, _37920_, _37913_);
  and (_37922_, _04566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_37924_, \oc8051_golden_model_1.IRAM[6] [7], _40552_);
  or (_37925_, _37924_, _37922_);
  nand (_37926_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_37927_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_37928_, _37927_, _37926_);
  or (_37929_, _37928_, _37925_);
  and (_37930_, _04942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_37931_, \oc8051_golden_model_1.IRAM[6] [4], _40536_);
  or (_37932_, _37931_, _37930_);
  and (_37933_, \oc8051_golden_model_1.IRAM[6] [5], _40539_);
  and (_37935_, _04836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_37936_, _37935_, _37933_);
  or (_37937_, _37936_, _37932_);
  or (_37938_, _37937_, _37929_);
  or (_37939_, _37938_, _37921_);
  and (_37940_, _03957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37941_, \oc8051_golden_model_1.IRAM[7] [1], _40575_);
  or (_37942_, _37941_, _37940_);
  and (_37943_, _03765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37944_, \oc8051_golden_model_1.IRAM[7] [0], _40564_);
  or (_37946_, _37944_, _37943_);
  or (_37947_, _37946_, _37942_);
  and (_37948_, _04389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_37949_, \oc8051_golden_model_1.IRAM[7] [2], _40586_);
  or (_37950_, _37949_, _37948_);
  nand (_37951_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_37952_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37953_, _37952_, _37951_);
  or (_37954_, _37953_, _37950_);
  or (_37955_, _37954_, _37947_);
  or (_37957_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_37958_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_37959_, _37958_, _37957_);
  or (_37960_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_37961_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_37962_, _37961_, _37960_);
  or (_37963_, _37962_, _37959_);
  and (_37964_, _04564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_37965_, \oc8051_golden_model_1.IRAM[7] [7], _40239_);
  or (_37966_, _37965_, _37964_);
  nand (_37968_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_37969_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_37970_, _37969_, _37968_);
  or (_37971_, _37970_, _37966_);
  or (_37972_, _37971_, _37963_);
  or (_37973_, _37972_, _37955_);
  or (_37974_, _37973_, _37939_);
  or (_37975_, _37974_, _37905_);
  or (_37976_, _37975_, _37836_);
  and (_37977_, \oc8051_golden_model_1.IRAM[8] [0], _40644_);
  and (_37979_, _03787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_37980_, _37979_, _37977_);
  and (_37981_, _03978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_37982_, \oc8051_golden_model_1.IRAM[8] [1], _40655_);
  or (_37983_, _37982_, _37981_);
  or (_37984_, _37983_, _37980_);
  or (_37985_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nand (_37986_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_37987_, _37986_, _37985_);
  or (_37988_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_37990_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_37991_, _37990_, _37988_);
  or (_37992_, _37991_, _37987_);
  or (_37993_, _37992_, _37984_);
  or (_37994_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand (_37995_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_37996_, _37995_, _37994_);
  or (_37997_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_37998_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_37999_, _37998_, _37997_);
  or (_38001_, _37999_, _37996_);
  or (_38002_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_38003_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_38004_, _38003_, _38002_);
  or (_38005_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nand (_38006_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_38007_, _38006_, _38005_);
  or (_38008_, _38007_, _38004_);
  or (_38009_, _38008_, _38001_);
  or (_38010_, _38009_, _37993_);
  or (_38012_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_38013_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_38014_, _38013_, _38012_);
  or (_38015_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nand (_38016_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_38017_, _38016_, _38015_);
  or (_38018_, _38017_, _38014_);
  or (_38019_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_38020_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_38021_, _38020_, _38019_);
  or (_38023_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_38024_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_38025_, _38024_, _38023_);
  or (_38026_, _38025_, _38021_);
  or (_38027_, _38026_, _38018_);
  or (_38028_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_38029_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_38030_, _38029_, _38028_);
  or (_38031_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nand (_38032_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38034_, _38032_, _38031_);
  or (_38035_, _38034_, _38030_);
  and (_38036_, \oc8051_golden_model_1.IRAM[9] [4], _40728_);
  and (_38037_, _04962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_38038_, _38037_, _38036_);
  and (_38039_, _04857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_38040_, \oc8051_golden_model_1.IRAM[9] [5], _40731_);
  or (_38041_, _38040_, _38039_);
  or (_38042_, _38041_, _38038_);
  or (_38043_, _38042_, _38035_);
  or (_38045_, _38043_, _38027_);
  or (_38046_, _38045_, _38010_);
  and (_38047_, _04409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_38048_, \oc8051_golden_model_1.IRAM[10] [2], _40744_);
  or (_38049_, _38048_, _38047_);
  nand (_38050_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_38051_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_38052_, _38051_, _38050_);
  or (_38053_, _38052_, _38049_);
  or (_38054_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand (_38056_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_38057_, _38056_, _38054_);
  or (_38058_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand (_38059_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_38060_, _38059_, _38058_);
  or (_38061_, _38060_, _38057_);
  or (_38062_, _38061_, _38053_);
  or (_38063_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nand (_38064_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38065_, _38064_, _38063_);
  and (_38067_, _04580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38068_, \oc8051_golden_model_1.IRAM[10] [7], _40253_);
  or (_38069_, _38068_, _38067_);
  or (_38070_, _38069_, _38065_);
  and (_38071_, \oc8051_golden_model_1.IRAM[10] [4], _40750_);
  and (_38072_, _04957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_38073_, _38072_, _38071_);
  and (_38074_, _04852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38075_, \oc8051_golden_model_1.IRAM[10] [5], _40753_);
  or (_38076_, _38075_, _38074_);
  or (_38078_, _38076_, _38073_);
  or (_38079_, _38078_, _38070_);
  or (_38080_, _38079_, _38062_);
  and (_38081_, _03782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_38082_, \oc8051_golden_model_1.IRAM[11] [0], _40761_);
  or (_38083_, _38082_, _38081_);
  and (_38084_, \oc8051_golden_model_1.IRAM[11] [1], _40764_);
  and (_38085_, _03973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_38086_, _38085_, _38084_);
  or (_38087_, _38086_, _38083_);
  and (_38089_, _04407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_38090_, \oc8051_golden_model_1.IRAM[11] [2], _40767_);
  or (_38091_, _38090_, _38089_);
  nand (_38092_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_38093_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_38094_, _38093_, _38092_);
  or (_38095_, _38094_, _38091_);
  or (_38096_, _38095_, _38087_);
  or (_38097_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_38098_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_38100_, _38098_, _38097_);
  or (_38101_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_38102_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_38103_, _38102_, _38101_);
  or (_38104_, _38103_, _38100_);
  and (_38105_, _04578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38106_, \oc8051_golden_model_1.IRAM[11] [7], _40779_);
  or (_38107_, _38106_, _38105_);
  or (_38108_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_38109_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_38111_, _38109_, _38108_);
  or (_38112_, _38111_, _38107_);
  or (_38113_, _38112_, _38104_);
  or (_38114_, _38113_, _38096_);
  or (_38115_, _38114_, _38080_);
  or (_38116_, _38115_, _38046_);
  or (_38117_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_38118_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_38119_, _38118_, _38117_);
  nand (_38120_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_38122_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_38123_, _38122_, _38120_);
  or (_38124_, _38123_, _38119_);
  and (_38125_, \oc8051_golden_model_1.IRAM[12] [0], _40783_);
  and (_38126_, _03799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_38127_, _38126_, _38125_);
  and (_38128_, _03990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_38129_, \oc8051_golden_model_1.IRAM[12] [1], _40786_);
  or (_38130_, _38129_, _38128_);
  or (_38131_, _38130_, _38127_);
  or (_38133_, _38131_, _38124_);
  or (_38134_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_38135_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38136_, _38135_, _38134_);
  nand (_38137_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_38138_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_38139_, _38138_, _38137_);
  or (_38140_, _38139_, _38136_);
  or (_38141_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_38142_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_38144_, _38142_, _38141_);
  or (_38145_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand (_38146_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_38147_, _38146_, _38145_);
  or (_38148_, _38147_, _38144_);
  or (_38149_, _38148_, _38140_);
  or (_38150_, _38149_, _38133_);
  or (_38151_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_38152_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_38153_, _38152_, _38151_);
  or (_38155_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_38156_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_38157_, _38156_, _38155_);
  or (_38158_, _38157_, _38153_);
  or (_38159_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_38160_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_38161_, _38160_, _38159_);
  nand (_38162_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_38163_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_38164_, _38163_, _38162_);
  or (_38166_, _38164_, _38161_);
  or (_38167_, _38166_, _38158_);
  and (_38168_, _04974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_38169_, \oc8051_golden_model_1.IRAM[13] [4], _40814_);
  or (_38170_, _38169_, _38168_);
  and (_38171_, _04869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_38172_, \oc8051_golden_model_1.IRAM[13] [5], _40817_);
  or (_38173_, _38172_, _38171_);
  or (_38174_, _38173_, _38170_);
  or (_38175_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_38177_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_38178_, _38177_, _38175_);
  nand (_38179_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_38180_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38181_, _38180_, _38179_);
  or (_38182_, _38181_, _38178_);
  or (_38183_, _38182_, _38174_);
  or (_38184_, _38183_, _38167_);
  or (_38185_, _38184_, _38150_);
  or (_38186_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand (_38188_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_38189_, _38188_, _38186_);
  or (_38190_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand (_38191_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_38192_, _38191_, _38190_);
  or (_38193_, _38192_, _38189_);
  nand (_38194_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_38195_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_38196_, _38195_, _38194_);
  and (_38197_, _04421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_38199_, \oc8051_golden_model_1.IRAM[14] [2], _40830_);
  or (_38200_, _38199_, _38197_);
  or (_38201_, _38200_, _38196_);
  or (_38202_, _38201_, _38193_);
  and (_38203_, _04969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38204_, \oc8051_golden_model_1.IRAM[14] [4], _40835_);
  or (_38205_, _38204_, _38203_);
  and (_38206_, \oc8051_golden_model_1.IRAM[14] [5], _40838_);
  and (_38207_, _04864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_38208_, _38207_, _38206_);
  or (_38210_, _38208_, _38205_);
  and (_38211_, _04592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38212_, \oc8051_golden_model_1.IRAM[14] [7], _40264_);
  or (_38213_, _38212_, _38211_);
  nand (_38214_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_38215_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38216_, _38215_, _38214_);
  or (_38217_, _38216_, _38213_);
  or (_38218_, _38217_, _38210_);
  or (_38219_, _38218_, _38202_);
  and (_38221_, _04419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_38222_, \oc8051_golden_model_1.IRAM[15] [2], _40852_);
  or (_38223_, _38222_, _38221_);
  nand (_38224_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_38225_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_38226_, _38225_, _38224_);
  or (_38227_, _38226_, _38223_);
  and (_38228_, _03794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_38229_, \oc8051_golden_model_1.IRAM[15] [0], _40846_);
  or (_38230_, _38229_, _38228_);
  and (_38232_, _03985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_38233_, \oc8051_golden_model_1.IRAM[15] [1], _40849_);
  or (_38234_, _38233_, _38232_);
  or (_38235_, _38234_, _38230_);
  or (_38236_, _38235_, _38227_);
  and (_38237_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38238_, \oc8051_golden_model_1.IRAM[15] [7], _40295_);
  or (_38239_, _38238_, _38237_);
  nand (_38240_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_38241_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38243_, _38241_, _38240_);
  or (_38244_, _38243_, _38239_);
  or (_38245_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_38246_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38247_, _38246_, _38245_);
  or (_38248_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_38249_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38250_, _38249_, _38248_);
  or (_38251_, _38250_, _38247_);
  or (_38252_, _38251_, _38244_);
  or (_38254_, _38252_, _38236_);
  or (_38255_, _38254_, _38219_);
  or (_38256_, _38255_, _38185_);
  or (_38257_, _38256_, _38116_);
  or (_38258_, _38257_, _37976_);
  and (property_invalid_iram, _38258_, _37493_);
  nand (_38259_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38260_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_38261_, _38260_, _38259_);
  and (_38262_, _17385_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_38264_, _17385_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38265_, _38264_, _38262_);
  or (_38266_, _38265_, _38261_);
  nor (_38267_, _17199_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38268_, _17199_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38269_, _38268_, _38267_);
  and (_38270_, _17289_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_38271_, _17289_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38272_, _38271_, _38270_);
  or (_38273_, _38272_, _38269_);
  or (_38275_, _38273_, _38266_);
  or (_38276_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_38277_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38278_, _38277_, _38276_);
  or (_38279_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_38280_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38281_, _38280_, _38279_);
  or (_38282_, _38281_, _38278_);
  and (_38283_, _08298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_38284_, _08298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38286_, _38284_, _38283_);
  nand (_38287_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38288_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_38289_, _38288_, _38287_);
  or (_38290_, _38289_, _38286_);
  or (_38291_, _38290_, _38282_);
  or (_38292_, _38291_, _38275_);
  and (property_invalid_dph, _38292_, _37493_);
  nand (_38293_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_38294_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38296_, _38294_, _38293_);
  and (_38297_, _16731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38298_, \oc8051_golden_model_1.DPL [2], _38887_);
  or (_38299_, _38298_, _38297_);
  or (_38300_, _38299_, _38296_);
  and (_38301_, \oc8051_golden_model_1.DPL [0], _38879_);
  and (_38302_, _16543_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_38303_, _38302_, _38301_);
  and (_38304_, _16632_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38305_, \oc8051_golden_model_1.DPL [1], _38883_);
  or (_38307_, _38305_, _38304_);
  or (_38308_, _38307_, _38303_);
  or (_38309_, _38308_, _38300_);
  or (_38310_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_38311_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38312_, _38311_, _38310_);
  or (_38313_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_38314_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38315_, _38314_, _38313_);
  or (_38316_, _38315_, _38312_);
  and (_38317_, _08201_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38318_, \oc8051_golden_model_1.DPL [7], _38599_);
  or (_38319_, _38318_, _38317_);
  nand (_38320_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_38321_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38322_, _38321_, _38320_);
  or (_38323_, _38322_, _38319_);
  or (_38324_, _38323_, _38316_);
  or (_38325_, _38324_, _38309_);
  and (property_invalid_dpl, _38325_, _37493_);
  nand (_38327_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_38328_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_38329_, _38328_, _38327_);
  and (_38330_, _06850_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_38331_, \oc8051_golden_model_1.B [2], _29796_);
  or (_38332_, _38331_, _38330_);
  or (_38333_, _38332_, _38329_);
  and (_38334_, \oc8051_golden_model_1.B [0], _28405_);
  and (_38335_, _06825_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_38336_, _38335_, _38334_);
  and (_38338_, _06796_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38339_, \oc8051_golden_model_1.B [1], _29119_);
  or (_38340_, _38339_, _38338_);
  or (_38341_, _38340_, _38336_);
  or (_38342_, _38341_, _38333_);
  or (_38343_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_38344_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38345_, _38344_, _38343_);
  or (_38346_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_38347_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38349_, _38347_, _38346_);
  or (_38350_, _38349_, _38345_);
  and (_38351_, _06210_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_38352_, \oc8051_golden_model_1.B [7], _27220_);
  or (_38353_, _38352_, _38351_);
  nand (_38354_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_38355_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_38356_, _38355_, _38354_);
  or (_38357_, _38356_, _38353_);
  or (_38358_, _38357_, _38350_);
  or (_38360_, _38358_, _38342_);
  and (property_invalid_b_reg, _38360_, _37493_);
  nand (_38361_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38362_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38363_, _38362_, _38361_);
  and (_38364_, _06964_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38365_, \oc8051_golden_model_1.ACC [2], _39095_);
  or (_38366_, _38365_, _38364_);
  or (_38367_, _38366_, _38363_);
  nor (_38368_, _02551_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38370_, _02551_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38371_, _38370_, _38368_);
  and (_38372_, _02667_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38373_, _02667_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_38374_, _38373_, _38372_);
  or (_38375_, _38374_, _38371_);
  or (_38376_, _38375_, _38367_);
  or (_38377_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38378_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38379_, _38378_, _38377_);
  or (_38381_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38382_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38383_, _38382_, _38381_);
  or (_38384_, _38383_, _38379_);
  and (_38385_, _06806_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38386_, _06806_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38387_, _38386_, _38385_);
  nand (_38388_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38389_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38390_, _38389_, _38388_);
  or (_38392_, _38390_, _38387_);
  or (_38393_, _38392_, _38384_);
  or (_38394_, _38393_, _38376_);
  and (property_invalid_acc, _38394_, _37493_);
  and (_38395_, _23300_, _42920_);
  nor (_38396_, _23300_, _42920_);
  and (_38397_, _25117_, _42891_);
  nor (_38398_, _25117_, _42891_);
  and (_38399_, _24394_, _42904_);
  nor (_38400_, _24394_, _42904_);
  and (_38402_, _24760_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_38403_, _24029_, _42909_);
  nor (_38404_, _24760_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_38405_, _38404_, _38403_);
  or (_38406_, _38405_, _38402_);
  nor (_38407_, _25478_, _42886_);
  and (_38408_, _25478_, _42886_);
  and (_38409_, _24029_, _42909_);
  nor (_38410_, _26154_, _38518_);
  and (_38411_, _26154_, _38518_);
  and (_38412_, _25822_, _38512_);
  nor (_38413_, _25822_, _38512_);
  nand (_38414_, _26478_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_38415_, _26478_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38416_, _38415_, _38414_);
  or (_38417_, _27102_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_38418_, _27102_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38419_, _38418_, _38417_);
  or (_38420_, _22909_, _42925_);
  nand (_38421_, _22909_, _42925_);
  and (_38423_, _38421_, _38420_);
  or (_38424_, _38423_, _38419_);
  and (_38425_, _09985_, _38540_);
  nor (_38426_, _09985_, _38540_);
  or (_38427_, _38426_, _38425_);
  or (_38428_, _38427_, _38424_);
  nor (_38429_, _27710_, _38535_);
  and (_38430_, _27710_, _38535_);
  or (_38431_, _38430_, _38429_);
  or (_38432_, _38431_, _38428_);
  and (_38434_, _26787_, _38508_);
  nor (_38435_, _26787_, _38508_);
  or (_38436_, _38435_, _38434_);
  or (_38437_, _38436_, _38432_);
  and (_38438_, _27409_, _38504_);
  nor (_38439_, _27409_, _38504_);
  or (_38440_, _38439_, _38438_);
  or (_38441_, _38440_, _38437_);
  or (_38442_, _38441_, _38416_);
  or (_38443_, _38442_, _38413_);
  or (_38445_, _38443_, _38412_);
  or (_38446_, _38445_, _38411_);
  or (_38447_, _38446_, _38410_);
  or (_38448_, _38447_, _38409_);
  or (_38449_, _38448_, _38408_);
  or (_38450_, _38449_, _38407_);
  or (_38451_, _38450_, _38406_);
  or (_38452_, _38451_, _38400_);
  or (_38453_, _38452_, _38399_);
  nor (_38454_, _23666_, _42915_);
  and (_38456_, _23666_, _42915_);
  or (_38457_, _38456_, _38454_);
  or (_38458_, _38457_, _38453_);
  or (_38459_, _38458_, _38398_);
  or (_38460_, _38459_, _38397_);
  or (_38461_, _38460_, _38396_);
  or (_38462_, _38461_, _38395_);
  and (property_invalid_pc, _38462_, _37143_);
  buf (_44045_, _43998_);
  buf (_44093_, _43998_);
  buf (_00033_, _43998_);
  buf (_00072_, _43998_);
  buf (_00114_, _43998_);
  buf (_00156_, _43998_);
  buf (_00199_, _43998_);
  buf (_00246_, _43998_);
  buf (_00290_, _43998_);
  buf (_00332_, _43998_);
  buf (_00381_, _43998_);
  buf (_00434_, _43998_);
  buf (_00487_, _43998_);
  buf (_00540_, _43998_);
  buf (_00593_, _43998_);
  buf (_38841_, _38736_);
  buf (_38843_, _38737_);
  buf (_38856_, _38736_);
  buf (_38857_, _38737_);
  buf (_39165_, _38757_);
  buf (_39166_, _38758_);
  buf (_39167_, _38759_);
  buf (_39168_, _38760_);
  buf (_39169_, _38761_);
  buf (_39170_, _38763_);
  buf (_39171_, _38764_);
  buf (_39172_, _38765_);
  buf (_39174_, _38766_);
  buf (_39175_, _38767_);
  buf (_39176_, _38769_);
  buf (_39177_, _38770_);
  buf (_39178_, _38771_);
  buf (_39179_, _38772_);
  buf (_39231_, _38757_);
  buf (_39232_, _38758_);
  buf (_39233_, _38759_);
  buf (_39234_, _38760_);
  buf (_39235_, _38761_);
  buf (_39236_, _38763_);
  buf (_39237_, _38764_);
  buf (_39238_, _38765_);
  buf (_39240_, _38766_);
  buf (_39241_, _38767_);
  buf (_39242_, _38769_);
  buf (_39243_, _38770_);
  buf (_39244_, _38771_);
  buf (_39245_, _38772_);
  buf (_39571_, _39538_);
  buf (_39683_, _39538_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _44001_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _44005_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _44009_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _44012_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _44016_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _44020_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _44023_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _43995_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _43998_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _44049_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _44053_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _44056_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _44060_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _44063_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _44067_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _44071_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _44043_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _44045_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00335_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00338_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00342_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00344_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00348_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00352_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00356_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00329_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00332_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00385_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00389_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00393_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00397_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00401_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00405_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00409_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00378_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00381_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00438_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00442_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00446_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00450_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00454_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00458_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00462_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00431_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00434_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00491_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00495_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00499_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00503_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00507_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00511_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00515_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00484_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00487_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00544_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00548_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00552_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00556_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00560_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00564_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00568_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00537_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00540_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00597_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00601_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00605_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00609_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00613_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00617_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00621_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00590_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00593_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _44097_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _44100_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _44104_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00008_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00009_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00010_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00013_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _44090_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _44093_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00036_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00039_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00042_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00045_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00046_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00050_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00053_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00030_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00033_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00075_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00079_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00082_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00085_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00088_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00092_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00095_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00070_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00072_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00117_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00121_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00124_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00127_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00130_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00134_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00137_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00112_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00114_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00159_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00163_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00166_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00169_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00172_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00176_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00179_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00154_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00156_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00203_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00206_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00210_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00213_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00217_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00221_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00224_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00196_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00199_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00249_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00253_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00256_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00260_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00263_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00266_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00270_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00243_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00246_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00293_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00296_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00300_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00303_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00306_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00309_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00313_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00287_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00290_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40710_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40711_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40712_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40713_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40714_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40715_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40716_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40484_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40699_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40700_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40702_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40703_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40704_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40705_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40706_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40707_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40688_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40689_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40691_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40692_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40693_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40694_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40695_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40697_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40678_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40679_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40680_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40681_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40682_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40683_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40684_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40685_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40667_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40668_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40669_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40670_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40672_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40673_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40674_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40675_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40656_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40657_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40658_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40659_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40660_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40662_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40663_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40664_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40645_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40646_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40647_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40648_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40649_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40651_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40652_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40653_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40633_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40634_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40635_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40636_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40637_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40638_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40640_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40641_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40622_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40623_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40624_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40625_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40627_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40628_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40629_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40630_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40611_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40612_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40613_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40614_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40615_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40617_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40618_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40619_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40600_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40601_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40602_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40603_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40604_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40606_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40607_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40608_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40588_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40590_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40591_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40592_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40593_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40594_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40596_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40597_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40577_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40578_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40579_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40580_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40582_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40583_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40584_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40585_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40566_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40567_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40568_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40569_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40570_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40571_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40573_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40574_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40554_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40555_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40556_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40557_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40559_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40560_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40561_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40562_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40542_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40543_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40545_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40546_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40547_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40548_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40549_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40550_);
  dff (\oc8051_golden_model_1.B [0], _43414_);
  dff (\oc8051_golden_model_1.B [1], _43415_);
  dff (\oc8051_golden_model_1.B [2], _43416_);
  dff (\oc8051_golden_model_1.B [3], _43417_);
  dff (\oc8051_golden_model_1.B [4], _43418_);
  dff (\oc8051_golden_model_1.B [5], _43419_);
  dff (\oc8051_golden_model_1.B [6], _43421_);
  dff (\oc8051_golden_model_1.B [7], _40486_);
  dff (\oc8051_golden_model_1.ACC [0], _43422_);
  dff (\oc8051_golden_model_1.ACC [1], _43423_);
  dff (\oc8051_golden_model_1.ACC [2], _43424_);
  dff (\oc8051_golden_model_1.ACC [3], _43425_);
  dff (\oc8051_golden_model_1.ACC [4], _43426_);
  dff (\oc8051_golden_model_1.ACC [5], _43427_);
  dff (\oc8051_golden_model_1.ACC [6], _43428_);
  dff (\oc8051_golden_model_1.ACC [7], _40487_);
  dff (\oc8051_golden_model_1.DPL [0], _43430_);
  dff (\oc8051_golden_model_1.DPL [1], _43431_);
  dff (\oc8051_golden_model_1.DPL [2], _43432_);
  dff (\oc8051_golden_model_1.DPL [3], _43433_);
  dff (\oc8051_golden_model_1.DPL [4], _43434_);
  dff (\oc8051_golden_model_1.DPL [5], _43435_);
  dff (\oc8051_golden_model_1.DPL [6], _43436_);
  dff (\oc8051_golden_model_1.DPL [7], _40488_);
  dff (\oc8051_golden_model_1.DPH [0], _43438_);
  dff (\oc8051_golden_model_1.DPH [1], _43439_);
  dff (\oc8051_golden_model_1.DPH [2], _43440_);
  dff (\oc8051_golden_model_1.DPH [3], _43441_);
  dff (\oc8051_golden_model_1.DPH [4], _43443_);
  dff (\oc8051_golden_model_1.DPH [5], _43444_);
  dff (\oc8051_golden_model_1.DPH [6], _43445_);
  dff (\oc8051_golden_model_1.DPH [7], _40489_);
  dff (\oc8051_golden_model_1.IE [0], _43446_);
  dff (\oc8051_golden_model_1.IE [1], _43447_);
  dff (\oc8051_golden_model_1.IE [2], _43448_);
  dff (\oc8051_golden_model_1.IE [3], _43449_);
  dff (\oc8051_golden_model_1.IE [4], _43450_);
  dff (\oc8051_golden_model_1.IE [5], _43451_);
  dff (\oc8051_golden_model_1.IE [6], _43452_);
  dff (\oc8051_golden_model_1.IE [7], _40490_);
  dff (\oc8051_golden_model_1.IP [0], _43454_);
  dff (\oc8051_golden_model_1.IP [1], _43455_);
  dff (\oc8051_golden_model_1.IP [2], _43456_);
  dff (\oc8051_golden_model_1.IP [3], _43457_);
  dff (\oc8051_golden_model_1.IP [4], _43458_);
  dff (\oc8051_golden_model_1.IP [5], _43459_);
  dff (\oc8051_golden_model_1.IP [6], _43461_);
  dff (\oc8051_golden_model_1.IP [7], _40491_);
  dff (\oc8051_golden_model_1.P0 [0], _43462_);
  dff (\oc8051_golden_model_1.P0 [1], _43463_);
  dff (\oc8051_golden_model_1.P0 [2], _43465_);
  dff (\oc8051_golden_model_1.P0 [3], _43466_);
  dff (\oc8051_golden_model_1.P0 [4], _43467_);
  dff (\oc8051_golden_model_1.P0 [5], _43468_);
  dff (\oc8051_golden_model_1.P0 [6], _43469_);
  dff (\oc8051_golden_model_1.P0 [7], _40492_);
  dff (\oc8051_golden_model_1.P1 [0], _43470_);
  dff (\oc8051_golden_model_1.P1 [1], _43471_);
  dff (\oc8051_golden_model_1.P1 [2], _43472_);
  dff (\oc8051_golden_model_1.P1 [3], _43473_);
  dff (\oc8051_golden_model_1.P1 [4], _43474_);
  dff (\oc8051_golden_model_1.P1 [5], _43475_);
  dff (\oc8051_golden_model_1.P1 [6], _43476_);
  dff (\oc8051_golden_model_1.P1 [7], _40493_);
  dff (\oc8051_golden_model_1.P2 [0], _43478_);
  dff (\oc8051_golden_model_1.P2 [1], _43479_);
  dff (\oc8051_golden_model_1.P2 [2], _43480_);
  dff (\oc8051_golden_model_1.P2 [3], _43481_);
  dff (\oc8051_golden_model_1.P2 [4], _43483_);
  dff (\oc8051_golden_model_1.P2 [5], _43484_);
  dff (\oc8051_golden_model_1.P2 [6], _43485_);
  dff (\oc8051_golden_model_1.P2 [7], _40494_);
  dff (\oc8051_golden_model_1.P3 [0], _43487_);
  dff (\oc8051_golden_model_1.P3 [1], _43488_);
  dff (\oc8051_golden_model_1.P3 [2], _43489_);
  dff (\oc8051_golden_model_1.P3 [3], _43490_);
  dff (\oc8051_golden_model_1.P3 [4], _43491_);
  dff (\oc8051_golden_model_1.P3 [5], _43492_);
  dff (\oc8051_golden_model_1.P3 [6], _43493_);
  dff (\oc8051_golden_model_1.P3 [7], _40495_);
  dff (\oc8051_golden_model_1.PC [0], _43495_);
  dff (\oc8051_golden_model_1.PC [1], _43496_);
  dff (\oc8051_golden_model_1.PC [2], _43497_);
  dff (\oc8051_golden_model_1.PC [3], _43498_);
  dff (\oc8051_golden_model_1.PC [4], _43499_);
  dff (\oc8051_golden_model_1.PC [5], _43500_);
  dff (\oc8051_golden_model_1.PC [6], _43501_);
  dff (\oc8051_golden_model_1.PC [7], _43502_);
  dff (\oc8051_golden_model_1.PC [8], _43504_);
  dff (\oc8051_golden_model_1.PC [9], _43505_);
  dff (\oc8051_golden_model_1.PC [10], _43506_);
  dff (\oc8051_golden_model_1.PC [11], _43507_);
  dff (\oc8051_golden_model_1.PC [12], _43508_);
  dff (\oc8051_golden_model_1.PC [13], _43509_);
  dff (\oc8051_golden_model_1.PC [14], _43510_);
  dff (\oc8051_golden_model_1.PC [15], _40497_);
  dff (\oc8051_golden_model_1.PSW [0], _43512_);
  dff (\oc8051_golden_model_1.PSW [1], _43513_);
  dff (\oc8051_golden_model_1.PSW [2], _43514_);
  dff (\oc8051_golden_model_1.PSW [3], _43515_);
  dff (\oc8051_golden_model_1.PSW [4], _43516_);
  dff (\oc8051_golden_model_1.PSW [5], _43517_);
  dff (\oc8051_golden_model_1.PSW [6], _43518_);
  dff (\oc8051_golden_model_1.PSW [7], _40498_);
  dff (\oc8051_golden_model_1.PCON [0], _43519_);
  dff (\oc8051_golden_model_1.PCON [1], _43520_);
  dff (\oc8051_golden_model_1.PCON [2], _43522_);
  dff (\oc8051_golden_model_1.PCON [3], _43523_);
  dff (\oc8051_golden_model_1.PCON [4], _43524_);
  dff (\oc8051_golden_model_1.PCON [5], _43525_);
  dff (\oc8051_golden_model_1.PCON [6], _43526_);
  dff (\oc8051_golden_model_1.PCON [7], _40499_);
  dff (\oc8051_golden_model_1.SBUF [0], _43528_);
  dff (\oc8051_golden_model_1.SBUF [1], _43529_);
  dff (\oc8051_golden_model_1.SBUF [2], _43530_);
  dff (\oc8051_golden_model_1.SBUF [3], _43531_);
  dff (\oc8051_golden_model_1.SBUF [4], _43532_);
  dff (\oc8051_golden_model_1.SBUF [5], _43533_);
  dff (\oc8051_golden_model_1.SBUF [6], _43534_);
  dff (\oc8051_golden_model_1.SBUF [7], _40500_);
  dff (\oc8051_golden_model_1.SCON [0], _43536_);
  dff (\oc8051_golden_model_1.SCON [1], _43537_);
  dff (\oc8051_golden_model_1.SCON [2], _43538_);
  dff (\oc8051_golden_model_1.SCON [3], _43539_);
  dff (\oc8051_golden_model_1.SCON [4], _43540_);
  dff (\oc8051_golden_model_1.SCON [5], _43541_);
  dff (\oc8051_golden_model_1.SCON [6], _43542_);
  dff (\oc8051_golden_model_1.SCON [7], _40501_);
  dff (\oc8051_golden_model_1.SP [0], _43544_);
  dff (\oc8051_golden_model_1.SP [1], _43545_);
  dff (\oc8051_golden_model_1.SP [2], _43546_);
  dff (\oc8051_golden_model_1.SP [3], _43547_);
  dff (\oc8051_golden_model_1.SP [4], _43548_);
  dff (\oc8051_golden_model_1.SP [5], _43549_);
  dff (\oc8051_golden_model_1.SP [6], _43550_);
  dff (\oc8051_golden_model_1.SP [7], _40503_);
  dff (\oc8051_golden_model_1.TCON [0], _43552_);
  dff (\oc8051_golden_model_1.TCON [1], _43553_);
  dff (\oc8051_golden_model_1.TCON [2], _43554_);
  dff (\oc8051_golden_model_1.TCON [3], _43555_);
  dff (\oc8051_golden_model_1.TCON [4], _43556_);
  dff (\oc8051_golden_model_1.TCON [5], _43557_);
  dff (\oc8051_golden_model_1.TCON [6], _43559_);
  dff (\oc8051_golden_model_1.TCON [7], _40504_);
  dff (\oc8051_golden_model_1.TH0 [0], _43560_);
  dff (\oc8051_golden_model_1.TH0 [1], _43561_);
  dff (\oc8051_golden_model_1.TH0 [2], _43562_);
  dff (\oc8051_golden_model_1.TH0 [3], _43563_);
  dff (\oc8051_golden_model_1.TH0 [4], _43564_);
  dff (\oc8051_golden_model_1.TH0 [5], _43565_);
  dff (\oc8051_golden_model_1.TH0 [6], _43566_);
  dff (\oc8051_golden_model_1.TH0 [7], _40505_);
  dff (\oc8051_golden_model_1.TH1 [0], _43568_);
  dff (\oc8051_golden_model_1.TH1 [1], _43569_);
  dff (\oc8051_golden_model_1.TH1 [2], _43570_);
  dff (\oc8051_golden_model_1.TH1 [3], _43571_);
  dff (\oc8051_golden_model_1.TH1 [4], _43572_);
  dff (\oc8051_golden_model_1.TH1 [5], _43573_);
  dff (\oc8051_golden_model_1.TH1 [6], _43574_);
  dff (\oc8051_golden_model_1.TH1 [7], _40506_);
  dff (\oc8051_golden_model_1.TL0 [0], _43576_);
  dff (\oc8051_golden_model_1.TL0 [1], _43577_);
  dff (\oc8051_golden_model_1.TL0 [2], _43578_);
  dff (\oc8051_golden_model_1.TL0 [3], _43579_);
  dff (\oc8051_golden_model_1.TL0 [4], _43581_);
  dff (\oc8051_golden_model_1.TL0 [5], _43582_);
  dff (\oc8051_golden_model_1.TL0 [6], _43583_);
  dff (\oc8051_golden_model_1.TL0 [7], _40507_);
  dff (\oc8051_golden_model_1.TL1 [0], _43584_);
  dff (\oc8051_golden_model_1.TL1 [1], _43585_);
  dff (\oc8051_golden_model_1.TL1 [2], _43586_);
  dff (\oc8051_golden_model_1.TL1 [3], _43587_);
  dff (\oc8051_golden_model_1.TL1 [4], _43588_);
  dff (\oc8051_golden_model_1.TL1 [5], _43589_);
  dff (\oc8051_golden_model_1.TL1 [6], _43590_);
  dff (\oc8051_golden_model_1.TL1 [7], _40508_);
  dff (\oc8051_golden_model_1.TMOD [0], _43592_);
  dff (\oc8051_golden_model_1.TMOD [1], _43593_);
  dff (\oc8051_golden_model_1.TMOD [2], _43594_);
  dff (\oc8051_golden_model_1.TMOD [3], _43595_);
  dff (\oc8051_golden_model_1.TMOD [4], _43596_);
  dff (\oc8051_golden_model_1.TMOD [5], _43597_);
  dff (\oc8051_golden_model_1.TMOD [6], _43599_);
  dff (\oc8051_golden_model_1.TMOD [7], _40509_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43600_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43601_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43603_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43604_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43605_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43606_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43607_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40510_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43608_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43609_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43610_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43611_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43612_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43613_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43614_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40511_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43616_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43617_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43618_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43619_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43621_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43622_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43623_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40512_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43625_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43626_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43627_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43628_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43629_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43630_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43631_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40514_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03050_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03061_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03082_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03104_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03125_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _01072_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03136_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _01042_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03147_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03158_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03169_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03180_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03191_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03202_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03213_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01082_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02688_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _24751_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02889_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03093_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03304_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03505_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03706_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03907_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _04108_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04309_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04423_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04536_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04637_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04738_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04839_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04940_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _05041_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _26945_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38749_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38750_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38751_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38752_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38753_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38754_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38755_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38734_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38757_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38758_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38759_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38760_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38761_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38763_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38764_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38736_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38765_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38766_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38767_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38769_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38770_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38771_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38772_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38737_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04369_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _28812_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04372_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _28814_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04375_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _28816_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _28818_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04378_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _28820_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _28822_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04381_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _28824_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04384_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _28826_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _28828_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _28830_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04387_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _28833_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04390_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _04393_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _04453_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _04455_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04357_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _04458_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _04461_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04360_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _04464_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _04363_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _04467_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _04470_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _04473_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _04476_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _04479_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _04482_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _04485_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _04366_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39538_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38926_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38934_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39119_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39127_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39133_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38844_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38846_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39219_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38852_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39225_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39230_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39231_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39235_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39237_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39241_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39243_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39245_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38858_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39246_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39249_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39251_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39252_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38862_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39254_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39256_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39257_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39258_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39260_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39262_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39263_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39265_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39266_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39268_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39269_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39270_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39271_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39272_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39273_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39277_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39283_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39284_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39289_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39290_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39292_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39294_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39296_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38866_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39299_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39305_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39308_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39311_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39312_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39313_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38870_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39314_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39316_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39317_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39318_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39320_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39321_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39322_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39323_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39324_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39325_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39327_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39328_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39329_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39330_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38875_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39681_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39699_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39700_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39702_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39703_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39704_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39705_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39706_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39682_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39683_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39707_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39708_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _41661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _41666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _41671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _41676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _41681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _41686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _41692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _41694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _41732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _41735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _41739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _41742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _41746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _41749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _41753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _41756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _41906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _41910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _41913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _41917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _41920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _41924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _41927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _41930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _41876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _41879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _41883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _41886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _41890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _41893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _41897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _41899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _41847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _41851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _41854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _41858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _41862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _41865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _41869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _41871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _41819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _41823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _41826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _41830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _41833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _41837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _41840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _41843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _41791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _41795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _41798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _41802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _41805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _41809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _41812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _41815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _41761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _41764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _41768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _41771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _41775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _41778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _41782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _41784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _41701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _41705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _41708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _41712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _41715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _41719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _41722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _41725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _41934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _41938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _41941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _41945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _41948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _41952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _41955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _41958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _42088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _42092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _42096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _42099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _42103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _42106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _42110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _42113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _42056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _42060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _42064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _42068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _42072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _42076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _42080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _42083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _42024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _42028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _42032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _42036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _42040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _42044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _42048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _42051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _41991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _41995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _41999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _42003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _42007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _42011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _42015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _42018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _41962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _41966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _41968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _41972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _41975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _41979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _41983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _41986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _42118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _42122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _42126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _42129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _42133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _42137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _42141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _41418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _43977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _43979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _43980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _43982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _43984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _43986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _43988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _41408_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39567_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39569_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39629_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39631_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39632_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39633_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39634_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39635_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39636_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39570_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24377_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22437_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08996_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _09007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _09018_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _09029_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41319_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10770_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10781_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09600_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1046 , \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1063 , \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1214 , \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1300 , \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1424 [8], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1425 , \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1430 [4], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1431 , \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1439 , \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1456 , \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1461 [8], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1462 , \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1475 , \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1496 [8], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1497 , \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1593 [8], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1594 , \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1597 [4], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1598 , \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1605 , \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1622 , \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1627 [8], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1630 [4], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1631 , \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1638 , \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1655 , \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1748 [0], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1748 [1], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1748 [2], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1748 [3], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1748 [4], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1748 [5], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1748 [6], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1821 , \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1879 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1879 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1879 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1879 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1879 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1879 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1879 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1880 [0], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1880 [1], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1880 [2], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1880 [3], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1880 [4], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1880 [5], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1880 [6], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1936 , \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1953 , \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2085 , \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2102 , \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2141 , \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2200 , \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2444 , \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2446 , \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2452 , \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [1], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 [5], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2484 [6], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [1], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 [5], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2514 [6], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2734 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2734 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2734 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2734 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2734 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2734 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2734 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2735 [0], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2752 , \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2753 , \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2754 , \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2755 , \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2756 , \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2757 , \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2758 , \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2759 , \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2853 , \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2875 , \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(PC_gm[0], \oc8051_golden_model_1.PC [0]);
  buf(PC_gm[1], \oc8051_golden_model_1.PC [1]);
  buf(PC_gm[2], \oc8051_golden_model_1.PC [2]);
  buf(PC_gm[3], \oc8051_golden_model_1.PC [3]);
  buf(PC_gm[4], \oc8051_golden_model_1.PC [4]);
  buf(PC_gm[5], \oc8051_golden_model_1.PC [5]);
  buf(PC_gm[6], \oc8051_golden_model_1.PC [6]);
  buf(PC_gm[7], \oc8051_golden_model_1.PC [7]);
  buf(PC_gm[8], \oc8051_golden_model_1.PC [8]);
  buf(PC_gm[9], \oc8051_golden_model_1.PC [9]);
  buf(PC_gm[10], \oc8051_golden_model_1.PC [10]);
  buf(PC_gm[11], \oc8051_golden_model_1.PC [11]);
  buf(PC_gm[12], \oc8051_golden_model_1.PC [12]);
  buf(PC_gm[13], \oc8051_golden_model_1.PC [13]);
  buf(PC_gm[14], \oc8051_golden_model_1.PC [14]);
  buf(PC_gm[15], \oc8051_golden_model_1.PC [15]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc_impl[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc_impl[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc_impl[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc_impl[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc_impl[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc_impl[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc_impl[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc_impl[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc_impl[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc_impl[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc_impl[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc_impl[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc_impl[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc_impl[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc_impl[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc_impl[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(property_invalid_dec_rom_pc, 1'b0);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
