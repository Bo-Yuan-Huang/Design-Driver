
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, property_invalid_jc, property_invalid_jnc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire [15:0] _28201_;
  wire [7:0] _28202_;
  wire [7:0] _28203_;
  wire [7:0] _28204_;
  wire [7:0] _28205_;
  wire [7:0] _28206_;
  wire [7:0] _28207_;
  wire [7:0] _28208_;
  wire [7:0] _28209_;
  wire [7:0] _28210_;
  wire [7:0] _28211_;
  wire [7:0] _28212_;
  wire [7:0] _28213_;
  wire [7:0] _28214_;
  wire [7:0] _28215_;
  wire [7:0] _28216_;
  wire [7:0] _28217_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_ajmp;
  output property_invalid_jc;
  output property_invalid_jnc;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [31:0] word_in;
  not _28218_ (_23914_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _28219_ (_23915_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _23914_);
  and _28220_ (_23916_, _23915_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _28221_ (_23917_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _23914_);
  and _28222_ (_23918_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _23914_);
  nor _28223_ (_23919_, _23918_, _23917_);
  and _28224_ (_23920_, _23919_, _23916_);
  not _28225_ (_23921_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _28226_ (_23922_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _23921_);
  not _28227_ (_23923_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _28228_ (_23924_, _23923_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nor _28229_ (_23925_, _23924_, _23922_);
  nand _28230_ (_23926_, _23925_, _23920_);
  not _28231_ (_27355_, rst);
  or _28232_ (_23927_, _23920_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _28233_ (_23928_, _23927_, _27355_);
  and _28234_ (_23530_, _23928_, _23926_);
  nor _28235_ (_23929_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _28236_ (_23930_, _23929_);
  and _28237_ (_23931_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not _28238_ (_23932_, _23931_);
  and _28239_ (_23933_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _28240_ (_23934_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _28241_ (_23935_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _28242_ (_23936_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _28243_ (_23937_, _23936_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _28244_ (_23938_, _23937_, _23935_);
  or _28245_ (_23939_, _23938_, _23934_);
  not _28246_ (_23940_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _28247_ (_23941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _28248_ (_23942_, _23941_, _23935_);
  or _28249_ (_23943_, _23942_, _23940_);
  and _28250_ (_23944_, _23943_, _23939_);
  or _28251_ (_23945_, _23937_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _28252_ (_23946_, _23945_);
  nand _28253_ (_23947_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _28254_ (_23948_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _28255_ (_23949_, _23948_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _28256_ (_23950_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _28257_ (_23951_, _23950_, _23947_);
  and _28258_ (_23952_, _23951_, _23944_);
  not _28259_ (_23953_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _28260_ (_23954_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23953_);
  or _28261_ (_23955_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not _28262_ (_23956_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _28263_ (_23957_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23956_);
  and _28264_ (_23958_, _23957_, _23955_);
  or _28265_ (_23959_, _23958_, _23954_);
  nand _28266_ (_23960_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23953_);
  or _28267_ (_23961_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _28268_ (_23962_, _23961_, _23959_);
  or _28269_ (_23963_, _23941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _28270_ (_23964_, _23963_, _23962_);
  not _28271_ (_23965_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _28272_ (_23966_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _28273_ (_23967_, _23966_, _23935_);
  or _28274_ (_23968_, _23967_, _23965_);
  and _28275_ (_23969_, _23966_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _28276_ (_23970_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _28277_ (_23971_, _23970_, _23968_);
  and _28278_ (_23972_, _23971_, _23964_);
  and _28279_ (_23973_, _23972_, _23952_);
  not _28280_ (_23974_, _23973_);
  or _28281_ (_23975_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or _28282_ (_23976_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or _28283_ (_23977_, _23956_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and _28284_ (_23978_, _23977_, _23976_);
  or _28285_ (_23979_, _23978_, _23954_);
  or _28286_ (_23980_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _28287_ (_23981_, _23980_, _23979_);
  or _28288_ (_23982_, _23981_, _23975_);
  and _28289_ (_23983_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _28290_ (_23984_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _28291_ (_23985_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _28292_ (_23986_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _28293_ (_23987_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _23986_);
  nor _28294_ (_23988_, _23987_, _23985_);
  nor _28295_ (_23989_, _23988_, _23984_);
  and _28296_ (_23990_, _23989_, _23982_);
  nand _28297_ (_23991_, _23990_, _23929_);
  not _28298_ (_23992_, _23922_);
  or _28299_ (_23993_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or _28300_ (_23994_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23956_);
  and _28301_ (_23995_, _23994_, _23993_);
  or _28302_ (_23996_, _23995_, _23954_);
  or _28303_ (_23997_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _28304_ (_23998_, _23997_, _23996_);
  or _28305_ (_23999_, _23998_, _23975_);
  nand _28306_ (_24000_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not _28307_ (_24001_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _28308_ (_24002_, _23987_, _24001_);
  and _28309_ (_24003_, _24002_, _24000_);
  and _28310_ (_24004_, _24003_, _23999_);
  or _28311_ (_24005_, _24004_, _23992_);
  not _28312_ (_24006_, _23924_);
  or _28313_ (_24007_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _28314_ (_24008_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23956_);
  and _28315_ (_24009_, _24008_, _24007_);
  or _28316_ (_24010_, _24009_, _23954_);
  or _28317_ (_24011_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _28318_ (_24012_, _24011_, _24010_);
  or _28319_ (_24013_, _24012_, _23975_);
  nand _28320_ (_24014_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not _28321_ (_24015_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _28322_ (_24016_, _23987_, _24015_);
  and _28323_ (_24017_, _24016_, _24014_);
  and _28324_ (_24018_, _24017_, _24013_);
  or _28325_ (_24019_, _24018_, _24006_);
  and _28326_ (_24020_, _24019_, _24005_);
  or _28327_ (_24021_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _28328_ (_24022_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23956_);
  and _28329_ (_24023_, _24022_, _24021_);
  or _28330_ (_24024_, _24023_, _23954_);
  or _28331_ (_24025_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _28332_ (_24026_, _24025_, _24024_);
  or _28333_ (_24027_, _24026_, _23975_);
  nand _28334_ (_24028_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not _28335_ (_24029_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _28336_ (_24030_, _23987_, _24029_);
  and _28337_ (_24031_, _24030_, _24028_);
  nand _28338_ (_24032_, _24031_, _24027_);
  or _28339_ (_24033_, _24032_, _23921_);
  nand _28340_ (_24034_, _24033_, _23925_);
  nand _28341_ (_24035_, _24034_, _24020_);
  and _28342_ (_24036_, _24035_, _23991_);
  and _28343_ (_24037_, _24036_, _23974_);
  or _28344_ (_24038_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or _28345_ (_24039_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23956_);
  and _28346_ (_24040_, _24039_, _24038_);
  or _28347_ (_24041_, _24040_, _23954_);
  or _28348_ (_24042_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _28349_ (_24043_, _24042_, _24041_);
  or _28350_ (_24044_, _24043_, _23975_);
  nand _28351_ (_24045_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not _28352_ (_24046_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _28353_ (_24047_, _23987_, _24046_);
  and _28354_ (_24048_, _24047_, _24045_);
  nand _28355_ (_24049_, _24048_, _24044_);
  or _28356_ (_24050_, _24049_, _23930_);
  or _28357_ (_24051_, _23962_, _23975_);
  nand _28358_ (_24052_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or _28359_ (_24053_, _23987_, _23965_);
  and _28360_ (_24054_, _24053_, _24052_);
  and _28361_ (_24055_, _24054_, _24051_);
  or _28362_ (_24056_, _24055_, _23992_);
  or _28363_ (_24057_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or _28364_ (_24058_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23956_);
  and _28365_ (_24059_, _24058_, _24057_);
  or _28366_ (_24060_, _24059_, _23954_);
  or _28367_ (_24061_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _28368_ (_24062_, _24061_, _24060_);
  or _28369_ (_24063_, _24062_, _23975_);
  nand _28370_ (_24064_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _28371_ (_24065_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _28372_ (_24066_, _23987_, _24065_);
  and _28373_ (_24067_, _24066_, _24064_);
  and _28374_ (_24068_, _24067_, _24063_);
  or _28375_ (_24069_, _24068_, _24006_);
  and _28376_ (_24070_, _24069_, _24056_);
  or _28377_ (_24071_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _28378_ (_24072_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23956_);
  and _28379_ (_24073_, _24072_, _24071_);
  or _28380_ (_24074_, _24073_, _23954_);
  or _28381_ (_24075_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _28382_ (_24076_, _24075_, _24074_);
  or _28383_ (_24077_, _24076_, _23975_);
  nand _28384_ (_24078_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not _28385_ (_24079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _28386_ (_24080_, _23987_, _24079_);
  and _28387_ (_24081_, _24080_, _24078_);
  nand _28388_ (_24082_, _24081_, _24077_);
  or _28389_ (_24083_, _24082_, _23921_);
  nand _28390_ (_24084_, _24083_, _23925_);
  nand _28391_ (_24085_, _24084_, _24070_);
  and _28392_ (_24086_, _24085_, _24050_);
  not _28393_ (_24087_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _28394_ (_24088_, _23938_, _24087_);
  not _28395_ (_24089_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _28396_ (_24090_, _23942_, _24089_);
  and _28397_ (_24091_, _24090_, _24088_);
  nand _28398_ (_24092_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nand _28399_ (_24093_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _28400_ (_24094_, _24093_, _24092_);
  and _28401_ (_24095_, _24094_, _24091_);
  or _28402_ (_24096_, _24012_, _23963_);
  or _28403_ (_24097_, _23967_, _24015_);
  nand _28404_ (_24098_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _28405_ (_24099_, _24098_, _24097_);
  and _28406_ (_24100_, _24099_, _24096_);
  and _28407_ (_24101_, _24100_, _24095_);
  not _28408_ (_24102_, _24101_);
  and _28409_ (_24103_, _24102_, _24086_);
  and _28410_ (_24104_, _24103_, _24037_);
  and _28411_ (_24105_, _23974_, _24086_);
  not _28412_ (_24106_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _28413_ (_24107_, _23938_, _24106_);
  not _28414_ (_24108_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _28415_ (_24109_, _23942_, _24108_);
  and _28416_ (_24110_, _24109_, _24107_);
  nand _28417_ (_24111_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nand _28418_ (_24112_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _28419_ (_24113_, _24112_, _24111_);
  and _28420_ (_24114_, _24113_, _24110_);
  or _28421_ (_24115_, _23998_, _23963_);
  nand _28422_ (_24116_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  or _28423_ (_24117_, _23967_, _24001_);
  and _28424_ (_24118_, _24117_, _24116_);
  and _28425_ (_24119_, _24118_, _24115_);
  nand _28426_ (_24120_, _24119_, _24114_);
  and _28427_ (_24121_, _24120_, _24036_);
  nand _28428_ (_24122_, _24121_, _24105_);
  and _28429_ (_24123_, _24120_, _24086_);
  or _28430_ (_24124_, _24123_, _24037_);
  and _28431_ (_24125_, _24124_, _24122_);
  and _28432_ (_24126_, _24125_, _24104_);
  not _28433_ (_24127_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _28434_ (_24128_, _23938_, _24127_);
  not _28435_ (_24129_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _28436_ (_24130_, _23942_, _24129_);
  and _28437_ (_24131_, _24130_, _24128_);
  nand _28438_ (_24132_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nand _28439_ (_24133_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and _28440_ (_24134_, _24133_, _24132_);
  and _28441_ (_24135_, _24134_, _24131_);
  or _28442_ (_24136_, _23963_, _24043_);
  or _28443_ (_24137_, _23967_, _24046_);
  nand _28444_ (_24138_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _28445_ (_24139_, _24138_, _24137_);
  and _28446_ (_24140_, _24139_, _24136_);
  and _28447_ (_24141_, _24140_, _24135_);
  or _28448_ (_24142_, _24141_, _24122_);
  not _28449_ (_24143_, _24141_);
  and _28450_ (_24144_, _24143_, _24086_);
  not _28451_ (_24145_, _24144_);
  nand _28452_ (_24146_, _24145_, _24122_);
  and _28453_ (_24147_, _24146_, _24142_);
  nand _28454_ (_24148_, _24147_, _24121_);
  or _28455_ (_24149_, _24144_, _24121_);
  and _28456_ (_24150_, _24149_, _24148_);
  nand _28457_ (_24151_, _24150_, _24126_);
  not _28458_ (_24152_, _24151_);
  not _28459_ (_24153_, _24142_);
  and _28460_ (_24154_, _24147_, _24121_);
  nand _28461_ (_24155_, _24035_, _23991_);
  or _28462_ (_24156_, _24141_, _24155_);
  nand _28463_ (_24157_, _24085_, _24050_);
  not _28464_ (_24158_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _28465_ (_24159_, _23942_, _24158_);
  not _28466_ (_24160_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or _28467_ (_24161_, _23938_, _24160_);
  and _28468_ (_24162_, _24161_, _24159_);
  or _28469_ (_24163_, _23967_, _23985_);
  nand _28470_ (_24164_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _28471_ (_24165_, _24164_, _24163_);
  and _28472_ (_24166_, _24165_, _24162_);
  or _28473_ (_24167_, _23981_, _23963_);
  nand _28474_ (_24168_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nand _28475_ (_24169_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and _28476_ (_24170_, _24169_, _24168_);
  and _28477_ (_24171_, _24170_, _24167_);
  and _28478_ (_24172_, _24171_, _24166_);
  or _28479_ (_24173_, _24172_, _24157_);
  or _28480_ (_24174_, _24173_, _24156_);
  nand _28481_ (_24175_, _24173_, _24156_);
  and _28482_ (_24176_, _24175_, _24174_);
  nand _28483_ (_24177_, _24176_, _24154_);
  or _28484_ (_24178_, _24176_, _24154_);
  and _28485_ (_24179_, _24178_, _24177_);
  nand _28486_ (_24180_, _24179_, _24153_);
  or _28487_ (_24181_, _24179_, _24153_);
  and _28488_ (_24182_, _24181_, _24180_);
  nand _28489_ (_24183_, _24182_, _24152_);
  or _28490_ (_24184_, _24182_, _24152_);
  nand _28491_ (_24185_, _24184_, _24183_);
  not _28492_ (_24186_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _28493_ (_24187_, _23938_, _24186_);
  not _28494_ (_24188_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _28495_ (_24189_, _23942_, _24188_);
  and _28496_ (_24190_, _24189_, _24187_);
  nand _28497_ (_24191_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand _28498_ (_24192_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _28499_ (_24193_, _24192_, _24191_);
  and _28500_ (_24194_, _24193_, _24190_);
  or _28501_ (_24195_, _24026_, _23963_);
  or _28502_ (_24196_, _23967_, _24029_);
  nand _28503_ (_24197_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _28504_ (_24198_, _24197_, _24196_);
  and _28505_ (_24199_, _24198_, _24195_);
  nand _28506_ (_24200_, _24199_, _24194_);
  and _28507_ (_24201_, _24200_, _24036_);
  not _28508_ (_24202_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _28509_ (_24203_, _23938_, _24202_);
  not _28510_ (_24204_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _28511_ (_24205_, _23942_, _24204_);
  and _28512_ (_24206_, _24205_, _24203_);
  nand _28513_ (_24207_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  or _28514_ (_24208_, _23967_, _24065_);
  and _28515_ (_24209_, _24208_, _24207_);
  and _28516_ (_24210_, _24209_, _24206_);
  or _28517_ (_24211_, _23963_, _24062_);
  nand _28518_ (_24212_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _28519_ (_24213_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _28520_ (_24214_, _24213_, _24212_);
  and _28521_ (_24215_, _24214_, _24211_);
  nand _28522_ (_24216_, _24215_, _24210_);
  and _28523_ (_24217_, _24216_, _24086_);
  and _28524_ (_24218_, _24217_, _24201_);
  not _28525_ (_24219_, _24218_);
  and _28526_ (_24220_, _24200_, _24086_);
  not _28527_ (_24221_, _24220_);
  and _28528_ (_24222_, _24216_, _24036_);
  and _28529_ (_24223_, _24222_, _24221_);
  nand _28530_ (_24224_, _24223_, _24103_);
  nand _28531_ (_24225_, _24224_, _24219_);
  not _28532_ (_24226_, _24104_);
  and _28533_ (_24227_, _24102_, _24036_);
  or _28534_ (_24228_, _24227_, _24105_);
  and _28535_ (_24229_, _24228_, _24226_);
  and _28536_ (_24230_, _24229_, _24225_);
  not _28537_ (_24231_, _24126_);
  or _28538_ (_24232_, _24125_, _24104_);
  and _28539_ (_24233_, _24232_, _24231_);
  and _28540_ (_24234_, _24233_, _24230_);
  or _28541_ (_24235_, _24150_, _24126_);
  and _28542_ (_24236_, _24235_, _24151_);
  nand _28543_ (_24237_, _24236_, _24234_);
  not _28544_ (_24238_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _28545_ (_24239_, _23938_, _24238_);
  not _28546_ (_24240_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _28547_ (_24241_, _23942_, _24240_);
  nor _28548_ (_24242_, _24241_, _24239_);
  and _28549_ (_24243_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _28550_ (_24244_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _28551_ (_24245_, _24244_, _24243_);
  and _28552_ (_24246_, _24245_, _24242_);
  nor _28553_ (_24247_, _23963_, _24076_);
  nor _28554_ (_24248_, _23967_, _24079_);
  and _28555_ (_24249_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _28556_ (_24250_, _24249_, _24248_);
  not _28557_ (_24251_, _24250_);
  nor _28558_ (_24252_, _24251_, _24247_);
  and _28559_ (_24253_, _24252_, _24246_);
  not _28560_ (_24254_, _24253_);
  and _28561_ (_24255_, _24254_, _24036_);
  and _28562_ (_24256_, _24255_, _24220_);
  or _28563_ (_24257_, _24217_, _24201_);
  and _28564_ (_24258_, _24257_, _24219_);
  and _28565_ (_24259_, _24258_, _24256_);
  or _28566_ (_24260_, _24223_, _24103_);
  and _28567_ (_24261_, _24260_, _24224_);
  nand _28568_ (_24262_, _24261_, _24259_);
  not _28569_ (_24263_, _24262_);
  nand _28570_ (_24264_, _24229_, _24225_);
  or _28571_ (_24265_, _24229_, _24225_);
  and _28572_ (_24266_, _24265_, _24264_);
  nand _28573_ (_24267_, _24266_, _24263_);
  nand _28574_ (_24268_, _24233_, _24230_);
  or _28575_ (_24269_, _24233_, _24230_);
  nand _28576_ (_24270_, _24269_, _24268_);
  or _28577_ (_24271_, _24270_, _24267_);
  or _28578_ (_24272_, _24236_, _24234_);
  nand _28579_ (_24273_, _24272_, _24237_);
  or _28580_ (_24274_, _24273_, _24271_);
  and _28581_ (_24275_, _24274_, _24237_);
  or _28582_ (_24276_, _24275_, _24185_);
  nand _28583_ (_24277_, _24276_, _24183_);
  not _28584_ (_24278_, _24172_);
  and _28585_ (_24279_, _24278_, _24036_);
  and _28586_ (_24280_, _24279_, _24145_);
  and _28587_ (_24281_, _24180_, _24177_);
  not _28588_ (_24282_, _24281_);
  nand _28589_ (_24283_, _24282_, _24280_);
  or _28590_ (_24284_, _24282_, _24280_);
  and _28591_ (_24285_, _24284_, _24283_);
  nand _28592_ (_24286_, _24285_, _24277_);
  and _28593_ (_24287_, _24283_, _24174_);
  nand _28594_ (_24288_, _24287_, _24286_);
  nand _28595_ (_24289_, _24288_, _23933_);
  or _28596_ (_24290_, _24288_, _23933_);
  nand _28597_ (_24291_, _24290_, _24289_);
  and _28598_ (_24292_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or _28599_ (_24293_, _24285_, _24277_);
  and _28600_ (_24294_, _24293_, _24286_);
  nand _28601_ (_24295_, _24294_, _24292_);
  or _28602_ (_24296_, _24295_, _24291_);
  nand _28603_ (_24297_, _24296_, _24289_);
  and _28604_ (_24298_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _28605_ (_24299_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _28606_ (_24300_, _24299_, _24298_);
  and _28607_ (_24301_, _24300_, _24297_);
  and _28608_ (_24302_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand _28609_ (_24303_, _24275_, _24185_);
  and _28610_ (_24304_, _24303_, _24276_);
  nand _28611_ (_24305_, _24304_, _24302_);
  or _28612_ (_24309_, _24304_, _24302_);
  and _28613_ (_24310_, _24309_, _24305_);
  and _28614_ (_24311_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand _28615_ (_24312_, _24273_, _24271_);
  and _28616_ (_24313_, _24312_, _24274_);
  nand _28617_ (_24314_, _24313_, _24311_);
  or _28618_ (_24315_, _24313_, _24311_);
  nand _28619_ (_24316_, _24315_, _24314_);
  and _28620_ (_24317_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand _28621_ (_24318_, _24270_, _24267_);
  and _28622_ (_24319_, _24318_, _24271_);
  nand _28623_ (_24326_, _24319_, _24317_);
  or _28624_ (_24332_, _24319_, _24317_);
  and _28625_ (_24338_, _24332_, _24326_);
  and _28626_ (_24344_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _28627_ (_24345_, _24266_, _24263_);
  and _28628_ (_24346_, _24345_, _24267_);
  nand _28629_ (_24347_, _24346_, _24344_);
  and _28630_ (_24348_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _28631_ (_24349_, _24261_, _24259_);
  and _28632_ (_24350_, _24349_, _24262_);
  nand _28633_ (_24351_, _24350_, _24348_);
  and _28634_ (_24352_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _28635_ (_24353_, _24258_, _24256_);
  or _28636_ (_24354_, _24258_, _24256_);
  and _28637_ (_24355_, _24354_, _24353_);
  and _28638_ (_24356_, _24355_, _24352_);
  not _28639_ (_24357_, _24356_);
  or _28640_ (_24358_, _24350_, _24348_);
  nand _28641_ (_24359_, _24358_, _24351_);
  or _28642_ (_24360_, _24359_, _24357_);
  nand _28643_ (_24361_, _24360_, _24351_);
  or _28644_ (_24362_, _24346_, _24344_);
  and _28645_ (_24363_, _24362_, _24347_);
  nand _28646_ (_24364_, _24363_, _24361_);
  nand _28647_ (_24365_, _24364_, _24347_);
  nand _28648_ (_24366_, _24365_, _24338_);
  and _28649_ (_24367_, _24366_, _24326_);
  or _28650_ (_24368_, _24367_, _24316_);
  nand _28651_ (_24369_, _24368_, _24314_);
  nand _28652_ (_24371_, _24369_, _24310_);
  and _28653_ (_24373_, _24371_, _24305_);
  and _28654_ (_24374_, _24290_, _24289_);
  or _28655_ (_24375_, _24294_, _24292_);
  and _28656_ (_24376_, _24375_, _24295_);
  and _28657_ (_24377_, _24376_, _24374_);
  nand _28658_ (_24378_, _24300_, _24377_);
  nor _28659_ (_24379_, _24378_, _24373_);
  or _28660_ (_24380_, _24379_, _24301_);
  and _28661_ (_24381_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _28662_ (_24382_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _28663_ (_24383_, _24382_, _24381_);
  nand _28664_ (_24384_, _24383_, _24380_);
  nor _28665_ (_24385_, _24384_, _23932_);
  not _28666_ (_24386_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or _28667_ (_24387_, _23929_, _24386_);
  nor _28668_ (_24388_, _24387_, _24385_);
  and _28669_ (_24389_, _24385_, _24386_);
  or _28670_ (_24390_, _24389_, _24388_);
  and _28671_ (_23899_, _24390_, _27355_);
  nor _28672_ (_24391_, _23920_, _23923_);
  and _28673_ (_24392_, _23920_, _23923_);
  or _28674_ (_24393_, _24392_, _24391_);
  and _28675_ (_02784_, _24393_, _27355_);
  and _28676_ (_24394_, _24254_, _24086_);
  and _28677_ (_02984_, _24394_, _27355_);
  nor _28678_ (_24395_, _24255_, _24220_);
  nor _28679_ (_24396_, _24395_, _24256_);
  and _28680_ (_03157_, _24396_, _27355_);
  nor _28681_ (_24397_, _24355_, _24352_);
  nor _28682_ (_24398_, _24397_, _24356_);
  and _28683_ (_03302_, _24398_, _27355_);
  and _28684_ (_24399_, _24359_, _24357_);
  not _28685_ (_24400_, _24399_);
  and _28686_ (_24401_, _24400_, _24360_);
  and _28687_ (_03443_, _24401_, _27355_);
  or _28688_ (_24402_, _24363_, _24361_);
  and _28689_ (_24403_, _24402_, _24364_);
  and _28690_ (_03584_, _24403_, _27355_);
  or _28691_ (_24408_, _24365_, _24338_);
  and _28692_ (_24413_, _24408_, _24366_);
  and _28693_ (_03782_, _24413_, _27355_);
  and _28694_ (_24425_, _24367_, _24316_);
  not _28695_ (_24432_, _24425_);
  and _28696_ (_24441_, _24432_, _24368_);
  and _28697_ (_03985_, _24441_, _27355_);
  or _28698_ (_24442_, _24369_, _24310_);
  and _28699_ (_24443_, _24442_, _24371_);
  and _28700_ (_04190_, _24443_, _27355_);
  not _28701_ (_24444_, _24376_);
  or _28702_ (_24445_, _24444_, _24373_);
  not _28703_ (_24446_, _24445_);
  and _28704_ (_24447_, _24444_, _24373_);
  nor _28705_ (_24448_, _24447_, _24446_);
  and _28706_ (_04293_, _24448_, _27355_);
  and _28707_ (_24449_, _24445_, _24295_);
  or _28708_ (_24450_, _24449_, _24291_);
  nand _28709_ (_24451_, _24449_, _24291_);
  and _28710_ (_24452_, _24451_, _24450_);
  and _28711_ (_04397_, _24452_, _27355_);
  nand _28712_ (_24453_, _24450_, _24289_);
  nand _28713_ (_24454_, _24453_, _24298_);
  or _28714_ (_24455_, _24453_, _24298_);
  and _28715_ (_24456_, _24455_, _24454_);
  and _28716_ (_04499_, _24456_, _27355_);
  not _28717_ (_24457_, _24380_);
  not _28718_ (_24458_, _24299_);
  nand _28719_ (_24459_, _24458_, _24454_);
  and _28720_ (_24460_, _24459_, _24457_);
  and _28721_ (_04604_, _24460_, _27355_);
  and _28722_ (_24461_, _24381_, _24380_);
  nor _28723_ (_24462_, _24381_, _24380_);
  nor _28724_ (_24463_, _24462_, _24461_);
  and _28725_ (_04707_, _24463_, _27355_);
  or _28726_ (_24464_, _24382_, _24461_);
  and _28727_ (_24465_, _24464_, _24384_);
  and _28728_ (_04810_, _24465_, _27355_);
  and _28729_ (_24466_, _24384_, _23932_);
  or _28730_ (_24467_, _24466_, _24385_);
  nor _28731_ (_04914_, _24467_, rst);
  and _28732_ (_24468_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _23914_);
  nor _28733_ (_24469_, _24468_, _23915_);
  not _28734_ (_24471_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _28735_ (_24482_, _23917_, _24471_);
  and _28736_ (_24487_, _24482_, _24469_);
  and _28737_ (_24488_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _28738_ (_24489_, _24488_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _28739_ (_24496_, _24488_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _28740_ (_24506_, _24496_, _24489_);
  and _28741_ (_00958_, _24506_, _27355_);
  and _28742_ (_00985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _27355_);
  nor _28743_ (_24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _28744_ (_24508_, _24507_, _24172_);
  nor _28745_ (_24509_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _28746_ (_24510_, _24509_);
  and _28747_ (_24511_, _24510_, _24508_);
  not _28748_ (_24512_, _24511_);
  or _28749_ (_24513_, _24082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _28750_ (_24514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _28751_ (_24515_, _24067_, _24063_);
  or _28752_ (_24516_, _24515_, _24514_);
  and _28753_ (_24517_, _24516_, _24513_);
  or _28754_ (_24518_, _24517_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _28755_ (_24519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _28756_ (_24520_, _24054_, _24051_);
  or _28757_ (_24521_, _24520_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _28758_ (_24522_, _24049_, _24514_);
  and _28759_ (_24523_, _24522_, _24521_);
  or _28760_ (_24524_, _24523_, _24519_);
  and _28761_ (_24525_, _24524_, _24518_);
  or _28762_ (_24526_, _24525_, _24512_);
  nand _28763_ (_24527_, _24507_, _24141_);
  nor _28764_ (_24528_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _28765_ (_24529_, _24528_);
  and _28766_ (_24530_, _24529_, _24527_);
  and _28767_ (_24531_, _24032_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _28768_ (_24532_, _24531_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _28769_ (_24533_, _24017_, _24013_);
  or _28770_ (_24534_, _24533_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _28771_ (_24535_, _24003_, _23999_);
  or _28772_ (_24536_, _24535_, _24514_);
  and _28773_ (_24537_, _24536_, _24534_);
  or _28774_ (_24538_, _24537_, _24519_);
  nand _28775_ (_24539_, _24538_, _24532_);
  nand _28776_ (_24540_, _24539_, _24530_);
  nand _28777_ (_24541_, _24524_, _24518_);
  or _28778_ (_24542_, _24541_, _24511_);
  and _28779_ (_24543_, _24542_, _24526_);
  not _28780_ (_24544_, _24543_);
  or _28781_ (_24545_, _24544_, _24540_);
  and _28782_ (_24546_, _24545_, _24526_);
  or _28783_ (_24547_, _24539_, _24530_);
  and _28784_ (_24548_, _24547_, _24540_);
  and _28785_ (_24549_, _24548_, _24543_);
  not _28786_ (_24550_, _24507_);
  or _28787_ (_24551_, _24550_, _24120_);
  nor _28788_ (_24552_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _28789_ (_24553_, _24552_);
  nand _28790_ (_24554_, _24553_, _24551_);
  and _28791_ (_24555_, _24082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _28792_ (_24556_, _24555_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _28793_ (_24557_, _24515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _28794_ (_24558_, _24520_, _24514_);
  and _28795_ (_24559_, _24558_, _24557_);
  or _28796_ (_24560_, _24559_, _24519_);
  and _28797_ (_24561_, _24560_, _24556_);
  or _28798_ (_24562_, _24561_, _24554_);
  or _28799_ (_24563_, _24032_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _28800_ (_24564_, _24533_, _24514_);
  and _28801_ (_24565_, _24564_, _24563_);
  and _28802_ (_24566_, _24565_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _28803_ (_24567_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _28804_ (_24568_, _24567_);
  nand _28805_ (_24569_, _24507_, _23973_);
  and _28806_ (_24570_, _24569_, _24568_);
  not _28807_ (_24571_, _24570_);
  or _28808_ (_24572_, _24571_, _24566_);
  and _28809_ (_24573_, _24553_, _24551_);
  nand _28810_ (_24574_, _24560_, _24556_);
  or _28811_ (_24575_, _24574_, _24573_);
  nand _28812_ (_24576_, _24575_, _24562_);
  or _28813_ (_24577_, _24576_, _24572_);
  nand _28814_ (_24578_, _24577_, _24562_);
  nand _28815_ (_24579_, _24578_, _24549_);
  and _28816_ (_24580_, _24579_, _24546_);
  and _28817_ (_24581_, _24517_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _28818_ (_24582_, _24581_);
  nand _28819_ (_24583_, _24507_, _24101_);
  nor _28820_ (_24584_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _28821_ (_24585_, _24584_);
  and _28822_ (_24586_, _24585_, _24583_);
  nand _28823_ (_24587_, _24586_, _24582_);
  or _28824_ (_24588_, _24586_, _24582_);
  nand _28825_ (_24589_, _24588_, _24587_);
  nand _28826_ (_24590_, _24531_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _28827_ (_24591_, _24550_, _24216_);
  nor _28828_ (_24592_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _28829_ (_24593_, _24592_);
  and _28830_ (_24594_, _24593_, _24591_);
  nand _28831_ (_24595_, _24594_, _24590_);
  and _28832_ (_24596_, _24555_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _28833_ (_24597_, _24550_, _24200_);
  nor _28834_ (_24598_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _28835_ (_24599_, _24598_);
  nand _28836_ (_24600_, _24599_, _24597_);
  and _28837_ (_24601_, _24600_, _24596_);
  or _28838_ (_24602_, _24594_, _24590_);
  nand _28839_ (_24603_, _24602_, _24595_);
  or _28840_ (_24604_, _24603_, _24601_);
  and _28841_ (_24605_, _24604_, _24595_);
  or _28842_ (_24606_, _24605_, _24589_);
  nand _28843_ (_24607_, _24606_, _24587_);
  not _28844_ (_24608_, _24566_);
  or _28845_ (_24609_, _24570_, _24608_);
  and _28846_ (_24610_, _24609_, _24572_);
  not _28847_ (_24611_, _24610_);
  nor _28848_ (_24612_, _24576_, _24611_);
  and _28849_ (_24613_, _24612_, _24549_);
  nand _28850_ (_24614_, _24613_, _24607_);
  nand _28851_ (_24615_, _24614_, _24580_);
  not _28852_ (_24616_, _24049_);
  and _28853_ (_24617_, _23990_, _24616_);
  nor _28854_ (_24618_, _24617_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _28855_ (_24619_, _24537_, _24523_);
  or _28856_ (_24620_, _24535_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _28857_ (_24621_, _23990_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _28858_ (_24622_, _24621_, _24620_);
  nor _28859_ (_24623_, _24622_, _24559_);
  nand _28860_ (_24624_, _24623_, _24619_);
  and _28861_ (_24625_, _24624_, _24519_);
  nor _28862_ (_24626_, _24625_, _24618_);
  nor _28863_ (_24627_, _24565_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _28864_ (_24628_, _24622_, _24519_);
  nor _28865_ (_24629_, _24628_, _24627_);
  not _28866_ (_24630_, _24629_);
  and _28867_ (_24631_, _24630_, _24626_);
  and _28868_ (_24632_, _24631_, _24615_);
  nor _28869_ (_24633_, _24632_, _24512_);
  not _28870_ (_24634_, _24633_);
  not _28871_ (_24635_, _24548_);
  and _28872_ (_24636_, _24577_, _24562_);
  nand _28873_ (_24637_, _24612_, _24607_);
  and _28874_ (_24638_, _24637_, _24636_);
  or _28875_ (_24639_, _24638_, _24635_);
  and _28876_ (_24640_, _24639_, _24540_);
  nand _28877_ (_24641_, _24640_, _24543_);
  or _28878_ (_24642_, _24640_, _24543_);
  nand _28879_ (_24643_, _24642_, _24641_);
  nand _28880_ (_24644_, _24643_, _24632_);
  and _28881_ (_24645_, _24644_, _24634_);
  and _28882_ (_24646_, _24645_, _24629_);
  nor _28883_ (_24647_, _24645_, _24629_);
  and _28884_ (_24648_, _24638_, _24635_);
  not _28885_ (_24649_, _24648_);
  nand _28886_ (_24650_, _24649_, _24639_);
  nand _28887_ (_24651_, _24650_, _24632_);
  nor _28888_ (_24652_, _24632_, _24530_);
  not _28889_ (_24653_, _24652_);
  and _28890_ (_24654_, _24653_, _24651_);
  and _28891_ (_24655_, _24654_, _24541_);
  nor _28892_ (_24656_, _24655_, _24647_);
  or _28893_ (_24657_, _24656_, _24646_);
  nor _28894_ (_24658_, _24647_, _24646_);
  not _28895_ (_24659_, _24655_);
  or _28896_ (_24660_, _24654_, _24541_);
  and _28897_ (_24661_, _24660_, _24659_);
  and _28898_ (_24662_, _24661_, _24658_);
  not _28899_ (_24663_, _24632_);
  nand _28900_ (_24664_, _24610_, _24607_);
  and _28901_ (_24665_, _24664_, _24572_);
  and _28902_ (_24666_, _24576_, _24665_);
  nor _28903_ (_24667_, _24576_, _24665_);
  nor _28904_ (_24668_, _24667_, _24666_);
  nor _28905_ (_24669_, _24668_, _24663_);
  nor _28906_ (_24670_, _24632_, _24573_);
  nor _28907_ (_24671_, _24670_, _24669_);
  and _28908_ (_24672_, _24671_, _24539_);
  not _28909_ (_24673_, _24672_);
  nor _28910_ (_24674_, _24671_, _24539_);
  nor _28911_ (_24675_, _24632_, _24571_);
  nor _28912_ (_24676_, _24610_, _24607_);
  not _28913_ (_24677_, _24676_);
  and _28914_ (_24678_, _24677_, _24664_);
  and _28915_ (_24679_, _24678_, _24632_);
  or _28916_ (_24680_, _24679_, _24675_);
  and _28917_ (_24681_, _24680_, _24574_);
  not _28918_ (_24682_, _24681_);
  and _28919_ (_24683_, _24605_, _24589_);
  not _28920_ (_24684_, _24683_);
  and _28921_ (_24685_, _24684_, _24606_);
  or _28922_ (_24686_, _24685_, _24663_);
  or _28923_ (_24687_, _24632_, _24586_);
  and _28924_ (_24688_, _24687_, _24686_);
  nor _28925_ (_24689_, _24688_, _24608_);
  or _28926_ (_24690_, _24632_, _24600_);
  not _28927_ (_24691_, _24596_);
  and _28928_ (_24694_, _24600_, _24691_);
  nor _28929_ (_24705_, _24600_, _24691_);
  nor _28930_ (_24716_, _24705_, _24694_);
  nand _28931_ (_24727_, _24632_, _24716_);
  nand _28932_ (_24734_, _24727_, _24690_);
  nand _28933_ (_24742_, _24734_, _24590_);
  or _28934_ (_24753_, _24734_, _24590_);
  nand _28935_ (_24764_, _24753_, _24742_);
  nor _28936_ (_24775_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _28937_ (_24786_, _24507_, _24253_);
  nor _28938_ (_24797_, _24786_, _24775_);
  nor _28939_ (_24808_, _24797_, _24691_);
  or _28940_ (_24819_, _24808_, _24764_);
  and _28941_ (_24830_, _24819_, _24742_);
  or _28942_ (_24841_, _24632_, _24594_);
  and _28943_ (_24852_, _24603_, _24601_);
  not _28944_ (_24863_, _24852_);
  and _28945_ (_24874_, _24863_, _24604_);
  or _28946_ (_24885_, _24874_, _24663_);
  and _28947_ (_24896_, _24885_, _24841_);
  nand _28948_ (_24906_, _24896_, _24582_);
  or _28949_ (_24907_, _24896_, _24582_);
  nand _28950_ (_24908_, _24907_, _24906_);
  or _28951_ (_24909_, _24908_, _24830_);
  and _28952_ (_24910_, _24688_, _24608_);
  not _28953_ (_24911_, _24910_);
  and _28954_ (_24912_, _24911_, _24906_);
  and _28955_ (_24913_, _24912_, _24909_);
  nor _28956_ (_24914_, _24913_, _24689_);
  nor _28957_ (_24915_, _24680_, _24574_);
  nor _28958_ (_24916_, _24915_, _24681_);
  nand _28959_ (_24917_, _24916_, _24914_);
  and _28960_ (_24918_, _24917_, _24682_);
  or _28961_ (_24919_, _24918_, _24674_);
  nand _28962_ (_24920_, _24919_, _24673_);
  nand _28963_ (_24921_, _24920_, _24662_);
  nand _28964_ (_24922_, _24921_, _24657_);
  and _28965_ (_24923_, _24922_, _24626_);
  nor _28966_ (_24924_, _24923_, _24645_);
  and _28967_ (_24925_, _24920_, _24661_);
  or _28968_ (_24926_, _24925_, _24655_);
  or _28969_ (_24927_, _24926_, _24658_);
  nand _28970_ (_24928_, _24926_, _24658_);
  and _28971_ (_24929_, _24928_, _24927_);
  and _28972_ (_24930_, _24929_, _24923_);
  or _28973_ (_24931_, _24930_, _24924_);
  and _28974_ (_01001_, _24931_, _27355_);
  and _28975_ (_03039_, _24923_, _27355_);
  and _28976_ (_03049_, _24632_, _27355_);
  and _28977_ (_03068_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _27355_);
  and _28978_ (_03084_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _27355_);
  and _28979_ (_03100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _27355_);
  or _28980_ (_24932_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _28981_ (_24933_, _24488_, rst);
  and _28982_ (_03108_, _24933_, _24932_);
  nand _28983_ (_24934_, _24923_, _24596_);
  and _28984_ (_24935_, _24934_, _24797_);
  nor _28985_ (_24936_, _24934_, _24797_);
  or _28986_ (_24937_, _24936_, _24935_);
  and _28987_ (_03117_, _24937_, _27355_);
  nand _28988_ (_24938_, _24922_, _24626_);
  and _28989_ (_24939_, _24808_, _24764_);
  not _28990_ (_24940_, _24939_);
  and _28991_ (_24941_, _24940_, _24819_);
  or _28992_ (_24942_, _24941_, _24938_);
  or _28993_ (_24943_, _24923_, _24734_);
  and _28994_ (_24944_, _24943_, _24942_);
  and _28995_ (_03125_, _24944_, _27355_);
  not _28996_ (_24945_, _24909_);
  and _28997_ (_24946_, _24908_, _24830_);
  nor _28998_ (_24947_, _24946_, _24945_);
  or _28999_ (_24948_, _24947_, _24938_);
  or _29000_ (_24949_, _24923_, _24896_);
  and _29001_ (_24950_, _24949_, _24948_);
  and _29002_ (_03132_, _24950_, _27355_);
  or _29003_ (_24951_, _24910_, _24689_);
  and _29004_ (_24952_, _24909_, _24906_);
  nor _29005_ (_24953_, _24952_, _24951_);
  and _29006_ (_24954_, _24952_, _24951_);
  nor _29007_ (_24955_, _24954_, _24953_);
  or _29008_ (_24956_, _24955_, _24938_);
  or _29009_ (_24957_, _24923_, _24688_);
  and _29010_ (_24958_, _24957_, _24956_);
  and _29011_ (_03141_, _24958_, _27355_);
  or _29012_ (_24959_, _24916_, _24914_);
  and _29013_ (_24960_, _24959_, _24917_);
  or _29014_ (_24961_, _24960_, _24938_);
  or _29015_ (_24962_, _24923_, _24680_);
  and _29016_ (_24963_, _24962_, _24961_);
  and _29017_ (_03149_, _24963_, _27355_);
  or _29018_ (_24964_, _24674_, _24672_);
  nand _29019_ (_24965_, _24964_, _24918_);
  or _29020_ (_24966_, _24964_, _24918_);
  and _29021_ (_24967_, _24966_, _24965_);
  or _29022_ (_24968_, _24967_, _24938_);
  or _29023_ (_24969_, _24923_, _24671_);
  and _29024_ (_24970_, _24969_, _24968_);
  and _29025_ (_03158_, _24970_, _27355_);
  nor _29026_ (_24971_, _24920_, _24661_);
  or _29027_ (_24972_, _24971_, _24925_);
  and _29028_ (_24973_, _24972_, _24923_);
  nor _29029_ (_24974_, _24923_, _24654_);
  or _29030_ (_24975_, _24974_, _24973_);
  nor _29031_ (_03166_, _24975_, rst);
  not _29032_ (_24976_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _29033_ (_24977_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _23914_);
  and _29034_ (_24978_, _24977_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _29035_ (_24979_, _24978_, _24976_);
  and _29036_ (_24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _29037_ (_24981_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _29038_ (_24982_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _29039_ (_24983_, _24982_, _24981_);
  and _29040_ (_24984_, _24983_, _24979_);
  not _29041_ (_24985_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _29042_ (_24986_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _23914_);
  and _29043_ (_24988_, _24986_, _24976_);
  and _29044_ (_24990_, _24988_, _24985_);
  and _29045_ (_24992_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _29046_ (_24994_, _24992_, _24984_);
  not _29047_ (_24996_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _29048_ (_24998_, _24977_, _24996_);
  and _29049_ (_25000_, _24998_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _29050_ (_25002_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _29051_ (_25004_, _24998_, _24976_);
  and _29052_ (_25006_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or _29053_ (_25008_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _29054_ (_25010_, _25008_, _23914_);
  nor _29055_ (_25012_, _25010_, _24977_);
  and _29056_ (_25014_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _29057_ (_25016_, _25014_, _25006_);
  nor _29058_ (_25018_, _25016_, _25002_);
  and _29059_ (_25020_, _25018_, _24994_);
  and _29060_ (_25022_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor _29061_ (_25024_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _29062_ (_25026_, _25024_, _24980_);
  and _29063_ (_25028_, _25026_, _24979_);
  nor _29064_ (_25030_, _25028_, _25022_);
  and _29065_ (_25032_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _29066_ (_25034_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _29067_ (_25036_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _29068_ (_25038_, _25036_, _25034_);
  nor _29069_ (_25040_, _25038_, _25032_);
  and _29070_ (_25042_, _25040_, _25030_);
  and _29071_ (_25043_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and _29072_ (_25044_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _29073_ (_25045_, _25044_, _25043_);
  not _29074_ (_25046_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _29075_ (_25047_, _24979_, _25046_);
  not _29076_ (_25048_, _25047_);
  and _29077_ (_25049_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _29078_ (_25050_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _29079_ (_25051_, _25050_, _25049_);
  and _29080_ (_25052_, _25051_, _25048_);
  and _29081_ (_25053_, _25052_, _25045_);
  and _29082_ (_25054_, _25053_, _25042_);
  and _29083_ (_25055_, _25054_, _25020_);
  and _29084_ (_25056_, _24981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _29085_ (_25057_, _25056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _29086_ (_25058_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _29087_ (_25059_, _25058_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _29088_ (_25060_, _25059_);
  not _29089_ (_25061_, _24979_);
  nor _29090_ (_25062_, _25058_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _29091_ (_25063_, _25062_, _25061_);
  and _29092_ (_25064_, _25063_, _25060_);
  not _29093_ (_25065_, _25064_);
  and _29094_ (_25066_, _24978_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _29095_ (_25067_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _29096_ (_25068_, _25067_, _25066_);
  and _29097_ (_25069_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _29098_ (_25070_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _29099_ (_25071_, _25070_, _25069_);
  and _29100_ (_25072_, _25071_, _25068_);
  and _29101_ (_25073_, _25072_, _25065_);
  nor _29102_ (_25074_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _29103_ (_25075_, _25074_);
  nor _29104_ (_25076_, _25058_, _25061_);
  and _29105_ (_25077_, _25076_, _25075_);
  not _29106_ (_25078_, _25077_);
  and _29107_ (_25079_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _29108_ (_25080_, _25079_, _25066_);
  and _29109_ (_25081_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _29110_ (_25082_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _29111_ (_25083_, _25082_, _25081_);
  and _29112_ (_25084_, _25083_, _25080_);
  and _29113_ (_25085_, _25084_, _25078_);
  nor _29114_ (_25086_, _25085_, _25073_);
  not _29115_ (_25087_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _29116_ (_25088_, _25059_, _25087_);
  and _29117_ (_25089_, _25059_, _25087_);
  nor _29118_ (_25090_, _25089_, _25088_);
  nor _29119_ (_25091_, _25090_, _25061_);
  not _29120_ (_25092_, _25091_);
  and _29121_ (_25093_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not _29122_ (_25094_, _25093_);
  not _29123_ (_25095_, _25066_);
  and _29124_ (_25096_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and _29125_ (_25097_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _29126_ (_25098_, _25097_, _25096_);
  and _29127_ (_25099_, _25098_, _25095_);
  and _29128_ (_25100_, _25099_, _25094_);
  and _29129_ (_25101_, _25100_, _25092_);
  not _29130_ (_25102_, _25101_);
  and _29131_ (_25103_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _29132_ (_25104_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _29133_ (_25105_, _25104_, _25103_);
  not _29134_ (_25106_, _25056_);
  nor _29135_ (_25107_, _24981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _29136_ (_25108_, _25107_, _25061_);
  and _29137_ (_25109_, _25108_, _25106_);
  and _29138_ (_25110_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _29139_ (_25111_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _29140_ (_25112_, _25111_, _25110_);
  not _29141_ (_25113_, _25112_);
  nor _29142_ (_25114_, _25113_, _25109_);
  and _29143_ (_25115_, _25114_, _25105_);
  not _29144_ (_25116_, _25115_);
  and _29145_ (_25117_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor _29146_ (_25118_, _25117_, _25066_);
  nor _29147_ (_25119_, _25056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _29148_ (_25120_, _25119_, _25061_);
  nor _29149_ (_25121_, _25120_, _25057_);
  and _29150_ (_25122_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _29151_ (_25123_, _25122_, _25121_);
  and _29152_ (_25124_, _25123_, _25118_);
  and _29153_ (_25125_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _29154_ (_25126_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _29155_ (_25127_, _25126_, _25125_);
  and _29156_ (_25128_, _25127_, _25124_);
  nor _29157_ (_25129_, _25128_, _25116_);
  and _29158_ (_25130_, _25129_, _25102_);
  and _29159_ (_25131_, _25130_, _25086_);
  nand _29160_ (_25132_, _25131_, _25055_);
  and _29161_ (_25133_, _24931_, _24487_);
  and _29162_ (_25134_, _24390_, _23920_);
  nor _29163_ (_25135_, _23973_, _24055_);
  and _29164_ (_25136_, _23973_, _24055_);
  nor _29165_ (_25137_, _25136_, _25135_);
  nor _29166_ (_25138_, _24101_, _24018_);
  and _29167_ (_25139_, _24101_, _24018_);
  nor _29168_ (_25140_, _25139_, _25138_);
  and _29169_ (_25141_, _24216_, _24515_);
  nor _29170_ (_25142_, _24216_, _24515_);
  nor _29171_ (_25143_, _25142_, _25141_);
  not _29172_ (_25144_, _25143_);
  and _29173_ (_25145_, _24200_, _24032_);
  not _29174_ (_25146_, _24082_);
  nor _29175_ (_25147_, _24253_, _25146_);
  nor _29176_ (_25148_, _24200_, _24032_);
  nor _29177_ (_25149_, _25148_, _25145_);
  and _29178_ (_25150_, _25149_, _25147_);
  nor _29179_ (_25151_, _25150_, _25145_);
  nor _29180_ (_25152_, _25151_, _25144_);
  nor _29181_ (_25153_, _25152_, _25141_);
  nor _29182_ (_25155_, _25153_, _25140_);
  and _29183_ (_25164_, _25153_, _25140_);
  nor _29184_ (_25165_, _25164_, _25155_);
  nor _29185_ (_25166_, _23960_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _29186_ (_25167_, _25166_);
  nor _29187_ (_25168_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _29188_ (_25169_, _25168_, _23958_);
  and _29189_ (_25170_, _25169_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _29190_ (_25171_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _29191_ (_25172_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25171_);
  nand _29192_ (_25173_, _25172_, _23995_);
  not _29193_ (_25174_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _29194_ (_25175_, _25174_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _29195_ (_25176_, _25175_, _24040_);
  and _29196_ (_25177_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _29197_ (_25178_, _25177_, _23978_);
  and _29198_ (_25179_, _25178_, _25176_);
  and _29199_ (_25180_, _25179_, _25173_);
  nand _29200_ (_25181_, _25180_, _25170_);
  not _29201_ (_25182_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _29202_ (_25183_, _25168_, _24073_);
  and _29203_ (_25184_, _25183_, _25182_);
  nand _29204_ (_25185_, _25177_, _24009_);
  nand _29205_ (_25186_, _25175_, _24059_);
  nand _29206_ (_25187_, _25172_, _24023_);
  and _29207_ (_25188_, _25187_, _25186_);
  and _29208_ (_25189_, _25188_, _25185_);
  nand _29209_ (_25190_, _25189_, _25184_);
  nand _29210_ (_25191_, _25190_, _25181_);
  nand _29211_ (_25192_, _25191_, _23960_);
  and _29212_ (_25193_, _25192_, _25167_);
  and _29213_ (_25194_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _29214_ (_25195_, _25194_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _29215_ (_25196_, _25195_);
  and _29216_ (_25197_, _25196_, _25193_);
  and _29217_ (_25198_, _25196_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _29218_ (_25199_, _25198_, _25197_);
  and _29219_ (_25200_, _24253_, _25146_);
  nor _29220_ (_25201_, _25200_, _25147_);
  not _29221_ (_25202_, _25201_);
  nor _29222_ (_25203_, _25202_, _25199_);
  and _29223_ (_25204_, _25203_, _25149_);
  and _29224_ (_25205_, _25151_, _25144_);
  nor _29225_ (_25206_, _25205_, _25152_);
  and _29226_ (_25207_, _25206_, _25204_);
  not _29227_ (_25208_, _25207_);
  nor _29228_ (_25209_, _25208_, _25165_);
  nor _29229_ (_25210_, _25153_, _25139_);
  or _29230_ (_25211_, _25210_, _25138_);
  or _29231_ (_25212_, _25211_, _25209_);
  and _29232_ (_25213_, _25212_, _25137_);
  and _29233_ (_25214_, _24120_, _24535_);
  nor _29234_ (_25215_, _24120_, _24535_);
  nor _29235_ (_25216_, _25215_, _25214_);
  and _29236_ (_25217_, _25216_, _25135_);
  nor _29237_ (_25218_, _25216_, _25135_);
  nor _29238_ (_25219_, _25218_, _25217_);
  and _29239_ (_25220_, _25219_, _25213_);
  nor _29240_ (_25221_, _24141_, _24616_);
  and _29241_ (_25222_, _24141_, _24616_);
  nor _29242_ (_25223_, _25222_, _25221_);
  not _29243_ (_25224_, _25223_);
  nor _29244_ (_25225_, _25217_, _25214_);
  nor _29245_ (_25226_, _25225_, _25224_);
  and _29246_ (_25227_, _25225_, _25224_);
  nor _29247_ (_25228_, _25227_, _25226_);
  and _29248_ (_25229_, _25228_, _25220_);
  nor _29249_ (_25230_, _25226_, _25221_);
  not _29250_ (_25231_, _25230_);
  nor _29251_ (_25232_, _25231_, _25229_);
  nor _29252_ (_25233_, _24172_, _23990_);
  and _29253_ (_25234_, _24172_, _23990_);
  nor _29254_ (_25235_, _25234_, _25233_);
  not _29255_ (_25236_, _25235_);
  nor _29256_ (_25237_, _25236_, _25232_);
  not _29257_ (_25238_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _29258_ (_25239_, _24468_, _25238_);
  and _29259_ (_25240_, _25239_, _23919_);
  nand _29260_ (_25241_, _25236_, _25232_);
  nand _29261_ (_25242_, _25241_, _25240_);
  nor _29262_ (_25243_, _25242_, _25237_);
  not _29263_ (_25244_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _29264_ (_25245_, _23915_, _25244_);
  and _29265_ (_25246_, _25245_, _23919_);
  not _29266_ (_25247_, _25246_);
  nor _29267_ (_25248_, _24141_, _24049_);
  and _29268_ (_25249_, _24120_, _24004_);
  and _29269_ (_25250_, _23973_, _24520_);
  nor _29270_ (_25251_, _25250_, _25216_);
  nor _29271_ (_25252_, _25251_, _25249_);
  nor _29272_ (_25253_, _25252_, _25223_);
  nor _29273_ (_25254_, _25253_, _25248_);
  and _29274_ (_25255_, _25252_, _25223_);
  nor _29275_ (_25256_, _25255_, _25253_);
  not _29276_ (_25257_, _25256_);
  and _29277_ (_25258_, _25250_, _25216_);
  nor _29278_ (_25259_, _25258_, _25251_);
  not _29279_ (_25260_, _25259_);
  not _29280_ (_25266_, _25137_);
  not _29281_ (_25277_, _25140_);
  and _29282_ (_25288_, _24253_, _24082_);
  nor _29283_ (_25299_, _25288_, _25149_);
  not _29284_ (_25310_, _24032_);
  and _29285_ (_25321_, _24200_, _25310_);
  nor _29286_ (_25323_, _25321_, _25299_);
  nor _29287_ (_25324_, _25323_, _25143_);
  and _29288_ (_25325_, _24216_, _24068_);
  nor _29289_ (_25326_, _25325_, _25324_);
  nor _29290_ (_25327_, _25326_, _25277_);
  and _29291_ (_25328_, _25326_, _25277_);
  nor _29292_ (_25329_, _25328_, _25327_);
  and _29293_ (_25330_, _25323_, _25143_);
  nor _29294_ (_25331_, _25330_, _25324_);
  not _29295_ (_25332_, _25331_);
  and _29296_ (_25333_, _25288_, _25149_);
  nor _29297_ (_25334_, _25333_, _25299_);
  not _29298_ (_25335_, _25334_);
  nor _29299_ (_25336_, _25201_, _25199_);
  and _29300_ (_25337_, _25336_, _25335_);
  and _29301_ (_25338_, _25337_, _25332_);
  and _29302_ (_25339_, _25338_, _25329_);
  or _29303_ (_25340_, _24101_, _24533_);
  and _29304_ (_25341_, _24101_, _24533_);
  or _29305_ (_25342_, _25326_, _25341_);
  and _29306_ (_25343_, _25342_, _25340_);
  or _29307_ (_25344_, _25343_, _25339_);
  and _29308_ (_25345_, _25344_, _25266_);
  and _29309_ (_25346_, _25345_, _25260_);
  and _29310_ (_25347_, _25346_, _25257_);
  nor _29311_ (_25348_, _25347_, _25254_);
  nor _29312_ (_25349_, _25348_, _25235_);
  and _29313_ (_25350_, _25348_, _25235_);
  nor _29314_ (_25351_, _25350_, _25349_);
  nor _29315_ (_25352_, _25351_, _25247_);
  and _29316_ (_25353_, _23918_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _29317_ (_25354_, _25353_, _25245_);
  not _29318_ (_25355_, _24200_);
  nor _29319_ (_25356_, _24253_, _25355_);
  and _29320_ (_25357_, _25356_, _24216_);
  and _29321_ (_25358_, _25357_, _24102_);
  and _29322_ (_25359_, _25358_, _23974_);
  and _29323_ (_25360_, _25359_, _24120_);
  and _29324_ (_25361_, _25360_, _24143_);
  and _29325_ (_25362_, _25361_, _25199_);
  not _29326_ (_25363_, _25199_);
  not _29327_ (_25364_, _24120_);
  and _29328_ (_25365_, _24141_, _25364_);
  nor _29329_ (_25366_, _24216_, _24200_);
  and _29330_ (_25367_, _25366_, _24253_);
  and _29331_ (_25368_, _25367_, _24101_);
  and _29332_ (_25369_, _25368_, _23973_);
  and _29333_ (_25370_, _25369_, _25365_);
  and _29334_ (_25371_, _25370_, _25363_);
  nor _29335_ (_25372_, _25371_, _25362_);
  and _29336_ (_25373_, _25372_, _24172_);
  nor _29337_ (_25374_, _25372_, _24172_);
  nor _29338_ (_25375_, _25374_, _25373_);
  and _29339_ (_25376_, _25375_, _25354_);
  not _29340_ (_25377_, _23990_);
  nor _29341_ (_25378_, _25199_, _25377_);
  not _29342_ (_25379_, _25378_);
  and _29343_ (_25380_, _25199_, _24172_);
  and _29344_ (_25381_, _25353_, _23916_);
  not _29345_ (_25382_, _25381_);
  nor _29346_ (_25383_, _25382_, _25380_);
  and _29347_ (_25384_, _25383_, _25379_);
  nor _29348_ (_25385_, _25384_, _25376_);
  not _29349_ (_25386_, _25365_);
  and _29350_ (_25390_, _25239_, _24482_);
  nor _29351_ (_25394_, _25366_, _24101_);
  and _29352_ (_25395_, _25394_, _25390_);
  and _29353_ (_25396_, _25395_, _23974_);
  nor _29354_ (_25397_, _25396_, _25386_);
  nor _29355_ (_25398_, _25365_, _24172_);
  nor _29356_ (_25399_, _25398_, _25395_);
  and _29357_ (_25400_, _25399_, _25199_);
  nor _29358_ (_25401_, _25400_, _25397_);
  nand _29359_ (_25402_, _25401_, _24278_);
  or _29360_ (_25403_, _25401_, _24278_);
  and _29361_ (_25404_, _25403_, _25390_);
  and _29362_ (_25405_, _25404_, _25402_);
  and _29363_ (_25406_, _25353_, _25239_);
  and _29364_ (_25407_, _25406_, _25363_);
  not _29365_ (_25408_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _29366_ (_25409_, _23918_, _25408_);
  and _29367_ (_25410_, _25409_, _25239_);
  not _29368_ (_25411_, _25410_);
  nor _29369_ (_25412_, _25411_, _25234_);
  and _29370_ (_25413_, _25409_, _24469_);
  and _29371_ (_25414_, _25413_, _25235_);
  nor _29372_ (_25415_, _25414_, _25412_);
  and _29373_ (_25416_, _24482_, _23916_);
  and _29374_ (_25417_, _25416_, _25233_);
  and _29375_ (_25418_, _25245_, _24482_);
  and _29376_ (_25419_, _25418_, _24172_);
  nor _29377_ (_25420_, _25419_, _25417_);
  and _29378_ (_25421_, _25353_, _24469_);
  and _29379_ (_25422_, _25421_, _24254_);
  and _29380_ (_25423_, _24469_, _23919_);
  not _29381_ (_25424_, _25423_);
  nor _29382_ (_25425_, _25424_, _24172_);
  and _29383_ (_25426_, _25409_, _23915_);
  not _29384_ (_25427_, _25426_);
  nor _29385_ (_25428_, _25427_, _24141_);
  or _29386_ (_25429_, _25428_, _25425_);
  nor _29387_ (_25430_, _25429_, _25422_);
  and _29388_ (_25431_, _25430_, _25420_);
  nand _29389_ (_25432_, _25431_, _25415_);
  or _29390_ (_25433_, _25432_, _25407_);
  nor _29391_ (_25434_, _25433_, _25405_);
  nand _29392_ (_25435_, _25434_, _25385_);
  or _29393_ (_25437_, _25435_, _25352_);
  or _29394_ (_25438_, _25437_, _25243_);
  or _29395_ (_25440_, _25438_, _25134_);
  or _29396_ (_25441_, _25440_, _25133_);
  or _29397_ (_25443_, _25441_, _25132_);
  not _29398_ (_25444_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _29399_ (_25446_, \oc8051_top_1.oc8051_decoder1.wr , _23914_);
  not _29400_ (_25447_, _25446_);
  nor _29401_ (_25449_, _25447_, _24988_);
  and _29402_ (_25450_, _25449_, _25444_);
  not _29403_ (_25452_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _29404_ (_25453_, _25132_, _25452_);
  and _29405_ (_25455_, _25453_, _25450_);
  and _29406_ (_25456_, _25455_, _25443_);
  nor _29407_ (_25458_, _25449_, _25452_);
  not _29408_ (_25459_, _25240_);
  nor _29409_ (_25461_, _25237_, _25233_);
  nor _29410_ (_25462_, _25461_, _25459_);
  not _29411_ (_25464_, _25462_);
  and _29412_ (_25465_, _24172_, _25377_);
  nor _29413_ (_25466_, _25465_, _25349_);
  nor _29414_ (_25467_, _25466_, _25247_);
  and _29415_ (_25468_, _25397_, _25199_);
  nor _29416_ (_25469_, _25468_, _25380_);
  not _29417_ (_25470_, _25390_);
  not _29418_ (_25471_, _25397_);
  nor _29419_ (_25472_, _25199_, _24172_);
  and _29420_ (_25473_, _25472_, _25471_);
  nor _29421_ (_25474_, _25473_, _25470_);
  and _29422_ (_25475_, _25474_, _25469_);
  and _29423_ (_25476_, _25195_, _25193_);
  and _29424_ (_25477_, _25409_, _25245_);
  and _29425_ (_25478_, _25416_, _25193_);
  nor _29426_ (_25479_, _25478_, _25477_);
  nor _29427_ (_25480_, _25479_, _25476_);
  nor _29428_ (_25481_, _25199_, _25193_);
  and _29429_ (_25482_, _25481_, _25421_);
  and _29430_ (_25483_, _25418_, _25199_);
  or _29431_ (_25484_, _25483_, _25482_);
  nor _29432_ (_25491_, _25198_, _25193_);
  not _29433_ (_25496_, _25413_);
  nor _29434_ (_25497_, _25496_, _25197_);
  nor _29435_ (_25498_, _25497_, _25410_);
  nor _29436_ (_25499_, _25498_, _25491_);
  nor _29437_ (_25500_, _25424_, _25199_);
  and _29438_ (_25501_, _25409_, _23916_);
  not _29439_ (_25502_, _25501_);
  nor _29440_ (_25503_, _25502_, _24172_);
  and _29441_ (_25504_, _25406_, _24254_);
  or _29442_ (_25505_, _25504_, _25395_);
  or _29443_ (_25506_, _25505_, _25503_);
  or _29444_ (_25507_, _25506_, _25500_);
  or _29445_ (_25508_, _25507_, _25499_);
  or _29446_ (_25509_, _25508_, _25484_);
  or _29447_ (_25510_, _25509_, _25480_);
  nor _29448_ (_25511_, _25510_, _25475_);
  not _29449_ (_25512_, _25511_);
  nor _29450_ (_25513_, _25512_, _25467_);
  and _29451_ (_25514_, _25513_, _25464_);
  not _29452_ (_25515_, _25020_);
  nor _29453_ (_25516_, _25053_, _25042_);
  and _29454_ (_25517_, _25516_, _25515_);
  and _29455_ (_25518_, _25517_, _25131_);
  nand _29456_ (_25519_, _25518_, _25514_);
  or _29457_ (_25520_, _25518_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _29458_ (_25521_, _25449_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _29459_ (_25522_, _25521_, _25520_);
  and _29460_ (_25523_, _25522_, _25519_);
  or _29461_ (_25524_, _25523_, _25458_);
  or _29462_ (_25525_, _25524_, _25456_);
  and _29463_ (_06524_, _25525_, _27355_);
  nand _29464_ (_25526_, _24937_, _24487_);
  and _29465_ (_25527_, _24448_, _23920_);
  and _29466_ (_25528_, _25202_, _25199_);
  nor _29467_ (_25529_, _25528_, _25203_);
  not _29468_ (_25530_, _25529_);
  nor _29469_ (_25531_, _25246_, _25240_);
  nor _29470_ (_25532_, _25531_, _25530_);
  nor _29471_ (_25533_, _25502_, _25199_);
  not _29472_ (_25534_, _25533_);
  and _29473_ (_25535_, _25413_, _25201_);
  not _29474_ (_25536_, _25535_);
  nor _29475_ (_25537_, _25411_, _25200_);
  not _29476_ (_25538_, _25537_);
  and _29477_ (_25539_, _25416_, _25147_);
  and _29478_ (_25540_, _25418_, _24253_);
  nor _29479_ (_25541_, _25540_, _25539_);
  and _29480_ (_25542_, _25541_, _25538_);
  and _29481_ (_25543_, _25542_, _25536_);
  and _29482_ (_25544_, _25381_, _24082_);
  and _29483_ (_25545_, _25354_, _24253_);
  nor _29484_ (_25546_, _25545_, _25544_);
  and _29485_ (_25547_, _25477_, _24278_);
  not _29486_ (_25548_, _25547_);
  and _29487_ (_25549_, _25353_, _25238_);
  and _29488_ (_25550_, _25549_, _24200_);
  nor _29489_ (_25551_, _25423_, _25390_);
  nor _29490_ (_25552_, _25551_, _24253_);
  nor _29491_ (_25553_, _25552_, _25550_);
  and _29492_ (_25554_, _25553_, _25548_);
  and _29493_ (_25555_, _25554_, _25546_);
  and _29494_ (_25556_, _25555_, _25543_);
  and _29495_ (_25557_, _25556_, _25534_);
  not _29496_ (_25558_, _25557_);
  nor _29497_ (_25559_, _25558_, _25532_);
  not _29498_ (_25560_, _25559_);
  nor _29499_ (_25561_, _25560_, _25527_);
  and _29500_ (_25562_, _25561_, _25526_);
  not _29501_ (_25563_, _25562_);
  or _29502_ (_25564_, _25563_, _25132_);
  not _29503_ (_25565_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _29504_ (_25566_, _25132_, _25565_);
  and _29505_ (_25570_, _25566_, _25450_);
  and _29506_ (_25572_, _25570_, _25564_);
  nor _29507_ (_25573_, _25449_, _25565_);
  not _29508_ (_25574_, _25514_);
  or _29509_ (_25575_, _25574_, _25132_);
  and _29510_ (_25576_, _25566_, _25521_);
  and _29511_ (_25577_, _25576_, _25575_);
  or _29512_ (_25578_, _25577_, _25573_);
  or _29513_ (_25579_, _25578_, _25572_);
  and _29514_ (_08841_, _25579_, _27355_);
  nand _29515_ (_25580_, _24944_, _24487_);
  nor _29516_ (_25581_, _25394_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _29517_ (_25582_, _25581_, _24200_);
  nor _29518_ (_25583_, _25581_, _24200_);
  nor _29519_ (_25584_, _25583_, _25582_);
  nor _29520_ (_25585_, _25584_, _25470_);
  not _29521_ (_25595_, _25585_);
  nor _29522_ (_25596_, _25427_, _24253_);
  and _29523_ (_25597_, _25423_, _24200_);
  and _29524_ (_25598_, _25549_, _24216_);
  or _29525_ (_25599_, _25598_, _25597_);
  nor _29526_ (_25600_, _25599_, _25596_);
  and _29527_ (_25601_, _25413_, _25149_);
  nor _29528_ (_25602_, _25411_, _25148_);
  not _29529_ (_25603_, _25602_);
  and _29530_ (_25604_, _25416_, _25145_);
  and _29531_ (_25605_, _25418_, _25355_);
  nor _29532_ (_25606_, _25605_, _25604_);
  nand _29533_ (_25607_, _25606_, _25603_);
  nor _29534_ (_25608_, _25607_, _25601_);
  and _29535_ (_25609_, _25608_, _25600_);
  and _29536_ (_25610_, _25609_, _25595_);
  nor _29537_ (_25611_, _25149_, _25147_);
  or _29538_ (_25612_, _25611_, _25150_);
  and _29539_ (_25613_, _25612_, _25203_);
  nor _29540_ (_25614_, _25612_, _25203_);
  or _29541_ (_25615_, _25614_, _25613_);
  and _29542_ (_25616_, _25615_, _25240_);
  nor _29543_ (_25617_, _25336_, _25335_);
  nor _29544_ (_25619_, _25617_, _25337_);
  nor _29545_ (_25620_, _25619_, _25247_);
  nor _29546_ (_25621_, _25620_, _25616_);
  and _29547_ (_25623_, _25621_, _25610_);
  nand _29548_ (_25624_, _24452_, _23920_);
  and _29549_ (_25626_, _25381_, _24032_);
  not _29550_ (_25627_, _25626_);
  and _29551_ (_25628_, _24253_, _25355_);
  nor _29552_ (_25630_, _25628_, _25356_);
  and _29553_ (_25631_, _25630_, _25363_);
  or _29554_ (_25632_, _25630_, _25363_);
  nand _29555_ (_25633_, _25632_, _25354_);
  or _29556_ (_25635_, _25633_, _25631_);
  and _29557_ (_25636_, _25635_, _25627_);
  and _29558_ (_25637_, _25636_, _25624_);
  and _29559_ (_25638_, _25637_, _25623_);
  nand _29560_ (_25639_, _25638_, _25580_);
  or _29561_ (_25641_, _25639_, _25132_);
  not _29562_ (_25642_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _29563_ (_25643_, _25132_, _25642_);
  and _29564_ (_25644_, _25643_, _25450_);
  and _29565_ (_25645_, _25644_, _25641_);
  nor _29566_ (_25646_, _25449_, _25642_);
  nand _29567_ (_25648_, _25131_, _25020_);
  not _29568_ (_25649_, _25053_);
  and _29569_ (_25650_, _25649_, _25042_);
  not _29570_ (_25651_, _25650_);
  nor _29571_ (_25652_, _25651_, _25648_);
  nand _29572_ (_25653_, _25652_, _25514_);
  or _29573_ (_25654_, _25652_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _29574_ (_25656_, _25654_, _25521_);
  and _29575_ (_25657_, _25656_, _25653_);
  or _29576_ (_25658_, _25657_, _25646_);
  or _29577_ (_25659_, _25658_, _25645_);
  and _29578_ (_08853_, _25659_, _27355_);
  nand _29579_ (_25660_, _24456_, _23920_);
  nand _29580_ (_25661_, _24950_, _24487_);
  and _29581_ (_25662_, _25381_, _24515_);
  not _29582_ (_25664_, _24216_);
  nand _29583_ (_25665_, _25356_, _25199_);
  nand _29584_ (_25666_, _25628_, _25363_);
  and _29585_ (_25667_, _25666_, _25665_);
  nand _29586_ (_25668_, _25667_, _25664_);
  or _29587_ (_25669_, _25667_, _25664_);
  and _29588_ (_25670_, _25669_, _25668_);
  and _29589_ (_25671_, _25670_, _25354_);
  nor _29590_ (_25672_, _25671_, _25662_);
  nor _29591_ (_25674_, _25337_, _25332_);
  nor _29592_ (_25675_, _25674_, _25338_);
  nor _29593_ (_25676_, _25675_, _25247_);
  not _29594_ (_25677_, _25676_);
  and _29595_ (_25678_, _25549_, _24102_);
  and _29596_ (_25679_, _25416_, _25141_);
  and _29597_ (_25680_, _25418_, _25664_);
  nor _29598_ (_25681_, _25680_, _25679_);
  nor _29599_ (_25682_, _25411_, _25142_);
  and _29600_ (_25684_, _25413_, _25143_);
  nor _29601_ (_25685_, _25684_, _25682_);
  and _29602_ (_25686_, _25423_, _24216_);
  and _29603_ (_25687_, _25426_, _24200_);
  nor _29604_ (_25688_, _25687_, _25686_);
  and _29605_ (_25689_, _25688_, _25685_);
  nand _29606_ (_25690_, _25689_, _25681_);
  nor _29607_ (_25691_, _25690_, _25678_);
  and _29608_ (_25692_, _25691_, _25677_);
  nor _29609_ (_25693_, _25206_, _25204_);
  nor _29610_ (_25694_, _25693_, _25459_);
  and _29611_ (_25695_, _25694_, _25208_);
  nor _29612_ (_25696_, _25583_, _25664_);
  and _29613_ (_25697_, _25366_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _29614_ (_25698_, _25697_, _25696_);
  nor _29615_ (_25699_, _25698_, _25470_);
  nor _29616_ (_25700_, _25699_, _25695_);
  and _29617_ (_25701_, _25700_, _25692_);
  and _29618_ (_25702_, _25701_, _25672_);
  and _29619_ (_25703_, _25702_, _25661_);
  and _29620_ (_25704_, _25703_, _25660_);
  not _29621_ (_25705_, _25704_);
  or _29622_ (_25706_, _25705_, _25132_);
  not _29623_ (_25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _29624_ (_25708_, _25132_, _25707_);
  and _29625_ (_25709_, _25708_, _25450_);
  and _29626_ (_25710_, _25709_, _25706_);
  nor _29627_ (_25711_, _25449_, _25707_);
  or _29628_ (_25712_, _25516_, _25648_);
  and _29629_ (_25713_, _25712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _29630_ (_25714_, _25042_);
  and _29631_ (_25715_, _25020_, _25053_);
  and _29632_ (_25716_, _25715_, _25714_);
  not _29633_ (_25717_, _25716_);
  nor _29634_ (_25718_, _25717_, _25514_);
  nand _29635_ (_25719_, _25020_, _25042_);
  nor _29636_ (_25720_, _25719_, _25707_);
  or _29637_ (_25721_, _25720_, _25718_);
  and _29638_ (_25722_, _25721_, _25131_);
  or _29639_ (_25723_, _25722_, _25713_);
  and _29640_ (_25724_, _25723_, _25521_);
  or _29641_ (_25725_, _25724_, _25711_);
  or _29642_ (_25726_, _25725_, _25710_);
  and _29643_ (_08864_, _25726_, _27355_);
  nand _29644_ (_25727_, _24460_, _23920_);
  nand _29645_ (_25728_, _24958_, _24487_);
  and _29646_ (_25729_, _25381_, _24533_);
  nand _29647_ (_25730_, _25357_, _25199_);
  nand _29648_ (_25731_, _25367_, _25363_);
  nand _29649_ (_25732_, _25731_, _25730_);
  and _29650_ (_25733_, _25732_, _24102_);
  or _29651_ (_25734_, _25732_, _24102_);
  nand _29652_ (_25735_, _25734_, _25354_);
  nor _29653_ (_25736_, _25735_, _25733_);
  nor _29654_ (_25737_, _25736_, _25729_);
  not _29655_ (_25738_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _29656_ (_25739_, _25366_, _25738_);
  nor _29657_ (_25740_, _25739_, _24102_);
  or _29658_ (_25741_, _25740_, _25470_);
  nor _29659_ (_25742_, _25741_, _25394_);
  not _29660_ (_25743_, _25742_);
  nor _29661_ (_25744_, _25411_, _25139_);
  and _29662_ (_25745_, _25413_, _25140_);
  nor _29663_ (_25746_, _25745_, _25744_);
  and _29664_ (_25747_, _25416_, _25138_);
  and _29665_ (_25748_, _25418_, _24101_);
  nor _29666_ (_25749_, _25748_, _25747_);
  and _29667_ (_25750_, _25549_, _23974_);
  not _29668_ (_25751_, _25750_);
  nor _29669_ (_25752_, _25424_, _24101_);
  and _29670_ (_25753_, _25426_, _24216_);
  nor _29671_ (_25754_, _25753_, _25752_);
  and _29672_ (_25755_, _25754_, _25751_);
  and _29673_ (_25756_, _25755_, _25749_);
  and _29674_ (_25757_, _25756_, _25746_);
  and _29675_ (_25758_, _25757_, _25743_);
  nor _29676_ (_25759_, _25338_, _25329_);
  nor _29677_ (_25760_, _25759_, _25339_);
  nor _29678_ (_25761_, _25760_, _25247_);
  and _29679_ (_25762_, _25208_, _25165_);
  or _29680_ (_25763_, _25762_, _25459_);
  nor _29681_ (_25764_, _25763_, _25209_);
  nor _29682_ (_25765_, _25764_, _25761_);
  and _29683_ (_25766_, _25765_, _25758_);
  and _29684_ (_25767_, _25766_, _25737_);
  and _29685_ (_25768_, _25767_, _25728_);
  and _29686_ (_25769_, _25768_, _25727_);
  not _29687_ (_25770_, _25769_);
  or _29688_ (_25771_, _25770_, _25132_);
  not _29689_ (_25772_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _29690_ (_25773_, _25132_, _25772_);
  and _29691_ (_25774_, _25773_, _25450_);
  and _29692_ (_25775_, _25774_, _25771_);
  nor _29693_ (_25776_, _25449_, _25772_);
  and _29694_ (_25777_, _25648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _29695_ (_25778_, _25516_, _25020_);
  and _29696_ (_25779_, _25778_, _25574_);
  or _29697_ (_25780_, _25516_, _25515_);
  nor _29698_ (_25781_, _25780_, _25772_);
  or _29699_ (_25782_, _25781_, _25779_);
  and _29700_ (_25783_, _25782_, _25131_);
  or _29701_ (_25784_, _25783_, _25777_);
  and _29702_ (_25785_, _25784_, _25521_);
  or _29703_ (_25786_, _25785_, _25776_);
  or _29704_ (_25787_, _25786_, _25775_);
  and _29705_ (_08876_, _25787_, _27355_);
  and _29706_ (_25788_, _24963_, _24487_);
  and _29707_ (_25789_, _24463_, _23920_);
  nor _29708_ (_25790_, _25344_, _25137_);
  and _29709_ (_25791_, _25344_, _25137_);
  nor _29710_ (_25792_, _25791_, _25790_);
  and _29711_ (_25793_, _25792_, _25246_);
  or _29712_ (_25794_, _25212_, _25137_);
  nor _29713_ (_25795_, _25459_, _25213_);
  and _29714_ (_25796_, _25795_, _25794_);
  nor _29715_ (_25797_, _25199_, _24055_);
  and _29716_ (_25798_, _25199_, _23974_);
  nor _29717_ (_25799_, _25798_, _25797_);
  nor _29718_ (_25800_, _25799_, _25382_);
  and _29719_ (_25801_, _25358_, _25199_);
  and _29720_ (_25802_, _25368_, _25363_);
  nor _29721_ (_25803_, _25802_, _25801_);
  and _29722_ (_25804_, _25803_, _23973_);
  nor _29723_ (_25805_, _25803_, _23973_);
  nor _29724_ (_25806_, _25805_, _25804_);
  and _29725_ (_25807_, _25806_, _25354_);
  nor _29726_ (_25808_, _25807_, _25800_);
  or _29727_ (_25809_, _25395_, _23974_);
  nor _29728_ (_25810_, _25424_, _23973_);
  nor _29729_ (_25811_, _25396_, _25470_);
  or _29730_ (_25812_, _25811_, _25810_);
  and _29731_ (_25813_, _25812_, _25809_);
  and _29732_ (_25814_, _25413_, _25137_);
  and _29733_ (_25815_, _25416_, _25135_);
  nor _29734_ (_25816_, _25411_, _25136_);
  and _29735_ (_25817_, _25418_, _23973_);
  or _29736_ (_25818_, _25817_, _25816_);
  or _29737_ (_25819_, _25818_, _25815_);
  nor _29738_ (_25820_, _25819_, _25814_);
  and _29739_ (_25821_, _25549_, _24120_);
  nor _29740_ (_25822_, _25427_, _24101_);
  nor _29741_ (_25823_, _25822_, _25821_);
  nand _29742_ (_25824_, _25823_, _25820_);
  nor _29743_ (_25825_, _25824_, _25813_);
  nand _29744_ (_25826_, _25825_, _25808_);
  or _29745_ (_25827_, _25826_, _25796_);
  or _29746_ (_25828_, _25827_, _25793_);
  or _29747_ (_25829_, _25828_, _25789_);
  or _29748_ (_25830_, _25829_, _25788_);
  or _29749_ (_25831_, _25830_, _25132_);
  not _29750_ (_25832_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _29751_ (_25833_, _25132_, _25832_);
  and _29752_ (_25834_, _25833_, _25450_);
  and _29753_ (_25835_, _25834_, _25831_);
  nor _29754_ (_25836_, _25449_, _25832_);
  not _29755_ (_25837_, _25131_);
  and _29756_ (_25838_, _25054_, _25515_);
  nor _29757_ (_25839_, _25054_, _25515_);
  nor _29758_ (_25840_, _25839_, _25838_);
  or _29759_ (_25841_, _25840_, _25837_);
  and _29760_ (_25842_, _25841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _29761_ (_25843_, _25838_, _25574_);
  and _29762_ (_25844_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _29763_ (_25845_, _25844_, _25843_);
  and _29764_ (_25846_, _25845_, _25131_);
  or _29765_ (_25847_, _25846_, _25842_);
  and _29766_ (_25848_, _25847_, _25521_);
  or _29767_ (_25849_, _25848_, _25836_);
  or _29768_ (_25850_, _25849_, _25835_);
  and _29769_ (_08887_, _25850_, _27355_);
  and _29770_ (_25851_, _24970_, _24487_);
  and _29771_ (_25852_, _24465_, _23920_);
  or _29772_ (_25853_, _25219_, _25213_);
  nor _29773_ (_25854_, _25459_, _25220_);
  and _29774_ (_25855_, _25854_, _25853_);
  nor _29775_ (_25856_, _25345_, _25260_);
  nor _29776_ (_25857_, _25856_, _25346_);
  nor _29777_ (_25858_, _25857_, _25247_);
  nor _29778_ (_25859_, _25199_, _24004_);
  and _29779_ (_25860_, _25199_, _24120_);
  nor _29780_ (_25861_, _25860_, _25859_);
  nor _29781_ (_25862_, _25861_, _25382_);
  and _29782_ (_25863_, _25359_, _25199_);
  and _29783_ (_25864_, _25369_, _25363_);
  nor _29784_ (_25865_, _25864_, _25863_);
  and _29785_ (_25866_, _25865_, _25364_);
  not _29786_ (_25867_, _25354_);
  nor _29787_ (_25868_, _25865_, _25364_);
  or _29788_ (_25869_, _25868_, _25867_);
  nor _29789_ (_25870_, _25869_, _25866_);
  nor _29790_ (_25871_, _25870_, _25862_);
  nor _29791_ (_25872_, _25396_, _24120_);
  not _29792_ (_25873_, _25400_);
  and _29793_ (_25874_, _25873_, _25872_);
  or _29794_ (_25875_, _25400_, _25396_);
  and _29795_ (_25876_, _25875_, _24120_);
  or _29796_ (_25877_, _25876_, _25874_);
  and _29797_ (_25878_, _25877_, _25390_);
  and _29798_ (_25879_, _25413_, _25216_);
  nor _29799_ (_25880_, _25411_, _25215_);
  not _29800_ (_25881_, _25880_);
  and _29801_ (_25882_, _25416_, _25214_);
  and _29802_ (_25883_, _25418_, _25364_);
  nor _29803_ (_25884_, _25883_, _25882_);
  nand _29804_ (_25885_, _25884_, _25881_);
  nor _29805_ (_25886_, _25885_, _25879_);
  and _29806_ (_25887_, _25549_, _24143_);
  and _29807_ (_25888_, _25423_, _24120_);
  nor _29808_ (_25889_, _25427_, _23973_);
  or _29809_ (_25890_, _25889_, _25888_);
  nor _29810_ (_25891_, _25890_, _25887_);
  nand _29811_ (_25892_, _25891_, _25886_);
  nor _29812_ (_25893_, _25892_, _25878_);
  nand _29813_ (_25894_, _25893_, _25871_);
  or _29814_ (_25895_, _25894_, _25858_);
  or _29815_ (_25896_, _25895_, _25855_);
  or _29816_ (_25897_, _25896_, _25852_);
  or _29817_ (_25898_, _25897_, _25851_);
  or _29818_ (_25899_, _25898_, _25132_);
  not _29819_ (_25900_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _29820_ (_25901_, _25132_, _25900_);
  and _29821_ (_25902_, _25901_, _25450_);
  and _29822_ (_25903_, _25902_, _25899_);
  nor _29823_ (_25904_, _25449_, _25900_);
  and _29824_ (_25905_, _25650_, _25515_);
  and _29825_ (_25906_, _25905_, _25131_);
  nand _29826_ (_25907_, _25906_, _25514_);
  or _29827_ (_25908_, _25906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _29828_ (_25909_, _25908_, _25521_);
  and _29829_ (_25910_, _25909_, _25907_);
  or _29830_ (_25911_, _25910_, _25904_);
  or _29831_ (_25912_, _25911_, _25903_);
  and _29832_ (_08898_, _25912_, _27355_);
  not _29833_ (_25913_, _24487_);
  or _29834_ (_25914_, _24975_, _25913_);
  not _29835_ (_25915_, _23920_);
  or _29836_ (_25916_, _24467_, _25915_);
  nor _29837_ (_25917_, _25346_, _25257_);
  nor _29838_ (_25918_, _25917_, _25347_);
  nor _29839_ (_25919_, _25918_, _25247_);
  not _29840_ (_25920_, _25919_);
  nor _29841_ (_25921_, _25228_, _25220_);
  not _29842_ (_25922_, _25921_);
  nor _29843_ (_25923_, _25459_, _25229_);
  and _29844_ (_25924_, _25923_, _25922_);
  and _29845_ (_25925_, _25199_, _24143_);
  nor _29846_ (_25926_, _25199_, _24616_);
  or _29847_ (_25927_, _25926_, _25925_);
  and _29848_ (_25928_, _25927_, _25381_);
  or _29849_ (_25929_, _25199_, _25364_);
  or _29850_ (_25930_, _25864_, _25360_);
  and _29851_ (_25931_, _25930_, _25929_);
  nor _29852_ (_25932_, _25931_, _24143_);
  and _29853_ (_25933_, _25931_, _24143_);
  or _29854_ (_25934_, _25933_, _25867_);
  nor _29855_ (_25935_, _25934_, _25932_);
  nor _29856_ (_25936_, _25935_, _25928_);
  nor _29857_ (_25937_, _25874_, _24141_);
  and _29858_ (_25938_, _25874_, _24141_);
  nor _29859_ (_25939_, _25938_, _25937_);
  nor _29860_ (_25940_, _25939_, _25470_);
  nor _29861_ (_25941_, _25424_, _24141_);
  not _29862_ (_25942_, _25941_);
  and _29863_ (_25943_, _25549_, _24278_);
  and _29864_ (_25944_, _25426_, _24120_);
  nor _29865_ (_25945_, _25944_, _25943_);
  and _29866_ (_25946_, _25945_, _25942_);
  and _29867_ (_25947_, _25413_, _25223_);
  nor _29868_ (_25948_, _25411_, _25222_);
  not _29869_ (_25949_, _25948_);
  and _29870_ (_25950_, _25416_, _25221_);
  and _29871_ (_25951_, _25418_, _24141_);
  nor _29872_ (_25952_, _25951_, _25950_);
  nand _29873_ (_25953_, _25952_, _25949_);
  nor _29874_ (_25954_, _25953_, _25947_);
  and _29875_ (_25955_, _25954_, _25946_);
  not _29876_ (_25956_, _25955_);
  nor _29877_ (_25957_, _25956_, _25940_);
  and _29878_ (_25958_, _25957_, _25936_);
  not _29879_ (_25959_, _25958_);
  nor _29880_ (_25960_, _25959_, _25924_);
  and _29881_ (_25961_, _25960_, _25920_);
  and _29882_ (_25962_, _25961_, _25916_);
  and _29883_ (_25963_, _25962_, _25914_);
  not _29884_ (_25964_, _25963_);
  or _29885_ (_25965_, _25964_, _25132_);
  not _29886_ (_25966_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _29887_ (_25967_, _25132_, _25966_);
  and _29888_ (_25968_, _25967_, _25450_);
  and _29889_ (_25969_, _25968_, _25965_);
  nor _29890_ (_25970_, _25449_, _25966_);
  nor _29891_ (_25971_, _25020_, _25042_);
  and _29892_ (_25972_, _25971_, _25053_);
  and _29893_ (_25973_, _25972_, _25131_);
  nand _29894_ (_25974_, _25973_, _25514_);
  or _29895_ (_25975_, _25973_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _29896_ (_25976_, _25975_, _25521_);
  and _29897_ (_25977_, _25976_, _25974_);
  or _29898_ (_25978_, _25977_, _25970_);
  or _29899_ (_25979_, _25978_, _25969_);
  and _29900_ (_08909_, _25979_, _27355_);
  and _29901_ (_25980_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29902_ (_25981_, _25980_);
  nor _29903_ (_25982_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _29904_ (_25983_, _25982_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29905_ (_25984_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _29906_ (_25985_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _29907_ (_25986_, _25985_, _25984_);
  and _29908_ (_25987_, _25982_, _23914_);
  and _29909_ (_25988_, _25987_, _25986_);
  and _29910_ (_25989_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _29911_ (_25990_, _25989_);
  not _29912_ (_25991_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _29913_ (_25992_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _29914_ (_25993_, _25992_);
  not _29915_ (_25994_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand _29916_ (_25995_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _29917_ (_25996_, _25995_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or _29918_ (_25997_, _25996_, _25994_);
  not _29919_ (_25998_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not _29920_ (_25999_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _29921_ (_26000_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _29922_ (_26001_, _26000_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _29923_ (_26002_, _26001_, _25999_);
  or _29924_ (_26003_, _26002_, _25998_);
  and _29925_ (_26004_, _26003_, _25997_);
  or _29926_ (_26005_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _29927_ (_26006_, _26005_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _29928_ (_26007_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  not _29929_ (_26008_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _29930_ (_26009_, _26005_, _25999_);
  or _29931_ (_26010_, _26009_, _26008_);
  and _29932_ (_26011_, _26010_, _26007_);
  nor _29933_ (_26012_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _29934_ (_26013_, _26012_, _25999_);
  nand _29935_ (_26014_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _29936_ (_26015_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not _29937_ (_26016_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _29938_ (_26017_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26016_);
  nand _29939_ (_26018_, _26017_, _25999_);
  or _29940_ (_26019_, _26018_, _26015_);
  and _29941_ (_26020_, _26019_, _26014_);
  and _29942_ (_26021_, _26020_, _26011_);
  nand _29943_ (_26022_, _26021_, _26004_);
  nand _29944_ (_26023_, _26022_, _25993_);
  nand _29945_ (_26024_, _26023_, _25991_);
  nor _29946_ (_26025_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _25991_);
  nor _29947_ (_26026_, _26025_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _29948_ (_26027_, _26026_, _26024_);
  and _29949_ (_26028_, _26027_, _25990_);
  nand _29950_ (_26029_, _26028_, _25988_);
  not _29951_ (_26030_, _25986_);
  nor _29952_ (_26031_, _25987_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _29953_ (_26032_, _26031_, _26030_);
  and _29954_ (_26033_, _26032_, _26029_);
  not _29955_ (_26034_, _26033_);
  not _29956_ (_26035_, _25988_);
  and _29957_ (_26036_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _29958_ (_26037_, _26036_);
  not _29959_ (_26038_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _29960_ (_26039_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand _29961_ (_26041_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not _29962_ (_26043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _29963_ (_26045_, _26018_, _26043_);
  and _29964_ (_26047_, _26045_, _26041_);
  nand _29965_ (_26049_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not _29966_ (_26051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _29967_ (_26053_, _26009_, _26051_);
  and _29968_ (_26055_, _26053_, _26049_);
  not _29969_ (_26057_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _29970_ (_26059_, _25996_, _26057_);
  not _29971_ (_26061_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _29972_ (_26063_, _26002_, _26061_);
  and _29973_ (_26065_, _26063_, _26059_);
  and _29974_ (_26067_, _26065_, _26055_);
  nand _29975_ (_26069_, _26067_, _26047_);
  nand _29976_ (_26071_, _26069_, _25993_);
  nor _29977_ (_26073_, _26071_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _29978_ (_26075_, _26073_, _26039_);
  nand _29979_ (_26077_, _26075_, _26038_);
  nand _29980_ (_26079_, _26077_, _26037_);
  or _29981_ (_26081_, _26079_, _26035_);
  nor _29982_ (_26083_, _25987_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _29983_ (_26085_, _26083_, _26030_);
  nand _29984_ (_26087_, _26085_, _26081_);
  and _29985_ (_26089_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _29986_ (_26091_, _26089_);
  not _29987_ (_26093_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _29988_ (_26095_, _26002_, _26093_);
  not _29989_ (_26097_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _29990_ (_26099_, _26018_, _26097_);
  and _29991_ (_26101_, _26099_, _26095_);
  nand _29992_ (_26103_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not _29993_ (_26105_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _29994_ (_26107_, _26009_, _26105_);
  and _29995_ (_26109_, _26107_, _26103_);
  nand _29996_ (_26110_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not _29997_ (_26111_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _29998_ (_26112_, _25996_, _26111_);
  and _29999_ (_26113_, _26112_, _26110_);
  and _30000_ (_26114_, _26113_, _26109_);
  and _30001_ (_26115_, _26114_, _26101_);
  or _30002_ (_26116_, _26115_, _25992_);
  nand _30003_ (_26117_, _26116_, _25991_);
  nor _30004_ (_26118_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _25991_);
  nor _30005_ (_26119_, _26118_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _30006_ (_26120_, _26119_, _26117_);
  and _30007_ (_26121_, _26120_, _26091_);
  nand _30008_ (_26122_, _26121_, _25988_);
  nor _30009_ (_26123_, _25987_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _30010_ (_26124_, _26123_, _26030_);
  and _30011_ (_26125_, _26124_, _26122_);
  not _30012_ (_26126_, _26125_);
  not _30013_ (_26127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _30014_ (_26128_, _26009_, _26127_);
  not _30015_ (_26129_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _30016_ (_26130_, _25996_, _26129_);
  and _30017_ (_26131_, _26130_, _26128_);
  not _30018_ (_26132_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _30019_ (_26133_, _26018_, _26132_);
  and _30020_ (_26134_, _26133_, _26131_);
  not _30021_ (_26135_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _30022_ (_26136_, _26002_, _26135_);
  and _30023_ (_26137_, _26136_, _25993_);
  nand _30024_ (_26138_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _30025_ (_26139_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _30026_ (_26140_, _26139_, _26138_);
  and _30027_ (_26141_, _26140_, _26137_);
  nand _30028_ (_26142_, _26141_, _26134_);
  nor _30029_ (_26143_, _26142_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _30030_ (_26144_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _25991_);
  or _30031_ (_26145_, _26144_, _26143_);
  nand _30032_ (_26146_, _26145_, _26038_);
  nor _30033_ (_26147_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _26038_);
  not _30034_ (_26148_, _26147_);
  and _30035_ (_26149_, _26148_, _26146_);
  or _30036_ (_26150_, _26149_, _26035_);
  nor _30037_ (_26151_, _25987_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _30038_ (_26152_, _26151_, _26030_);
  and _30039_ (_26153_, _26152_, _26150_);
  and _30040_ (_26154_, _26153_, _26126_);
  and _30041_ (_26155_, _26154_, _26087_);
  and _30042_ (_26156_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not _30043_ (_26157_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _30044_ (_26158_, _26009_, _26157_);
  not _30045_ (_26159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _30046_ (_26160_, _25996_, _26159_);
  nand _30047_ (_26161_, _26160_, _26158_);
  nor _30048_ (_26162_, _26161_, _26156_);
  not _30049_ (_26163_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _30050_ (_26164_, _26002_, _26163_);
  and _30051_ (_26165_, _26164_, _25993_);
  nand _30052_ (_26166_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not _30053_ (_26167_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _30054_ (_26168_, _26018_, _26167_);
  and _30055_ (_26169_, _26168_, _26166_);
  and _30056_ (_26170_, _26169_, _26165_);
  nand _30057_ (_26171_, _26170_, _26162_);
  or _30058_ (_26172_, _26171_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _30059_ (_26173_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _25991_);
  nor _30060_ (_26174_, _26173_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _30061_ (_26175_, _26174_, _26172_);
  and _30062_ (_26176_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _30063_ (_26177_, _26176_, _26175_);
  or _30064_ (_26178_, _26177_, _26035_);
  nor _30065_ (_26179_, _25987_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _30066_ (_26180_, _26179_, _26030_);
  and _30067_ (_26181_, _26180_, _26178_);
  and _30068_ (_26182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not _30069_ (_26183_, _26182_);
  and _30070_ (_26184_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nand _30071_ (_26185_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not _30072_ (_26186_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _30073_ (_26187_, _26018_, _26186_);
  and _30074_ (_26188_, _26187_, _26185_);
  nand _30075_ (_26189_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not _30076_ (_26190_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _30077_ (_26191_, _26009_, _26190_);
  and _30078_ (_26192_, _26191_, _26189_);
  not _30079_ (_26193_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _30080_ (_26194_, _25996_, _26193_);
  not _30081_ (_26195_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _30082_ (_26196_, _26002_, _26195_);
  and _30083_ (_26197_, _26196_, _26194_);
  and _30084_ (_26198_, _26197_, _26192_);
  nand _30085_ (_26199_, _26198_, _26188_);
  nand _30086_ (_26200_, _26199_, _25993_);
  nor _30087_ (_26201_, _26200_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _30088_ (_26202_, _26201_, _26184_);
  nand _30089_ (_26203_, _26202_, _26038_);
  nand _30090_ (_26204_, _26203_, _26183_);
  or _30091_ (_26205_, _26204_, _26035_);
  nor _30092_ (_26206_, _25987_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _30093_ (_26207_, _26206_, _26030_);
  nand _30094_ (_26208_, _26207_, _26205_);
  not _30095_ (_26209_, _26208_);
  and _30096_ (_26210_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _30097_ (_26211_, _26210_);
  not _30098_ (_26212_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _30099_ (_26213_, _25996_, _26212_);
  not _30100_ (_26214_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _30101_ (_26215_, _26002_, _26214_);
  and _30102_ (_26216_, _26215_, _26213_);
  nand _30103_ (_26217_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not _30104_ (_26218_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _30105_ (_26219_, _26009_, _26218_);
  and _30106_ (_26220_, _26219_, _26217_);
  nand _30107_ (_26221_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _30108_ (_26222_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _30109_ (_26223_, _26018_, _26222_);
  and _30110_ (_26224_, _26223_, _26221_);
  and _30111_ (_26225_, _26224_, _26220_);
  nand _30112_ (_26226_, _26225_, _26216_);
  and _30113_ (_26227_, _26226_, _25993_);
  or _30114_ (_26228_, _26227_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _30115_ (_26229_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _25991_);
  nor _30116_ (_26230_, _26229_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _30117_ (_26231_, _26230_, _26228_);
  nand _30118_ (_26232_, _26231_, _26211_);
  or _30119_ (_26233_, _26232_, _26035_);
  nor _30120_ (_26234_, _25987_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _30121_ (_26235_, _26234_, _26030_);
  and _30122_ (_26236_, _26235_, _26233_);
  and _30123_ (_26237_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _30124_ (_26238_, _26237_);
  and _30125_ (_26239_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _30126_ (_26240_, _25992_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand _30127_ (_26241_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  not _30128_ (_26242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _30129_ (_26243_, _26002_, _26242_);
  and _30130_ (_26244_, _26243_, _26241_);
  not _30131_ (_26245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _30132_ (_26246_, _25996_, _26245_);
  not _30133_ (_26247_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _30134_ (_26248_, _26018_, _26247_);
  and _30135_ (_26249_, _26248_, _26246_);
  nand _30136_ (_26250_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not _30137_ (_26251_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _30138_ (_26252_, _26009_, _26251_);
  and _30139_ (_26253_, _26252_, _26250_);
  and _30140_ (_26254_, _26253_, _26249_);
  and _30141_ (_26255_, _26254_, _26244_);
  nor _30142_ (_26256_, _26255_, _26240_);
  or _30143_ (_26257_, _26256_, _26239_);
  nand _30144_ (_26258_, _26257_, _26038_);
  nand _30145_ (_26259_, _26258_, _26238_);
  or _30146_ (_26260_, _26259_, _26035_);
  nor _30147_ (_26261_, _25987_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _30148_ (_26262_, _26261_, _26030_);
  nand _30149_ (_26263_, _26262_, _26260_);
  and _30150_ (_26264_, _26263_, _26236_);
  and _30151_ (_26265_, _26264_, _26209_);
  and _30152_ (_26266_, _26265_, _26181_);
  and _30153_ (_26267_, _26266_, _26155_);
  and _30154_ (_26268_, _26267_, _26034_);
  not _30155_ (_26269_, _26181_);
  nor _30156_ (_26270_, _26263_, _26236_);
  and _30157_ (_26271_, _26270_, _26209_);
  and _30158_ (_26272_, _26271_, _26269_);
  and _30159_ (_26273_, _26155_, _26034_);
  and _30160_ (_26274_, _26273_, _26272_);
  or _30161_ (_26275_, _26274_, _26268_);
  not _30162_ (_26276_, _26275_);
  and _30163_ (_26277_, _26125_, _26087_);
  not _30164_ (_26278_, _26153_);
  and _30165_ (_26279_, _26278_, _26033_);
  and _30166_ (_26280_, _26279_, _26277_);
  and _30167_ (_26281_, _26270_, _26208_);
  and _30168_ (_26282_, _26281_, _26269_);
  and _30169_ (_26283_, _26282_, _26280_);
  and _30170_ (_26284_, _26126_, _26087_);
  nor _30171_ (_26285_, _26153_, _26033_);
  and _30172_ (_26286_, _26285_, _26284_);
  and _30173_ (_26287_, _26286_, _26265_);
  or _30174_ (_26288_, _26287_, _26283_);
  and _30175_ (_26289_, _26271_, _26181_);
  and _30176_ (_26290_, _26289_, _26280_);
  nand _30177_ (_26291_, _26235_, _26233_);
  and _30178_ (_26292_, _26263_, _26291_);
  and _30179_ (_26293_, _26292_, _26208_);
  and _30180_ (_26294_, _26293_, _26181_);
  and _30181_ (_26295_, _26294_, _26280_);
  nor _30182_ (_26296_, _26295_, _26290_);
  nor _30183_ (_26297_, _26263_, _26291_);
  and _30184_ (_26298_, _26297_, _26208_);
  and _30185_ (_26299_, _26298_, _26181_);
  and _30186_ (_26300_, _26299_, _26273_);
  and _30187_ (_26301_, _26282_, _26155_);
  nor _30188_ (_26302_, _26301_, _26300_);
  nand _30189_ (_26303_, _26302_, _26296_);
  nor _30190_ (_26304_, _26303_, _26288_);
  and _30191_ (_26305_, _26304_, _26276_);
  and _30192_ (_26306_, _26289_, _26155_);
  and _30193_ (_26307_, _26306_, _26034_);
  and _30194_ (_26308_, _26265_, _26269_);
  and _30195_ (_26309_, _26308_, _26273_);
  nor _30196_ (_26310_, _26309_, _26307_);
  and _30197_ (_26311_, _26264_, _26208_);
  and _30198_ (_26312_, _26311_, _26181_);
  and _30199_ (_26313_, _26312_, _26286_);
  and _30200_ (_26314_, _26311_, _26269_);
  and _30201_ (_26315_, _26314_, _26286_);
  and _30202_ (_26316_, _26294_, _26286_);
  or _30203_ (_26317_, _26316_, _26315_);
  or _30204_ (_26318_, _26317_, _26313_);
  not _30205_ (_26319_, _26318_);
  and _30206_ (_26320_, _26293_, _26269_);
  nand _30207_ (_26321_, _26320_, _26280_);
  not _30208_ (_26322_, _26087_);
  and _30209_ (_26323_, _26308_, _26322_);
  not _30210_ (_26324_, _26323_);
  and _30211_ (_26325_, _26153_, _26125_);
  and _30212_ (_26326_, _26325_, _26087_);
  and _30213_ (_26327_, _26326_, _26269_);
  nand _30214_ (_26328_, _26327_, _26265_);
  and _30215_ (_26329_, _26328_, _26324_);
  and _30216_ (_26330_, _26329_, _26321_);
  and _30217_ (_26331_, _26330_, _26319_);
  and _30218_ (_26332_, _26331_, _26310_);
  and _30219_ (_26333_, _26281_, _26181_);
  and _30220_ (_26334_, _26333_, _26155_);
  and _30221_ (_26335_, _26292_, _26209_);
  and _30222_ (_26336_, _26335_, _26269_);
  and _30223_ (_26337_, _26336_, _26273_);
  nor _30224_ (_26338_, _26337_, _26334_);
  or _30225_ (_26339_, _26333_, _26311_);
  and _30226_ (_26340_, _26339_, _26280_);
  and _30227_ (_26341_, _26298_, _26269_);
  and _30228_ (_26342_, _26341_, _26155_);
  and _30229_ (_26343_, _26286_, _26271_);
  or _30230_ (_26344_, _26343_, _26342_);
  nor _30231_ (_26345_, _26344_, _26340_);
  and _30232_ (_26346_, _26345_, _26338_);
  and _30233_ (_26347_, _26341_, _26280_);
  and _30234_ (_26348_, _26280_, _26272_);
  nor _30235_ (_26349_, _26348_, _26347_);
  and _30236_ (_26350_, _26297_, _26209_);
  and _30237_ (_26351_, _26350_, _26269_);
  nand _30238_ (_26352_, _26351_, _26280_);
  and _30239_ (_26353_, _26311_, _26273_);
  not _30240_ (_26354_, _26353_);
  and _30241_ (_26355_, _26354_, _26352_);
  and _30242_ (_26356_, _26355_, _26349_);
  and _30243_ (_26357_, _26336_, _26280_);
  not _30244_ (_26358_, _26357_);
  and _30245_ (_26359_, _26335_, _26181_);
  nand _30246_ (_26360_, _26359_, _26273_);
  and _30247_ (_26361_, _26360_, _26358_);
  or _30248_ (_26362_, _26359_, _26266_);
  nand _30249_ (_26363_, _26362_, _26280_);
  and _30250_ (_26364_, _26363_, _26361_);
  and _30251_ (_26365_, _26364_, _26356_);
  and _30252_ (_26366_, _26365_, _26346_);
  and _30253_ (_26367_, _26366_, _26332_);
  nand _30254_ (_26368_, _26367_, _26305_);
  nand _30255_ (_26369_, _26368_, _25983_);
  not _30256_ (_26370_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _30257_ (_26371_, _23914_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _30258_ (_26372_, _26371_, _26370_);
  not _30259_ (_26373_, _26263_);
  and _30260_ (_26374_, _26373_, _26208_);
  and _30261_ (_26375_, _26286_, _26374_);
  and _30262_ (_26376_, _26375_, _26372_);
  and _30263_ (_26377_, _26153_, _26034_);
  and _30264_ (_26378_, _26377_, _26284_);
  and _30265_ (_26379_, _26378_, _26312_);
  and _30266_ (_26380_, _26378_, _26314_);
  nor _30267_ (_26381_, _26380_, _26379_);
  and _30268_ (_26382_, \oc8051_top_1.oc8051_decoder1.state [0], _23914_);
  and _30269_ (_26383_, _26382_, \oc8051_top_1.oc8051_decoder1.state [1]);
  not _30270_ (_26384_, _26383_);
  nor _30271_ (_26385_, _26384_, _26381_);
  nor _30272_ (_26386_, _26385_, _26376_);
  nand _30273_ (_26387_, _26386_, _26369_);
  nand _30274_ (_26388_, _26387_, _23914_);
  and _30275_ (_26389_, _26388_, _25981_);
  not _30276_ (_26390_, _26389_);
  and _30277_ (_26391_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _30278_ (_26392_, _26391_);
  not _30279_ (_26393_, _25983_);
  nand _30280_ (_26394_, _26289_, _26286_);
  and _30281_ (_26395_, _26354_, _26394_);
  and _30282_ (_26396_, _26181_, _26087_);
  and _30283_ (_26397_, _26396_, _26325_);
  and _30284_ (_26398_, _26397_, _26265_);
  and _30285_ (_26399_, _26326_, _26293_);
  nor _30286_ (_26400_, _26399_, _26398_);
  and _30287_ (_26401_, _26400_, _26395_);
  and _30288_ (_26402_, _26397_, _26281_);
  and _30289_ (_26403_, _26326_, _26311_);
  or _30290_ (_26404_, _26403_, _26402_);
  and _30291_ (_26405_, _26326_, _26271_);
  not _30292_ (_26406_, _26405_);
  nand _30293_ (_26407_, _26359_, _26326_);
  and _30294_ (_26408_, _26407_, _26406_);
  not _30295_ (_26409_, _26408_);
  nor _30296_ (_26410_, _26409_, _26404_);
  and _30297_ (_26411_, _26410_, _26401_);
  and _30298_ (_26412_, _26154_, _26033_);
  and _30299_ (_26413_, _26412_, _26087_);
  and _30300_ (_26414_, _26308_, _26413_);
  not _30301_ (_26415_, _26414_);
  nand _30302_ (_26416_, _26359_, _26413_);
  nand _30303_ (_26417_, _26299_, _26413_);
  and _30304_ (_26418_, _26417_, _26416_);
  and _30305_ (_26419_, _26418_, _26415_);
  and _30306_ (_26420_, _26336_, _26326_);
  not _30307_ (_26421_, _26420_);
  not _30308_ (_26422_, _26327_);
  nor _30309_ (_26423_, _26350_, _26281_);
  or _30310_ (_26424_, _26423_, _26422_);
  nand _30311_ (_26425_, _26341_, _26326_);
  and _30312_ (_26426_, _26425_, _26424_);
  and _30313_ (_26427_, _26426_, _26421_);
  and _30314_ (_26428_, _26427_, _26419_);
  and _30315_ (_26429_, _26428_, _26411_);
  or _30316_ (_26430_, _26429_, _26393_);
  and _30317_ (_26431_, _26298_, _26286_);
  and _30318_ (_26432_, _26431_, _26372_);
  nor _30319_ (_26433_, _26432_, _26385_);
  and _30320_ (_26434_, _26433_, _26430_);
  or _30321_ (_26435_, _26434_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _30322_ (_26436_, _26435_, _26392_);
  and _30323_ (_26437_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _30324_ (_26438_, _26285_, _26277_);
  and _30325_ (_26439_, _26438_, _26336_);
  and _30326_ (_26440_, _26438_, _26308_);
  nor _30327_ (_26441_, _26440_, _26439_);
  and _30328_ (_26442_, _26441_, _26419_);
  nor _30329_ (_26443_, _26442_, _26393_);
  not _30330_ (_26444_, _26443_);
  and _30331_ (_26445_, _26372_, _26286_);
  and _30332_ (_26446_, _26445_, _26374_);
  and _30333_ (_26447_, _26440_, _23914_);
  and _30334_ (_26448_, _26439_, _23914_);
  nor _30335_ (_26449_, _26448_, _26447_);
  nor _30336_ (_26450_, _26449_, _25982_);
  nor _30337_ (_26451_, _26450_, _26446_);
  and _30338_ (_26452_, _26451_, _26444_);
  nor _30339_ (_26453_, _26452_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _30340_ (_26454_, _26453_, _26437_);
  nand _30341_ (_26455_, _26454_, _27355_);
  nor _30342_ (_24440_, _26455_, _26436_);
  and _30343_ (_09474_, _24440_, _26390_);
  and _30344_ (_26456_, _25450_, _25115_);
  and _30345_ (_26457_, _25128_, _25085_);
  not _30346_ (_26458_, _25073_);
  nor _30347_ (_26459_, _26458_, _25101_);
  and _30348_ (_26460_, _26459_, _26457_);
  and _30349_ (_26461_, _26460_, _25650_);
  and _30350_ (_26462_, _26461_, _25020_);
  and _30351_ (_26463_, _26462_, _26456_);
  not _30352_ (_26464_, _26463_);
  and _30353_ (_26465_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _30354_ (_26466_, _25239_, _24471_);
  nor _30355_ (_26467_, _26466_, _24487_);
  and _30356_ (_26468_, _26467_, _25915_);
  and _30357_ (_26469_, _26468_, _25424_);
  nor _30358_ (_26470_, _25426_, _25549_);
  and _30359_ (_26471_, _26470_, _26469_);
  nor _30360_ (_26472_, _26471_, _24141_);
  not _30361_ (_26473_, _26472_);
  and _30362_ (_26474_, _26473_, _25954_);
  and _30363_ (_26475_, _26474_, _25936_);
  nor _30364_ (_26476_, _26475_, _26464_);
  nor _30365_ (_26477_, _26476_, _26465_);
  and _30366_ (_26478_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _30367_ (_26479_, _26471_, _25364_);
  not _30368_ (_26480_, _26479_);
  and _30369_ (_26481_, _26480_, _25886_);
  and _30370_ (_26482_, _26481_, _25871_);
  nor _30371_ (_26483_, _26482_, _26464_);
  nor _30372_ (_26484_, _26483_, _26478_);
  and _30373_ (_26485_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _30374_ (_26486_, _26471_, _23973_);
  not _30375_ (_26487_, _26486_);
  and _30376_ (_26488_, _26487_, _25820_);
  and _30377_ (_26489_, _26488_, _25808_);
  nor _30378_ (_26490_, _26489_, _26464_);
  nor _30379_ (_26491_, _26490_, _26485_);
  and _30380_ (_26492_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _30381_ (_26493_, _26471_, _24101_);
  not _30382_ (_26494_, _26493_);
  and _30383_ (_26495_, _26494_, _25749_);
  and _30384_ (_26496_, _26495_, _25746_);
  and _30385_ (_26497_, _26496_, _25737_);
  nor _30386_ (_26498_, _26497_, _26464_);
  nor _30387_ (_26499_, _26498_, _26492_);
  and _30388_ (_26500_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _30389_ (_26501_, _26471_, _25664_);
  not _30390_ (_26502_, _26501_);
  and _30391_ (_26503_, _26502_, _25681_);
  and _30392_ (_26504_, _26503_, _25685_);
  and _30393_ (_26505_, _26504_, _25672_);
  nor _30394_ (_26506_, _26505_, _26464_);
  nor _30395_ (_26507_, _26506_, _26500_);
  and _30396_ (_26508_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _30397_ (_26509_, _26471_, _25355_);
  not _30398_ (_26510_, _26509_);
  and _30399_ (_26511_, _26510_, _25608_);
  and _30400_ (_26512_, _26511_, _25636_);
  nor _30401_ (_26513_, _26512_, _26464_);
  nor _30402_ (_26514_, _26513_, _26508_);
  and _30403_ (_26515_, _26456_, _25020_);
  and _30404_ (_26516_, _26515_, _26461_);
  nor _30405_ (_26517_, _26516_, _25046_);
  nor _30406_ (_26518_, _26471_, _24253_);
  not _30407_ (_26519_, _26518_);
  and _30408_ (_26520_, _26519_, _25546_);
  and _30409_ (_26521_, _26520_, _25543_);
  not _30410_ (_26522_, _26521_);
  and _30411_ (_26523_, _26522_, _26516_);
  nor _30412_ (_26524_, _26523_, _26517_);
  and _30413_ (_26525_, _26524_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _30414_ (_26526_, _26525_, _26514_);
  and _30415_ (_26527_, _26526_, _26507_);
  and _30416_ (_26528_, _26527_, _26499_);
  and _30417_ (_26529_, _26528_, _26491_);
  and _30418_ (_26530_, _26529_, _26484_);
  and _30419_ (_26531_, _26530_, _26477_);
  nor _30420_ (_26532_, _26516_, _25087_);
  nand _30421_ (_26533_, _26532_, _26531_);
  or _30422_ (_26534_, _26532_, _26531_);
  and _30423_ (_26535_, _26534_, _25061_);
  nand _30424_ (_26536_, _26535_, _26533_);
  nor _30425_ (_26537_, _26516_, _25091_);
  and _30426_ (_26538_, _26537_, _26536_);
  nor _30427_ (_26539_, _26471_, _24172_);
  not _30428_ (_26540_, _26539_);
  and _30429_ (_26541_, _26540_, _25420_);
  and _30430_ (_26542_, _26541_, _25415_);
  and _30431_ (_26543_, _26542_, _25385_);
  and _30432_ (_26544_, _26543_, _26463_);
  nor _30433_ (_26545_, _26544_, _26538_);
  and _30434_ (_09496_, _26545_, _27355_);
  not _30435_ (_26546_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _30436_ (_26547_, _26524_, _26546_);
  nor _30437_ (_26548_, _26524_, _26546_);
  nor _30438_ (_26549_, _26548_, _26547_);
  and _30439_ (_26550_, _26549_, _25061_);
  nor _30440_ (_26551_, _26550_, _25047_);
  nor _30441_ (_26552_, _26551_, _26463_);
  nor _30442_ (_26553_, _26552_, _26523_);
  nand _30443_ (_10718_, _26553_, _27355_);
  nor _30444_ (_26554_, _26525_, _26514_);
  nor _30445_ (_26555_, _26554_, _26526_);
  nor _30446_ (_26556_, _26555_, _24979_);
  nor _30447_ (_26557_, _26556_, _25028_);
  nor _30448_ (_26558_, _26557_, _26463_);
  nor _30449_ (_26559_, _26558_, _26513_);
  nand _30450_ (_10729_, _26559_, _27355_);
  nor _30451_ (_26560_, _26526_, _26507_);
  nor _30452_ (_26561_, _26560_, _26527_);
  nor _30453_ (_26562_, _26561_, _24979_);
  nor _30454_ (_26563_, _26562_, _24984_);
  nor _30455_ (_26564_, _26563_, _26463_);
  nor _30456_ (_26565_, _26564_, _26506_);
  nand _30457_ (_10740_, _26565_, _27355_);
  nor _30458_ (_26566_, _26527_, _26499_);
  nor _30459_ (_26567_, _26566_, _26528_);
  nor _30460_ (_26568_, _26567_, _24979_);
  nor _30461_ (_26569_, _26568_, _25109_);
  nor _30462_ (_26570_, _26569_, _26463_);
  nor _30463_ (_26571_, _26570_, _26498_);
  nor _30464_ (_10751_, _26571_, rst);
  nor _30465_ (_26572_, _26528_, _26491_);
  nor _30466_ (_26573_, _26572_, _26529_);
  nor _30467_ (_26574_, _26573_, _24979_);
  nor _30468_ (_26575_, _26574_, _25121_);
  nor _30469_ (_26576_, _26575_, _26463_);
  nor _30470_ (_26577_, _26576_, _26490_);
  nor _30471_ (_10762_, _26577_, rst);
  nor _30472_ (_26578_, _26529_, _26484_);
  nor _30473_ (_26579_, _26578_, _26530_);
  nor _30474_ (_26580_, _26579_, _24979_);
  nor _30475_ (_26581_, _26580_, _25077_);
  nor _30476_ (_26582_, _26581_, _26463_);
  nor _30477_ (_26583_, _26582_, _26483_);
  nor _30478_ (_10773_, _26583_, rst);
  nor _30479_ (_26584_, _26530_, _26477_);
  nor _30480_ (_26585_, _26584_, _26531_);
  nor _30481_ (_26586_, _26585_, _24979_);
  nor _30482_ (_26587_, _26586_, _25064_);
  nor _30483_ (_26588_, _26587_, _26463_);
  nor _30484_ (_26589_, _26588_, _26476_);
  nor _30485_ (_10784_, _26589_, rst);
  and _30486_ (_26590_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _23914_);
  and _30487_ (_26591_, _26590_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _30488_ (_26592_, _26460_, _25778_);
  nand _30489_ (_26593_, _26592_, _26456_);
  and _30490_ (_26594_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _30491_ (_26595_, _25020_, _25115_);
  and _30492_ (_26596_, _25516_, _26595_);
  and _30493_ (_26597_, _26596_, _26460_);
  and _30494_ (_26598_, _26597_, _25449_);
  and _30495_ (_26599_, _26598_, _25444_);
  and _30496_ (_26600_, _26599_, _25441_);
  or _30497_ (_26601_, _26600_, _26594_);
  or _30498_ (_26602_, _26601_, _26591_);
  not _30499_ (_26603_, _26591_);
  nor _30500_ (_26604_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _30501_ (_26605_, _24108_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30502_ (_26606_, _26605_, _26604_);
  nor _30503_ (_26607_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _30504_ (_26608_, _24089_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30505_ (_26609_, _26608_, _26607_);
  nor _30506_ (_26610_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _30507_ (_26611_, _24240_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30508_ (_26612_, _26611_, _26610_);
  not _30509_ (_26613_, _26612_);
  nor _30510_ (_26614_, _26613_, _25461_);
  nor _30511_ (_26615_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _30512_ (_26616_, _24188_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30513_ (_26617_, _26616_, _26615_);
  and _30514_ (_26618_, _26617_, _26614_);
  nor _30515_ (_26619_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _30516_ (_26620_, _24204_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30517_ (_26621_, _26620_, _26619_);
  and _30518_ (_26622_, _26621_, _26618_);
  and _30519_ (_26623_, _26622_, _26609_);
  nor _30520_ (_26624_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _30521_ (_26625_, _23940_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30522_ (_26626_, _26625_, _26624_);
  and _30523_ (_26627_, _26626_, _26623_);
  and _30524_ (_26628_, _26627_, _26606_);
  nor _30525_ (_26629_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _30526_ (_26630_, _24129_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30527_ (_26631_, _26630_, _26629_);
  and _30528_ (_26632_, _26631_, _26628_);
  nor _30529_ (_26633_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _30530_ (_26634_, _24158_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _30531_ (_26635_, _26634_, _26633_);
  or _30532_ (_26636_, _26635_, _26632_);
  nand _30533_ (_26637_, _26635_, _26632_);
  and _30534_ (_26638_, _26637_, _26636_);
  and _30535_ (_26639_, _26638_, _25240_);
  and _30536_ (_26640_, _24443_, _23920_);
  and _30537_ (_26641_, _25361_, _24278_);
  and _30538_ (_26642_, _26641_, _24082_);
  and _30539_ (_26643_, _26642_, _24032_);
  and _30540_ (_26644_, _26643_, _24515_);
  and _30541_ (_26645_, _26644_, _24533_);
  and _30542_ (_26646_, _26645_, _24520_);
  or _30543_ (_26647_, _26646_, _25363_);
  and _30544_ (_26648_, _25370_, _24172_);
  and _30545_ (_26649_, _24018_, _24068_);
  nor _30546_ (_26650_, _24032_, _24082_);
  and _30547_ (_26651_, _26650_, _26649_);
  and _30548_ (_26652_, _26651_, _26648_);
  and _30549_ (_26653_, _24004_, _24055_);
  and _30550_ (_26654_, _26653_, _26652_);
  nor _30551_ (_26655_, _26654_, _25199_);
  not _30552_ (_26656_, _26655_);
  nand _30553_ (_26657_, _25199_, _24004_);
  and _30554_ (_26658_, _26657_, _26656_);
  and _30555_ (_26659_, _26658_, _26647_);
  and _30556_ (_26660_, _25199_, _24616_);
  nor _30557_ (_26661_, _26660_, _25926_);
  and _30558_ (_26662_, _26661_, _26659_);
  or _30559_ (_26663_, _26662_, _25377_);
  nand _30560_ (_26664_, _26662_, _25377_);
  and _30561_ (_26665_, _26664_, _26663_);
  and _30562_ (_26666_, _26665_, _25354_);
  and _30563_ (_26667_, _25199_, _25377_);
  or _30564_ (_26668_, _26667_, _25472_);
  and _30565_ (_26669_, _26668_, _25381_);
  nor _30566_ (_26670_, _25502_, _24101_);
  nor _30567_ (_26671_, _25424_, _23990_);
  and _30568_ (_26672_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or _30569_ (_26673_, _26672_, _26671_);
  or _30570_ (_26674_, _26673_, _26670_);
  or _30571_ (_26675_, _26674_, _26669_);
  or _30572_ (_26676_, _26675_, _26666_);
  or _30573_ (_26677_, _26676_, _26640_);
  or _30574_ (_26678_, _26677_, _26639_);
  or _30575_ (_26679_, _26678_, _26603_);
  and _30576_ (_26680_, _26679_, _27355_);
  and _30577_ (_12743_, _26680_, _26602_);
  and _30578_ (_26681_, _26456_, _25716_);
  and _30579_ (_26682_, _26681_, _26460_);
  nor _30580_ (_26683_, _26682_, _26591_);
  or _30581_ (_26684_, _26683_, _25441_);
  not _30582_ (_26685_, _26683_);
  or _30583_ (_26686_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _30584_ (_26687_, _26686_, _27355_);
  and _30585_ (_12764_, _26687_, _26684_);
  nor _30586_ (_26688_, _26593_, _25562_);
  and _30587_ (_26689_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _30588_ (_26690_, _26689_, _26591_);
  or _30589_ (_26691_, _26690_, _26688_);
  and _30590_ (_26692_, _26613_, _25461_);
  nor _30591_ (_26693_, _26692_, _26614_);
  and _30592_ (_26694_, _26693_, _25240_);
  nand _30593_ (_26695_, _24923_, _24487_);
  nor _30594_ (_26696_, _25472_, _25380_);
  not _30595_ (_26697_, _26696_);
  nor _30596_ (_26698_, _26697_, _25372_);
  nor _30597_ (_26699_, _26698_, _24082_);
  and _30598_ (_26700_, _26698_, _24082_);
  nor _30599_ (_26701_, _26700_, _26699_);
  and _30600_ (_26702_, _26701_, _25354_);
  and _30601_ (_26703_, _25423_, _24082_);
  and _30602_ (_26704_, _24394_, _23920_);
  nor _30603_ (_26705_, _25502_, _23973_);
  nor _30604_ (_26706_, _25382_, _24253_);
  or _30605_ (_26707_, _26706_, _26705_);
  or _30606_ (_26708_, _26707_, _26704_);
  nor _30607_ (_26709_, _26708_, _26703_);
  not _30608_ (_26710_, _26709_);
  nor _30609_ (_26711_, _26710_, _26702_);
  nand _30610_ (_26712_, _26711_, _26695_);
  or _30611_ (_26713_, _26712_, _26694_);
  or _30612_ (_26714_, _26713_, _26603_);
  and _30613_ (_26715_, _26714_, _27355_);
  and _30614_ (_13683_, _26715_, _26691_);
  and _30615_ (_26716_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _30616_ (_26717_, _26599_, _25639_);
  or _30617_ (_26718_, _26717_, _26716_);
  or _30618_ (_26719_, _26718_, _26591_);
  nor _30619_ (_26720_, _26617_, _26614_);
  not _30620_ (_26721_, _26720_);
  nor _30621_ (_26722_, _26618_, _25459_);
  and _30622_ (_26723_, _26722_, _26721_);
  not _30623_ (_26724_, _26723_);
  and _30624_ (_26725_, _24632_, _24487_);
  not _30625_ (_26726_, _26725_);
  and _30626_ (_26727_, _25423_, _24032_);
  nor _30627_ (_26728_, _26642_, _25363_);
  and _30628_ (_26729_, _26648_, _25146_);
  nor _30629_ (_26730_, _26729_, _25199_);
  or _30630_ (_26731_, _26730_, _26728_);
  and _30631_ (_26732_, _26731_, _25310_);
  not _30632_ (_26733_, _26732_);
  nor _30633_ (_26734_, _26731_, _25310_);
  nor _30634_ (_26735_, _26734_, _25867_);
  and _30635_ (_26736_, _26735_, _26733_);
  and _30636_ (_26737_, _24396_, _23920_);
  and _30637_ (_26738_, _25501_, _24120_);
  and _30638_ (_26739_, _25381_, _24200_);
  or _30639_ (_26740_, _26739_, _26738_);
  or _30640_ (_26741_, _26740_, _26737_);
  or _30641_ (_26742_, _26741_, _26736_);
  nor _30642_ (_26743_, _26742_, _26727_);
  and _30643_ (_26744_, _26743_, _26726_);
  and _30644_ (_26745_, _26744_, _26724_);
  nand _30645_ (_26746_, _26745_, _26591_);
  and _30646_ (_26747_, _26746_, _27355_);
  and _30647_ (_13694_, _26747_, _26719_);
  nor _30648_ (_26748_, _26593_, _25704_);
  and _30649_ (_26749_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _30650_ (_26750_, _26749_, _26591_);
  or _30651_ (_26751_, _26750_, _26748_);
  nor _30652_ (_26752_, _26621_, _26618_);
  nor _30653_ (_26753_, _26752_, _26622_);
  and _30654_ (_26754_, _26753_, _25240_);
  not _30655_ (_26755_, _26754_);
  and _30656_ (_26756_, _26729_, _25310_);
  and _30657_ (_26757_, _26756_, _25363_);
  and _30658_ (_26758_, _26643_, _25199_);
  nor _30659_ (_26759_, _26758_, _26757_);
  and _30660_ (_26760_, _26759_, _24068_);
  nor _30661_ (_26761_, _26759_, _24068_);
  nor _30662_ (_26762_, _26761_, _26760_);
  and _30663_ (_26763_, _26762_, _25354_);
  and _30664_ (_26764_, _25381_, _24216_);
  and _30665_ (_26765_, _25423_, _24515_);
  nor _30666_ (_26766_, _26765_, _26764_);
  and _30667_ (_26767_, _24398_, _23920_);
  nor _30668_ (_26768_, _25502_, _24141_);
  and _30669_ (_26769_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _30670_ (_26770_, _26769_, _26768_);
  nor _30671_ (_26771_, _26770_, _26767_);
  and _30672_ (_26772_, _26771_, _26766_);
  not _30673_ (_26773_, _26772_);
  nor _30674_ (_26774_, _26773_, _26763_);
  and _30675_ (_26775_, _26774_, _26755_);
  nand _30676_ (_26776_, _26775_, _26591_);
  and _30677_ (_26777_, _26776_, _27355_);
  and _30678_ (_13705_, _26777_, _26751_);
  nor _30679_ (_26778_, _26593_, _25769_);
  and _30680_ (_26779_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _30681_ (_26780_, _26779_, _26591_);
  or _30682_ (_26781_, _26780_, _26778_);
  nor _30683_ (_26782_, _26622_, _26609_);
  not _30684_ (_26783_, _26782_);
  nor _30685_ (_26784_, _26623_, _25459_);
  and _30686_ (_26785_, _26784_, _26783_);
  not _30687_ (_26786_, _26785_);
  and _30688_ (_26787_, _24401_, _23920_);
  not _30689_ (_26788_, _26787_);
  nor _30690_ (_26789_, _26645_, _25363_);
  nor _30691_ (_26790_, _26644_, _24533_);
  not _30692_ (_26791_, _26790_);
  and _30693_ (_26792_, _26791_, _26789_);
  and _30694_ (_26793_, _26756_, _24068_);
  nor _30695_ (_26794_, _26793_, _24018_);
  nor _30696_ (_26795_, _26794_, _26652_);
  nor _30697_ (_26796_, _26795_, _25199_);
  nor _30698_ (_26797_, _26796_, _26792_);
  nor _30699_ (_26798_, _26797_, _25867_);
  and _30700_ (_26799_, _25423_, _24533_);
  nor _30701_ (_26800_, _25382_, _24101_);
  and _30702_ (_26801_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _30703_ (_26802_, _26801_, _26800_);
  or _30704_ (_26803_, _26802_, _25503_);
  nor _30705_ (_26804_, _26803_, _26799_);
  not _30706_ (_26805_, _26804_);
  nor _30707_ (_26806_, _26805_, _26798_);
  and _30708_ (_26807_, _26806_, _26788_);
  and _30709_ (_26808_, _26807_, _26786_);
  nand _30710_ (_26809_, _26808_, _26591_);
  and _30711_ (_26810_, _26809_, _27355_);
  and _30712_ (_13716_, _26810_, _26781_);
  and _30713_ (_26811_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _30714_ (_26812_, _26599_, _25830_);
  or _30715_ (_26813_, _26812_, _26811_);
  or _30716_ (_26814_, _26813_, _26591_);
  or _30717_ (_26815_, _26626_, _26623_);
  nor _30718_ (_26816_, _26627_, _25459_);
  and _30719_ (_26817_, _26816_, _26815_);
  nor _30720_ (_26818_, _26652_, _25199_);
  nor _30721_ (_26819_, _26818_, _26789_);
  or _30722_ (_26820_, _26819_, _24520_);
  nand _30723_ (_26821_, _26819_, _24520_);
  and _30724_ (_26822_, _26821_, _26820_);
  and _30725_ (_26823_, _26822_, _25354_);
  and _30726_ (_26824_, _24403_, _23920_);
  or _30727_ (_26825_, _25199_, _23974_);
  nand _30728_ (_26826_, _25199_, _24055_);
  and _30729_ (_26827_, _26826_, _25381_);
  and _30730_ (_26828_, _26827_, _26825_);
  nor _30731_ (_26829_, _25502_, _24253_);
  and _30732_ (_26830_, _25423_, _24520_);
  and _30733_ (_26831_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _30734_ (_26832_, _26831_, _26830_);
  or _30735_ (_26833_, _26832_, _26829_);
  or _30736_ (_26834_, _26833_, _26828_);
  or _30737_ (_26835_, _26834_, _26824_);
  or _30738_ (_26836_, _26835_, _26823_);
  or _30739_ (_26837_, _26836_, _26817_);
  or _30740_ (_26838_, _26837_, _26603_);
  and _30741_ (_26839_, _26838_, _27355_);
  and _30742_ (_13727_, _26839_, _26814_);
  and _30743_ (_26840_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _30744_ (_26841_, _26599_, _25898_);
  or _30745_ (_26842_, _26841_, _26840_);
  or _30746_ (_26843_, _26842_, _26591_);
  or _30747_ (_26844_, _26627_, _26606_);
  nor _30748_ (_26845_, _26628_, _25459_);
  and _30749_ (_26846_, _26845_, _26844_);
  and _30750_ (_26847_, _24413_, _23920_);
  and _30751_ (_26848_, _26652_, _24055_);
  nor _30752_ (_26849_, _26848_, _25199_);
  not _30753_ (_26850_, _26849_);
  and _30754_ (_26851_, _26850_, _26647_);
  and _30755_ (_26852_, _26851_, _24004_);
  nor _30756_ (_26853_, _26851_, _24004_);
  or _30757_ (_26854_, _26853_, _26852_);
  and _30758_ (_26855_, _26854_, _25354_);
  or _30759_ (_26856_, _25199_, _24120_);
  and _30760_ (_26857_, _26657_, _25381_);
  and _30761_ (_26858_, _26857_, _26856_);
  and _30762_ (_26859_, _25501_, _24200_);
  and _30763_ (_26860_, _25423_, _24535_);
  and _30764_ (_26861_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _30765_ (_26862_, _26861_, _26860_);
  or _30766_ (_26863_, _26862_, _26859_);
  or _30767_ (_26864_, _26863_, _26858_);
  or _30768_ (_26865_, _26864_, _26855_);
  or _30769_ (_26866_, _26865_, _26847_);
  or _30770_ (_26867_, _26866_, _26846_);
  or _30771_ (_26868_, _26867_, _26603_);
  and _30772_ (_26869_, _26868_, _27355_);
  and _30773_ (_13738_, _26869_, _26843_);
  nor _30774_ (_26870_, _26593_, _25963_);
  and _30775_ (_26871_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _30776_ (_26872_, _26871_, _26591_);
  or _30777_ (_26873_, _26872_, _26870_);
  nor _30778_ (_26874_, _26631_, _26628_);
  nor _30779_ (_26875_, _26874_, _26632_);
  and _30780_ (_26876_, _26875_, _25240_);
  not _30781_ (_26877_, _26876_);
  and _30782_ (_26878_, _24441_, _23920_);
  nor _30783_ (_26879_, _26659_, _24616_);
  and _30784_ (_26880_, _26659_, _24616_);
  nor _30785_ (_26881_, _26880_, _26879_);
  nor _30786_ (_26882_, _26881_, _25867_);
  nor _30787_ (_26883_, _25199_, _24143_);
  not _30788_ (_26884_, _26883_);
  nor _30789_ (_26885_, _26660_, _25382_);
  and _30790_ (_26886_, _26885_, _26884_);
  and _30791_ (_26887_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  and _30792_ (_26888_, _25501_, _24216_);
  and _30793_ (_26889_, _25423_, _24049_);
  or _30794_ (_26890_, _26889_, _26888_);
  nor _30795_ (_26891_, _26890_, _26887_);
  not _30796_ (_26892_, _26891_);
  nor _30797_ (_26893_, _26892_, _26886_);
  not _30798_ (_26894_, _26893_);
  nor _30799_ (_26895_, _26894_, _26882_);
  not _30800_ (_26896_, _26895_);
  nor _30801_ (_26897_, _26896_, _26878_);
  and _30802_ (_26898_, _26897_, _26877_);
  nand _30803_ (_26899_, _26898_, _26591_);
  and _30804_ (_26900_, _26899_, _27355_);
  and _30805_ (_13749_, _26900_, _26873_);
  nand _30806_ (_26901_, _26685_, _25562_);
  or _30807_ (_26902_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _30808_ (_26903_, _26902_, _27355_);
  and _30809_ (_13760_, _26903_, _26901_);
  or _30810_ (_26904_, _26683_, _25639_);
  or _30811_ (_26905_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _30812_ (_26906_, _26905_, _27355_);
  and _30813_ (_13771_, _26906_, _26904_);
  nand _30814_ (_26907_, _26685_, _25704_);
  or _30815_ (_26908_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _30816_ (_26909_, _26908_, _27355_);
  and _30817_ (_13782_, _26909_, _26907_);
  nand _30818_ (_26910_, _26685_, _25769_);
  or _30819_ (_26911_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _30820_ (_26912_, _26911_, _27355_);
  and _30821_ (_13793_, _26912_, _26910_);
  or _30822_ (_26913_, _26683_, _25830_);
  or _30823_ (_26914_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _30824_ (_26915_, _26914_, _27355_);
  and _30825_ (_13804_, _26915_, _26913_);
  or _30826_ (_26916_, _26683_, _25898_);
  or _30827_ (_26917_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _30828_ (_26918_, _26917_, _27355_);
  and _30829_ (_13815_, _26918_, _26916_);
  nand _30830_ (_26919_, _26685_, _25963_);
  or _30831_ (_26920_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _30832_ (_26921_, _26920_, _27355_);
  and _30833_ (_13826_, _26921_, _26919_);
  not _30834_ (_26922_, _25085_);
  nor _30835_ (_26923_, _26922_, _25073_);
  and _30836_ (_26924_, _26923_, _25521_);
  and _30837_ (_26925_, _26924_, _25130_);
  not _30838_ (_26926_, _25517_);
  nor _30839_ (_26927_, _26926_, _25514_);
  not _30840_ (_26928_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _30841_ (_26929_, _25517_, _26928_);
  or _30842_ (_26930_, _26929_, _26927_);
  and _30843_ (_26931_, _26930_, _26925_);
  nor _30844_ (_26932_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _30845_ (_26933_, _26932_);
  nand _30846_ (_26934_, _26933_, _25514_);
  and _30847_ (_26935_, _26932_, _26928_);
  nor _30848_ (_26936_, _26935_, _26925_);
  and _30849_ (_26937_, _26936_, _26934_);
  nor _30850_ (_26938_, _25128_, _26922_);
  nor _30851_ (_26939_, _25073_, _25101_);
  and _30852_ (_26940_, _26456_, _25055_);
  and _30853_ (_26941_, _26940_, _26939_);
  and _30854_ (_26942_, _26941_, _26938_);
  or _30855_ (_26943_, _26942_, _26937_);
  or _30856_ (_26944_, _26943_, _26931_);
  nand _30857_ (_26945_, _26942_, _26543_);
  and _30858_ (_26946_, _26945_, _27355_);
  and _30859_ (_15222_, _26946_, _26944_);
  and _30860_ (_26947_, _25650_, _25020_);
  and _30861_ (_26948_, _26925_, _26947_);
  nand _30862_ (_26949_, _26948_, _25514_);
  not _30863_ (_26950_, _26942_);
  or _30864_ (_26951_, _26948_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _30865_ (_26952_, _26951_, _26950_);
  and _30866_ (_26953_, _26952_, _26949_);
  nor _30867_ (_26954_, _26950_, _26512_);
  or _30868_ (_26955_, _26954_, _26953_);
  and _30869_ (_17288_, _26955_, _27355_);
  or _30870_ (_26956_, _24452_, _24448_);
  or _30871_ (_26957_, _26956_, _24456_);
  or _30872_ (_26958_, _26957_, _24460_);
  nor _30873_ (_26959_, _26958_, _24465_);
  nand _30874_ (_26960_, _26959_, _24467_);
  and _30875_ (_26961_, _26960_, _23920_);
  and _30876_ (_26962_, _25465_, _25348_);
  not _30877_ (_26963_, _25348_);
  and _30878_ (_26964_, _25466_, _26963_);
  or _30879_ (_26965_, _26964_, _26962_);
  and _30880_ (_26966_, _26965_, _25246_);
  not _30881_ (_26967_, _25233_);
  nand _30882_ (_26968_, _25232_, _26967_);
  or _30883_ (_26969_, _25234_, _25232_);
  and _30884_ (_26970_, _25240_, _26969_);
  and _30885_ (_26971_, _26970_, _26968_);
  and _30886_ (_26972_, _26653_, _24617_);
  and _30887_ (_26973_, _26651_, _24487_);
  nand _30888_ (_26974_, _26973_, _26972_);
  nand _30889_ (_26975_, _26974_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _30890_ (_26976_, _26975_, _26971_);
  or _30891_ (_26977_, _26976_, _26966_);
  or _30892_ (_26978_, _26977_, _25789_);
  or _30893_ (_26979_, _26978_, _25134_);
  or _30894_ (_26980_, _26979_, _26961_);
  nor _30895_ (_26981_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _30896_ (_26982_, _26981_, _26925_);
  and _30897_ (_26983_, _26982_, _26980_);
  and _30898_ (_26984_, _25717_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _30899_ (_26985_, _26984_, _25718_);
  and _30900_ (_26986_, _26985_, _26925_);
  or _30901_ (_26987_, _26986_, _26942_);
  or _30902_ (_26988_, _26987_, _26983_);
  nand _30903_ (_26989_, _26942_, _26505_);
  and _30904_ (_26990_, _26989_, _27355_);
  and _30905_ (_17297_, _26990_, _26988_);
  and _30906_ (_26991_, _26925_, _25778_);
  nand _30907_ (_26992_, _26991_, _25514_);
  or _30908_ (_26993_, _26991_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _30909_ (_26994_, _26993_, _26950_);
  and _30910_ (_26995_, _26994_, _26992_);
  nor _30911_ (_26996_, _26950_, _26497_);
  or _30912_ (_26997_, _26996_, _26995_);
  and _30913_ (_17306_, _26997_, _27355_);
  not _30914_ (_26998_, _26925_);
  or _30915_ (_26999_, _26998_, _25840_);
  and _30916_ (_27000_, _26999_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _30917_ (_27001_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _30918_ (_27002_, _27001_, _25843_);
  and _30919_ (_27003_, _27002_, _26925_);
  or _30920_ (_27004_, _27003_, _27000_);
  and _30921_ (_27005_, _27004_, _26950_);
  nor _30922_ (_27006_, _26950_, _26489_);
  or _30923_ (_27007_, _27006_, _27005_);
  and _30924_ (_17315_, _27007_, _27355_);
  and _30925_ (_27008_, _26925_, _25905_);
  nand _30926_ (_27009_, _27008_, _25514_);
  or _30927_ (_27010_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _30928_ (_27011_, _27010_, _26950_);
  and _30929_ (_27012_, _27011_, _27009_);
  nor _30930_ (_27013_, _26950_, _26482_);
  or _30931_ (_27014_, _27013_, _27012_);
  and _30932_ (_17324_, _27014_, _27355_);
  and _30933_ (_27015_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _30934_ (_27016_, _25240_, _25212_);
  and _30935_ (_27017_, _25344_, _25246_);
  or _30936_ (_27018_, _27017_, _27016_);
  and _30937_ (_27019_, _27018_, _27015_);
  nand _30938_ (_27020_, _27015_, _25424_);
  and _30939_ (_27021_, _27020_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _30940_ (_27022_, _27021_, _26925_);
  or _30941_ (_27023_, _27022_, _27019_);
  not _30942_ (_27024_, _25972_);
  nor _30943_ (_27025_, _27024_, _25514_);
  or _30944_ (_27026_, _25972_, _25738_);
  nand _30945_ (_27027_, _27026_, _26925_);
  or _30946_ (_27028_, _27027_, _27025_);
  and _30947_ (_27029_, _27028_, _27023_);
  or _30948_ (_27030_, _27029_, _26942_);
  nand _30949_ (_27031_, _26942_, _26475_);
  and _30950_ (_27032_, _27031_, _27355_);
  and _30951_ (_17332_, _27032_, _27030_);
  nor _30952_ (_27033_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _30953_ (_27034_, _27033_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _30954_ (_27035_, _25055_, _25115_);
  and _30955_ (_27036_, _25128_, _26922_);
  and _30956_ (_27037_, _27036_, _26939_);
  and _30957_ (_27038_, _27037_, _27035_);
  and _30958_ (_27039_, _27038_, _25450_);
  nor _30959_ (_27040_, _27039_, _27034_);
  not _30960_ (_27041_, _27040_);
  and _30961_ (_27042_, _27041_, _25441_);
  not _30962_ (_27043_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _30963_ (_27044_, _26590_, _27043_);
  and _30964_ (_27045_, _25128_, _25115_);
  and _30965_ (_27046_, _27045_, _25086_);
  not _30966_ (_27047_, _25521_);
  nor _30967_ (_27048_, _27047_, _25101_);
  and _30968_ (_27049_, _27048_, _27046_);
  and _30969_ (_27050_, _27049_, _25517_);
  or _30970_ (_27051_, _27050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _30971_ (_27052_, _27044_);
  and _30972_ (_27053_, _27052_, _27040_);
  nand _30973_ (_27054_, _27050_, _25514_);
  and _30974_ (_27055_, _27054_, _27053_);
  and _30975_ (_27056_, _27055_, _27051_);
  or _30976_ (_27057_, _27056_, _27044_);
  or _30977_ (_27058_, _27057_, _27042_);
  or _30978_ (_27059_, _27052_, _26678_);
  and _30979_ (_27060_, _27059_, _27058_);
  and _30980_ (_17824_, _27060_, _27355_);
  or _30981_ (_27061_, _27040_, _25562_);
  and _30982_ (_27062_, _27049_, _25055_);
  nor _30983_ (_27063_, _27062_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not _30984_ (_27064_, _27063_);
  not _30985_ (_27065_, _27053_);
  and _30986_ (_27066_, _27062_, _25514_);
  nor _30987_ (_27067_, _27066_, _27065_);
  and _30988_ (_27068_, _27067_, _27064_);
  nor _30989_ (_27069_, _27068_, _27044_);
  nand _30990_ (_27070_, _27069_, _27061_);
  or _30991_ (_27071_, _27052_, _26713_);
  and _30992_ (_27072_, _27071_, _27070_);
  and _30993_ (_19498_, _27072_, _27355_);
  nor _30994_ (_27073_, _27052_, _26745_);
  not _30995_ (_27074_, _27073_);
  or _30996_ (_27075_, _27040_, _25639_);
  nor _30997_ (_27076_, _27049_, _24029_);
  not _30998_ (_27077_, _27076_);
  not _30999_ (_27078_, _27049_);
  not _31000_ (_27079_, _26947_);
  nor _31001_ (_27080_, _27079_, _25514_);
  nor _31002_ (_27081_, _26947_, _24029_);
  nor _31003_ (_27082_, _27081_, _27080_);
  or _31004_ (_27083_, _27082_, _27078_);
  and _31005_ (_27084_, _27083_, _27040_);
  and _31006_ (_27085_, _27084_, _27077_);
  nor _31007_ (_27086_, _27085_, _27044_);
  nand _31008_ (_27087_, _27086_, _27075_);
  nand _31009_ (_27088_, _27087_, _27074_);
  and _31010_ (_19508_, _27088_, _27355_);
  or _31011_ (_27089_, _27040_, _25704_);
  and _31012_ (_27090_, _27049_, _25716_);
  and _31013_ (_27091_, _27090_, _25514_);
  nor _31014_ (_27092_, _27090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _31015_ (_27093_, _27092_, _27065_);
  not _31016_ (_27094_, _27093_);
  nor _31017_ (_27095_, _27094_, _27091_);
  nor _31018_ (_27096_, _27095_, _27044_);
  nand _31019_ (_27097_, _27096_, _27089_);
  and _31020_ (_27098_, _27044_, _26775_);
  not _31021_ (_27099_, _27098_);
  and _31022_ (_27100_, _27099_, _27097_);
  and _31023_ (_19518_, _27100_, _27355_);
  or _31024_ (_27101_, _27040_, _25769_);
  and _31025_ (_27102_, _27053_, _27078_);
  and _31026_ (_27103_, _27102_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _31027_ (_27104_, _25778_, _24015_);
  nor _31028_ (_27105_, _27104_, _25779_);
  and _31029_ (_27106_, _27049_, _27052_);
  not _31030_ (_27107_, _27106_);
  nor _31031_ (_27108_, _27107_, _27105_);
  and _31032_ (_27109_, _27108_, _27053_);
  nor _31033_ (_27110_, _27109_, _27103_);
  and _31034_ (_27111_, _27110_, _27052_);
  nand _31035_ (_27112_, _27111_, _27101_);
  and _31036_ (_27113_, _27044_, _26808_);
  not _31037_ (_27114_, _27113_);
  and _31038_ (_27115_, _27114_, _27112_);
  and _31039_ (_19528_, _27115_, _27355_);
  and _31040_ (_27116_, _27041_, _25830_);
  and _31041_ (_27117_, _27049_, _25838_);
  or _31042_ (_27118_, _27117_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _31043_ (_27119_, _27117_, _25514_);
  and _31044_ (_27120_, _27119_, _27053_);
  and _31045_ (_27121_, _27120_, _27118_);
  or _31046_ (_27122_, _27121_, _27044_);
  or _31047_ (_27123_, _27122_, _27116_);
  or _31048_ (_27124_, _27052_, _26837_);
  and _31049_ (_27125_, _27124_, _27123_);
  and _31050_ (_19539_, _27125_, _27355_);
  and _31051_ (_27126_, _27041_, _25898_);
  and _31052_ (_27127_, _27049_, _25905_);
  or _31053_ (_27128_, _27127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _31054_ (_27129_, _27127_, _25514_);
  and _31055_ (_27130_, _27129_, _27053_);
  and _31056_ (_27131_, _27130_, _27128_);
  or _31057_ (_27132_, _27131_, _27044_);
  or _31058_ (_27133_, _27132_, _27126_);
  or _31059_ (_27134_, _27052_, _26867_);
  and _31060_ (_27135_, _27134_, _27133_);
  and _31061_ (_19549_, _27135_, _27355_);
  or _31062_ (_27136_, _27040_, _25963_);
  and _31063_ (_27137_, _27049_, _25972_);
  nor _31064_ (_27138_, _27137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _31065_ (_27139_, _27138_);
  and _31066_ (_27140_, _27137_, _25514_);
  nor _31067_ (_27141_, _27140_, _27065_);
  and _31068_ (_27142_, _27141_, _27139_);
  nor _31069_ (_27143_, _27142_, _27044_);
  and _31070_ (_27144_, _27143_, _27136_);
  and _31071_ (_27145_, _27044_, _26898_);
  or _31072_ (_27146_, _27145_, _27144_);
  nor _31073_ (_19559_, _27146_, rst);
  and _31074_ (_27147_, _25085_, _25073_);
  and _31075_ (_27148_, _27045_, _25102_);
  and _31076_ (_27149_, _27148_, _27147_);
  and _31077_ (_27150_, _27149_, _25517_);
  nand _31078_ (_27151_, _27150_, _25514_);
  or _31079_ (_27152_, _27150_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _31080_ (_27153_, _27152_, _25521_);
  and _31081_ (_27154_, _27153_, _27151_);
  and _31082_ (_27155_, _26460_, _27035_);
  nand _31083_ (_27156_, _27155_, _26543_);
  or _31084_ (_27157_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _31085_ (_27158_, _27157_, _25450_);
  and _31086_ (_27159_, _27158_, _27156_);
  not _31087_ (_27160_, _25449_);
  and _31088_ (_27161_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _31089_ (_27162_, _27161_, rst);
  or _31090_ (_27163_, _27162_, _27159_);
  or _31091_ (_23900_, _27163_, _27154_);
  and _31092_ (_27164_, _27147_, _25130_);
  and _31093_ (_27165_, _27164_, _25517_);
  nand _31094_ (_27166_, _27165_, _25514_);
  or _31095_ (_27167_, _27165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _31096_ (_27168_, _27167_, _25521_);
  and _31097_ (_27169_, _27168_, _27166_);
  and _31098_ (_27170_, _26938_, _26459_);
  and _31099_ (_27171_, _27170_, _27035_);
  nand _31100_ (_27172_, _27171_, _26543_);
  or _31101_ (_27173_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _31102_ (_27174_, _27173_, _25450_);
  and _31103_ (_27175_, _27174_, _27172_);
  and _31104_ (_27176_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _31105_ (_27177_, _27176_, rst);
  or _31106_ (_27178_, _27177_, _27175_);
  or _31107_ (_23901_, _27178_, _27169_);
  and _31108_ (_27179_, _26922_, _25073_);
  and _31109_ (_27180_, _27179_, _27148_);
  and _31110_ (_27181_, _27180_, _25517_);
  nand _31111_ (_27182_, _27181_, _25514_);
  or _31112_ (_27183_, _27181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _31113_ (_27184_, _27183_, _25521_);
  and _31114_ (_27185_, _27184_, _27182_);
  and _31115_ (_27186_, _27036_, _26459_);
  and _31116_ (_27187_, _27186_, _27035_);
  not _31117_ (_27188_, _27187_);
  nor _31118_ (_27189_, _27188_, _26543_);
  and _31119_ (_27190_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _31120_ (_27191_, _27190_, _27189_);
  and _31121_ (_27192_, _27191_, _25450_);
  and _31122_ (_27193_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _31123_ (_27194_, _27193_, rst);
  or _31124_ (_27195_, _27194_, _27192_);
  or _31125_ (_23902_, _27195_, _27185_);
  and _31126_ (_27196_, _27179_, _25130_);
  and _31127_ (_27197_, _27196_, _25517_);
  nand _31128_ (_27198_, _27197_, _25514_);
  or _31129_ (_27199_, _27197_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _31130_ (_27200_, _27199_, _25521_);
  and _31131_ (_27201_, _27200_, _27198_);
  nor _31132_ (_27202_, _25128_, _25085_);
  and _31133_ (_27203_, _26459_, _27202_);
  and _31134_ (_27204_, _27203_, _27035_);
  not _31135_ (_27205_, _27204_);
  nor _31136_ (_27206_, _27205_, _26543_);
  and _31137_ (_27207_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _31138_ (_27208_, _27207_, _27206_);
  and _31139_ (_27209_, _27208_, _25450_);
  and _31140_ (_27210_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _31141_ (_27211_, _27210_, rst);
  or _31142_ (_27212_, _27211_, _27209_);
  or _31143_ (_23903_, _27212_, _27201_);
  or _31144_ (_27213_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _31145_ (_27214_, _27213_, _25521_);
  nand _31146_ (_27215_, _27155_, _25514_);
  and _31147_ (_27216_, _27215_, _27214_);
  nand _31148_ (_27217_, _27155_, _26521_);
  and _31149_ (_27218_, _27217_, _25450_);
  and _31150_ (_27219_, _27218_, _27213_);
  not _31151_ (_27220_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _31152_ (_27221_, _25449_, _27220_);
  or _31153_ (_27222_, _27221_, rst);
  or _31154_ (_27223_, _27222_, _27219_);
  or _31155_ (_24987_, _27223_, _27216_);
  and _31156_ (_27224_, _25650_, _26595_);
  and _31157_ (_27225_, _27224_, _26460_);
  nand _31158_ (_27226_, _27225_, _25514_);
  or _31159_ (_27227_, _27225_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _31160_ (_27228_, _27227_, _25521_);
  and _31161_ (_27229_, _27228_, _27226_);
  nand _31162_ (_27230_, _27155_, _26512_);
  or _31163_ (_27231_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _31164_ (_27232_, _27231_, _25450_);
  and _31165_ (_27233_, _27232_, _27230_);
  and _31166_ (_27234_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _31167_ (_27235_, _27234_, rst);
  or _31168_ (_27236_, _27235_, _27233_);
  or _31169_ (_24989_, _27236_, _27229_);
  not _31170_ (_27237_, _25780_);
  nand _31171_ (_27238_, _27149_, _27237_);
  and _31172_ (_27239_, _27238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not _31173_ (_27240_, _25719_);
  and _31174_ (_27241_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _31175_ (_27242_, _27241_, _25718_);
  and _31176_ (_27243_, _27242_, _27149_);
  or _31177_ (_27244_, _27243_, _27239_);
  and _31178_ (_27245_, _27244_, _25521_);
  nand _31179_ (_27246_, _27155_, _26505_);
  or _31180_ (_27247_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _31181_ (_27248_, _27247_, _25450_);
  and _31182_ (_27249_, _27248_, _27246_);
  and _31183_ (_27250_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _31184_ (_27251_, _27250_, rst);
  or _31185_ (_27252_, _27251_, _27249_);
  or _31186_ (_24991_, _27252_, _27245_);
  nand _31187_ (_27253_, _27149_, _25020_);
  and _31188_ (_27254_, _27253_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _31189_ (_27255_, _27237_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _31190_ (_27256_, _27255_, _25779_);
  and _31191_ (_27257_, _27256_, _27149_);
  or _31192_ (_27258_, _27257_, _27254_);
  and _31193_ (_27259_, _27258_, _25521_);
  nand _31194_ (_27260_, _27155_, _26497_);
  or _31195_ (_27261_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _31196_ (_27262_, _27261_, _25450_);
  and _31197_ (_27263_, _27262_, _27260_);
  and _31198_ (_27264_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _31199_ (_27265_, _27264_, rst);
  or _31200_ (_27266_, _27265_, _27263_);
  or _31201_ (_24993_, _27266_, _27259_);
  not _31202_ (_27267_, _27149_);
  or _31203_ (_27268_, _27267_, _25840_);
  and _31204_ (_27269_, _27268_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _31205_ (_27270_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _31206_ (_27271_, _27270_, _25843_);
  and _31207_ (_27272_, _27271_, _27149_);
  or _31208_ (_27273_, _27272_, _27269_);
  and _31209_ (_27274_, _27273_, _25521_);
  nand _31210_ (_27275_, _27155_, _26489_);
  or _31211_ (_27276_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _31212_ (_27277_, _27276_, _25450_);
  and _31213_ (_27278_, _27277_, _27275_);
  and _31214_ (_27279_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _31215_ (_27280_, _27279_, rst);
  or _31216_ (_27281_, _27280_, _27278_);
  or _31217_ (_24995_, _27281_, _27274_);
  and _31218_ (_27282_, _27149_, _25905_);
  nand _31219_ (_27283_, _27282_, _25514_);
  or _31220_ (_27284_, _27282_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _31221_ (_27285_, _27284_, _25521_);
  and _31222_ (_27286_, _27285_, _27283_);
  nand _31223_ (_27287_, _27155_, _26482_);
  or _31224_ (_27288_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _31225_ (_27289_, _27288_, _25450_);
  and _31226_ (_27290_, _27289_, _27287_);
  and _31227_ (_27291_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _31228_ (_27292_, _27291_, rst);
  or _31229_ (_27293_, _27292_, _27290_);
  or _31230_ (_24997_, _27293_, _27286_);
  and _31231_ (_27295_, _27149_, _25972_);
  nand _31232_ (_27297_, _27295_, _25514_);
  or _31233_ (_27299_, _27295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _31234_ (_27300_, _27299_, _25521_);
  and _31235_ (_27302_, _27300_, _27297_);
  nand _31236_ (_27304_, _27155_, _26475_);
  or _31237_ (_27306_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _31238_ (_27308_, _27306_, _25450_);
  and _31239_ (_27309_, _27308_, _27304_);
  and _31240_ (_27310_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _31241_ (_27311_, _27310_, rst);
  or _31242_ (_27312_, _27311_, _27309_);
  or _31243_ (_24999_, _27312_, _27302_);
  and _31244_ (_27313_, _27164_, _25055_);
  nand _31245_ (_27314_, _27313_, _25514_);
  or _31246_ (_27315_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _31247_ (_27316_, _27315_, _25521_);
  and _31248_ (_27317_, _27316_, _27314_);
  nand _31249_ (_27318_, _27171_, _26521_);
  and _31250_ (_27319_, _27318_, _25450_);
  and _31251_ (_27320_, _27319_, _27315_);
  not _31252_ (_27321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _31253_ (_27322_, _25449_, _27321_);
  or _31254_ (_27323_, _27322_, rst);
  or _31255_ (_27324_, _27323_, _27320_);
  or _31256_ (_25001_, _27324_, _27317_);
  and _31257_ (_27325_, _27164_, _26947_);
  nand _31258_ (_27326_, _27325_, _25514_);
  or _31259_ (_27327_, _27325_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _31260_ (_27328_, _27327_, _25521_);
  and _31261_ (_27329_, _27328_, _27326_);
  nand _31262_ (_27330_, _27171_, _26512_);
  or _31263_ (_27331_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _31264_ (_27332_, _27331_, _25450_);
  and _31265_ (_27333_, _27332_, _27330_);
  and _31266_ (_27334_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _31267_ (_27335_, _27334_, rst);
  or _31268_ (_27336_, _27335_, _27333_);
  or _31269_ (_25003_, _27336_, _27329_);
  and _31270_ (_27337_, _27164_, _25716_);
  nand _31271_ (_27338_, _27337_, _25514_);
  or _31272_ (_27339_, _27337_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _31273_ (_27340_, _27339_, _25521_);
  and _31274_ (_27342_, _27340_, _27338_);
  nand _31275_ (_27344_, _27171_, _26505_);
  or _31276_ (_27346_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _31277_ (_27348_, _27346_, _25450_);
  and _31278_ (_27350_, _27348_, _27344_);
  and _31279_ (_27352_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _31280_ (_27354_, _27352_, rst);
  or _31281_ (_27356_, _27354_, _27350_);
  or _31282_ (_25005_, _27356_, _27342_);
  and _31283_ (_27358_, _27164_, _25778_);
  nand _31284_ (_27360_, _27358_, _25514_);
  or _31285_ (_27361_, _27358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _31286_ (_27362_, _27361_, _25521_);
  and _31287_ (_27363_, _27362_, _27360_);
  nand _31288_ (_27364_, _27171_, _26497_);
  or _31289_ (_27365_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _31290_ (_27366_, _27365_, _25450_);
  and _31291_ (_27367_, _27366_, _27364_);
  and _31292_ (_27368_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _31293_ (_27369_, _27368_, rst);
  or _31294_ (_27370_, _27369_, _27367_);
  or _31295_ (_25007_, _27370_, _27363_);
  and _31296_ (_27371_, _27164_, _25838_);
  nand _31297_ (_27372_, _27371_, _25514_);
  or _31298_ (_27373_, _27371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _31299_ (_27374_, _27373_, _25521_);
  and _31300_ (_27375_, _27374_, _27372_);
  nand _31301_ (_27376_, _27171_, _26489_);
  or _31302_ (_27377_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _31303_ (_27378_, _27377_, _25450_);
  and _31304_ (_27379_, _27378_, _27376_);
  and _31305_ (_27380_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _31306_ (_27381_, _27380_, rst);
  or _31307_ (_27382_, _27381_, _27379_);
  or _31308_ (_25009_, _27382_, _27375_);
  and _31309_ (_27383_, _27164_, _25905_);
  nand _31310_ (_27384_, _27383_, _25514_);
  or _31311_ (_27385_, _27383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _31312_ (_27386_, _27385_, _25521_);
  and _31313_ (_27387_, _27386_, _27384_);
  nand _31314_ (_27388_, _27171_, _26482_);
  or _31315_ (_27389_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _31316_ (_27390_, _27389_, _25450_);
  and _31317_ (_27391_, _27390_, _27388_);
  and _31318_ (_27392_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _31319_ (_27393_, _27392_, rst);
  or _31320_ (_27394_, _27393_, _27391_);
  or _31321_ (_25011_, _27394_, _27387_);
  and _31322_ (_27395_, _27164_, _25972_);
  nand _31323_ (_27396_, _27395_, _25514_);
  or _31324_ (_27397_, _27395_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _31325_ (_27398_, _27397_, _25521_);
  and _31326_ (_27399_, _27398_, _27396_);
  nand _31327_ (_27400_, _27171_, _26475_);
  or _31328_ (_27401_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _31329_ (_27402_, _27401_, _25450_);
  and _31330_ (_27403_, _27402_, _27400_);
  and _31331_ (_27404_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _31332_ (_27405_, _27404_, rst);
  or _31333_ (_27406_, _27405_, _27403_);
  or _31334_ (_25013_, _27406_, _27399_);
  and _31335_ (_27407_, _27180_, _25055_);
  nand _31336_ (_27408_, _27407_, _25514_);
  or _31337_ (_27409_, _27187_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _31338_ (_27410_, _27409_, _25521_);
  and _31339_ (_27411_, _27410_, _27408_);
  nand _31340_ (_27412_, _27187_, _26521_);
  and _31341_ (_27413_, _27412_, _25450_);
  and _31342_ (_27414_, _27413_, _27409_);
  not _31343_ (_27415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _31344_ (_27416_, _25449_, _27415_);
  or _31345_ (_27417_, _27416_, rst);
  or _31346_ (_27418_, _27417_, _27414_);
  or _31347_ (_25015_, _27418_, _27411_);
  and _31348_ (_27419_, _27180_, _26947_);
  nand _31349_ (_27420_, _27419_, _25514_);
  or _31350_ (_27421_, _27419_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _31351_ (_27422_, _27421_, _25521_);
  and _31352_ (_27423_, _27422_, _27420_);
  nor _31353_ (_27424_, _27188_, _26512_);
  and _31354_ (_27425_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _31355_ (_27426_, _27425_, _27424_);
  and _31356_ (_27427_, _27426_, _25450_);
  and _31357_ (_27428_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _31358_ (_27429_, _27428_, rst);
  or _31359_ (_27430_, _27429_, _27427_);
  or _31360_ (_25017_, _27430_, _27423_);
  and _31361_ (_27431_, _27180_, _25716_);
  nand _31362_ (_27432_, _27431_, _25514_);
  or _31363_ (_27433_, _27431_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _31364_ (_27434_, _27433_, _25521_);
  and _31365_ (_27435_, _27434_, _27432_);
  nor _31366_ (_27436_, _27188_, _26505_);
  and _31367_ (_27437_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _31368_ (_27438_, _27437_, _27436_);
  and _31369_ (_27439_, _27438_, _25450_);
  and _31370_ (_27440_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _31371_ (_27441_, _27440_, rst);
  or _31372_ (_27442_, _27441_, _27439_);
  or _31373_ (_25019_, _27442_, _27435_);
  and _31374_ (_27443_, _27180_, _25778_);
  nand _31375_ (_27444_, _27443_, _25514_);
  or _31376_ (_27445_, _27443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _31377_ (_27446_, _27445_, _25521_);
  and _31378_ (_27447_, _27446_, _27444_);
  nor _31379_ (_27448_, _27188_, _26497_);
  and _31380_ (_27449_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _31381_ (_27450_, _27449_, _27448_);
  and _31382_ (_27451_, _27450_, _25450_);
  and _31383_ (_27452_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _31384_ (_27453_, _27452_, rst);
  or _31385_ (_27454_, _27453_, _27451_);
  or _31386_ (_25021_, _27454_, _27447_);
  and _31387_ (_27455_, _27180_, _25838_);
  nand _31388_ (_27456_, _27455_, _25514_);
  or _31389_ (_27457_, _27455_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _31390_ (_27458_, _27457_, _25521_);
  and _31391_ (_27459_, _27458_, _27456_);
  nor _31392_ (_27460_, _27188_, _26489_);
  and _31393_ (_27461_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _31394_ (_27462_, _27461_, _27460_);
  and _31395_ (_27463_, _27462_, _25450_);
  and _31396_ (_27464_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _31397_ (_27465_, _27464_, rst);
  or _31398_ (_27466_, _27465_, _27463_);
  or _31399_ (_25023_, _27466_, _27459_);
  and _31400_ (_27467_, _27180_, _25905_);
  nand _31401_ (_27468_, _27467_, _25514_);
  or _31402_ (_27469_, _27467_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _31403_ (_27470_, _27469_, _25521_);
  and _31404_ (_27471_, _27470_, _27468_);
  nor _31405_ (_27472_, _27188_, _26482_);
  and _31406_ (_27473_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _31407_ (_27474_, _27473_, _27472_);
  and _31408_ (_27475_, _27474_, _25450_);
  and _31409_ (_27476_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _31410_ (_27477_, _27476_, rst);
  or _31411_ (_27478_, _27477_, _27475_);
  or _31412_ (_25025_, _27478_, _27471_);
  and _31413_ (_27479_, _27180_, _25972_);
  nand _31414_ (_27480_, _27479_, _25514_);
  or _31415_ (_27481_, _27479_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _31416_ (_27482_, _27481_, _25521_);
  and _31417_ (_27483_, _27482_, _27480_);
  nor _31418_ (_27484_, _27188_, _26475_);
  and _31419_ (_27485_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _31420_ (_27486_, _27485_, _27484_);
  and _31421_ (_27487_, _27486_, _25450_);
  and _31422_ (_27488_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _31423_ (_27489_, _27488_, rst);
  or _31424_ (_27490_, _27489_, _27487_);
  or _31425_ (_25027_, _27490_, _27483_);
  and _31426_ (_27491_, _27196_, _25055_);
  nand _31427_ (_27492_, _27491_, _25514_);
  or _31428_ (_27493_, _27204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _31429_ (_27494_, _27493_, _25521_);
  and _31430_ (_27495_, _27494_, _27492_);
  nand _31431_ (_27496_, _27204_, _26521_);
  and _31432_ (_27497_, _27496_, _25450_);
  and _31433_ (_27498_, _27497_, _27493_);
  not _31434_ (_27499_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _31435_ (_27500_, _25449_, _27499_);
  or _31436_ (_27501_, _27500_, rst);
  or _31437_ (_27502_, _27501_, _27498_);
  or _31438_ (_25029_, _27502_, _27495_);
  and _31439_ (_27503_, _27196_, _26947_);
  nand _31440_ (_27504_, _27503_, _25514_);
  or _31441_ (_27505_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _31442_ (_27506_, _27505_, _25521_);
  and _31443_ (_27507_, _27506_, _27504_);
  nor _31444_ (_27508_, _27205_, _26512_);
  and _31445_ (_27509_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _31446_ (_27510_, _27509_, _27508_);
  and _31447_ (_27511_, _27510_, _25450_);
  and _31448_ (_27512_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _31449_ (_27513_, _27512_, rst);
  or _31450_ (_27514_, _27513_, _27511_);
  or _31451_ (_25031_, _27514_, _27507_);
  and _31452_ (_27515_, _27196_, _25716_);
  nand _31453_ (_27516_, _27515_, _25514_);
  or _31454_ (_27517_, _27515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _31455_ (_27518_, _27517_, _25521_);
  and _31456_ (_27519_, _27518_, _27516_);
  nor _31457_ (_27520_, _27205_, _26505_);
  and _31458_ (_27521_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _31459_ (_27522_, _27521_, _27520_);
  and _31460_ (_27523_, _27522_, _25450_);
  and _31461_ (_27524_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _31462_ (_27525_, _27524_, rst);
  or _31463_ (_27526_, _27525_, _27523_);
  or _31464_ (_25033_, _27526_, _27519_);
  and _31465_ (_27527_, _27196_, _25778_);
  nand _31466_ (_27528_, _27527_, _25514_);
  or _31467_ (_27529_, _27527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _31468_ (_27530_, _27529_, _25521_);
  and _31469_ (_27531_, _27530_, _27528_);
  nor _31470_ (_27532_, _27205_, _26497_);
  and _31471_ (_27533_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _31472_ (_27534_, _27533_, _27532_);
  and _31473_ (_27535_, _27534_, _25450_);
  and _31474_ (_27536_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _31475_ (_27537_, _27536_, rst);
  or _31476_ (_27538_, _27537_, _27535_);
  or _31477_ (_25035_, _27538_, _27531_);
  and _31478_ (_27539_, _27196_, _25838_);
  nand _31479_ (_27540_, _27539_, _25514_);
  or _31480_ (_27541_, _27539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _31481_ (_27542_, _27541_, _25521_);
  and _31482_ (_27543_, _27542_, _27540_);
  nor _31483_ (_27544_, _27205_, _26489_);
  and _31484_ (_27545_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _31485_ (_27546_, _27545_, _27544_);
  and _31486_ (_27547_, _27546_, _25450_);
  and _31487_ (_27548_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _31488_ (_27549_, _27548_, rst);
  or _31489_ (_27550_, _27549_, _27547_);
  or _31490_ (_25037_, _27550_, _27543_);
  and _31491_ (_27551_, _27196_, _25905_);
  nand _31492_ (_27552_, _27551_, _25514_);
  or _31493_ (_27553_, _27551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _31494_ (_27554_, _27553_, _25521_);
  and _31495_ (_27555_, _27554_, _27552_);
  nor _31496_ (_27556_, _27205_, _26482_);
  and _31497_ (_27557_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _31498_ (_27558_, _27557_, _27556_);
  and _31499_ (_27559_, _27558_, _25450_);
  and _31500_ (_27560_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _31501_ (_27561_, _27560_, rst);
  or _31502_ (_27562_, _27561_, _27559_);
  or _31503_ (_25039_, _27562_, _27555_);
  and _31504_ (_27563_, _27196_, _25972_);
  nand _31505_ (_27564_, _27563_, _25514_);
  or _31506_ (_27565_, _27563_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _31507_ (_27566_, _27565_, _25521_);
  and _31508_ (_27567_, _27566_, _27564_);
  nor _31509_ (_27568_, _27205_, _26475_);
  and _31510_ (_27569_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _31511_ (_27570_, _27569_, _27568_);
  and _31512_ (_27571_, _27570_, _25450_);
  and _31513_ (_27572_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _31514_ (_27573_, _27572_, rst);
  or _31515_ (_27574_, _27573_, _27571_);
  or _31516_ (_25041_, _27574_, _27567_);
  and _31517_ (_25436_, t0_i, _27355_);
  and _31518_ (_25439_, t1_i, _27355_);
  not _31519_ (_27575_, _25450_);
  nor _31520_ (_27576_, _27575_, _25115_);
  and _31521_ (_27577_, _27576_, _25778_);
  and _31522_ (_27578_, _27577_, _26460_);
  nand _31523_ (_27579_, _27578_, _26543_);
  not _31524_ (_27580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _31525_ (_27581_, _27580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _31526_ (_27582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _31527_ (_27583_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _27582_);
  nor _31528_ (_27584_, _27583_, _27581_);
  nor _31529_ (_27585_, _25020_, _25115_);
  and _31530_ (_27586_, _27585_, _26461_);
  and _31531_ (_27587_, _27586_, _25450_);
  nor _31532_ (_27588_, _27587_, _27584_);
  not _31533_ (_27589_, _27588_);
  and _31534_ (_27590_, _27589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _31535_ (_27591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _31536_ (_27592_, t1_i);
  and _31537_ (_27593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _27592_);
  nor _31538_ (_27594_, _27593_, _27591_);
  not _31539_ (_27595_, _27594_);
  not _31540_ (_27596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _31541_ (_27597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _27596_);
  nor _31542_ (_27598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _31543_ (_27599_, _27598_);
  and _31544_ (_27600_, _27599_, _27597_);
  and _31545_ (_27601_, _27600_, _27595_);
  and _31546_ (_27602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _31547_ (_27603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _31548_ (_27604_, _27603_, _27602_);
  and _31549_ (_27605_, _27604_, _27601_);
  and _31550_ (_27606_, _27605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _31551_ (_27607_, _27606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _31552_ (_27608_, _27607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _31553_ (_27609_, _27608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _31554_ (_27610_, _27604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _31555_ (_27611_, _27610_, _27601_);
  and _31556_ (_27612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _31557_ (_27613_, _27612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _31558_ (_27614_, _27613_, _27611_);
  nor _31559_ (_27615_, _27614_, _27584_);
  and _31560_ (_27616_, _27615_, _27609_);
  and _31561_ (_27617_, _27614_, _27581_);
  and _31562_ (_27618_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _31563_ (_27619_, _27618_, _27616_);
  nor _31564_ (_27620_, _27619_, _27587_);
  or _31565_ (_27621_, _27620_, _27590_);
  or _31566_ (_27622_, _27621_, _27578_);
  and _31567_ (_27623_, _27622_, _27355_);
  and _31568_ (_25442_, _27623_, _27579_);
  and _31569_ (_27624_, _27578_, _27355_);
  and _31570_ (_27625_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _31571_ (_27626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _31572_ (_27627_, _27626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _31573_ (_27628_, _27627_, _27611_);
  and _31574_ (_27629_, _27628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _31575_ (_27630_, _27629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _31576_ (_27631_, _27630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _31577_ (_27632_, _27631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _31578_ (_27633_, _27632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _31579_ (_27634_, _27632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _31580_ (_27635_, _27634_, _27613_);
  not _31581_ (_27636_, _27583_);
  nor _31582_ (_27637_, _27613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _31583_ (_27638_, _27637_, _27636_);
  nor _31584_ (_27639_, _27638_, _27635_);
  and _31585_ (_27640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _31586_ (_27641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _31587_ (_27642_, _27641_);
  nor _31588_ (_27643_, _27634_, _27642_);
  or _31589_ (_27644_, _27643_, _27640_);
  or _31590_ (_27645_, _27644_, _27639_);
  nand _31591_ (_27646_, _27645_, _27633_);
  nor _31592_ (_27647_, _27646_, _27587_);
  not _31593_ (_27648_, _27587_);
  nor _31594_ (_27649_, _27648_, _26543_);
  or _31595_ (_27650_, _27649_, _27647_);
  nor _31596_ (_27651_, _27578_, rst);
  and _31597_ (_27652_, _27651_, _27650_);
  or _31598_ (_25445_, _27652_, _27625_);
  not _31599_ (_27653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _31600_ (_27654_, _27601_, _27653_);
  or _31601_ (_27655_, _27654_, _27635_);
  and _31602_ (_27656_, _27655_, _27583_);
  or _31603_ (_27657_, _27654_, _27634_);
  and _31604_ (_27658_, _27657_, _27641_);
  nand _31605_ (_27659_, _27601_, _27580_);
  and _31606_ (_27660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _31607_ (_27661_, _27660_, _27659_);
  or _31608_ (_27662_, _27661_, _27617_);
  or _31609_ (_27663_, _27662_, _27658_);
  nor _31610_ (_27664_, _27663_, _27656_);
  nor _31611_ (_27665_, _27664_, _27587_);
  and _31612_ (_25448_, _27665_, _27651_);
  and _31613_ (_27666_, _27576_, _25716_);
  and _31614_ (_27667_, _27666_, _26460_);
  not _31615_ (_27668_, _27667_);
  and _31616_ (_27669_, _27576_, _25838_);
  and _31617_ (_27670_, _27669_, _26460_);
  nor _31618_ (_27671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _31619_ (_27672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _31620_ (_27673_, t0_i);
  and _31621_ (_27674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _27673_);
  nor _31622_ (_27675_, _27674_, _27672_);
  not _31623_ (_27676_, _27675_);
  not _31624_ (_27677_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _31625_ (_27678_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _31626_ (_27679_, _27678_, _27677_);
  and _31627_ (_27680_, _27679_, _27676_);
  not _31628_ (_27681_, _27680_);
  and _31629_ (_27682_, _27681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _31630_ (_27683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _31631_ (_27684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _31632_ (_27685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _31633_ (_27686_, _27685_, _27684_);
  and _31634_ (_27687_, _27686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _31635_ (_27688_, _27687_, _27680_);
  and _31636_ (_27689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _31637_ (_27690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _31638_ (_27691_, _27690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _31639_ (_27692_, _27691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _31640_ (_27693_, _27692_, _27689_);
  and _31641_ (_27694_, _27693_, _27688_);
  and _31642_ (_27695_, _27694_, _27683_);
  or _31643_ (_27696_, _27695_, _27682_);
  and _31644_ (_27697_, _27696_, _27671_);
  and _31645_ (_27698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _31646_ (_27699_, _27698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _31647_ (_27700_, _27699_, _27688_);
  not _31648_ (_27701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _31649_ (_27702_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _27701_);
  and _31650_ (_27703_, _27693_, _27683_);
  and _31651_ (_27704_, _27703_, _27702_);
  or _31652_ (_27705_, _27704_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _31653_ (_27706_, _27705_, _27700_);
  not _31654_ (_27707_, _27671_);
  and _31655_ (_27708_, _27682_, _27707_);
  or _31656_ (_27709_, _27708_, _27706_);
  or _31657_ (_27710_, _27709_, _27697_);
  nand _31658_ (_27711_, _27710_, _27355_);
  nor _31659_ (_27712_, _27711_, _27670_);
  and _31660_ (_25451_, _27712_, _27668_);
  nand _31661_ (_27713_, _27667_, _26543_);
  not _31662_ (_27714_, _27670_);
  or _31663_ (_27715_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _31664_ (_27716_, _27671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _31665_ (_27717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _31666_ (_27718_, _27717_, _27688_);
  or _31667_ (_27719_, _27718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _31668_ (_27720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _31669_ (_27721_, _27720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _31670_ (_27722_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _31671_ (_27723_, _27722_, _27700_);
  and _31672_ (_27724_, _27723_, _27707_);
  or _31673_ (_27725_, _27724_, _27670_);
  and _31674_ (_27726_, _27725_, _27719_);
  or _31675_ (_27727_, _27726_, _27716_);
  and _31676_ (_27728_, _27727_, _27715_);
  or _31677_ (_27729_, _27728_, _27667_);
  and _31678_ (_27730_, _27729_, _27355_);
  and _31679_ (_25454_, _27730_, _27713_);
  nand _31680_ (_27731_, _27670_, _26543_);
  or _31681_ (_27732_, _27721_, _27702_);
  not _31682_ (_27733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _31683_ (_27734_, _27699_, _27687_);
  and _31684_ (_27735_, _27680_, _27701_);
  and _31685_ (_27736_, _27735_, _27734_);
  and _31686_ (_27737_, _27736_, _27693_);
  and _31687_ (_27738_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _31688_ (_27739_, _27738_, _27733_);
  and _31689_ (_27740_, _27738_, _27733_);
  or _31690_ (_27741_, _27740_, _27739_);
  and _31691_ (_27742_, _27741_, _27732_);
  and _31692_ (_27743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _31693_ (_27744_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _31694_ (_27745_, _27744_, _27692_);
  and _31695_ (_27746_, _27745_, _27689_);
  and _31696_ (_27747_, _27746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _31697_ (_27748_, _27747_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _31698_ (_27749_, _27744_, _27703_);
  and _31699_ (_27750_, _27749_, _27748_);
  and _31700_ (_27751_, _27750_, _27743_);
  and _31701_ (_27752_, _27694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _31702_ (_27753_, _27752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _31703_ (_27754_, _27695_, _27707_);
  and _31704_ (_27755_, _27754_, _27753_);
  or _31705_ (_27756_, _27755_, _27751_);
  or _31706_ (_27757_, _27756_, _27742_);
  or _31707_ (_27758_, _27757_, _27670_);
  and _31708_ (_27759_, _27758_, _27668_);
  and _31709_ (_27760_, _27759_, _27731_);
  and _31710_ (_27761_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _31711_ (_27762_, _27761_, _27760_);
  and _31712_ (_25457_, _27762_, _27355_);
  or _31713_ (_27763_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _31714_ (_27764_, _27743_, _27355_);
  and _31715_ (_27765_, _27764_, _27763_);
  not _31716_ (_27766_, _27744_);
  or _31717_ (_27767_, _27766_, _27703_);
  nand _31718_ (_27768_, _27767_, _27765_);
  nor _31719_ (_27769_, _27768_, _27670_);
  and _31720_ (_25460_, _27769_, _27668_);
  and _31721_ (_27770_, _27576_, _26462_);
  or _31722_ (_27771_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _31723_ (_27772_, _27771_, _27355_);
  nand _31724_ (_27773_, _27770_, _26543_);
  and _31725_ (_25463_, _27773_, _27772_);
  nor _31726_ (_27774_, _26521_, rst);
  or _31727_ (_27775_, _27774_, _27651_);
  and _31728_ (_27776_, _27601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _31729_ (_27777_, _27601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _31730_ (_27778_, _27777_, _27776_);
  and _31731_ (_27779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _31732_ (_27780_, _27779_, _27587_);
  and _31733_ (_27781_, _27780_, _27778_);
  and _31734_ (_27782_, _27613_, _27610_);
  and _31735_ (_27783_, _27782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _31736_ (_27784_, _27783_, _27581_);
  nor _31737_ (_27785_, _27784_, _27587_);
  or _31738_ (_27786_, _27785_, _27578_);
  not _31739_ (_27787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _31740_ (_27788_, _27780_, _27787_);
  or _31741_ (_27789_, _27788_, _27786_);
  or _31742_ (_27790_, _27789_, _27781_);
  and _31743_ (_26040_, _27790_, _27775_);
  and _31744_ (_27791_, _27776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _31745_ (_27792_, _27776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _31746_ (_27793_, _27792_, _27791_);
  nand _31747_ (_27794_, _27793_, _27780_);
  or _31748_ (_27795_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _31749_ (_27796_, _27795_, _27794_);
  and _31750_ (_27797_, _27608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _31751_ (_27798_, _27797_, _27581_);
  nand _31752_ (_27799_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _31753_ (_27800_, _27799_, _27587_);
  or _31754_ (_27801_, _27800_, _27578_);
  or _31755_ (_27802_, _27801_, _27796_);
  nand _31756_ (_27803_, _27578_, _26512_);
  and _31757_ (_27804_, _27803_, _27355_);
  and _31758_ (_26042_, _27804_, _27802_);
  not _31759_ (_27805_, _26505_);
  and _31760_ (_27806_, _27624_, _27805_);
  nor _31761_ (_27807_, _27791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _31762_ (_27808_, _27776_, _27602_);
  or _31763_ (_27809_, _27808_, _27807_);
  nand _31764_ (_27810_, _27809_, _27780_);
  or _31765_ (_27811_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _31766_ (_27812_, _27811_, _27810_);
  nand _31767_ (_27813_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _31768_ (_27814_, _27813_, _27587_);
  or _31769_ (_27815_, _27814_, _27812_);
  and _31770_ (_27816_, _27815_, _27651_);
  or _31771_ (_26044_, _27816_, _27806_);
  not _31772_ (_27817_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _31773_ (_27818_, _27780_, _27817_);
  or _31774_ (_27819_, _27808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _31775_ (_27820_, _27779_, _27605_);
  and _31776_ (_27821_, _27820_, _27819_);
  and _31777_ (_27822_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _31778_ (_27823_, _27822_, _27821_);
  nor _31779_ (_27824_, _27823_, _27587_);
  or _31780_ (_27825_, _27824_, _27818_);
  and _31781_ (_27826_, _27825_, _27651_);
  not _31782_ (_27827_, _26497_);
  and _31783_ (_27828_, _27624_, _27827_);
  or _31784_ (_26046_, _27828_, _27826_);
  not _31785_ (_27829_, _26489_);
  and _31786_ (_27830_, _27624_, _27829_);
  and _31787_ (_27831_, _27617_, _27648_);
  and _31788_ (_27832_, _27831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _31789_ (_27833_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _31790_ (_27834_, _27605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _31791_ (_27835_, _27834_, _27611_);
  nand _31792_ (_27836_, _27835_, _27780_);
  and _31793_ (_27837_, _27836_, _27833_);
  or _31794_ (_27838_, _27837_, _27832_);
  and _31795_ (_27839_, _27838_, _27651_);
  or _31796_ (_26048_, _27839_, _27830_);
  not _31797_ (_27840_, _26482_);
  and _31798_ (_27841_, _27624_, _27840_);
  and _31799_ (_27842_, _27589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _31800_ (_27843_, _27611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _31801_ (_27844_, _27611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _31802_ (_27845_, _27844_, _27584_);
  and _31803_ (_27846_, _27845_, _27843_);
  and _31804_ (_27847_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _31805_ (_27848_, _27847_, _27846_);
  nor _31806_ (_27849_, _27848_, _27587_);
  or _31807_ (_27850_, _27849_, _27842_);
  and _31808_ (_27851_, _27850_, _27651_);
  or _31809_ (_26050_, _27851_, _27841_);
  not _31810_ (_27852_, _26475_);
  and _31811_ (_27853_, _27624_, _27852_);
  and _31812_ (_27854_, _27782_, _27601_);
  and _31813_ (_27855_, _27581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _31814_ (_27856_, _27855_, _27854_);
  nor _31815_ (_27857_, _27856_, _27587_);
  or _31816_ (_27858_, _27588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _31817_ (_27859_, _27844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _31818_ (_27860_, _27859_, _27608_);
  nand _31819_ (_27861_, _27860_, _27588_);
  and _31820_ (_27862_, _27861_, _27858_);
  or _31821_ (_27863_, _27862_, _27857_);
  and _31822_ (_27864_, _27863_, _27651_);
  or _31823_ (_26052_, _27864_, _27853_);
  and _31824_ (_27865_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _31825_ (_27866_, _27641_, _27611_);
  and _31826_ (_27867_, _27854_, _27583_);
  nor _31827_ (_27868_, _27867_, _27866_);
  and _31828_ (_27869_, _27868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _31829_ (_27870_, _27868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _31830_ (_27871_, _27870_, _27869_);
  or _31831_ (_27872_, _27871_, _27587_);
  nand _31832_ (_27873_, _27587_, _26521_);
  and _31833_ (_27874_, _27873_, _27651_);
  and _31834_ (_27875_, _27874_, _27872_);
  or _31835_ (_26054_, _27875_, _27865_);
  and _31836_ (_27876_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _31837_ (_27877_, _27587_, _26512_);
  and _31838_ (_27878_, _27783_, _27601_);
  nor _31839_ (_27879_, _27878_, _27636_);
  and _31840_ (_27880_, _27582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _31841_ (_27881_, _27880_, _27611_);
  nor _31842_ (_27882_, _27881_, _27583_);
  nor _31843_ (_27883_, _27882_, _27879_);
  or _31844_ (_27884_, _27883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _31845_ (_27885_, _27883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _31846_ (_27886_, _27885_, _27884_);
  or _31847_ (_27887_, _27886_, _27587_);
  and _31848_ (_27888_, _27887_, _27651_);
  and _31849_ (_27889_, _27888_, _27877_);
  or _31850_ (_26056_, _27889_, _27876_);
  and _31851_ (_27890_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _31852_ (_27891_, _27587_, _26505_);
  and _31853_ (_27892_, _27626_, _27610_);
  and _31854_ (_27893_, _27892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _31855_ (_27894_, _27893_, _27601_);
  nor _31856_ (_27895_, _27894_, _27642_);
  or _31857_ (_27896_, _27895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand _31858_ (_27897_, _27628_, _27613_);
  and _31859_ (_27898_, _27897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or _31860_ (_27899_, _27898_, _27896_);
  and _31861_ (_27900_, _27899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _31862_ (_27901_, _27867_, _27626_);
  and _31863_ (_27902_, _27626_, _27641_);
  and _31864_ (_27903_, _27902_, _27611_);
  nor _31865_ (_27904_, _27903_, _27901_);
  nor _31866_ (_27905_, _27904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _31867_ (_27906_, _27905_, _27900_);
  or _31868_ (_27907_, _27906_, _27587_);
  and _31869_ (_27908_, _27907_, _27651_);
  and _31870_ (_27909_, _27908_, _27891_);
  or _31871_ (_26058_, _27909_, _27890_);
  and _31872_ (_27910_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _31873_ (_27911_, _27587_, _26497_);
  and _31874_ (_27912_, _27783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _31875_ (_27913_, _27912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _31876_ (_27914_, _27913_, _27601_);
  and _31877_ (_27915_, _27914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _31878_ (_27916_, _27914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _31879_ (_27917_, _27916_, _27583_);
  nor _31880_ (_27918_, _27917_, _27915_);
  and _31881_ (_27919_, _27896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _31882_ (_27920_, _27894_, _27641_);
  nor _31883_ (_27921_, _27920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _31884_ (_27922_, _27921_, _27919_);
  or _31885_ (_27923_, _27922_, _27918_);
  or _31886_ (_27924_, _27923_, _27587_);
  and _31887_ (_27925_, _27924_, _27651_);
  and _31888_ (_27926_, _27925_, _27911_);
  or _31889_ (_26060_, _27926_, _27910_);
  and _31890_ (_27927_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _31891_ (_27928_, _27587_, _26489_);
  and _31892_ (_27929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _31893_ (_27930_, _27914_, _27929_);
  or _31894_ (_27931_, _27915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _31895_ (_27932_, _27931_, _27583_);
  nor _31896_ (_27933_, _27932_, _27930_);
  and _31897_ (_27934_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _31898_ (_27935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _31899_ (_27936_, _27894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _31900_ (_27937_, _27936_, _27935_);
  or _31901_ (_27938_, _27936_, _27935_);
  and _31902_ (_27939_, _27938_, _27937_);
  and _31903_ (_27940_, _27939_, _27641_);
  or _31904_ (_27941_, _27940_, _27934_);
  or _31905_ (_27942_, _27941_, _27933_);
  or _31906_ (_27943_, _27942_, _27587_);
  and _31907_ (_27944_, _27943_, _27651_);
  and _31908_ (_27945_, _27944_, _27928_);
  or _31909_ (_26062_, _27945_, _27927_);
  and _31910_ (_27946_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _31911_ (_27947_, _27587_, _26482_);
  not _31912_ (_27948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _31913_ (_27949_, _27630_, _27641_);
  and _31914_ (_27950_, _27930_, _27583_);
  nor _31915_ (_27951_, _27950_, _27949_);
  and _31916_ (_27952_, _27951_, _27948_);
  nor _31917_ (_27953_, _27951_, _27948_);
  nor _31918_ (_27954_, _27953_, _27952_);
  or _31919_ (_27955_, _27954_, _27587_);
  and _31920_ (_27956_, _27955_, _27651_);
  and _31921_ (_27957_, _27956_, _27947_);
  or _31922_ (_26064_, _27957_, _27946_);
  and _31923_ (_27958_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _31924_ (_27959_, _27587_, _26475_);
  not _31925_ (_27960_, _27953_);
  nor _31926_ (_27961_, _27960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _31927_ (_27962_, _27960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _31928_ (_27963_, _27962_, _27961_);
  or _31929_ (_27964_, _27963_, _27587_);
  and _31930_ (_27965_, _27964_, _27651_);
  and _31931_ (_27966_, _27965_, _27959_);
  or _31932_ (_26066_, _27966_, _27958_);
  nor _31933_ (_27967_, _27681_, _27670_);
  or _31934_ (_27968_, _27967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _31935_ (_27969_, _27680_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _31936_ (_27970_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _31937_ (_27971_, _27970_, _27734_);
  nand _31938_ (_27972_, _27971_, _27969_);
  or _31939_ (_27973_, _27972_, _27670_);
  and _31940_ (_27974_, _27973_, _27968_);
  or _31941_ (_27975_, _27974_, _27667_);
  nand _31942_ (_27976_, _27667_, _26521_);
  and _31943_ (_27977_, _27976_, _27355_);
  and _31944_ (_26068_, _27977_, _27975_);
  nor _31945_ (_27978_, _27969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _31946_ (_27979_, _27969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _31947_ (_27980_, _27979_, _27978_);
  and _31948_ (_27981_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _31949_ (_27982_, _27981_, _27700_);
  nor _31950_ (_27983_, _27982_, _27980_);
  nor _31951_ (_27984_, _27983_, _27670_);
  and _31952_ (_27985_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _31953_ (_27986_, _27985_, _27984_);
  and _31954_ (_27987_, _27986_, _27668_);
  nor _31955_ (_27988_, _27668_, _26512_);
  or _31956_ (_27989_, _27988_, _27987_);
  and _31957_ (_26070_, _27989_, _27355_);
  nand _31958_ (_27990_, _27667_, _26505_);
  nor _31959_ (_27991_, _27979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _31960_ (_27992_, _27969_, _27684_);
  nor _31961_ (_27993_, _27992_, _27991_);
  and _31962_ (_27994_, _27721_, _27700_);
  and _31963_ (_27995_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _31964_ (_27996_, _27995_, _27993_);
  nor _31965_ (_27997_, _27996_, _27670_);
  and _31966_ (_27998_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _31967_ (_27999_, _27998_, _27997_);
  or _31968_ (_28000_, _27999_, _27667_);
  and _31969_ (_28001_, _28000_, _27355_);
  and _31970_ (_26072_, _28001_, _27990_);
  nand _31971_ (_28002_, _27667_, _26497_);
  and _31972_ (_28003_, _27686_, _27680_);
  nor _31973_ (_28004_, _27992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _31974_ (_28005_, _28004_, _28003_);
  and _31975_ (_28006_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _31976_ (_28007_, _28006_, _28005_);
  nor _31977_ (_28008_, _28007_, _27670_);
  and _31978_ (_28009_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _31979_ (_28010_, _28009_, _28008_);
  or _31980_ (_28011_, _28010_, _27667_);
  and _31981_ (_28012_, _28011_, _27355_);
  and _31982_ (_26074_, _28012_, _28002_);
  nor _31983_ (_28013_, _28003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _31984_ (_28014_, _28013_, _27688_);
  and _31985_ (_28015_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _31986_ (_28016_, _28015_, _28014_);
  or _31987_ (_28017_, _28016_, _27670_);
  or _31988_ (_28018_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _31989_ (_28019_, _28018_, _27668_);
  and _31990_ (_28020_, _28019_, _28017_);
  nor _31991_ (_28021_, _27668_, _26489_);
  or _31992_ (_28022_, _28021_, _28020_);
  and _31993_ (_26076_, _28022_, _27355_);
  nand _31994_ (_28023_, _27667_, _26482_);
  or _31995_ (_28024_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _31996_ (_28025_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _31997_ (_28026_, _27688_, _27707_);
  or _31998_ (_28027_, _28026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _31999_ (_28028_, _28026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _32000_ (_28029_, _28028_);
  or _32001_ (_28030_, _28029_, _27670_);
  and _32002_ (_28031_, _28030_, _28027_);
  or _32003_ (_28032_, _28031_, _28025_);
  and _32004_ (_28033_, _28032_, _28024_);
  or _32005_ (_28034_, _28033_, _27667_);
  and _32006_ (_28035_, _28034_, _27355_);
  and _32007_ (_26078_, _28035_, _28023_);
  and _32008_ (_28036_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _32009_ (_28037_, _28036_, _27680_);
  and _32010_ (_28038_, _28037_, _27734_);
  nor _32011_ (_28039_, _28029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _32012_ (_28040_, _28039_, _28038_);
  nor _32013_ (_28041_, _28040_, _27670_);
  and _32014_ (_28042_, _28030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _32015_ (_28043_, _28042_, _28041_);
  and _32016_ (_28044_, _28043_, _27668_);
  nor _32017_ (_28045_, _27668_, _26475_);
  or _32018_ (_28046_, _28045_, _28044_);
  and _32019_ (_26080_, _28046_, _27355_);
  nor _32020_ (_28047_, _27736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _32021_ (_28048_, _27736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _32022_ (_28049_, _28048_, _28047_);
  and _32023_ (_28050_, _28049_, _27732_);
  and _32024_ (_28051_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _32025_ (_28052_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _32026_ (_28053_, _28052_, _27743_);
  nor _32027_ (_28054_, _28053_, _28051_);
  and _32028_ (_28055_, _27688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _32029_ (_28056_, _27688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _32030_ (_28057_, _28056_, _27671_);
  nor _32031_ (_28058_, _28057_, _28055_);
  or _32032_ (_28059_, _28058_, _28054_);
  nor _32033_ (_28060_, _28059_, _28050_);
  nand _32034_ (_28061_, _28060_, _27714_);
  nand _32035_ (_28062_, _27670_, _26521_);
  and _32036_ (_28063_, _28062_, _27668_);
  and _32037_ (_28064_, _28063_, _28061_);
  and _32038_ (_28065_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _32039_ (_28066_, _28065_, _28064_);
  and _32040_ (_26082_, _28066_, _27355_);
  nand _32041_ (_28067_, _27670_, _26512_);
  or _32042_ (_28068_, _28048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _32043_ (_28069_, _27734_, _27680_);
  and _32044_ (_28070_, _28069_, _27690_);
  not _32045_ (_28071_, _28070_);
  or _32046_ (_28072_, _28071_, _27721_);
  and _32047_ (_28073_, _28072_, _27732_);
  and _32048_ (_28074_, _28073_, _28068_);
  and _32049_ (_28075_, _27744_, _27690_);
  or _32050_ (_28076_, _28051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _32051_ (_28077_, _28076_, _27743_);
  nor _32052_ (_28078_, _28077_, _28075_);
  and _32053_ (_28079_, _28055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _32054_ (_28080_, _28055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _32055_ (_28081_, _28080_, _27671_);
  nor _32056_ (_28082_, _28081_, _28079_);
  or _32057_ (_28083_, _28082_, _28078_);
  or _32058_ (_28084_, _28083_, _28074_);
  or _32059_ (_28085_, _28084_, _27670_);
  and _32060_ (_28086_, _28085_, _27668_);
  and _32061_ (_28087_, _28086_, _28067_);
  and _32062_ (_28088_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _32063_ (_28089_, _28088_, _28087_);
  and _32064_ (_26084_, _28089_, _27355_);
  nand _32065_ (_28090_, _27670_, _26505_);
  or _32066_ (_28091_, _28070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _32067_ (_28092_, _28069_, _27691_);
  not _32068_ (_28093_, _28092_);
  and _32069_ (_28094_, _28093_, _27702_);
  and _32070_ (_28095_, _28094_, _28091_);
  or _32071_ (_28096_, _28079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _32072_ (_28097_, _27691_, _27688_);
  nor _32073_ (_28098_, _28097_, _27707_);
  and _32074_ (_28099_, _28098_, _28096_);
  and _32075_ (_28100_, _28075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _32076_ (_28101_, _28100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _32077_ (_28102_, _27744_, _27691_);
  nand _32078_ (_28103_, _28102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _32079_ (_28104_, _28103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _32080_ (_28105_, _28104_, _28101_);
  or _32081_ (_28106_, _28105_, _28099_);
  or _32082_ (_28107_, _28106_, _28095_);
  or _32083_ (_28108_, _28107_, _27670_);
  and _32084_ (_28109_, _28108_, _27668_);
  and _32085_ (_28110_, _28109_, _28090_);
  and _32086_ (_28111_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _32087_ (_28112_, _28111_, _28110_);
  and _32088_ (_26086_, _28112_, _27355_);
  nand _32089_ (_28113_, _27670_, _26497_);
  not _32090_ (_28114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _32091_ (_28115_, _28092_, _27701_);
  nor _32092_ (_28116_, _28115_, _28114_);
  and _32093_ (_28117_, _28115_, _28114_);
  or _32094_ (_28118_, _28117_, _28116_);
  and _32095_ (_28119_, _28118_, _27732_);
  or _32096_ (_28120_, _28102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _32097_ (_28121_, _27745_);
  and _32098_ (_28122_, _28121_, _27743_);
  and _32099_ (_28123_, _28122_, _28120_);
  or _32100_ (_28124_, _28097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _32101_ (_28125_, _27692_, _27688_);
  nor _32102_ (_28126_, _28125_, _27707_);
  and _32103_ (_28127_, _28126_, _28124_);
  or _32104_ (_28128_, _28127_, _28123_);
  or _32105_ (_28129_, _28128_, _28119_);
  or _32106_ (_28130_, _28129_, _27670_);
  and _32107_ (_28131_, _28130_, _27668_);
  and _32108_ (_28132_, _28131_, _28113_);
  and _32109_ (_28133_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _32110_ (_28134_, _28133_, _28132_);
  and _32111_ (_26088_, _28134_, _27355_);
  nand _32112_ (_28135_, _27670_, _26489_);
  or _32113_ (_28136_, _28125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _32114_ (_28137_, _28079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _32115_ (_28138_, _28137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _32116_ (_28139_, _28138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _32117_ (_28140_, _28139_, _27707_);
  and _32118_ (_28141_, _28140_, _28136_);
  and _32119_ (_28142_, _28069_, _27692_);
  nand _32120_ (_28143_, _28142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _32121_ (_28144_, _28142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _32122_ (_28145_, _28144_, _27702_);
  and _32123_ (_28146_, _28145_, _28143_);
  and _32124_ (_28147_, _27745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _32125_ (_28148_, _28147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _32126_ (_28149_, _28148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _32127_ (_28150_, _27745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _32128_ (_28151_, _28150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _32129_ (_28152_, _28151_, _28149_);
  or _32130_ (_28153_, _28152_, _28146_);
  or _32131_ (_28154_, _28153_, _28141_);
  or _32132_ (_28155_, _28154_, _27670_);
  and _32133_ (_28156_, _28155_, _27668_);
  and _32134_ (_28157_, _28156_, _28135_);
  and _32135_ (_28158_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _32136_ (_28159_, _28158_, _28157_);
  and _32137_ (_26090_, _28159_, _27355_);
  nand _32138_ (_28160_, _27670_, _26482_);
  nor _32139_ (_28161_, _28143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _32140_ (_28162_, _28161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _32141_ (_28163_, _28161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _32142_ (_28164_, _28163_, _27732_);
  and _32143_ (_28165_, _28164_, _28162_);
  not _32144_ (_28166_, _27746_);
  and _32145_ (_28167_, _28166_, _27743_);
  or _32146_ (_28168_, _28150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _32147_ (_28169_, _28168_, _28167_);
  not _32148_ (_28170_, _28139_);
  nor _32149_ (_28171_, _28170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _32150_ (_28172_, _28170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _32151_ (_28173_, _28172_, _28171_);
  and _32152_ (_28174_, _28173_, _27671_);
  or _32153_ (_28175_, _28174_, _28169_);
  or _32154_ (_28176_, _28175_, _28165_);
  or _32155_ (_28177_, _28176_, _27670_);
  and _32156_ (_28178_, _28177_, _27668_);
  and _32157_ (_28179_, _28178_, _28160_);
  and _32158_ (_28180_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _32159_ (_28181_, _28180_, _28179_);
  and _32160_ (_26092_, _28181_, _27355_);
  nand _32161_ (_28182_, _27670_, _26475_);
  or _32162_ (_28183_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _32163_ (_28184_, _28183_, _27732_);
  nor _32164_ (_28185_, _28184_, _27738_);
  or _32165_ (_28186_, _27746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _32166_ (_28187_, _27747_);
  and _32167_ (_28188_, _28187_, _27743_);
  and _32168_ (_28189_, _28188_, _28186_);
  or _32169_ (_28190_, _27694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _32170_ (_28191_, _27752_, _27707_);
  and _32171_ (_28192_, _28191_, _28190_);
  or _32172_ (_28193_, _28192_, _28189_);
  or _32173_ (_28194_, _28193_, _28185_);
  or _32174_ (_28195_, _28194_, _27670_);
  and _32175_ (_28196_, _28195_, _27668_);
  and _32176_ (_28197_, _28196_, _28182_);
  and _32177_ (_28198_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _32178_ (_28199_, _28198_, _28197_);
  and _32179_ (_26094_, _28199_, _27355_);
  nor _32180_ (_28200_, _27770_, _27720_);
  and _32181_ (_00002_, _27770_, _26522_);
  or _32182_ (_00003_, _00002_, _28200_);
  and _32183_ (_26096_, _00003_, _27355_);
  or _32184_ (_00004_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _32185_ (_00005_, _00004_, _27355_);
  nand _32186_ (_00006_, _27770_, _26512_);
  and _32187_ (_26098_, _00006_, _00005_);
  or _32188_ (_00007_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _32189_ (_00008_, _00007_, _27355_);
  nand _32190_ (_00009_, _27770_, _26505_);
  and _32191_ (_26100_, _00009_, _00008_);
  or _32192_ (_00010_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _32193_ (_00011_, _00010_, _27355_);
  nand _32194_ (_00012_, _27770_, _26497_);
  and _32195_ (_26102_, _00012_, _00011_);
  or _32196_ (_00013_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _32197_ (_00014_, _00013_, _27355_);
  nand _32198_ (_00015_, _27770_, _26489_);
  and _32199_ (_26104_, _00015_, _00014_);
  or _32200_ (_00016_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _32201_ (_00017_, _00016_, _27355_);
  nand _32202_ (_00018_, _27770_, _26482_);
  and _32203_ (_26106_, _00018_, _00017_);
  or _32204_ (_00019_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _32205_ (_00020_, _00019_, _27355_);
  nand _32206_ (_00021_, _27770_, _26475_);
  and _32207_ (_26108_, _00021_, _00020_);
  nor _32208_ (_00022_, _25128_, _25115_);
  and _32209_ (_00023_, _00022_, _27048_);
  and _32210_ (_00024_, _00023_, _27179_);
  and _32211_ (_00025_, _00024_, _25517_);
  nand _32212_ (_00026_, _00025_, _25514_);
  and _32213_ (_00027_, _26456_, _25517_);
  and _32214_ (_00028_, _00027_, _27203_);
  not _32215_ (_00029_, _00028_);
  or _32216_ (_00030_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _32217_ (_00031_, _00030_, _00029_);
  and _32218_ (_00032_, _00031_, _00026_);
  nor _32219_ (_00033_, _00029_, _26543_);
  or _32220_ (_00034_, _00033_, _00032_);
  and _32221_ (_27294_, _00034_, _27355_);
  and _32222_ (_00035_, _27576_, _25055_);
  and _32223_ (_00036_, _00035_, _27186_);
  and _32224_ (_00037_, _25128_, _25116_);
  and _32225_ (_00038_, _00037_, _27048_);
  and _32226_ (_00039_, _00038_, _27179_);
  and _32227_ (_00040_, _00039_, _25517_);
  nand _32228_ (_00041_, _00040_, _25514_);
  or _32229_ (_00042_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _32230_ (_00043_, _00042_, _00041_);
  or _32231_ (_00044_, _00043_, _00036_);
  nand _32232_ (_00045_, _00036_, _26543_);
  and _32233_ (_00046_, _00045_, _27355_);
  and _32234_ (_27296_, _00046_, _00044_);
  and _32235_ (_00047_, _00035_, _26460_);
  and _32236_ (_00048_, _00038_, _27147_);
  nand _32237_ (_00049_, _00048_, _25053_);
  and _32238_ (_00050_, _00049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _32239_ (_00051_, _00050_, _00047_);
  nor _32240_ (_00052_, _27047_, _25115_);
  and _32241_ (_00053_, _00052_, _25128_);
  and _32242_ (_00054_, _00053_, _25102_);
  and _32243_ (_00055_, _00054_, _27147_);
  or _32244_ (_00056_, _25054_, _25715_);
  and _32245_ (_00057_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _32246_ (_00058_, _00057_, _27025_);
  and _32247_ (_00059_, _00058_, _00055_);
  or _32248_ (_00060_, _00059_, _00051_);
  nand _32249_ (_00061_, _00047_, _26475_);
  and _32250_ (_00062_, _00061_, _27355_);
  and _32251_ (_27298_, _00062_, _00060_);
  not _32252_ (_00063_, _00047_);
  nor _32253_ (_00064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _32254_ (_00065_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _32255_ (_00066_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _32256_ (_00067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _32257_ (_00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _32258_ (_00069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00068_);
  and _32259_ (_00070_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _32260_ (_00071_, _00070_, _00069_);
  nor _32261_ (_00072_, _00071_, _00067_);
  or _32262_ (_00073_, _00072_, _00066_);
  and _32263_ (_00074_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _32264_ (_00075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _32265_ (_00076_, _00075_, _00074_);
  nor _32266_ (_00077_, _00076_, _00067_);
  and _32267_ (_00078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00068_);
  and _32268_ (_00079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _32269_ (_00080_, _00079_, _00078_);
  nand _32270_ (_00081_, _00080_, _00077_);
  or _32271_ (_00082_, _00081_, _00073_);
  and _32272_ (_00083_, _00082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _32273_ (_00084_, _00083_, _00065_);
  and _32274_ (_00085_, _26460_, _25517_);
  and _32275_ (_00086_, _00085_, _00052_);
  or _32276_ (_00087_, _00086_, _00084_);
  and _32277_ (_00088_, _00087_, _00063_);
  nand _32278_ (_00089_, _00086_, _25514_);
  and _32279_ (_00090_, _00089_, _00088_);
  nor _32280_ (_00091_, _00063_, _26543_);
  or _32281_ (_00092_, _00091_, _00090_);
  and _32282_ (_27301_, _00092_, _27355_);
  and _32283_ (_00093_, _27586_, _25521_);
  nand _32284_ (_00094_, _00093_, _25514_);
  not _32285_ (_00095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _32286_ (_00096_, _00095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _32287_ (_00097_, _00080_, _00067_);
  not _32288_ (_00098_, _00097_);
  or _32289_ (_00099_, _00098_, _00077_);
  or _32290_ (_00100_, _00099_, _00073_);
  and _32291_ (_00101_, _00100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _32292_ (_00102_, _00101_, _00096_);
  or _32293_ (_00103_, _00102_, _00093_);
  and _32294_ (_00104_, _00103_, _00063_);
  and _32295_ (_00105_, _00104_, _00094_);
  nor _32296_ (_00106_, _00063_, _26482_);
  or _32297_ (_00107_, _00106_, _00105_);
  and _32298_ (_27303_, _00107_, _27355_);
  not _32299_ (_00108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _32300_ (_00109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _00108_);
  nand _32301_ (_00110_, _00072_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _32302_ (_00111_, _00097_, _00077_);
  or _32303_ (_00112_, _00111_, _00110_);
  and _32304_ (_00113_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _32305_ (_00114_, _00113_, _00109_);
  and _32306_ (_00115_, _00052_, _26462_);
  or _32307_ (_00116_, _00115_, _00114_);
  and _32308_ (_00117_, _00116_, _00063_);
  nand _32309_ (_00118_, _00115_, _25514_);
  and _32310_ (_00119_, _00118_, _00117_);
  nor _32311_ (_00120_, _00063_, _26512_);
  or _32312_ (_00121_, _00120_, _00119_);
  and _32313_ (_27305_, _00121_, _27355_);
  and _32314_ (_00122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _32315_ (_00123_, _00110_, _00099_);
  and _32316_ (_00124_, _00123_, _00122_);
  and _32317_ (_00125_, _00052_, _26592_);
  or _32318_ (_00126_, _00125_, _00124_);
  and _32319_ (_00127_, _00126_, _00063_);
  nand _32320_ (_00128_, _00125_, _25514_);
  and _32321_ (_00129_, _00128_, _00127_);
  nor _32322_ (_00130_, _00063_, _26497_);
  or _32323_ (_00131_, _00130_, _00129_);
  and _32324_ (_27307_, _00131_, _27355_);
  nand _32325_ (_00132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _32326_ (_00133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00068_);
  and _32327_ (_00134_, _00133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _32328_ (_00135_, _00134_, _00132_);
  or _32329_ (_00136_, _00135_, _00067_);
  and _32330_ (_00137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _32331_ (_00138_, _00137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _32332_ (_00139_, _00138_);
  and _32333_ (_00140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _32334_ (_00141_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _32335_ (_00143_, _00141_);
  and _32336_ (_00145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _32337_ (_00147_, _00145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _32338_ (_00149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _32339_ (_00151_, _00149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _32340_ (_00153_, _00151_, _00147_);
  and _32341_ (_00155_, _00153_, _00143_);
  and _32342_ (_00157_, _00155_, _00139_);
  not _32343_ (_00159_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _32344_ (_00161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _32345_ (_00163_, _00161_, _00159_);
  nand _32346_ (_00165_, _00163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _32347_ (_00167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _32348_ (_00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _32349_ (_00171_, _00169_, _00167_);
  and _32350_ (_00173_, _00171_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _32351_ (_00175_, _00173_);
  and _32352_ (_00177_, _00175_, _00165_);
  nand _32353_ (_00179_, _00177_, _00157_);
  and _32354_ (_00181_, _00179_, _00136_);
  and _32355_ (_00183_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _32356_ (_00185_, _00183_, _00068_);
  and _32357_ (_00187_, _00185_, _00181_);
  not _32358_ (_00189_, _00187_);
  not _32359_ (_00191_, _00185_);
  and _32360_ (_00193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _00067_);
  not _32361_ (_00195_, _00193_);
  not _32362_ (_00197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _32363_ (_00199_, _00140_, _00197_);
  not _32364_ (_00201_, _00199_);
  not _32365_ (_00203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _32366_ (_00204_, _00145_, _00203_);
  not _32367_ (_00205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _32368_ (_00206_, _00149_, _00205_);
  nor _32369_ (_00207_, _00206_, _00204_);
  and _32370_ (_00208_, _00207_, _00201_);
  nor _32371_ (_00209_, _00208_, _00195_);
  not _32372_ (_00210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _32373_ (_00211_, _00163_, _00210_);
  not _32374_ (_00212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _32375_ (_00213_, _00171_, _00212_);
  nor _32376_ (_00214_, _00213_, _00211_);
  not _32377_ (_00215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _32378_ (_00216_, _00137_, _00215_);
  not _32379_ (_00217_, _00216_);
  and _32380_ (_00218_, _00217_, _00214_);
  nor _32381_ (_00219_, _00218_, _00195_);
  nor _32382_ (_00220_, _00219_, _00209_);
  or _32383_ (_00221_, _00220_, _00191_);
  and _32384_ (_00222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27355_);
  and _32385_ (_00223_, _00222_, _00221_);
  and _32386_ (_27341_, _00223_, _00189_);
  nor _32387_ (_00224_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _32388_ (_00225_, _00224_);
  not _32389_ (_00226_, _00181_);
  and _32390_ (_00227_, _00220_, _00226_);
  nor _32391_ (_00228_, _00227_, _00225_);
  nand _32392_ (_00229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27355_);
  nor _32393_ (_27343_, _00229_, _00228_);
  and _32394_ (_00230_, _00177_, _00139_);
  nand _32395_ (_00231_, _00230_, _00181_);
  or _32396_ (_00232_, _00219_, _00181_);
  and _32397_ (_00233_, _00232_, _00185_);
  and _32398_ (_00234_, _00233_, _00231_);
  or _32399_ (_00235_, _00234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _32400_ (_00236_, _00189_, _00155_);
  nor _32401_ (_00237_, _00191_, _00181_);
  nand _32402_ (_00238_, _00237_, _00209_);
  and _32403_ (_00239_, _00238_, _27355_);
  and _32404_ (_00240_, _00239_, _00236_);
  and _32405_ (_27345_, _00240_, _00235_);
  and _32406_ (_00241_, _00231_, _00224_);
  or _32407_ (_00242_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _32408_ (_00243_, _00224_, _00181_);
  not _32409_ (_00244_, _00243_);
  or _32410_ (_00245_, _00244_, _00155_);
  or _32411_ (_00246_, _00219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _32412_ (_00247_, _00224_, _00209_);
  and _32413_ (_00248_, _00247_, _00246_);
  or _32414_ (_00249_, _00248_, _00181_);
  and _32415_ (_00250_, _00249_, _27355_);
  and _32416_ (_00251_, _00250_, _00245_);
  and _32417_ (_27347_, _00251_, _00242_);
  nand _32418_ (_00252_, _00227_, _00067_);
  nor _32419_ (_00253_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _32420_ (_00254_, _00253_, _00183_);
  and _32421_ (_00255_, _00254_, _27355_);
  and _32422_ (_27349_, _00255_, _00252_);
  and _32423_ (_00256_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _32424_ (_00257_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _32425_ (_00258_, _00257_, _00253_);
  nor _32426_ (_00259_, _00258_, _00226_);
  or _32427_ (_00260_, _00259_, _00183_);
  or _32428_ (_00261_, _00260_, _00256_);
  not _32429_ (_00262_, _00183_);
  or _32430_ (_00263_, _00258_, _00262_);
  and _32431_ (_00264_, _00263_, _27355_);
  and _32432_ (_27351_, _00264_, _00261_);
  and _32433_ (_00265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27355_);
  and _32434_ (_27353_, _00265_, _00183_);
  nor _32435_ (_27357_, _00064_, rst);
  and _32436_ (_27359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _27355_);
  nor _32437_ (_00266_, _00227_, _00183_);
  and _32438_ (_00267_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _32439_ (_00268_, _00267_, _00266_);
  and _32440_ (_00142_, _00268_, _27355_);
  and _32441_ (_00269_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _32442_ (_00270_, _00269_, _00266_);
  and _32443_ (_00144_, _00270_, _27355_);
  and _32444_ (_00271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _27355_);
  and _32445_ (_00146_, _00271_, _00183_);
  nor _32446_ (_00272_, _00220_, _00181_);
  not _32447_ (_00273_, _00206_);
  nor _32448_ (_00274_, _00213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _32449_ (_00275_, _00274_, _00211_);
  or _32450_ (_00276_, _00275_, _00216_);
  and _32451_ (_00277_, _00276_, _00273_);
  or _32452_ (_00278_, _00277_, _00204_);
  and _32453_ (_00279_, _00278_, _00201_);
  and _32454_ (_00280_, _00279_, _00272_);
  not _32455_ (_00281_, _00151_);
  or _32456_ (_00282_, _00173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _32457_ (_00283_, _00282_, _00165_);
  or _32458_ (_00284_, _00283_, _00138_);
  and _32459_ (_00285_, _00284_, _00281_);
  or _32460_ (_00286_, _00285_, _00147_);
  and _32461_ (_00287_, _00181_, _00143_);
  and _32462_ (_00288_, _00287_, _00286_);
  or _32463_ (_00289_, _00288_, _00183_);
  or _32464_ (_00290_, _00289_, _00280_);
  or _32465_ (_00291_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _32466_ (_00292_, _00291_, _27355_);
  and _32467_ (_00148_, _00292_, _00290_);
  nor _32468_ (_00293_, _00204_, _00199_);
  or _32469_ (_00294_, _00216_, _00206_);
  and _32470_ (_00295_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _32471_ (_00296_, _00295_, _00294_);
  and _32472_ (_00297_, _00296_, _00293_);
  and _32473_ (_00298_, _00297_, _00272_);
  not _32474_ (_00299_, _00147_);
  or _32475_ (_00300_, _00151_, _00138_);
  and _32476_ (_00301_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _32477_ (_00302_, _00301_, _00300_);
  and _32478_ (_00303_, _00302_, _00299_);
  and _32479_ (_00304_, _00303_, _00287_);
  or _32480_ (_00305_, _00304_, _00183_);
  or _32481_ (_00306_, _00305_, _00298_);
  or _32482_ (_00307_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _32483_ (_00308_, _00307_, _27355_);
  and _32484_ (_00150_, _00308_, _00306_);
  and _32485_ (_00309_, _00217_, _00193_);
  nand _32486_ (_00310_, _00309_, _00208_);
  or _32487_ (_00311_, _00310_, _00214_);
  nor _32488_ (_00312_, _00311_, _00181_);
  nand _32489_ (_00313_, _00157_, _00136_);
  nor _32490_ (_00314_, _00313_, _00177_);
  or _32491_ (_00315_, _00314_, _00183_);
  or _32492_ (_00316_, _00315_, _00312_);
  or _32493_ (_00317_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _32494_ (_00318_, _00317_, _27355_);
  and _32495_ (_00152_, _00318_, _00316_);
  and _32496_ (_00319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _27355_);
  and _32497_ (_00154_, _00319_, _00183_);
  and _32498_ (_00320_, _00183_, _00068_);
  or _32499_ (_00321_, _00320_, _00228_);
  or _32500_ (_00322_, _00321_, _00237_);
  and _32501_ (_00156_, _00322_, _27355_);
  not _32502_ (_00323_, _00266_);
  and _32503_ (_00324_, _00323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _32504_ (_00325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00068_);
  or _32505_ (_00326_, _00325_, _00143_);
  and _32506_ (_00327_, _00326_, _00181_);
  not _32507_ (_00328_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _32508_ (_00329_, _00173_, _00068_);
  or _32509_ (_00330_, _00329_, _00328_);
  nor _32510_ (_00331_, _00165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _32511_ (_00332_, _00331_, _00138_);
  nand _32512_ (_00333_, _00332_, _00330_);
  or _32513_ (_00334_, _00139_, _00070_);
  and _32514_ (_00335_, _00334_, _00333_);
  or _32515_ (_00336_, _00335_, _00151_);
  or _32516_ (_00337_, _00325_, _00281_);
  and _32517_ (_00338_, _00337_, _00299_);
  and _32518_ (_00339_, _00338_, _00336_);
  and _32519_ (_00340_, _00147_, _00070_);
  or _32520_ (_00341_, _00340_, _00141_);
  or _32521_ (_00342_, _00341_, _00339_);
  and _32522_ (_00343_, _00342_, _00327_);
  or _32523_ (_00344_, _00325_, _00201_);
  and _32524_ (_00345_, _00213_, _00068_);
  or _32525_ (_00346_, _00345_, _00328_);
  and _32526_ (_00347_, _00211_, _00068_);
  nor _32527_ (_00348_, _00347_, _00216_);
  nand _32528_ (_00349_, _00348_, _00346_);
  or _32529_ (_00350_, _00217_, _00070_);
  and _32530_ (_00351_, _00350_, _00349_);
  or _32531_ (_00352_, _00351_, _00206_);
  not _32532_ (_00353_, _00204_);
  or _32533_ (_00354_, _00325_, _00273_);
  and _32534_ (_00355_, _00354_, _00353_);
  and _32535_ (_00356_, _00355_, _00352_);
  and _32536_ (_00357_, _00204_, _00070_);
  or _32537_ (_00358_, _00357_, _00199_);
  or _32538_ (_00359_, _00358_, _00356_);
  and _32539_ (_00360_, _00359_, _00272_);
  and _32540_ (_00361_, _00360_, _00344_);
  or _32541_ (_00362_, _00361_, _00343_);
  and _32542_ (_00363_, _00362_, _00262_);
  or _32543_ (_00364_, _00363_, _00324_);
  and _32544_ (_00158_, _00364_, _27355_);
  or _32545_ (_00365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00068_);
  and _32546_ (_00366_, _00365_, _00143_);
  or _32547_ (_00367_, _00366_, _00155_);
  or _32548_ (_00368_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _32549_ (_00369_, _00368_, _00332_);
  nand _32550_ (_00370_, _00138_, _00079_);
  nand _32551_ (_00371_, _00370_, _00153_);
  or _32552_ (_00372_, _00371_, _00369_);
  and _32553_ (_00373_, _00372_, _00367_);
  nand _32554_ (_00374_, _00141_, _00079_);
  nand _32555_ (_00375_, _00374_, _00181_);
  or _32556_ (_00376_, _00375_, _00373_);
  or _32557_ (_00377_, _00345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _32558_ (_00378_, _00377_, _00348_);
  and _32559_ (_00379_, _00216_, _00079_);
  or _32560_ (_00380_, _00379_, _00378_);
  and _32561_ (_00381_, _00380_, _00207_);
  not _32562_ (_00382_, _00207_);
  and _32563_ (_00383_, _00365_, _00382_);
  or _32564_ (_00384_, _00383_, _00199_);
  or _32565_ (_00385_, _00384_, _00381_);
  or _32566_ (_00386_, _00201_, _00079_);
  nand _32567_ (_00387_, _00386_, _00385_);
  nand _32568_ (_00388_, _00387_, _00272_);
  and _32569_ (_00389_, _00388_, _00376_);
  or _32570_ (_00390_, _00389_, _00183_);
  or _32571_ (_00391_, _00266_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _32572_ (_00392_, _00391_, _27355_);
  and _32573_ (_00160_, _00392_, _00390_);
  and _32574_ (_00393_, _00323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _32575_ (_00394_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _32576_ (_00395_, _00394_, _00143_);
  and _32577_ (_00396_, _00395_, _00181_);
  not _32578_ (_00397_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _32579_ (_00398_, _00173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _32580_ (_00399_, _00398_, _00397_);
  nor _32581_ (_00400_, _00165_, _00068_);
  nor _32582_ (_00401_, _00400_, _00138_);
  nand _32583_ (_00402_, _00401_, _00399_);
  or _32584_ (_00403_, _00139_, _00069_);
  and _32585_ (_00404_, _00403_, _00402_);
  or _32586_ (_00405_, _00404_, _00151_);
  or _32587_ (_00406_, _00394_, _00281_);
  and _32588_ (_00407_, _00406_, _00299_);
  and _32589_ (_00408_, _00407_, _00405_);
  and _32590_ (_00409_, _00147_, _00069_);
  or _32591_ (_00410_, _00409_, _00141_);
  or _32592_ (_00411_, _00410_, _00408_);
  and _32593_ (_00412_, _00411_, _00396_);
  or _32594_ (_00413_, _00394_, _00201_);
  and _32595_ (_00414_, _00213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _32596_ (_00415_, _00414_, _00397_);
  and _32597_ (_00416_, _00211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _32598_ (_00417_, _00416_, _00216_);
  nand _32599_ (_00418_, _00417_, _00415_);
  or _32600_ (_00419_, _00217_, _00069_);
  and _32601_ (_00420_, _00419_, _00418_);
  or _32602_ (_00421_, _00420_, _00206_);
  or _32603_ (_00422_, _00394_, _00273_);
  and _32604_ (_00423_, _00422_, _00353_);
  and _32605_ (_00424_, _00423_, _00421_);
  and _32606_ (_00425_, _00204_, _00069_);
  or _32607_ (_00426_, _00425_, _00199_);
  or _32608_ (_00427_, _00426_, _00424_);
  and _32609_ (_00428_, _00427_, _00272_);
  and _32610_ (_00429_, _00428_, _00413_);
  or _32611_ (_00430_, _00429_, _00412_);
  and _32612_ (_00431_, _00430_, _00262_);
  or _32613_ (_00432_, _00431_, _00393_);
  and _32614_ (_00162_, _00432_, _27355_);
  and _32615_ (_00433_, _00199_, _00078_);
  or _32616_ (_00434_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _32617_ (_00435_, _00434_, _00201_);
  or _32618_ (_00436_, _00435_, _00208_);
  and _32619_ (_00437_, _00216_, _00078_);
  or _32620_ (_00438_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _32621_ (_00439_, _00438_, _00417_);
  or _32622_ (_00440_, _00439_, _00382_);
  or _32623_ (_00441_, _00440_, _00437_);
  and _32624_ (_00442_, _00441_, _00436_);
  or _32625_ (_00443_, _00442_, _00433_);
  and _32626_ (_00444_, _00443_, _00272_);
  or _32627_ (_00445_, _00398_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _32628_ (_00446_, _00445_, _00401_);
  and _32629_ (_00447_, _00138_, _00078_);
  or _32630_ (_00448_, _00447_, _00446_);
  and _32631_ (_00449_, _00448_, _00153_);
  not _32632_ (_00450_, _00153_);
  and _32633_ (_00451_, _00434_, _00450_);
  or _32634_ (_00452_, _00451_, _00141_);
  or _32635_ (_00453_, _00452_, _00449_);
  or _32636_ (_00454_, _00143_, _00078_);
  and _32637_ (_00455_, _00454_, _00181_);
  and _32638_ (_00456_, _00455_, _00453_);
  and _32639_ (_00457_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _32640_ (_00458_, _00457_, _00183_);
  or _32641_ (_00459_, _00458_, _00456_);
  or _32642_ (_00460_, _00459_, _00444_);
  or _32643_ (_00461_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _32644_ (_00462_, _00461_, _27355_);
  and _32645_ (_00164_, _00462_, _00460_);
  or _32646_ (_00463_, _00225_, _00220_);
  and _32647_ (_00464_, _00463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _32648_ (_00465_, _00464_, _00243_);
  and _32649_ (_00166_, _00465_, _27355_);
  and _32650_ (_00466_, _00221_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _32651_ (_00467_, _00466_, _00187_);
  and _32652_ (_00168_, _00467_, _27355_);
  or _32653_ (_00468_, _00049_, _25719_);
  or _32654_ (_00469_, _00468_, _25574_);
  nand _32655_ (_00470_, _00468_, _00108_);
  and _32656_ (_00471_, _00470_, _00063_);
  and _32657_ (_00472_, _00471_, _00469_);
  nor _32658_ (_00473_, _00063_, _26521_);
  or _32659_ (_00474_, _00473_, _00472_);
  and _32660_ (_00170_, _00474_, _27355_);
  nand _32661_ (_00475_, _00055_, _25716_);
  nor _32662_ (_00476_, _00475_, _25514_);
  and _32663_ (_00477_, _00475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _32664_ (_00478_, _00477_, _00047_);
  or _32665_ (_00479_, _00478_, _00476_);
  nand _32666_ (_00480_, _00047_, _26505_);
  and _32667_ (_00481_, _00480_, _27355_);
  and _32668_ (_00172_, _00481_, _00479_);
  and _32669_ (_00482_, _00055_, _25838_);
  or _32670_ (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _32671_ (_00484_, _00483_, _00063_);
  nand _32672_ (_00485_, _00482_, _25514_);
  and _32673_ (_00486_, _00485_, _00484_);
  nor _32674_ (_00487_, _00063_, _26489_);
  or _32675_ (_00488_, _00487_, _00486_);
  and _32676_ (_00174_, _00488_, _27355_);
  and _32677_ (_00489_, _00039_, _25055_);
  nand _32678_ (_00490_, _00489_, _25514_);
  not _32679_ (_00491_, _00036_);
  or _32680_ (_00492_, _00489_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _32681_ (_00493_, _00492_, _00491_);
  and _32682_ (_00494_, _00493_, _00490_);
  nor _32683_ (_00495_, _00491_, _26521_);
  or _32684_ (_00496_, _00495_, _00494_);
  and _32685_ (_00176_, _00496_, _27355_);
  and _32686_ (_00497_, _00039_, _26947_);
  or _32687_ (_00498_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _32688_ (_00499_, _00498_, _00491_);
  nand _32689_ (_00500_, _00497_, _25514_);
  and _32690_ (_00501_, _00500_, _00499_);
  nor _32691_ (_00502_, _00491_, _26512_);
  or _32692_ (_00503_, _00502_, _00501_);
  and _32693_ (_00178_, _00503_, _27355_);
  nand _32694_ (_00504_, _00039_, _27237_);
  and _32695_ (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _32696_ (_00506_, _00505_, _00036_);
  and _32697_ (_00507_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _32698_ (_00508_, _00507_, _25718_);
  and _32699_ (_00509_, _00508_, _00039_);
  or _32700_ (_00510_, _00509_, _00506_);
  nand _32701_ (_00511_, _00036_, _26505_);
  and _32702_ (_00512_, _00511_, _27355_);
  and _32703_ (_00180_, _00512_, _00510_);
  and _32704_ (_00513_, _00039_, _25778_);
  or _32705_ (_00514_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _32706_ (_00515_, _00514_, _00491_);
  nand _32707_ (_00516_, _00513_, _25514_);
  and _32708_ (_00517_, _00516_, _00515_);
  nor _32709_ (_00518_, _00491_, _26497_);
  or _32710_ (_00519_, _00518_, _00517_);
  and _32711_ (_00182_, _00519_, _27355_);
  and _32712_ (_00520_, _00039_, _25838_);
  nand _32713_ (_00521_, _00520_, _25514_);
  or _32714_ (_00522_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _32715_ (_00523_, _00522_, _00521_);
  or _32716_ (_00524_, _00523_, _00036_);
  nand _32717_ (_00525_, _00036_, _26489_);
  and _32718_ (_00526_, _00525_, _27355_);
  and _32719_ (_00184_, _00526_, _00524_);
  and _32720_ (_00527_, _00039_, _25905_);
  or _32721_ (_00528_, _00527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _32722_ (_00529_, _00528_, _00491_);
  nand _32723_ (_00530_, _00527_, _25514_);
  and _32724_ (_00531_, _00530_, _00529_);
  nor _32725_ (_00532_, _00491_, _26482_);
  or _32726_ (_00533_, _00532_, _00531_);
  and _32727_ (_00186_, _00533_, _27355_);
  and _32728_ (_00534_, _00039_, _25972_);
  or _32729_ (_00535_, _00534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _32730_ (_00536_, _00535_, _00491_);
  nand _32731_ (_00537_, _00534_, _25514_);
  and _32732_ (_00538_, _00537_, _00536_);
  nor _32733_ (_00539_, _00491_, _26475_);
  or _32734_ (_00540_, _00539_, _00538_);
  and _32735_ (_00188_, _00540_, _27355_);
  and _32736_ (_00541_, _00024_, _25055_);
  nand _32737_ (_00542_, _00541_, _25514_);
  or _32738_ (_00543_, _00541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor _32739_ (_00544_, _00028_, rst);
  and _32740_ (_00545_, _00544_, _00543_);
  and _32741_ (_00546_, _00545_, _00542_);
  and _32742_ (_00547_, _00028_, _27774_);
  or _32743_ (_00190_, _00547_, _00546_);
  and _32744_ (_00548_, _00024_, _26947_);
  nand _32745_ (_00549_, _00548_, _25514_);
  or _32746_ (_00550_, _00548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _32747_ (_00551_, _00550_, _00029_);
  and _32748_ (_00552_, _00551_, _00549_);
  nor _32749_ (_00553_, _00029_, _26512_);
  or _32750_ (_00554_, _00553_, _00552_);
  and _32751_ (_00192_, _00554_, _27355_);
  nor _32752_ (_00555_, _25719_, _00205_);
  or _32753_ (_00556_, _00555_, _25718_);
  and _32754_ (_00557_, _00556_, _00024_);
  nand _32755_ (_00558_, _00024_, _27237_);
  and _32756_ (_00559_, _00558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _32757_ (_00560_, _00559_, _00028_);
  or _32758_ (_00561_, _00560_, _00557_);
  nand _32759_ (_00562_, _00028_, _26505_);
  and _32760_ (_00563_, _00562_, _27355_);
  and _32761_ (_00194_, _00563_, _00561_);
  and _32762_ (_00564_, _00024_, _25778_);
  nand _32763_ (_00565_, _00564_, _25514_);
  or _32764_ (_00566_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _32765_ (_00567_, _00566_, _00565_);
  or _32766_ (_00568_, _00567_, _00028_);
  nand _32767_ (_00569_, _00028_, _26497_);
  and _32768_ (_00570_, _00569_, _27355_);
  and _32769_ (_00196_, _00570_, _00568_);
  and _32770_ (_00571_, _00024_, _25838_);
  nand _32771_ (_00572_, _00571_, _25514_);
  or _32772_ (_00573_, _00571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _32773_ (_00574_, _00573_, _00572_);
  or _32774_ (_00575_, _00574_, _00028_);
  nand _32775_ (_00576_, _00028_, _26489_);
  and _32776_ (_00577_, _00576_, _27355_);
  and _32777_ (_00198_, _00577_, _00575_);
  and _32778_ (_00578_, _00024_, _25905_);
  nand _32779_ (_00579_, _00578_, _25514_);
  or _32780_ (_00580_, _00578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _32781_ (_00581_, _00580_, _00579_);
  or _32782_ (_00582_, _00581_, _00028_);
  nand _32783_ (_00583_, _00028_, _26482_);
  and _32784_ (_00584_, _00583_, _27355_);
  and _32785_ (_00200_, _00584_, _00582_);
  and _32786_ (_00585_, _00024_, _25972_);
  nand _32787_ (_00586_, _00585_, _25514_);
  or _32788_ (_00588_, _00585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _32789_ (_00589_, _00588_, _00029_);
  and _32790_ (_00591_, _00589_, _00586_);
  nor _32791_ (_00592_, _00029_, _26475_);
  or _32792_ (_00594_, _00592_, _00591_);
  and _32793_ (_00202_, _00594_, _27355_);
  and _32794_ (_00596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _32795_ (_00597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _32796_ (_00599_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _32797_ (_00600_, _00599_, _00597_);
  not _32798_ (_00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _32799_ (_00603_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _32800_ (_00605_, _00603_, _00600_);
  nor _32801_ (_00606_, _00605_, _00596_);
  or _32802_ (_00608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _32803_ (_00609_, _00608_, _27355_);
  nor _32804_ (_00590_, _00609_, _00606_);
  nor _32805_ (_00611_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _32806_ (_00613_, _00611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _32807_ (_00614_, _00611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _32808_ (_00616_, _00614_, _27355_);
  and _32809_ (_00593_, _00616_, _00613_);
  not _32810_ (_00618_, rxd_i);
  and _32811_ (_00619_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00618_);
  nor _32812_ (_00621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _32813_ (_00622_, _00621_);
  and _32814_ (_00624_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _32815_ (_00625_, _00624_, _00622_);
  and _32816_ (_00627_, _00625_, _00619_);
  not _32817_ (_00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _32818_ (_00630_, _00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _32819_ (_00631_, _00630_, _00621_);
  or _32820_ (_00633_, _00631_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _32821_ (_00634_, _00633_, _00627_);
  and _32822_ (_00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _27355_);
  and _32823_ (_00595_, _00636_, _00634_);
  and _32824_ (_00638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _32825_ (_00639_, _00638_, _00622_);
  nor _32826_ (_00640_, _00621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _32827_ (_00641_, _00640_, _00628_);
  nor _32828_ (_00642_, _00641_, _00639_);
  not _32829_ (_00643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _32830_ (_00644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _00643_);
  not _32831_ (_00645_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _32832_ (_00646_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _00645_);
  and _32833_ (_00647_, _00646_, _00644_);
  not _32834_ (_00648_, _00647_);
  or _32835_ (_00649_, _00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _32836_ (_00650_, _00647_, _00639_);
  and _32837_ (_00651_, _00639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _32838_ (_00652_, _00651_, _00650_);
  and _32839_ (_00653_, _00652_, _00649_);
  or _32840_ (_00654_, _00653_, _00642_);
  and _32841_ (_00655_, _00621_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _32842_ (_00656_, _00655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _32843_ (_00657_, _00656_);
  or _32844_ (_00658_, _00657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _32845_ (_00659_, _00658_, _00654_);
  nand _32846_ (_00598_, _00659_, _00636_);
  not _32847_ (_00660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _32848_ (_00661_, _00639_);
  nor _32849_ (_00662_, _00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _32850_ (_00663_, _00662_);
  not _32851_ (_00664_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _32852_ (_00665_, _00621_, _00664_);
  and _32853_ (_00666_, _00665_, _00663_);
  and _32854_ (_00667_, _00666_, _00661_);
  nor _32855_ (_00668_, _00667_, _00660_);
  and _32856_ (_00669_, _00667_, rxd_i);
  or _32857_ (_00670_, _00669_, rst);
  or _32858_ (_00601_, _00670_, _00668_);
  nor _32859_ (_00671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _32860_ (_00672_, _00671_, _00644_);
  and _32861_ (_00673_, _00672_, _00651_);
  nand _32862_ (_00674_, _00673_, _00618_);
  or _32863_ (_00675_, _00673_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _32864_ (_00676_, _00675_, _27355_);
  and _32865_ (_00604_, _00676_, _00674_);
  and _32866_ (_00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _32867_ (_00678_, _00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _32868_ (_00679_, _00678_, _00643_);
  and _32869_ (_00680_, _00679_, _00651_);
  and _32870_ (_00681_, _00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _32871_ (_00682_, _00681_, _00651_);
  nor _32872_ (_00683_, _00678_, _00661_);
  or _32873_ (_00684_, _00683_, _00682_);
  and _32874_ (_00685_, _00684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _32875_ (_00686_, _00685_, _00680_);
  and _32876_ (_00607_, _00686_, _27355_);
  and _32877_ (_00687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _27355_);
  nand _32878_ (_00688_, _00687_, _00664_);
  nand _32879_ (_00689_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _32880_ (_00610_, _00689_, _00688_);
  and _32881_ (_00690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00664_);
  not _32882_ (_00691_, _00625_);
  not _32883_ (_00692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _32884_ (_00693_, _00631_, _00692_);
  and _32885_ (_00694_, _00693_, _00691_);
  and _32886_ (_00695_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _32887_ (_00696_, _00695_, _00639_);
  or _32888_ (_00697_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _32889_ (_00698_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _32890_ (_00699_, _00698_, _00650_);
  and _32891_ (_00700_, _00699_, _00697_);
  and _32892_ (_00701_, _00700_, _00696_);
  or _32893_ (_00702_, _00701_, _00656_);
  nand _32894_ (_00703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _32895_ (_00704_, _00703_, _00639_);
  or _32896_ (_00705_, _00704_, _00648_);
  and _32897_ (_00706_, _00705_, _00657_);
  or _32898_ (_00707_, _00706_, rxd_i);
  and _32899_ (_00708_, _00707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _32900_ (_00709_, _00708_, _00702_);
  or _32901_ (_00710_, _00709_, _00690_);
  and _32902_ (_00612_, _00710_, _27355_);
  and _32903_ (_00711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _32904_ (_00712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _32905_ (_00713_, _00599_, _00712_);
  or _32906_ (_00714_, _00713_, _00603_);
  nor _32907_ (_00715_, _00714_, _00711_);
  or _32908_ (_00716_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _32909_ (_00717_, _00716_, _27355_);
  nor _32910_ (_00615_, _00717_, _00715_);
  nor _32911_ (_00718_, _00715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _32912_ (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _32913_ (_00720_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _32914_ (_00721_, _00720_, _27355_);
  and _32915_ (_00617_, _00721_, _00719_);
  and _32916_ (_00722_, _00655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _32917_ (_00723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _32918_ (_00724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _32919_ (_00725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _32920_ (_00726_, _00725_, _00724_);
  and _32921_ (_00727_, _00726_, _00723_);
  not _32922_ (_00728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _32923_ (_00729_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _32924_ (_00730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _32925_ (_00731_, _00730_, _00729_);
  and _32926_ (_00732_, _00731_, _00728_);
  and _32927_ (_00733_, _00732_, _00727_);
  or _32928_ (_00734_, _00733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _32929_ (_00735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _32930_ (_00736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _32931_ (_00737_, _00736_, _00735_);
  and _32932_ (_00738_, _00622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _32933_ (_00739_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _32934_ (_00740_, _00739_, _00737_);
  not _32935_ (_00741_, _00740_);
  or _32936_ (_00742_, _00741_, _00734_);
  and _32937_ (_00743_, _00737_, _00738_);
  not _32938_ (_00744_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _32939_ (_00745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00744_);
  or _32940_ (_00746_, _00745_, _00743_);
  and _32941_ (_00747_, _00746_, _00742_);
  or _32942_ (_00748_, _00747_, _00722_);
  not _32943_ (_00749_, _00722_);
  not _32944_ (_00750_, _00733_);
  or _32945_ (_00751_, _00750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _32946_ (_00752_, _00751_, _00734_);
  or _32947_ (_00753_, _00752_, _00749_);
  nand _32948_ (_00754_, _00753_, _00748_);
  nand _32949_ (_00755_, _26947_, _25116_);
  nor _32950_ (_00756_, _00755_, _27575_);
  and _32951_ (_00757_, _00756_, _27170_);
  nor _32952_ (_00758_, _00757_, rst);
  nand _32953_ (_00759_, _00758_, _00754_);
  not _32954_ (_00760_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _32955_ (_00761_, _00757_, _27355_);
  nand _32956_ (_00762_, _00761_, _00760_);
  and _32957_ (_00620_, _00762_, _00759_);
  nor _32958_ (_00763_, _00750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _32959_ (_00764_, _00743_, _00763_);
  and _32960_ (_00765_, _00733_, _00722_);
  or _32961_ (_00766_, _00744_, rst);
  nor _32962_ (_00767_, _00766_, _00765_);
  and _32963_ (_00768_, _00767_, _00764_);
  or _32964_ (_00623_, _00768_, _00761_);
  or _32965_ (_00769_, _00741_, _00763_);
  or _32966_ (_00770_, _00743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _32967_ (_00771_, _00655_, _00744_);
  and _32968_ (_00772_, _00771_, _00770_);
  and _32969_ (_00773_, _00772_, _00769_);
  or _32970_ (_00774_, _00773_, _00765_);
  and _32971_ (_00626_, _00774_, _00758_);
  and _32972_ (_00775_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _32973_ (_00776_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _32974_ (_00777_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _32975_ (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _32976_ (_00779_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _32977_ (_00780_, _00779_, _00778_);
  and _32978_ (_00629_, _00780_, _00758_);
  nor _32979_ (_00781_, _00740_, _00722_);
  and _32980_ (_00782_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _32981_ (_00783_, _00782_, _00758_);
  and _32982_ (_00784_, _00761_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _32983_ (_00632_, _00784_, _00783_);
  and _32984_ (_00785_, _00027_, _26460_);
  or _32985_ (_00786_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _32986_ (_00787_, _00786_, _27355_);
  nand _32987_ (_00788_, _00785_, _26543_);
  and _32988_ (_00635_, _00788_, _00787_);
  and _32989_ (_00789_, _00023_, _27147_);
  and _32990_ (_00790_, _00789_, _25517_);
  nand _32991_ (_00791_, _00790_, _25514_);
  and _32992_ (_00792_, _00035_, _27170_);
  not _32993_ (_00793_, _00792_);
  or _32994_ (_00794_, _00790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _32995_ (_00795_, _00794_, _00793_);
  and _32996_ (_00796_, _00795_, _00791_);
  nor _32997_ (_00797_, _00793_, _26543_);
  or _32998_ (_00798_, _00797_, _00796_);
  and _32999_ (_00637_, _00798_, _27355_);
  nor _33000_ (_00799_, _00656_, _00650_);
  not _33001_ (_00800_, _00799_);
  nor _33002_ (_00801_, _00694_, _00639_);
  nor _33003_ (_00802_, _00801_, _00800_);
  nor _33004_ (_00803_, _00802_, _00664_);
  or _33005_ (_00804_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _33006_ (_00805_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _00664_);
  or _33007_ (_00806_, _00805_, _00799_);
  and _33008_ (_00807_, _00806_, _27355_);
  and _33009_ (_01239_, _00807_, _00804_);
  or _33010_ (_00808_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _33011_ (_00809_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _00664_);
  or _33012_ (_00810_, _00809_, _00799_);
  and _33013_ (_00811_, _00810_, _27355_);
  and _33014_ (_01241_, _00811_, _00808_);
  or _33015_ (_00812_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _33016_ (_00813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _00664_);
  or _33017_ (_00814_, _00813_, _00799_);
  and _33018_ (_00815_, _00814_, _27355_);
  and _33019_ (_01243_, _00815_, _00812_);
  or _33020_ (_00816_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _33021_ (_00817_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _00664_);
  or _33022_ (_00818_, _00817_, _00799_);
  and _33023_ (_00819_, _00818_, _27355_);
  and _33024_ (_01245_, _00819_, _00816_);
  or _33025_ (_00820_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _33026_ (_00821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _00664_);
  or _33027_ (_00822_, _00821_, _00799_);
  and _33028_ (_00823_, _00822_, _27355_);
  and _33029_ (_01247_, _00823_, _00820_);
  or _33030_ (_00824_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _33031_ (_00825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _00664_);
  or _33032_ (_00826_, _00825_, _00799_);
  and _33033_ (_00827_, _00826_, _27355_);
  and _33034_ (_01248_, _00827_, _00824_);
  or _33035_ (_00828_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _33036_ (_00829_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _00664_);
  or _33037_ (_00830_, _00829_, _00799_);
  and _33038_ (_00831_, _00830_, _27355_);
  and _33039_ (_01250_, _00831_, _00828_);
  or _33040_ (_00832_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _33041_ (_00833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _00664_);
  or _33042_ (_00834_, _00833_, _00799_);
  and _33043_ (_00835_, _00834_, _27355_);
  and _33044_ (_01252_, _00835_, _00832_);
  nor _33045_ (_00836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _33046_ (_00837_, _00836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _33047_ (_00838_, _00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _33048_ (_00839_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _33049_ (_00840_, _00839_, _00639_);
  and _33050_ (_00841_, _00840_, _00838_);
  or _33051_ (_00842_, _00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _33052_ (_00843_, _00842_, _00693_);
  and _33053_ (_00844_, _00843_, _00661_);
  or _33054_ (_00845_, _00844_, _00841_);
  or _33055_ (_00846_, _00845_, _00656_);
  or _33056_ (_00847_, _00657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _33057_ (_00848_, _00847_, _00636_);
  and _33058_ (_00849_, _00848_, _00846_);
  or _33059_ (_01254_, _00849_, _00837_);
  and _33060_ (_00850_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _33061_ (_00851_, _00850_, _00694_);
  or _33062_ (_00852_, _00851_, _00802_);
  and _33063_ (_00853_, _00852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _33064_ (_00854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _00664_);
  nand _33065_ (_00855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _33066_ (_00856_, _00855_, _00799_);
  or _33067_ (_00857_, _00856_, _00854_);
  or _33068_ (_00858_, _00857_, _00853_);
  and _33069_ (_01256_, _00858_, _27355_);
  not _33070_ (_00859_, _00803_);
  and _33071_ (_00860_, _00859_, _00687_);
  or _33072_ (_00861_, _00851_, _00800_);
  and _33073_ (_00862_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _33074_ (_00863_, _00862_, _00861_);
  or _33075_ (_01258_, _00863_, _00860_);
  or _33076_ (_00864_, _00680_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _33077_ (_00865_, _00680_, _00618_);
  and _33078_ (_00866_, _00865_, _27355_);
  and _33079_ (_01260_, _00866_, _00864_);
  or _33080_ (_00867_, _00682_, _00645_);
  or _33081_ (_00868_, _00651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _33082_ (_00869_, _00868_, _27355_);
  and _33083_ (_01262_, _00869_, _00867_);
  and _33084_ (_00870_, _00682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _33085_ (_00871_, _00671_, _00677_);
  and _33086_ (_00872_, _00871_, _00651_);
  or _33087_ (_00873_, _00872_, _00870_);
  and _33088_ (_01264_, _00873_, _27355_);
  and _33089_ (_00874_, _00684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _33090_ (_00875_, _00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _33091_ (_00876_, _00875_, _00683_);
  or _33092_ (_00877_, _00876_, _00874_);
  and _33093_ (_01266_, _00877_, _27355_);
  and _33094_ (_00878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _00664_);
  and _33095_ (_00879_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33096_ (_00880_, _00879_, _00878_);
  and _33097_ (_01267_, _00880_, _27355_);
  and _33098_ (_00881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _00664_);
  and _33099_ (_00882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33100_ (_00883_, _00882_, _00881_);
  and _33101_ (_01269_, _00883_, _27355_);
  and _33102_ (_00884_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _00664_);
  and _33103_ (_00885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33104_ (_00886_, _00885_, _00884_);
  and _33105_ (_01271_, _00886_, _27355_);
  and _33106_ (_00887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _00664_);
  and _33107_ (_00888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33108_ (_00889_, _00888_, _00887_);
  and _33109_ (_01273_, _00889_, _27355_);
  and _33110_ (_00890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _00664_);
  and _33111_ (_00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33112_ (_00892_, _00891_, _00890_);
  and _33113_ (_01275_, _00892_, _27355_);
  and _33114_ (_00893_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _33115_ (_01277_, _00893_, _00837_);
  and _33116_ (_00894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _33117_ (_00895_, _00894_, _00854_);
  and _33118_ (_01279_, _00895_, _27355_);
  nor _33119_ (_00896_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _33120_ (_00897_, _00896_, _00775_);
  and _33121_ (_01281_, _00897_, _00758_);
  nor _33122_ (_00898_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _33123_ (_00899_, _00898_, _00776_);
  and _33124_ (_01282_, _00899_, _00758_);
  nor _33125_ (_00900_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _33126_ (_00901_, _00900_, _00777_);
  and _33127_ (_01284_, _00901_, _00758_);
  or _33128_ (_00902_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _33129_ (_00903_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _33130_ (_00904_, _00903_, _00902_);
  and _33131_ (_00905_, _00904_, _00749_);
  and _33132_ (_00906_, _00733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _33133_ (_00907_, _00906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _33134_ (_00908_, _00907_, _00722_);
  or _33135_ (_00909_, _00908_, _00905_);
  and _33136_ (_00910_, _00909_, _00758_);
  nor _33137_ (_00911_, _00622_, _26521_);
  and _33138_ (_00912_, _00911_, _00761_);
  or _33139_ (_01286_, _00912_, _00910_);
  not _33140_ (_00913_, _00781_);
  and _33141_ (_00914_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _33142_ (_00915_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _33143_ (_00916_, _00915_, _00914_);
  and _33144_ (_00917_, _00916_, _00758_);
  nand _33145_ (_00918_, _00621_, _26512_);
  nand _33146_ (_00919_, _00622_, _26521_);
  and _33147_ (_00920_, _00919_, _00761_);
  and _33148_ (_00921_, _00920_, _00918_);
  or _33149_ (_01288_, _00921_, _00917_);
  nor _33150_ (_00922_, _00781_, _00728_);
  and _33151_ (_00923_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _33152_ (_00924_, _00923_, _00922_);
  and _33153_ (_00925_, _00924_, _00758_);
  nand _33154_ (_00926_, _00621_, _26505_);
  nand _33155_ (_00927_, _00622_, _26512_);
  and _33156_ (_00928_, _00927_, _00761_);
  and _33157_ (_00929_, _00928_, _00926_);
  or _33158_ (_01290_, _00929_, _00925_);
  nor _33159_ (_00930_, _00781_, _00724_);
  and _33160_ (_00931_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _33161_ (_00932_, _00931_, _00930_);
  and _33162_ (_00933_, _00932_, _00758_);
  nand _33163_ (_00934_, _00622_, _26505_);
  nand _33164_ (_00935_, _00621_, _26497_);
  and _33165_ (_00936_, _00935_, _00761_);
  and _33166_ (_00937_, _00936_, _00934_);
  or _33167_ (_01292_, _00937_, _00933_);
  and _33168_ (_00938_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _33169_ (_00939_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _33170_ (_00940_, _00939_, _00938_);
  and _33171_ (_00941_, _00940_, _00758_);
  nand _33172_ (_00942_, _00621_, _26489_);
  nand _33173_ (_00943_, _00622_, _26497_);
  and _33174_ (_00944_, _00943_, _00761_);
  and _33175_ (_00945_, _00944_, _00942_);
  or _33176_ (_01294_, _00945_, _00941_);
  and _33177_ (_00946_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _33178_ (_00947_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _33179_ (_00948_, _00947_, _00946_);
  and _33180_ (_00949_, _00948_, _00758_);
  nand _33181_ (_00950_, _00622_, _26489_);
  nand _33182_ (_00951_, _00621_, _26482_);
  and _33183_ (_00952_, _00951_, _00761_);
  and _33184_ (_00953_, _00952_, _00950_);
  or _33185_ (_01296_, _00953_, _00949_);
  and _33186_ (_00954_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _33187_ (_00955_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _33188_ (_00956_, _00955_, _00954_);
  and _33189_ (_00957_, _00956_, _00758_);
  nand _33190_ (_00959_, _00621_, _26475_);
  nand _33191_ (_00960_, _00622_, _26482_);
  and _33192_ (_00961_, _00960_, _00761_);
  and _33193_ (_00962_, _00961_, _00959_);
  or _33194_ (_01297_, _00962_, _00957_);
  and _33195_ (_00963_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _33196_ (_00964_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _33197_ (_00965_, _00964_, _00963_);
  and _33198_ (_00966_, _00965_, _00758_);
  nand _33199_ (_00967_, _00621_, _26543_);
  nand _33200_ (_00968_, _00622_, _26475_);
  and _33201_ (_00969_, _00968_, _00761_);
  and _33202_ (_00970_, _00969_, _00967_);
  or _33203_ (_01299_, _00970_, _00966_);
  and _33204_ (_00971_, _00757_, _00622_);
  nand _33205_ (_00972_, _00971_, _26543_);
  and _33206_ (_00973_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _33207_ (_00974_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _33208_ (_00975_, _00974_, _00973_);
  or _33209_ (_00976_, _00975_, _00757_);
  and _33210_ (_00977_, _00976_, _27355_);
  and _33211_ (_01301_, _00977_, _00972_);
  and _33212_ (_00978_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _33213_ (_00979_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _33214_ (_00980_, _00979_, _00978_);
  and _33215_ (_00981_, _00980_, _00758_);
  or _33216_ (_00982_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _33217_ (_00983_, _00982_, _00622_);
  and _33218_ (_00984_, _00983_, _00761_);
  or _33219_ (_01303_, _00984_, _00981_);
  nand _33220_ (_00986_, _00785_, _26521_);
  or _33221_ (_00987_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _33222_ (_00988_, _00987_, _27355_);
  and _33223_ (_01305_, _00988_, _00986_);
  or _33224_ (_00989_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _33225_ (_00990_, _00989_, _27355_);
  nand _33226_ (_00991_, _00785_, _26512_);
  and _33227_ (_01307_, _00991_, _00990_);
  or _33228_ (_00992_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _33229_ (_00993_, _00992_, _27355_);
  nand _33230_ (_00994_, _00785_, _26505_);
  and _33231_ (_01309_, _00994_, _00993_);
  or _33232_ (_00995_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _33233_ (_00996_, _00995_, _27355_);
  nand _33234_ (_00997_, _00785_, _26497_);
  and _33235_ (_01310_, _00997_, _00996_);
  or _33236_ (_00998_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _33237_ (_00999_, _00998_, _27355_);
  nand _33238_ (_01000_, _00785_, _26489_);
  and _33239_ (_01312_, _01000_, _00999_);
  or _33240_ (_01002_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _33241_ (_01003_, _01002_, _27355_);
  nand _33242_ (_01004_, _00785_, _26482_);
  and _33243_ (_01314_, _01004_, _01003_);
  or _33244_ (_01005_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _33245_ (_01006_, _01005_, _27355_);
  nand _33246_ (_01007_, _00785_, _26475_);
  and _33247_ (_01316_, _01007_, _01006_);
  nand _33248_ (_01008_, _25514_, _25055_);
  or _33249_ (_01009_, _25055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _33250_ (_01010_, _01009_, _00789_);
  and _33251_ (_01011_, _01010_, _01008_);
  not _33252_ (_01012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _33253_ (_01013_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01012_);
  or _33254_ (_01014_, _01013_, _00621_);
  nor _33255_ (_01015_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _33256_ (_01016_, _01015_, _01014_);
  nor _33257_ (_01017_, _01016_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _33258_ (_01018_, _01017_, _00789_);
  or _33259_ (_01019_, _01018_, _00792_);
  or _33260_ (_01020_, _01019_, _01011_);
  nand _33261_ (_01021_, _00792_, _26521_);
  and _33262_ (_01022_, _01021_, _27355_);
  and _33263_ (_01318_, _01022_, _01020_);
  or _33264_ (_01023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _33265_ (_01024_, _01023_, _00789_);
  nand _33266_ (_01025_, _27079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _33267_ (_01026_, _01025_, _00789_);
  or _33268_ (_01027_, _01026_, _27080_);
  and _33269_ (_01028_, _01027_, _01024_);
  or _33270_ (_01029_, _01028_, _00792_);
  nand _33271_ (_01030_, _00792_, _26512_);
  and _33272_ (_01031_, _01030_, _27355_);
  and _33273_ (_01320_, _01031_, _01029_);
  not _33274_ (_01032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _33275_ (_01033_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _33276_ (_01034_, _00640_, _01033_);
  nor _33277_ (_01035_, _01034_, _01032_);
  and _33278_ (_01036_, _01034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _33279_ (_01037_, _01036_, _01035_);
  or _33280_ (_01038_, _01037_, _00789_);
  or _33281_ (_01039_, _25716_, _01032_);
  nand _33282_ (_01040_, _01039_, _00789_);
  or _33283_ (_01041_, _01040_, _25718_);
  and _33284_ (_01042_, _01041_, _01038_);
  or _33285_ (_01043_, _01042_, _00792_);
  nand _33286_ (_01044_, _00792_, _26505_);
  and _33287_ (_01045_, _01044_, _27355_);
  and _33288_ (_01322_, _01045_, _01043_);
  and _33289_ (_01046_, _00789_, _25778_);
  nand _33290_ (_01047_, _01046_, _25514_);
  or _33291_ (_01048_, _01046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _33292_ (_01049_, _01048_, _00793_);
  and _33293_ (_01050_, _01049_, _01047_);
  nor _33294_ (_01051_, _00793_, _26497_);
  or _33295_ (_01052_, _01051_, _01050_);
  and _33296_ (_01323_, _01052_, _27355_);
  and _33297_ (_01053_, _00789_, _25838_);
  nand _33298_ (_01054_, _01053_, _25514_);
  or _33299_ (_01055_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _33300_ (_01056_, _01055_, _00793_);
  and _33301_ (_01057_, _01056_, _01054_);
  nor _33302_ (_01058_, _00793_, _26489_);
  or _33303_ (_01059_, _01058_, _01057_);
  and _33304_ (_01325_, _01059_, _27355_);
  and _33305_ (_01060_, _00789_, _25905_);
  nand _33306_ (_01061_, _01060_, _25514_);
  or _33307_ (_01062_, _01060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _33308_ (_01063_, _01062_, _01061_);
  or _33309_ (_01064_, _01063_, _00792_);
  nand _33310_ (_01065_, _00792_, _26482_);
  and _33311_ (_01066_, _01065_, _27355_);
  and _33312_ (_01327_, _01066_, _01064_);
  and _33313_ (_01067_, _00789_, _25972_);
  nand _33314_ (_01068_, _01067_, _25514_);
  or _33315_ (_01069_, _01067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _33316_ (_01070_, _01069_, _00793_);
  and _33317_ (_01071_, _01070_, _01068_);
  nor _33318_ (_01072_, _00793_, _26475_);
  or _33319_ (_01073_, _01072_, _01071_);
  and _33320_ (_01329_, _01073_, _27355_);
  and _33321_ (_01640_, t2_i, _27355_);
  nor _33322_ (_01074_, t2_i, rst);
  and _33323_ (_01643_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _33324_ (_01075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _27355_);
  nor _33325_ (_01646_, _01075_, t2ex_i);
  and _33326_ (_01649_, t2ex_i, _27355_);
  and _33327_ (_01076_, _26457_, _26939_);
  and _33328_ (_01077_, _01076_, _27666_);
  nand _33329_ (_01078_, _01077_, _26543_);
  and _33330_ (_01079_, _01076_, _27577_);
  not _33331_ (_01080_, _01079_);
  and _33332_ (_01081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _33333_ (_01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _33334_ (_01083_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _33335_ (_01084_, _01083_, _01081_);
  not _33336_ (_01085_, _01084_);
  and _33337_ (_01086_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _33338_ (_01087_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _33339_ (_01088_, _01087_, _01086_);
  or _33340_ (_01089_, _01077_, _01088_);
  and _33341_ (_01090_, _01089_, _01080_);
  and _33342_ (_01091_, _01090_, _01078_);
  and _33343_ (_01092_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _33344_ (_01093_, _01092_, _01091_);
  and _33345_ (_01652_, _01093_, _27355_);
  nand _33346_ (_01094_, _01079_, _26543_);
  nor _33347_ (_01095_, _01077_, _01085_);
  or _33348_ (_01096_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _33349_ (_01097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _33350_ (_01098_, _01095_, _01097_);
  and _33351_ (_01099_, _01098_, _01096_);
  or _33352_ (_01100_, _01099_, _01079_);
  and _33353_ (_01101_, _01100_, _27355_);
  and _33354_ (_01655_, _01101_, _01094_);
  not _33355_ (_01102_, _01082_);
  or _33356_ (_01103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _33357_ (_01104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _33358_ (_01105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01104_);
  and _33359_ (_01106_, _01105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _33360_ (_01107_, _01106_, _01103_);
  and _33361_ (_01108_, _01076_, _25905_);
  and _33362_ (_01109_, _01108_, _27576_);
  and _33363_ (_01110_, _01076_, _27669_);
  nor _33364_ (_01111_, _01110_, _01109_);
  and _33365_ (_01112_, _01111_, _01107_);
  and _33366_ (_01113_, _01112_, _01102_);
  and _33367_ (_01114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _33368_ (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _33369_ (_01116_, _01115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _33370_ (_01117_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _33371_ (_01118_, _01117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _33372_ (_01119_, _01118_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _33373_ (_01120_, _01119_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _33374_ (_01121_, _01120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _33375_ (_01122_, _01121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _33376_ (_01123_, _01122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _33377_ (_01124_, _01123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _33378_ (_01125_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _33379_ (_01126_, _01125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _33380_ (_01127_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _33381_ (_01128_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _33382_ (_01129_, _01128_);
  nand _33383_ (_01130_, _01129_, _01113_);
  or _33384_ (_01131_, _01113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _33385_ (_01132_, _01131_, _27355_);
  and _33386_ (_01658_, _01132_, _01130_);
  nand _33387_ (_01133_, _01110_, _26543_);
  not _33388_ (_01134_, _01109_);
  not _33389_ (_01135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _33390_ (_01136_, _01081_, _01135_);
  and _33391_ (_01137_, _01136_, _01082_);
  and _33392_ (_01138_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _33393_ (_01139_, _01137_);
  not _33394_ (_01140_, _01083_);
  and _33395_ (_01141_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _33396_ (_01142_, _01128_, _01107_);
  and _33397_ (_01143_, _01142_, _01141_);
  and _33398_ (_01144_, _01119_, _01107_);
  or _33399_ (_01145_, _01144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _33400_ (_01146_, _01144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _33401_ (_01147_, _01146_, _01145_);
  or _33402_ (_01148_, _01147_, _01143_);
  and _33403_ (_01149_, _01148_, _01139_);
  or _33404_ (_01150_, _01149_, _01138_);
  or _33405_ (_01151_, _01150_, _01110_);
  and _33406_ (_01152_, _01151_, _01134_);
  and _33407_ (_01153_, _01152_, _01133_);
  and _33408_ (_01154_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _33409_ (_01155_, _01154_, _01153_);
  and _33410_ (_01661_, _01155_, _27355_);
  nand _33411_ (_01156_, _01109_, _26543_);
  nor _33412_ (_01157_, _01137_, _01097_);
  and _33413_ (_01158_, _01139_, _01107_);
  and _33414_ (_01159_, _01158_, _01127_);
  or _33415_ (_01160_, _01159_, _01157_);
  nand _33416_ (_01161_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _33417_ (_01162_, _01161_, _01142_);
  and _33418_ (_01163_, _01162_, _01160_);
  nand _33419_ (_01164_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _33420_ (_01165_, _01164_, _01111_);
  or _33421_ (_01166_, _01165_, _01163_);
  nand _33422_ (_01167_, _01110_, _01097_);
  and _33423_ (_01168_, _01167_, _27355_);
  and _33424_ (_01169_, _01168_, _01166_);
  and _33425_ (_01664_, _01169_, _01156_);
  not _33426_ (_01170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor _33427_ (_01171_, _01111_, _01170_);
  and _33428_ (_01172_, _01158_, _01082_);
  and _33429_ (_01173_, _01172_, _01111_);
  and _33430_ (_01174_, _01173_, _01128_);
  or _33431_ (_01175_, _01174_, _01171_);
  and _33432_ (_01667_, _01175_, _27355_);
  or _33433_ (_01176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _33434_ (_01177_, _00038_, _26923_);
  or _33435_ (_01178_, _01177_, _01176_);
  nand _33436_ (_01179_, _26926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _33437_ (_01180_, _01179_, _01177_);
  or _33438_ (_01181_, _01180_, _26927_);
  and _33439_ (_01182_, _01181_, _01178_);
  and _33440_ (_01183_, _01076_, _00035_);
  or _33441_ (_01184_, _01183_, _01182_);
  nand _33442_ (_01185_, _01183_, _26543_);
  and _33443_ (_01186_, _01185_, _27355_);
  and _33444_ (_01670_, _01186_, _01184_);
  or _33445_ (_01187_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _33446_ (_01188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _33447_ (_01189_, _01084_, _01188_);
  and _33448_ (_01190_, _01189_, _01187_);
  or _33449_ (_01191_, _01190_, _01077_);
  nand _33450_ (_01192_, _01077_, _26521_);
  and _33451_ (_01193_, _01192_, _01191_);
  or _33452_ (_01194_, _01193_, _01079_);
  not _33453_ (_01195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _33454_ (_01196_, _01079_, _01195_);
  and _33455_ (_01197_, _01196_, _27355_);
  and _33456_ (_02203_, _01197_, _01194_);
  nand _33457_ (_01198_, _01077_, _26512_);
  and _33458_ (_01199_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _33459_ (_01200_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _33460_ (_01201_, _01200_, _01199_);
  or _33461_ (_01202_, _01201_, _01077_);
  and _33462_ (_01203_, _01202_, _01080_);
  and _33463_ (_01204_, _01203_, _01198_);
  and _33464_ (_01205_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _33465_ (_01206_, _01205_, _01204_);
  and _33466_ (_02205_, _01206_, _27355_);
  nand _33467_ (_01207_, _01077_, _26505_);
  and _33468_ (_01208_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _33469_ (_01209_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _33470_ (_01210_, _01209_, _01208_);
  or _33471_ (_01211_, _01210_, _01077_);
  and _33472_ (_01212_, _01211_, _01080_);
  and _33473_ (_01213_, _01212_, _01207_);
  and _33474_ (_01214_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _33475_ (_01215_, _01214_, _01213_);
  and _33476_ (_02207_, _01215_, _27355_);
  nand _33477_ (_01216_, _01077_, _26497_);
  and _33478_ (_01217_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _33479_ (_01218_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _33480_ (_01219_, _01218_, _01217_);
  or _33481_ (_01220_, _01219_, _01077_);
  and _33482_ (_01221_, _01220_, _01080_);
  and _33483_ (_01222_, _01221_, _01216_);
  and _33484_ (_01223_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _33485_ (_01224_, _01223_, _01222_);
  and _33486_ (_02209_, _01224_, _27355_);
  nand _33487_ (_01225_, _01077_, _26489_);
  and _33488_ (_01226_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _33489_ (_01227_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _33490_ (_01228_, _01227_, _01226_);
  or _33491_ (_01229_, _01228_, _01077_);
  and _33492_ (_01230_, _01229_, _01080_);
  and _33493_ (_01231_, _01230_, _01225_);
  and _33494_ (_01232_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _33495_ (_01233_, _01232_, _01231_);
  and _33496_ (_02211_, _01233_, _27355_);
  nand _33497_ (_01234_, _01077_, _26482_);
  and _33498_ (_01235_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _33499_ (_01236_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _33500_ (_01237_, _01236_, _01235_);
  or _33501_ (_01238_, _01237_, _01077_);
  and _33502_ (_01240_, _01238_, _01080_);
  and _33503_ (_01242_, _01240_, _01234_);
  and _33504_ (_01244_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _33505_ (_01246_, _01244_, _01242_);
  and _33506_ (_02213_, _01246_, _27355_);
  nand _33507_ (_01249_, _01077_, _26475_);
  and _33508_ (_01251_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _33509_ (_01253_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _33510_ (_01255_, _01253_, _01251_);
  or _33511_ (_01257_, _01255_, _01077_);
  and _33512_ (_01259_, _01257_, _01080_);
  and _33513_ (_01261_, _01259_, _01249_);
  and _33514_ (_01263_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _33515_ (_01265_, _01263_, _01261_);
  and _33516_ (_02215_, _01265_, _27355_);
  and _33517_ (_01268_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  not _33518_ (_01270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _33519_ (_01272_, _01095_, _01270_);
  or _33520_ (_01274_, _01272_, _01268_);
  or _33521_ (_01276_, _01274_, _01079_);
  nand _33522_ (_01278_, _01079_, _26521_);
  and _33523_ (_01280_, _01278_, _27355_);
  and _33524_ (_02217_, _01280_, _01276_);
  nand _33525_ (_01283_, _01079_, _26512_);
  and _33526_ (_01285_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not _33527_ (_01287_, _01095_);
  and _33528_ (_01289_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _33529_ (_01291_, _01289_, _01285_);
  or _33530_ (_01293_, _01291_, _01079_);
  and _33531_ (_01295_, _01293_, _27355_);
  and _33532_ (_02219_, _01295_, _01283_);
  nand _33533_ (_01298_, _01079_, _26505_);
  and _33534_ (_01300_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _33535_ (_01302_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _33536_ (_01304_, _01302_, _01300_);
  or _33537_ (_01306_, _01304_, _01079_);
  and _33538_ (_01308_, _01306_, _27355_);
  and _33539_ (_02221_, _01308_, _01298_);
  nand _33540_ (_01311_, _01079_, _26497_);
  and _33541_ (_01313_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _33542_ (_01315_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _33543_ (_01317_, _01315_, _01313_);
  or _33544_ (_01319_, _01317_, _01079_);
  and _33545_ (_01321_, _01319_, _27355_);
  and _33546_ (_02223_, _01321_, _01311_);
  nand _33547_ (_01324_, _01079_, _26489_);
  and _33548_ (_01326_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _33549_ (_01328_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _33550_ (_01330_, _01328_, _01326_);
  or _33551_ (_01331_, _01330_, _01079_);
  and _33552_ (_01332_, _01331_, _27355_);
  and _33553_ (_02225_, _01332_, _01324_);
  nand _33554_ (_01333_, _01079_, _26482_);
  and _33555_ (_01334_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _33556_ (_01335_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _33557_ (_01336_, _01335_, _01334_);
  or _33558_ (_01337_, _01336_, _01079_);
  and _33559_ (_01338_, _01337_, _27355_);
  and _33560_ (_02227_, _01338_, _01333_);
  nand _33561_ (_01339_, _01079_, _26475_);
  and _33562_ (_01340_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _33563_ (_01341_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _33564_ (_01342_, _01341_, _01340_);
  or _33565_ (_01343_, _01342_, _01079_);
  and _33566_ (_01344_, _01343_, _27355_);
  and _33567_ (_02229_, _01344_, _01339_);
  and _33568_ (_01345_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _33569_ (_01346_, _01083_, _01195_);
  nand _33570_ (_01347_, _01346_, _01128_);
  nand _33571_ (_01348_, _01347_, _01345_);
  or _33572_ (_01349_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _33573_ (_01350_, _01349_, _01139_);
  and _33574_ (_01351_, _01350_, _01348_);
  nand _33575_ (_01352_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _33576_ (_01353_, _01352_, _01111_);
  or _33577_ (_01354_, _01353_, _01351_);
  nand _33578_ (_01355_, _01109_, _01188_);
  nand _33579_ (_01356_, _01110_, _26521_);
  and _33580_ (_01357_, _01356_, _27355_);
  and _33581_ (_01358_, _01357_, _01355_);
  and _33582_ (_02231_, _01358_, _01354_);
  and _33583_ (_01359_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _33584_ (_01360_, _01359_, _01158_);
  and _33585_ (_01361_, _01360_, _01128_);
  and _33586_ (_01362_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _33587_ (_01363_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _33588_ (_01364_, _01114_, _01107_);
  nor _33589_ (_01365_, _01364_, _01137_);
  and _33590_ (_01366_, _01365_, _01363_);
  nor _33591_ (_01367_, _01366_, _01362_);
  nand _33592_ (_01368_, _01367_, _01111_);
  or _33593_ (_01369_, _01368_, _01361_);
  nand _33594_ (_01370_, _01110_, _26512_);
  or _33595_ (_01371_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _33596_ (_01372_, _01371_, _27355_);
  and _33597_ (_01373_, _01372_, _01370_);
  and _33598_ (_02233_, _01373_, _01369_);
  and _33599_ (_01374_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _33600_ (_01375_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _33601_ (_01376_, _01375_, _01142_);
  not _33602_ (_01377_, _01364_);
  nor _33603_ (_01378_, _01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _33604_ (_01379_, _01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _33605_ (_01380_, _01379_, _01378_);
  or _33606_ (_01381_, _01380_, _01376_);
  and _33607_ (_01382_, _01381_, _01139_);
  or _33608_ (_01383_, _01382_, _01374_);
  or _33609_ (_01384_, _01383_, _01110_);
  nand _33610_ (_01385_, _01110_, _26505_);
  and _33611_ (_01386_, _01385_, _01134_);
  and _33612_ (_01387_, _01386_, _01384_);
  and _33613_ (_01388_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _33614_ (_01389_, _01388_, _01387_);
  and _33615_ (_02235_, _01389_, _27355_);
  not _33616_ (_01390_, _01110_);
  nor _33617_ (_01391_, _01390_, _26497_);
  and _33618_ (_01392_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _33619_ (_01393_, _01392_, _01142_);
  nand _33620_ (_01394_, _01115_, _01107_);
  and _33621_ (_01395_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _33622_ (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _33623_ (_01397_, _01396_, _01137_);
  or _33624_ (_01398_, _01397_, _01395_);
  or _33625_ (_01399_, _01398_, _01393_);
  or _33626_ (_01400_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _33627_ (_01401_, _01400_, _01111_);
  and _33628_ (_01402_, _01401_, _01399_);
  and _33629_ (_01403_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _33630_ (_01404_, _01403_, _01402_);
  or _33631_ (_01405_, _01404_, _01391_);
  and _33632_ (_02237_, _01405_, _27355_);
  and _33633_ (_01406_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _33634_ (_01407_, _01406_, _01142_);
  nand _33635_ (_01408_, _01116_, _01107_);
  and _33636_ (_01409_, _01408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _33637_ (_01410_, _01408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _33638_ (_01411_, _01410_, _01137_);
  or _33639_ (_01412_, _01411_, _01409_);
  or _33640_ (_01413_, _01412_, _01407_);
  nor _33641_ (_01414_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _33642_ (_01415_, _01414_, _01110_);
  and _33643_ (_01416_, _01415_, _01413_);
  nor _33644_ (_01417_, _01390_, _26489_);
  or _33645_ (_01418_, _01417_, _01416_);
  or _33646_ (_01419_, _01418_, _01109_);
  or _33647_ (_01420_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _33648_ (_01421_, _01420_, _27355_);
  and _33649_ (_02239_, _01421_, _01419_);
  and _33650_ (_01422_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _33651_ (_01423_, _01422_, _01142_);
  nand _33652_ (_01424_, _01117_, _01107_);
  and _33653_ (_01425_, _01424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _33654_ (_01426_, _01424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _33655_ (_01427_, _01426_, _01137_);
  or _33656_ (_01428_, _01427_, _01425_);
  or _33657_ (_01429_, _01428_, _01423_);
  nor _33658_ (_01430_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _33659_ (_01431_, _01430_, _01110_);
  and _33660_ (_01432_, _01431_, _01429_);
  nor _33661_ (_01433_, _01390_, _26482_);
  or _33662_ (_01434_, _01433_, _01432_);
  or _33663_ (_01435_, _01434_, _01109_);
  or _33664_ (_01436_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _33665_ (_01437_, _01436_, _27355_);
  and _33666_ (_02241_, _01437_, _01435_);
  nor _33667_ (_01438_, _01390_, _26475_);
  and _33668_ (_01439_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _33669_ (_01440_, _01439_, _01142_);
  and _33670_ (_01441_, _01118_, _01107_);
  nor _33671_ (_01442_, _01441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _33672_ (_01443_, _01442_, _01144_);
  or _33673_ (_01444_, _01443_, _01137_);
  or _33674_ (_01445_, _01444_, _01440_);
  nor _33675_ (_01446_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _33676_ (_01447_, _01446_, _01110_);
  and _33677_ (_01448_, _01447_, _01445_);
  or _33678_ (_01449_, _01448_, _01109_);
  or _33679_ (_01450_, _01449_, _01438_);
  or _33680_ (_01451_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _33681_ (_01452_, _01451_, _27355_);
  and _33682_ (_02243_, _01452_, _01450_);
  nor _33683_ (_01453_, _01083_, _01270_);
  and _33684_ (_01454_, _01453_, _01142_);
  and _33685_ (_01455_, _01120_, _01107_);
  or _33686_ (_01456_, _01455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _33687_ (_01457_, _01455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _33688_ (_01458_, _01457_, _01456_);
  or _33689_ (_01459_, _01458_, _01137_);
  or _33690_ (_01460_, _01459_, _01454_);
  and _33691_ (_01461_, _01137_, _01270_);
  nor _33692_ (_01462_, _01461_, _01110_);
  and _33693_ (_01463_, _01462_, _01460_);
  and _33694_ (_01464_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _33695_ (_01465_, _01464_, _01109_);
  or _33696_ (_01466_, _01465_, _01463_);
  nand _33697_ (_01467_, _01109_, _26521_);
  and _33698_ (_01468_, _01467_, _27355_);
  and _33699_ (_02245_, _01468_, _01466_);
  and _33700_ (_01469_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _33701_ (_01470_, _01469_, _01142_);
  and _33702_ (_01471_, _01121_, _01107_);
  or _33703_ (_01472_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _33704_ (_01473_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _33705_ (_01474_, _01473_, _01472_);
  or _33706_ (_01475_, _01474_, _01137_);
  or _33707_ (_01476_, _01475_, _01470_);
  nor _33708_ (_01477_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _33709_ (_01478_, _01477_, _01110_);
  and _33710_ (_01479_, _01478_, _01476_);
  and _33711_ (_01480_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _33712_ (_01481_, _01480_, _01109_);
  or _33713_ (_01482_, _01481_, _01479_);
  nand _33714_ (_01483_, _01109_, _26512_);
  and _33715_ (_01484_, _01483_, _27355_);
  and _33716_ (_02247_, _01484_, _01482_);
  and _33717_ (_01485_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _33718_ (_01486_, _01485_, _01142_);
  nand _33719_ (_01487_, _01122_, _01107_);
  and _33720_ (_01488_, _01487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _33721_ (_01489_, _01487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _33722_ (_01490_, _01489_, _01137_);
  or _33723_ (_01491_, _01490_, _01488_);
  or _33724_ (_01492_, _01491_, _01486_);
  nor _33725_ (_01493_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _33726_ (_01494_, _01493_, _01110_);
  and _33727_ (_01495_, _01494_, _01492_);
  and _33728_ (_01496_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _33729_ (_01497_, _01496_, _01109_);
  or _33730_ (_01498_, _01497_, _01495_);
  nand _33731_ (_01499_, _01109_, _26505_);
  and _33732_ (_01500_, _01499_, _27355_);
  and _33733_ (_02249_, _01500_, _01498_);
  and _33734_ (_01501_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _33735_ (_01502_, _01501_, _01142_);
  nand _33736_ (_01503_, _01123_, _01107_);
  and _33737_ (_01504_, _01503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor _33738_ (_01505_, _01503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _33739_ (_01506_, _01505_, _01137_);
  or _33740_ (_01507_, _01506_, _01504_);
  or _33741_ (_01508_, _01507_, _01502_);
  nor _33742_ (_01509_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _33743_ (_01510_, _01509_, _01110_);
  and _33744_ (_01511_, _01510_, _01508_);
  and _33745_ (_01512_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _33746_ (_01513_, _01512_, _01109_);
  or _33747_ (_01514_, _01513_, _01511_);
  nand _33748_ (_01515_, _01109_, _26497_);
  and _33749_ (_01516_, _01515_, _27355_);
  and _33750_ (_02251_, _01516_, _01514_);
  nand _33751_ (_01517_, _01109_, _26489_);
  and _33752_ (_01518_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _33753_ (_01519_, _01518_, _01142_);
  nand _33754_ (_01520_, _01124_, _01107_);
  and _33755_ (_01521_, _01520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _33756_ (_01522_, _01520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _33757_ (_01523_, _01522_, _01137_);
  or _33758_ (_01524_, _01523_, _01521_);
  or _33759_ (_01525_, _01524_, _01519_);
  nor _33760_ (_01526_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _33761_ (_01527_, _01526_, _01110_);
  and _33762_ (_01528_, _01527_, _01525_);
  and _33763_ (_01529_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _33764_ (_01530_, _01529_, _01109_);
  or _33765_ (_01531_, _01530_, _01528_);
  and _33766_ (_01532_, _01531_, _27355_);
  and _33767_ (_02253_, _01532_, _01517_);
  and _33768_ (_01533_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _33769_ (_01534_, _01533_, _01142_);
  nand _33770_ (_01535_, _01125_, _01107_);
  and _33771_ (_01536_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _33772_ (_01537_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _33773_ (_01538_, _01537_, _01137_);
  or _33774_ (_01539_, _01538_, _01536_);
  or _33775_ (_01540_, _01539_, _01534_);
  nor _33776_ (_01541_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _33777_ (_01542_, _01541_, _01110_);
  and _33778_ (_01543_, _01542_, _01540_);
  and _33779_ (_01544_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _33780_ (_01545_, _01544_, _01109_);
  or _33781_ (_01546_, _01545_, _01543_);
  nand _33782_ (_01547_, _01109_, _26482_);
  and _33783_ (_01548_, _01547_, _27355_);
  and _33784_ (_02255_, _01548_, _01546_);
  and _33785_ (_01549_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _33786_ (_01550_, _01549_, _01142_);
  nand _33787_ (_01551_, _01126_, _01107_);
  and _33788_ (_01552_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _33789_ (_01553_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _33790_ (_01554_, _01553_, _01137_);
  or _33791_ (_01555_, _01554_, _01552_);
  or _33792_ (_01556_, _01555_, _01550_);
  nor _33793_ (_01557_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _33794_ (_01558_, _01557_, _01110_);
  and _33795_ (_01559_, _01558_, _01556_);
  and _33796_ (_01560_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _33797_ (_01561_, _01560_, _01109_);
  or _33798_ (_01562_, _01561_, _01559_);
  nand _33799_ (_01563_, _01109_, _26475_);
  and _33800_ (_01564_, _01563_, _27355_);
  and _33801_ (_02257_, _01564_, _01562_);
  and _33802_ (_01565_, _01177_, _25055_);
  nand _33803_ (_01566_, _01565_, _25514_);
  not _33804_ (_01567_, _01183_);
  or _33805_ (_01568_, _01565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _33806_ (_01569_, _01568_, _01567_);
  and _33807_ (_01570_, _01569_, _01566_);
  nor _33808_ (_01571_, _01567_, _26521_);
  or _33809_ (_01572_, _01571_, _01570_);
  and _33810_ (_02259_, _01572_, _27355_);
  and _33811_ (_01573_, _01177_, _26947_);
  nand _33812_ (_01574_, _01573_, _25514_);
  or _33813_ (_01575_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _33814_ (_01576_, _01575_, _01574_);
  or _33815_ (_01577_, _01576_, _01183_);
  nand _33816_ (_01578_, _01183_, _26512_);
  and _33817_ (_01579_, _01578_, _27355_);
  and _33818_ (_02261_, _01579_, _01577_);
  nand _33819_ (_01580_, _01177_, _27237_);
  and _33820_ (_01581_, _01580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _33821_ (_01582_, _01581_, _01183_);
  and _33822_ (_01583_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _33823_ (_01584_, _01583_, _25718_);
  and _33824_ (_01585_, _01584_, _01177_);
  or _33825_ (_01586_, _01585_, _01582_);
  nand _33826_ (_01587_, _01183_, _26505_);
  and _33827_ (_01588_, _01587_, _27355_);
  and _33828_ (_02263_, _01588_, _01586_);
  and _33829_ (_01589_, _01177_, _25778_);
  or _33830_ (_01590_, _01589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _33831_ (_01591_, _01590_, _01567_);
  nand _33832_ (_01592_, _01589_, _25514_);
  and _33833_ (_01593_, _01592_, _01591_);
  nor _33834_ (_01594_, _01567_, _26497_);
  or _33835_ (_01595_, _01594_, _01593_);
  and _33836_ (_02265_, _01595_, _27355_);
  and _33837_ (_01596_, _01177_, _25838_);
  or _33838_ (_01597_, _01596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _33839_ (_01598_, _01597_, _01567_);
  nand _33840_ (_01599_, _01596_, _25514_);
  and _33841_ (_01600_, _01599_, _01598_);
  nor _33842_ (_01601_, _01567_, _26489_);
  or _33843_ (_01602_, _01601_, _01600_);
  and _33844_ (_02267_, _01602_, _27355_);
  and _33845_ (_01603_, _01177_, _25905_);
  or _33846_ (_01604_, _01603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _33847_ (_01605_, _01604_, _01567_);
  nand _33848_ (_01606_, _01603_, _25514_);
  and _33849_ (_01607_, _01606_, _01605_);
  nor _33850_ (_01608_, _01567_, _26482_);
  or _33851_ (_01609_, _01608_, _01607_);
  and _33852_ (_02269_, _01609_, _27355_);
  and _33853_ (_01610_, _01081_, _01170_);
  or _33854_ (_01611_, _01610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _33855_ (_01612_, _01611_, _01177_);
  nand _33856_ (_01613_, _27024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _33857_ (_01614_, _01613_, _01177_);
  or _33858_ (_01615_, _01614_, _27025_);
  and _33859_ (_01616_, _01615_, _01612_);
  or _33860_ (_01617_, _01616_, _01183_);
  nand _33861_ (_01618_, _01183_, _26475_);
  and _33862_ (_01619_, _01618_, _27355_);
  and _33863_ (_02271_, _01619_, _01617_);
  and _33864_ (_01620_, _25101_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _33865_ (_01621_, _01620_, _25116_);
  nor _33866_ (_01622_, _25053_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _33867_ (_01623_, _01622_, _01621_);
  nor _33868_ (_01624_, _26436_, _26389_);
  and _33869_ (_01625_, _01624_, _26454_);
  nand _33870_ (_01626_, _26545_, _01625_);
  nor _33871_ (_01627_, _26436_, _26390_);
  and _33872_ (_01628_, _26938_, _26939_);
  and _33873_ (_01629_, _01628_, _26940_);
  not _33874_ (_01630_, _01629_);
  and _33875_ (_01631_, _01630_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _33876_ (_01632_, _01631_, _26996_);
  and _33877_ (_01633_, _01632_, _25116_);
  nor _33878_ (_01634_, _01632_, _25116_);
  or _33879_ (_01635_, _01634_, _01633_);
  not _33880_ (_01636_, _01635_);
  not _33881_ (_01637_, _25128_);
  and _33882_ (_01638_, _01630_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _33883_ (_01639_, _01638_, _27006_);
  nor _33884_ (_01641_, _01639_, _01637_);
  and _33885_ (_01642_, _01639_, _01637_);
  nor _33886_ (_01644_, _01642_, _01641_);
  and _33887_ (_01645_, _26033_, _25053_);
  not _33888_ (_01647_, _01645_);
  nor _33889_ (_01648_, _26033_, _25053_);
  and _33890_ (_01650_, _25073_, _25101_);
  and _33891_ (_01651_, _01650_, _26938_);
  not _33892_ (_01653_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _33893_ (_01654_, _25446_, _01653_);
  not _33894_ (_01656_, _01654_);
  nor _33895_ (_01657_, _01656_, _00755_);
  and _33896_ (_01659_, _01657_, _01651_);
  not _33897_ (_01660_, _01659_);
  and _33898_ (_01662_, _25055_, _25116_);
  and _33899_ (_01663_, _01651_, _01662_);
  not _33900_ (_01665_, _01663_);
  and _33901_ (_01666_, _01650_, _26457_);
  and _33902_ (_01668_, _01666_, _01662_);
  not _33903_ (_01669_, _01668_);
  and _33904_ (_01671_, _01666_, _27035_);
  and _33905_ (_01672_, _01666_, _27224_);
  nor _33906_ (_01673_, _01672_, _01671_);
  and _33907_ (_01674_, _01673_, _01669_);
  not _33908_ (_01675_, _01666_);
  nor _33909_ (_01676_, _01675_, _00755_);
  not _33910_ (_01677_, _01676_);
  and _33911_ (_01678_, _01651_, _27035_);
  and _33912_ (_01679_, _01651_, _27224_);
  nor _33913_ (_01680_, _01679_, _01678_);
  and _33914_ (_01681_, _01680_, _01677_);
  and _33915_ (_01682_, _01681_, _01674_);
  and _33916_ (_01683_, _01682_, _01665_);
  or _33917_ (_01684_, _01683_, _01656_);
  and _33918_ (_01685_, _01684_, _01660_);
  nor _33919_ (_01686_, _01685_, _01648_);
  and _33920_ (_01687_, _01686_, _01647_);
  and _33921_ (_01688_, _01687_, _01644_);
  and _33922_ (_01689_, _01688_, _01636_);
  and _33923_ (_01690_, _01689_, _26543_);
  not _33924_ (_01691_, _01639_);
  and _33925_ (_01692_, _01632_, _26034_);
  and _33926_ (_01693_, _01692_, _01691_);
  and _33927_ (_01694_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _33928_ (_01695_, _01632_, _26033_);
  and _33929_ (_01696_, _01695_, _01639_);
  and _33930_ (_01697_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _33931_ (_01698_, _01697_, _01694_);
  nor _33932_ (_01699_, _01632_, _26034_);
  and _33933_ (_01700_, _01699_, _01691_);
  and _33934_ (_01701_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _33935_ (_01702_, _01632_, _26033_);
  and _33936_ (_01703_, _01702_, _01639_);
  and _33937_ (_01704_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _33938_ (_01705_, _01704_, _01701_);
  and _33939_ (_01706_, _01705_, _01698_);
  not _33940_ (_01707_, _01689_);
  and _33941_ (_01708_, _01702_, _01691_);
  nand _33942_ (_01709_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _33943_ (_01710_, _01692_, _01639_);
  nand _33944_ (_01711_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _33945_ (_01712_, _01711_, _01709_);
  and _33946_ (_01713_, _01695_, _01691_);
  nand _33947_ (_01714_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _33948_ (_01715_, _01699_, _01639_);
  nand _33949_ (_01716_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _33950_ (_01717_, _01716_, _01714_);
  and _33951_ (_01718_, _01717_, _01712_);
  and _33952_ (_01719_, _01718_, _01707_);
  and _33953_ (_01720_, _01719_, _01706_);
  nor _33954_ (_01721_, _01720_, _01690_);
  nand _33955_ (_01722_, _01721_, _01627_);
  and _33956_ (_01723_, _26454_, _26436_);
  not _33957_ (_01724_, _01723_);
  nor _33958_ (_01725_, _01724_, _26389_);
  not _33959_ (_01726_, _25987_);
  and _33960_ (_01727_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  nor _33961_ (_01728_, _25996_, _26190_);
  nor _33962_ (_01729_, _26018_, _26193_);
  nor _33963_ (_01730_, _01729_, _01728_);
  and _33964_ (_01731_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _33965_ (_01732_, _26002_, _26186_);
  nor _33966_ (_01733_, _01732_, _01731_);
  and _33967_ (_01734_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _33968_ (_01735_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _33969_ (_01736_, _26009_, _01735_);
  nor _33970_ (_01737_, _01736_, _01734_);
  and _33971_ (_01738_, _01737_, _01733_);
  and _33972_ (_01739_, _01738_, _01730_);
  and _33973_ (_01740_, _25993_, _25987_);
  not _33974_ (_01741_, _01740_);
  nor _33975_ (_01742_, _01741_, _01739_);
  nor _33976_ (_01743_, _01742_, _01727_);
  not _33977_ (_01744_, _01743_);
  nand _33978_ (_01745_, _01744_, _01725_);
  and _33979_ (_01746_, _01745_, _26454_);
  and _33980_ (_01747_, _01746_, _01722_);
  and _33981_ (_01748_, _01747_, _01626_);
  and _33982_ (_01749_, _26286_, _26266_);
  or _33983_ (_01750_, _01749_, _26337_);
  and _33984_ (_01751_, _26359_, _26273_);
  and _33985_ (_01752_, _26287_, _26269_);
  or _33986_ (_01753_, _01752_, _26300_);
  or _33987_ (_01754_, _01753_, _01751_);
  nor _33988_ (_01755_, _01754_, _01750_);
  nor _33989_ (_01756_, _26318_, _26275_);
  and _33990_ (_01757_, _01756_, _26310_);
  and _33991_ (_01758_, _01757_, _01755_);
  nor _33992_ (_01759_, _01758_, _26393_);
  or _33993_ (_01760_, _26316_, _26313_);
  and _33994_ (_01761_, _26372_, _01760_);
  nor _33995_ (_01762_, _01761_, _01759_);
  not _33996_ (_01763_, _01762_);
  and _33997_ (_01764_, _01763_, _01748_);
  not _33998_ (_01765_, _01764_);
  and _33999_ (_01766_, _01627_, _26454_);
  and _34000_ (_01767_, _01689_, _26497_);
  and _34001_ (_01768_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _34002_ (_01769_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _34003_ (_01770_, _01769_, _01768_);
  and _34004_ (_01771_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _34005_ (_01772_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _34006_ (_01773_, _01772_, _01771_);
  and _34007_ (_01774_, _01773_, _01770_);
  and _34008_ (_01775_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _34009_ (_01776_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _34010_ (_01777_, _01776_, _01775_);
  and _34011_ (_01778_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _34012_ (_01779_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _34013_ (_01780_, _01779_, _01778_);
  and _34014_ (_01781_, _01780_, _01777_);
  and _34015_ (_01782_, _01781_, _01707_);
  and _34016_ (_01783_, _01782_, _01774_);
  nor _34017_ (_01784_, _01783_, _01767_);
  and _34018_ (_01785_, _01784_, _01766_);
  not _34019_ (_01786_, _01785_);
  not _34020_ (_01787_, _01625_);
  or _34021_ (_01788_, _26571_, _01787_);
  not _34022_ (_01789_, _01632_);
  and _34023_ (_01790_, _01723_, _26389_);
  nand _34024_ (_01791_, _01790_, _01789_);
  and _34025_ (_01792_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _34026_ (_01793_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not _34027_ (_01794_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _34028_ (_01795_, _26009_, _01794_);
  nor _34029_ (_01796_, _01795_, _01793_);
  and _34030_ (_01797_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _34031_ (_01798_, _26018_, _26057_);
  nor _34032_ (_01799_, _01798_, _01797_);
  nor _34033_ (_01800_, _25996_, _26051_);
  nor _34034_ (_01801_, _26002_, _26043_);
  nor _34035_ (_01802_, _01801_, _01800_);
  and _34036_ (_01803_, _01802_, _01799_);
  and _34037_ (_01804_, _01803_, _01796_);
  nor _34038_ (_01805_, _01804_, _01741_);
  nor _34039_ (_01806_, _01805_, _01792_);
  not _34040_ (_01807_, _01806_);
  nand _34041_ (_01808_, _01807_, _01725_);
  and _34042_ (_01809_, _01808_, _01791_);
  and _34043_ (_01810_, _01809_, _01788_);
  and _34044_ (_01811_, _01810_, _01786_);
  or _34045_ (_01812_, _01811_, _01765_);
  and _34046_ (_01813_, _01689_, _26521_);
  and _34047_ (_01814_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _34048_ (_01815_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor _34049_ (_01816_, _01815_, _01814_);
  and _34050_ (_01817_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _34051_ (_01818_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _34052_ (_01819_, _01818_, _01817_);
  and _34053_ (_01820_, _01819_, _01816_);
  and _34054_ (_01821_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _34055_ (_01822_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _34056_ (_01823_, _01822_, _01821_);
  and _34057_ (_01824_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _34058_ (_01825_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _34059_ (_01826_, _01825_, _01824_);
  and _34060_ (_01827_, _01826_, _01823_);
  and _34061_ (_01828_, _01827_, _01707_);
  and _34062_ (_01829_, _01828_, _01820_);
  nor _34063_ (_01830_, _01829_, _01813_);
  and _34064_ (_01831_, _01830_, _01766_);
  not _34065_ (_01832_, _01831_);
  and _34066_ (_01833_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  nor _34067_ (_01834_, _25996_, _26008_);
  nor _34068_ (_01835_, _26018_, _25994_);
  nor _34069_ (_01836_, _01835_, _01834_);
  and _34070_ (_01837_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _34071_ (_01838_, _26002_, _26015_);
  nor _34072_ (_01839_, _01838_, _01837_);
  and _34073_ (_01840_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not _34074_ (_01841_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _34075_ (_01842_, _26009_, _01841_);
  nor _34076_ (_01843_, _01842_, _01840_);
  and _34077_ (_01844_, _01843_, _01839_);
  and _34078_ (_01845_, _01844_, _01836_);
  nor _34079_ (_01846_, _01845_, _01741_);
  nor _34080_ (_01847_, _01846_, _01833_);
  not _34081_ (_01848_, _01847_);
  and _34082_ (_01849_, _01848_, _01725_);
  or _34083_ (_01850_, _26553_, _01787_);
  nand _34084_ (_01851_, _01790_, _26033_);
  nand _34085_ (_01852_, _01851_, _01850_);
  nor _34086_ (_01853_, _01852_, _01849_);
  and _34087_ (_01854_, _01853_, _01832_);
  or _34088_ (_01855_, _01854_, _01763_);
  nand _34089_ (_01856_, _01855_, _01812_);
  and _34090_ (_01857_, _01856_, _01623_);
  nor _34091_ (_01858_, _01856_, _01623_);
  nor _34092_ (_01859_, _01858_, _01857_);
  and _34093_ (_01860_, _01620_, _01637_);
  nor _34094_ (_01861_, _25042_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _34095_ (_01862_, _01861_, _01860_);
  and _34096_ (_01863_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _34097_ (_01864_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _34098_ (_01865_, _01864_, _01863_);
  and _34099_ (_01866_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _34100_ (_01867_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _34101_ (_01868_, _01867_, _01866_);
  and _34102_ (_01869_, _01868_, _01865_);
  and _34103_ (_01870_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _34104_ (_01871_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _34105_ (_01872_, _01871_, _01870_);
  and _34106_ (_01873_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _34107_ (_01874_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _34108_ (_01875_, _01874_, _01873_);
  and _34109_ (_01876_, _01875_, _01872_);
  and _34110_ (_01877_, _01876_, _01707_);
  and _34111_ (_01878_, _01877_, _01869_);
  and _34112_ (_01879_, _01689_, _26489_);
  nor _34113_ (_01880_, _01879_, _01878_);
  and _34114_ (_01881_, _01880_, _01766_);
  not _34115_ (_01882_, _01881_);
  not _34116_ (_01883_, _26454_);
  and _34117_ (_01884_, _01883_, _26436_);
  nor _34118_ (_01885_, _26577_, _01787_);
  nor _34119_ (_01886_, _01885_, _01884_);
  and _34120_ (_01887_, _01790_, _01691_);
  and _34121_ (_01888_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  nor _34122_ (_01889_, _25996_, _26157_);
  nor _34123_ (_01890_, _26018_, _26159_);
  nor _34124_ (_01891_, _01890_, _01889_);
  not _34125_ (_01892_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _34126_ (_01893_, _26009_, _01892_);
  nor _34127_ (_01894_, _26002_, _26167_);
  nor _34128_ (_01895_, _01894_, _01893_);
  and _34129_ (_01896_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _34130_ (_01897_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _34131_ (_01898_, _01897_, _01896_);
  and _34132_ (_01899_, _01898_, _01895_);
  and _34133_ (_01900_, _01899_, _01891_);
  nor _34134_ (_01901_, _01900_, _01741_);
  nor _34135_ (_01902_, _01901_, _01888_);
  not _34136_ (_01903_, _01902_);
  and _34137_ (_01904_, _01903_, _01725_);
  nor _34138_ (_01905_, _01904_, _01887_);
  and _34139_ (_01906_, _01905_, _01886_);
  and _34140_ (_01907_, _01906_, _01882_);
  or _34141_ (_01908_, _01907_, _01765_);
  and _34142_ (_01909_, _01689_, _26512_);
  and _34143_ (_01910_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _34144_ (_01911_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _34145_ (_01912_, _01911_, _01910_);
  and _34146_ (_01913_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _34147_ (_01914_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _34148_ (_01915_, _01914_, _01913_);
  and _34149_ (_01916_, _01915_, _01912_);
  and _34150_ (_01917_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _34151_ (_01918_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _34152_ (_01919_, _01918_, _01917_);
  and _34153_ (_01920_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _34154_ (_01921_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _34155_ (_01922_, _01921_, _01920_);
  and _34156_ (_01923_, _01922_, _01919_);
  and _34157_ (_01924_, _01923_, _01707_);
  and _34158_ (_01925_, _01924_, _01916_);
  nor _34159_ (_01926_, _01925_, _01909_);
  and _34160_ (_01927_, _01926_, _01766_);
  not _34161_ (_01928_, _01927_);
  and _34162_ (_01929_, _01627_, _01883_);
  nor _34163_ (_01930_, _26559_, _01787_);
  nor _34164_ (_01931_, _01930_, _01929_);
  and _34165_ (_01932_, _01790_, _26153_);
  and _34166_ (_01933_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _34167_ (_01934_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not _34168_ (_01935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _34169_ (_01936_, _26009_, _01935_);
  nor _34170_ (_01937_, _01936_, _01934_);
  nor _34171_ (_01938_, _25996_, _26127_);
  nor _34172_ (_01939_, _26002_, _26132_);
  nor _34173_ (_01940_, _01939_, _01938_);
  and _34174_ (_01941_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _34175_ (_01942_, _26018_, _26129_);
  nor _34176_ (_01943_, _01942_, _01941_);
  and _34177_ (_01944_, _01943_, _01940_);
  and _34178_ (_01945_, _01944_, _01937_);
  nor _34179_ (_01946_, _01945_, _01741_);
  nor _34180_ (_01947_, _01946_, _01933_);
  not _34181_ (_01948_, _01947_);
  and _34182_ (_01949_, _01948_, _01725_);
  nor _34183_ (_01950_, _01949_, _01932_);
  and _34184_ (_01951_, _01950_, _01931_);
  and _34185_ (_01952_, _01951_, _01928_);
  or _34186_ (_01953_, _01952_, _01763_);
  and _34187_ (_01954_, _01953_, _01908_);
  and _34188_ (_01955_, _01954_, _01862_);
  nor _34189_ (_01956_, _01954_, _01862_);
  or _34190_ (_01957_, _01956_, _01955_);
  and _34191_ (_01958_, _01957_, _01859_);
  nor _34192_ (_01959_, _01620_, _26922_);
  not _34193_ (_01960_, _01959_);
  and _34194_ (_01961_, _01884_, _26389_);
  nor _34195_ (_01962_, _26583_, _01787_);
  nor _34196_ (_01963_, _01962_, _01961_);
  and _34197_ (_01964_, _01624_, _01883_);
  not _34198_ (_01965_, _01964_);
  and _34199_ (_01966_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  nor _34200_ (_01967_, _25996_, _26218_);
  nor _34201_ (_01968_, _26018_, _26212_);
  nor _34202_ (_01969_, _01968_, _01967_);
  and _34203_ (_01970_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not _34204_ (_01971_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _34205_ (_01972_, _26009_, _01971_);
  nor _34206_ (_01973_, _01972_, _01970_);
  and _34207_ (_01974_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _34208_ (_01975_, _26002_, _26222_);
  nor _34209_ (_01976_, _01975_, _01974_);
  and _34210_ (_01977_, _01976_, _01973_);
  and _34211_ (_01978_, _01977_, _01969_);
  nor _34212_ (_01979_, _01978_, _01741_);
  nor _34213_ (_01980_, _01979_, _01966_);
  not _34214_ (_01981_, _01980_);
  and _34215_ (_01982_, _01981_, _01725_);
  and _34216_ (_01983_, _01689_, _26482_);
  and _34217_ (_01984_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _34218_ (_01985_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _34219_ (_01986_, _01985_, _01984_);
  and _34220_ (_01987_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _34221_ (_01988_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _34222_ (_01989_, _01988_, _01987_);
  and _34223_ (_01990_, _01989_, _01986_);
  and _34224_ (_01991_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _34225_ (_01992_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _34226_ (_01993_, _01992_, _01991_);
  and _34227_ (_01994_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _34228_ (_01995_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _34229_ (_01996_, _01995_, _01994_);
  and _34230_ (_01997_, _01996_, _01993_);
  and _34231_ (_01998_, _01997_, _01707_);
  and _34232_ (_01999_, _01998_, _01990_);
  nor _34233_ (_02000_, _01999_, _01983_);
  and _34234_ (_02001_, _02000_, _01766_);
  nor _34235_ (_02002_, _02001_, _01982_);
  and _34236_ (_02003_, _02002_, _01965_);
  and _34237_ (_02004_, _02003_, _01963_);
  and _34238_ (_02005_, _02004_, _01765_);
  nor _34239_ (_02006_, _02005_, _01960_);
  not _34240_ (_02007_, _02006_);
  nor _34241_ (_02008_, _01620_, _25073_);
  not _34242_ (_02009_, _02008_);
  nor _34243_ (_02010_, _26589_, _01787_);
  not _34244_ (_02011_, _02010_);
  and _34245_ (_02012_, _01689_, _26475_);
  and _34246_ (_02013_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _34247_ (_02014_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _34248_ (_02015_, _02014_, _02013_);
  and _34249_ (_02016_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _34250_ (_02017_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _34251_ (_02018_, _02017_, _02016_);
  and _34252_ (_02019_, _02018_, _02015_);
  and _34253_ (_02020_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _34254_ (_02021_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _34255_ (_02022_, _02021_, _02020_);
  and _34256_ (_02023_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _34257_ (_02024_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor _34258_ (_02025_, _02024_, _02023_);
  and _34259_ (_02026_, _02025_, _02022_);
  and _34260_ (_02027_, _02026_, _01707_);
  and _34261_ (_02028_, _02027_, _02019_);
  nor _34262_ (_02029_, _02028_, _02012_);
  and _34263_ (_02030_, _02029_, _01766_);
  not _34264_ (_02031_, _02030_);
  and _34265_ (_02032_, _26436_, _26390_);
  and _34266_ (_02033_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _34267_ (_02034_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not _34268_ (_02035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _34269_ (_02036_, _26009_, _02035_);
  nor _34270_ (_02037_, _02036_, _02034_);
  nor _34271_ (_02038_, _25996_, _26251_);
  nor _34272_ (_02039_, _26002_, _26247_);
  nor _34273_ (_02040_, _02039_, _02038_);
  and _34274_ (_02041_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _34275_ (_02042_, _26018_, _26245_);
  nor _34276_ (_02043_, _02042_, _02041_);
  and _34277_ (_02044_, _02043_, _02040_);
  and _34278_ (_02045_, _02044_, _02037_);
  nor _34279_ (_02046_, _02045_, _01741_);
  nor _34280_ (_02047_, _02046_, _02033_);
  not _34281_ (_02048_, _02047_);
  and _34282_ (_02049_, _02048_, _02032_);
  nor _34283_ (_02050_, _01627_, _26454_);
  nor _34284_ (_02051_, _02050_, _02049_);
  and _34285_ (_02052_, _02051_, _02031_);
  and _34286_ (_02053_, _02052_, _02011_);
  nor _34287_ (_02054_, _02053_, _01764_);
  nor _34288_ (_02055_, _02054_, _02009_);
  and _34289_ (_02056_, _02054_, _02009_);
  nor _34290_ (_02057_, _02056_, _02055_);
  and _34291_ (_02058_, _02057_, _02007_);
  nor _34292_ (_02059_, _01748_, _25101_);
  and _34293_ (_02060_, _01748_, _25101_);
  nor _34294_ (_02061_, _02060_, _02059_);
  not _34295_ (_02062_, _02061_);
  nor _34296_ (_02063_, _01620_, _25128_);
  not _34297_ (_02064_, _02063_);
  nor _34298_ (_02065_, _01907_, _01764_);
  and _34299_ (_02066_, _02065_, _02064_);
  and _34300_ (_02067_, _02005_, _01960_);
  nor _34301_ (_02068_, _02067_, _02066_);
  and _34302_ (_02069_, _02068_, _02062_);
  and _34303_ (_02070_, _02069_, _02058_);
  and _34304_ (_02071_, _02070_, _01958_);
  and _34305_ (_02072_, _01620_, _26458_);
  nor _34306_ (_02073_, _01620_, _25115_);
  nor _34307_ (_02074_, _02073_, _02072_);
  and _34308_ (_02075_, _02053_, _01764_);
  and _34309_ (_02076_, _01811_, _01765_);
  nor _34310_ (_02077_, _02076_, _02075_);
  and _34311_ (_02078_, _02077_, _02074_);
  nor _34312_ (_02079_, _02077_, _02074_);
  or _34313_ (_02080_, _02079_, _02078_);
  not _34314_ (_02081_, _02080_);
  and _34315_ (_02082_, _01620_, _26922_);
  nor _34316_ (_02083_, _25020_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _34317_ (_02084_, _02083_, _02082_);
  not _34318_ (_02085_, _02084_);
  nor _34319_ (_02086_, _02004_, _01765_);
  and _34320_ (_02087_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _34321_ (_02088_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _34322_ (_02089_, _02088_, _02087_);
  and _34323_ (_02090_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _34324_ (_02091_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _34325_ (_02092_, _02091_, _02090_);
  and _34326_ (_02093_, _02092_, _02089_);
  and _34327_ (_02094_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _34328_ (_02095_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _34329_ (_02096_, _02095_, _02094_);
  and _34330_ (_02097_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _34331_ (_02098_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _34332_ (_02099_, _02098_, _02097_);
  and _34333_ (_02100_, _02099_, _02096_);
  and _34334_ (_02101_, _02100_, _01707_);
  and _34335_ (_02102_, _02101_, _02093_);
  and _34336_ (_02103_, _01689_, _26505_);
  nor _34337_ (_02104_, _02103_, _02102_);
  and _34338_ (_02105_, _02104_, _01766_);
  not _34339_ (_02106_, _02105_);
  and _34340_ (_02107_, _01790_, _26125_);
  not _34341_ (_02108_, _26565_);
  and _34342_ (_02109_, _02108_, _01625_);
  and _34343_ (_02110_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _34344_ (_02111_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not _34345_ (_02112_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _34346_ (_02113_, _26009_, _02112_);
  nor _34347_ (_02114_, _02113_, _02111_);
  nor _34348_ (_02115_, _26018_, _26111_);
  nor _34349_ (_02116_, _26002_, _26097_);
  nor _34350_ (_02117_, _02116_, _02115_);
  and _34351_ (_02118_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _34352_ (_02119_, _25996_, _26105_);
  nor _34353_ (_02120_, _02119_, _02118_);
  and _34354_ (_02121_, _02120_, _02117_);
  and _34355_ (_02122_, _02121_, _02114_);
  nor _34356_ (_02123_, _02122_, _01741_);
  nor _34357_ (_02124_, _02123_, _02110_);
  not _34358_ (_02125_, _02124_);
  and _34359_ (_02126_, _02125_, _01725_);
  or _34360_ (_02127_, _02126_, _02109_);
  nor _34361_ (_02128_, _02127_, _02107_);
  and _34362_ (_02129_, _02128_, _02106_);
  nor _34363_ (_02130_, _02129_, _01763_);
  nor _34364_ (_02131_, _02130_, _02086_);
  nor _34365_ (_02132_, _02131_, _02085_);
  and _34366_ (_02133_, _02131_, _02085_);
  nor _34367_ (_02134_, _02133_, _02132_);
  and _34368_ (_02135_, _02134_, _02081_);
  nor _34369_ (_02136_, _02065_, _02064_);
  and _34370_ (_02137_, _25446_, _25099_);
  not _34371_ (_02138_, _02137_);
  nor _34372_ (_02139_, _02138_, _02136_);
  and _34373_ (_02140_, _02139_, _02135_);
  and _34374_ (_02141_, _02140_, _02071_);
  not _34375_ (_02142_, _01748_);
  not _34376_ (_02143_, _02005_);
  not _34377_ (_02144_, _02131_);
  and _34378_ (_02145_, _01855_, _01812_);
  and _34379_ (_02146_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _34380_ (_02147_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _34381_ (_02148_, _02147_, _02146_);
  and _34382_ (_02149_, _02148_, _01954_);
  not _34383_ (_02150_, _01954_);
  and _34384_ (_02151_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _34385_ (_02152_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _34386_ (_02153_, _02152_, _02151_);
  and _34387_ (_02154_, _02153_, _02150_);
  or _34388_ (_02155_, _02154_, _02149_);
  or _34389_ (_02156_, _02155_, _02144_);
  not _34390_ (_02157_, _02077_);
  and _34391_ (_02158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and _34392_ (_02159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _34393_ (_02160_, _02159_, _02158_);
  and _34394_ (_02161_, _02160_, _01954_);
  and _34395_ (_02162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _34396_ (_02163_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _34397_ (_02164_, _02163_, _02162_);
  and _34398_ (_02165_, _02164_, _02150_);
  or _34399_ (_02166_, _02165_, _02161_);
  or _34400_ (_02167_, _02166_, _02131_);
  and _34401_ (_02168_, _02167_, _02157_);
  and _34402_ (_02169_, _02168_, _02156_);
  or _34403_ (_02170_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _34404_ (_02171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _34405_ (_02172_, _02171_, _02170_);
  and _34406_ (_02173_, _02172_, _01954_);
  or _34407_ (_02174_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _34408_ (_02175_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _34409_ (_02176_, _02175_, _02174_);
  and _34410_ (_02177_, _02176_, _02150_);
  or _34411_ (_02178_, _02177_, _02173_);
  or _34412_ (_02179_, _02178_, _02144_);
  or _34413_ (_02180_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _34414_ (_02181_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _34415_ (_02182_, _02181_, _02180_);
  and _34416_ (_02183_, _02182_, _01954_);
  or _34417_ (_02184_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _34418_ (_02185_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and _34419_ (_02186_, _02185_, _02184_);
  and _34420_ (_02187_, _02186_, _02150_);
  or _34421_ (_02188_, _02187_, _02183_);
  or _34422_ (_02189_, _02188_, _02131_);
  and _34423_ (_02190_, _02189_, _02077_);
  and _34424_ (_02191_, _02190_, _02179_);
  or _34425_ (_02192_, _02191_, _02169_);
  and _34426_ (_02193_, _02192_, _02065_);
  not _34427_ (_02194_, _02065_);
  and _34428_ (_02195_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _34429_ (_02196_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _34430_ (_02197_, _02196_, _02195_);
  and _34431_ (_02198_, _02197_, _01954_);
  and _34432_ (_02199_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _34433_ (_02200_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _34434_ (_02201_, _02200_, _02199_);
  and _34435_ (_02202_, _02201_, _02150_);
  or _34436_ (_02204_, _02202_, _02198_);
  or _34437_ (_02206_, _02204_, _02144_);
  and _34438_ (_02208_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _34439_ (_02210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _34440_ (_02212_, _02210_, _02208_);
  and _34441_ (_02214_, _02212_, _01954_);
  and _34442_ (_02216_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _34443_ (_02218_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _34444_ (_02220_, _02218_, _02216_);
  and _34445_ (_02222_, _02220_, _02150_);
  or _34446_ (_02224_, _02222_, _02214_);
  or _34447_ (_02226_, _02224_, _02131_);
  and _34448_ (_02228_, _02226_, _02157_);
  and _34449_ (_02230_, _02228_, _02206_);
  or _34450_ (_02232_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _34451_ (_02234_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _34452_ (_02236_, _02234_, _02150_);
  and _34453_ (_02238_, _02236_, _02232_);
  or _34454_ (_02240_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _34455_ (_02242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _34456_ (_02244_, _02242_, _01954_);
  and _34457_ (_02246_, _02244_, _02240_);
  or _34458_ (_02248_, _02246_, _02238_);
  or _34459_ (_02250_, _02248_, _02144_);
  or _34460_ (_02252_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _34461_ (_02254_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and _34462_ (_02256_, _02254_, _02150_);
  and _34463_ (_02258_, _02256_, _02252_);
  or _34464_ (_02260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _34465_ (_02262_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and _34466_ (_02264_, _02262_, _01954_);
  and _34467_ (_02266_, _02264_, _02260_);
  or _34468_ (_02268_, _02266_, _02258_);
  or _34469_ (_02270_, _02268_, _02131_);
  and _34470_ (_02272_, _02270_, _02077_);
  and _34471_ (_02273_, _02272_, _02250_);
  or _34472_ (_02274_, _02273_, _02230_);
  and _34473_ (_02275_, _02274_, _02194_);
  or _34474_ (_02276_, _02275_, _02193_);
  and _34475_ (_02277_, _02276_, _02143_);
  and _34476_ (_02278_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _34477_ (_02279_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _34478_ (_02280_, _02279_, _02278_);
  and _34479_ (_02281_, _02280_, _01954_);
  and _34480_ (_02282_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _34481_ (_02283_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _34482_ (_02284_, _02283_, _02282_);
  and _34483_ (_02285_, _02284_, _02150_);
  or _34484_ (_02286_, _02285_, _02281_);
  and _34485_ (_02287_, _02286_, _02131_);
  and _34486_ (_02288_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _34487_ (_02289_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _34488_ (_02290_, _02289_, _02288_);
  and _34489_ (_02291_, _02290_, _01954_);
  and _34490_ (_02292_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and _34491_ (_02293_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _34492_ (_02294_, _02293_, _02292_);
  and _34493_ (_02295_, _02294_, _02150_);
  or _34494_ (_02296_, _02295_, _02291_);
  and _34495_ (_02297_, _02296_, _02144_);
  or _34496_ (_02298_, _02297_, _02287_);
  and _34497_ (_02299_, _02298_, _02157_);
  or _34498_ (_02300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _34499_ (_02301_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _34500_ (_02302_, _02301_, _02150_);
  and _34501_ (_02303_, _02302_, _02300_);
  or _34502_ (_02304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _34503_ (_02305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _34504_ (_02306_, _02305_, _01954_);
  and _34505_ (_02307_, _02306_, _02304_);
  or _34506_ (_02308_, _02307_, _02303_);
  and _34507_ (_02309_, _02308_, _02131_);
  or _34508_ (_02310_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _34509_ (_02311_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _34510_ (_02312_, _02311_, _02150_);
  and _34511_ (_02313_, _02312_, _02310_);
  or _34512_ (_02314_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _34513_ (_02315_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _34514_ (_02316_, _02315_, _01954_);
  and _34515_ (_02317_, _02316_, _02314_);
  or _34516_ (_02318_, _02317_, _02313_);
  and _34517_ (_02319_, _02318_, _02144_);
  or _34518_ (_02320_, _02319_, _02309_);
  and _34519_ (_02321_, _02320_, _02077_);
  or _34520_ (_02322_, _02321_, _02299_);
  and _34521_ (_02323_, _02322_, _02194_);
  and _34522_ (_02324_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _34523_ (_02325_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _34524_ (_02326_, _02325_, _02324_);
  and _34525_ (_02327_, _02326_, _01954_);
  and _34526_ (_02328_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _34527_ (_02329_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _34528_ (_02330_, _02329_, _02328_);
  and _34529_ (_02331_, _02330_, _02150_);
  or _34530_ (_02332_, _02331_, _02327_);
  and _34531_ (_02333_, _02332_, _02131_);
  and _34532_ (_02334_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and _34533_ (_02335_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _34534_ (_02336_, _02335_, _02334_);
  and _34535_ (_02337_, _02336_, _01954_);
  and _34536_ (_02338_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _34537_ (_02339_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _34538_ (_02340_, _02339_, _02338_);
  and _34539_ (_02341_, _02340_, _02150_);
  or _34540_ (_02342_, _02341_, _02337_);
  and _34541_ (_02343_, _02342_, _02144_);
  or _34542_ (_02344_, _02343_, _02333_);
  and _34543_ (_02345_, _02344_, _02157_);
  or _34544_ (_02346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _34545_ (_02347_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _34546_ (_02348_, _02347_, _02346_);
  and _34547_ (_02349_, _02348_, _01954_);
  or _34548_ (_02350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _34549_ (_02351_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _34550_ (_02352_, _02351_, _02350_);
  and _34551_ (_02353_, _02352_, _02150_);
  or _34552_ (_02354_, _02353_, _02349_);
  and _34553_ (_02355_, _02354_, _02131_);
  or _34554_ (_02356_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _34555_ (_02357_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _34556_ (_02358_, _02357_, _02356_);
  and _34557_ (_02359_, _02358_, _01954_);
  or _34558_ (_02360_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _34559_ (_02361_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _34560_ (_02362_, _02361_, _02360_);
  and _34561_ (_02363_, _02362_, _02150_);
  or _34562_ (_02364_, _02363_, _02359_);
  and _34563_ (_02365_, _02364_, _02144_);
  or _34564_ (_02366_, _02365_, _02355_);
  and _34565_ (_02367_, _02366_, _02077_);
  or _34566_ (_02368_, _02367_, _02345_);
  and _34567_ (_02369_, _02368_, _02065_);
  or _34568_ (_02370_, _02369_, _02323_);
  and _34569_ (_02371_, _02370_, _02005_);
  or _34570_ (_02372_, _02371_, _02277_);
  or _34571_ (_02373_, _02372_, _02054_);
  not _34572_ (_02374_, _02054_);
  and _34573_ (_02375_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and _34574_ (_02376_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _34575_ (_02377_, _02376_, _02375_);
  and _34576_ (_02378_, _02377_, _01954_);
  and _34577_ (_02379_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _34578_ (_02380_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _34579_ (_02381_, _02380_, _02379_);
  and _34580_ (_02382_, _02381_, _02150_);
  or _34581_ (_02383_, _02382_, _02378_);
  or _34582_ (_02384_, _02383_, _02144_);
  and _34583_ (_02385_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and _34584_ (_02386_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _34585_ (_02387_, _02386_, _02385_);
  and _34586_ (_02388_, _02387_, _01954_);
  and _34587_ (_02389_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _34588_ (_02390_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _34589_ (_02391_, _02390_, _02389_);
  and _34590_ (_02392_, _02391_, _02150_);
  or _34591_ (_02393_, _02392_, _02388_);
  or _34592_ (_02394_, _02393_, _02131_);
  and _34593_ (_02395_, _02394_, _02157_);
  and _34594_ (_02396_, _02395_, _02384_);
  or _34595_ (_02397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _34596_ (_02398_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _34597_ (_02399_, _02398_, _02150_);
  and _34598_ (_02400_, _02399_, _02397_);
  or _34599_ (_02401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _34600_ (_02402_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and _34601_ (_02403_, _02402_, _01954_);
  and _34602_ (_02404_, _02403_, _02401_);
  or _34603_ (_02405_, _02404_, _02400_);
  or _34604_ (_02406_, _02405_, _02144_);
  or _34605_ (_02407_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _34606_ (_02408_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _34607_ (_02409_, _02408_, _02150_);
  and _34608_ (_02410_, _02409_, _02407_);
  or _34609_ (_02411_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _34610_ (_02412_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and _34611_ (_02413_, _02412_, _01954_);
  and _34612_ (_02414_, _02413_, _02411_);
  or _34613_ (_02415_, _02414_, _02410_);
  or _34614_ (_02416_, _02415_, _02131_);
  and _34615_ (_02417_, _02416_, _02077_);
  and _34616_ (_02418_, _02417_, _02406_);
  or _34617_ (_02419_, _02418_, _02396_);
  and _34618_ (_02420_, _02419_, _02194_);
  and _34619_ (_02421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _34620_ (_02422_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _34621_ (_02423_, _02422_, _02421_);
  and _34622_ (_02424_, _02423_, _01954_);
  and _34623_ (_02425_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _34624_ (_02426_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _34625_ (_02427_, _02426_, _02425_);
  and _34626_ (_02428_, _02427_, _02150_);
  or _34627_ (_02429_, _02428_, _02424_);
  or _34628_ (_02430_, _02429_, _02144_);
  and _34629_ (_02431_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _34630_ (_02432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _34631_ (_02433_, _02432_, _02431_);
  and _34632_ (_02434_, _02433_, _01954_);
  and _34633_ (_02435_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _34634_ (_02436_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _34635_ (_02437_, _02436_, _02435_);
  and _34636_ (_02438_, _02437_, _02150_);
  or _34637_ (_02439_, _02438_, _02434_);
  or _34638_ (_02440_, _02439_, _02131_);
  and _34639_ (_02441_, _02440_, _02157_);
  and _34640_ (_02442_, _02441_, _02430_);
  or _34641_ (_02443_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _34642_ (_02444_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _34643_ (_02445_, _02444_, _02443_);
  and _34644_ (_02446_, _02445_, _01954_);
  or _34645_ (_02447_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _34646_ (_02448_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _34647_ (_02449_, _02448_, _02447_);
  and _34648_ (_02450_, _02449_, _02150_);
  or _34649_ (_02451_, _02450_, _02446_);
  or _34650_ (_02452_, _02451_, _02144_);
  or _34651_ (_02453_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _34652_ (_02454_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _34653_ (_02455_, _02454_, _02453_);
  and _34654_ (_02456_, _02455_, _01954_);
  or _34655_ (_02457_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _34656_ (_02458_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _34657_ (_02459_, _02458_, _02457_);
  and _34658_ (_02460_, _02459_, _02150_);
  or _34659_ (_02461_, _02460_, _02456_);
  or _34660_ (_02462_, _02461_, _02131_);
  and _34661_ (_02463_, _02462_, _02077_);
  and _34662_ (_02464_, _02463_, _02452_);
  or _34663_ (_02465_, _02464_, _02442_);
  and _34664_ (_02466_, _02465_, _02065_);
  or _34665_ (_02467_, _02466_, _02420_);
  and _34666_ (_02468_, _02467_, _02143_);
  or _34667_ (_02469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _34668_ (_02470_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _34669_ (_02471_, _02470_, _02469_);
  and _34670_ (_02472_, _02471_, _01954_);
  or _34671_ (_02473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _34672_ (_02474_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and _34673_ (_02475_, _02474_, _02473_);
  and _34674_ (_02476_, _02475_, _02150_);
  or _34675_ (_02477_, _02476_, _02472_);
  and _34676_ (_02478_, _02477_, _02144_);
  or _34677_ (_02479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _34678_ (_02480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _34679_ (_02481_, _02480_, _02479_);
  and _34680_ (_02482_, _02481_, _01954_);
  or _34681_ (_02483_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _34682_ (_02484_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _34683_ (_02485_, _02484_, _02483_);
  and _34684_ (_02486_, _02485_, _02150_);
  or _34685_ (_02487_, _02486_, _02482_);
  and _34686_ (_02488_, _02487_, _02131_);
  or _34687_ (_02489_, _02488_, _02478_);
  and _34688_ (_02490_, _02489_, _02077_);
  and _34689_ (_02491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _34690_ (_02492_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _34691_ (_02493_, _02492_, _02491_);
  and _34692_ (_02494_, _02493_, _01954_);
  and _34693_ (_02495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _34694_ (_02496_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _34695_ (_02497_, _02496_, _02495_);
  and _34696_ (_02498_, _02497_, _02150_);
  or _34697_ (_02499_, _02498_, _02494_);
  and _34698_ (_02500_, _02499_, _02144_);
  and _34699_ (_02501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and _34700_ (_02502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _34701_ (_02503_, _02502_, _02501_);
  and _34702_ (_02504_, _02503_, _01954_);
  and _34703_ (_02505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and _34704_ (_02506_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _34705_ (_02507_, _02506_, _02505_);
  and _34706_ (_02508_, _02507_, _02150_);
  or _34707_ (_02509_, _02508_, _02504_);
  and _34708_ (_02510_, _02509_, _02131_);
  or _34709_ (_02511_, _02510_, _02500_);
  and _34710_ (_02512_, _02511_, _02157_);
  or _34711_ (_02513_, _02512_, _02490_);
  and _34712_ (_02514_, _02513_, _02065_);
  or _34713_ (_02515_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _34714_ (_02516_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _34715_ (_02517_, _02516_, _02150_);
  and _34716_ (_02518_, _02517_, _02515_);
  or _34717_ (_02519_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _34718_ (_02520_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _34719_ (_02521_, _02520_, _01954_);
  and _34720_ (_02522_, _02521_, _02519_);
  or _34721_ (_02523_, _02522_, _02518_);
  and _34722_ (_02524_, _02523_, _02144_);
  or _34723_ (_02525_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _34724_ (_02526_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and _34725_ (_02527_, _02526_, _02150_);
  and _34726_ (_02528_, _02527_, _02525_);
  or _34727_ (_02529_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _34728_ (_02530_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _34729_ (_02531_, _02530_, _01954_);
  and _34730_ (_02532_, _02531_, _02529_);
  or _34731_ (_02533_, _02532_, _02528_);
  and _34732_ (_02534_, _02533_, _02131_);
  or _34733_ (_02535_, _02534_, _02524_);
  and _34734_ (_02536_, _02535_, _02077_);
  and _34735_ (_02537_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and _34736_ (_02538_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _34737_ (_02539_, _02538_, _02537_);
  and _34738_ (_02540_, _02539_, _01954_);
  and _34739_ (_02541_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _34740_ (_02542_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _34741_ (_02543_, _02542_, _02541_);
  and _34742_ (_02544_, _02543_, _02150_);
  or _34743_ (_02545_, _02544_, _02540_);
  and _34744_ (_02546_, _02545_, _02144_);
  and _34745_ (_02547_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _34746_ (_02548_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _34747_ (_02549_, _02548_, _02547_);
  and _34748_ (_02550_, _02549_, _01954_);
  and _34749_ (_02551_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _34750_ (_02552_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _34751_ (_02553_, _02552_, _02551_);
  and _34752_ (_02554_, _02553_, _02150_);
  or _34753_ (_02555_, _02554_, _02550_);
  and _34754_ (_02556_, _02555_, _02131_);
  or _34755_ (_02557_, _02556_, _02546_);
  and _34756_ (_02558_, _02557_, _02157_);
  or _34757_ (_02559_, _02558_, _02536_);
  and _34758_ (_02560_, _02559_, _02194_);
  or _34759_ (_02561_, _02560_, _02514_);
  and _34760_ (_02562_, _02561_, _02005_);
  or _34761_ (_02563_, _02562_, _02468_);
  or _34762_ (_02564_, _02563_, _02374_);
  and _34763_ (_02565_, _02564_, _02373_);
  or _34764_ (_02566_, _02565_, _02142_);
  and _34765_ (_02567_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _34766_ (_02568_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _34767_ (_02569_, _02568_, _02567_);
  and _34768_ (_02570_, _02569_, _01954_);
  and _34769_ (_02571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _34770_ (_02572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _34771_ (_02573_, _02572_, _02571_);
  and _34772_ (_02574_, _02573_, _02150_);
  or _34773_ (_02575_, _02574_, _02570_);
  and _34774_ (_02576_, _02575_, _02131_);
  and _34775_ (_02577_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _34776_ (_02578_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _34777_ (_02579_, _02578_, _02577_);
  and _34778_ (_02580_, _02579_, _01954_);
  and _34779_ (_02581_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _34780_ (_02582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _34781_ (_02583_, _02582_, _02581_);
  and _34782_ (_02584_, _02583_, _02150_);
  or _34783_ (_02585_, _02584_, _02580_);
  and _34784_ (_02586_, _02585_, _02144_);
  or _34785_ (_02587_, _02586_, _02576_);
  and _34786_ (_02588_, _02587_, _02157_);
  or _34787_ (_02589_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _34788_ (_02590_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _34789_ (_02591_, _02590_, _02150_);
  and _34790_ (_02592_, _02591_, _02589_);
  or _34791_ (_02593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _34792_ (_02594_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _34793_ (_02595_, _02594_, _01954_);
  and _34794_ (_02596_, _02595_, _02593_);
  or _34795_ (_02597_, _02596_, _02592_);
  and _34796_ (_02598_, _02597_, _02131_);
  or _34797_ (_02599_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _34798_ (_02600_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _34799_ (_02601_, _02600_, _02150_);
  and _34800_ (_02602_, _02601_, _02599_);
  or _34801_ (_02603_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _34802_ (_02604_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _34803_ (_02605_, _02604_, _01954_);
  and _34804_ (_02606_, _02605_, _02603_);
  or _34805_ (_02607_, _02606_, _02602_);
  and _34806_ (_02608_, _02607_, _02144_);
  or _34807_ (_02609_, _02608_, _02598_);
  and _34808_ (_02610_, _02609_, _02077_);
  or _34809_ (_02611_, _02610_, _02588_);
  and _34810_ (_02612_, _02611_, _02194_);
  and _34811_ (_02613_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _34812_ (_02614_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _34813_ (_02615_, _02614_, _02613_);
  and _34814_ (_02616_, _02615_, _01954_);
  and _34815_ (_02617_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _34816_ (_02618_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _34817_ (_02619_, _02618_, _02617_);
  and _34818_ (_02620_, _02619_, _02150_);
  or _34819_ (_02621_, _02620_, _02616_);
  and _34820_ (_02622_, _02621_, _02131_);
  and _34821_ (_02623_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _34822_ (_02624_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _34823_ (_02625_, _02624_, _02623_);
  and _34824_ (_02626_, _02625_, _01954_);
  and _34825_ (_02627_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _34826_ (_02628_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _34827_ (_02629_, _02628_, _02627_);
  and _34828_ (_02630_, _02629_, _02150_);
  or _34829_ (_02631_, _02630_, _02626_);
  and _34830_ (_02632_, _02631_, _02144_);
  or _34831_ (_02633_, _02632_, _02622_);
  and _34832_ (_02634_, _02633_, _02157_);
  or _34833_ (_02635_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _34834_ (_02636_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _34835_ (_02637_, _02636_, _02635_);
  and _34836_ (_02638_, _02637_, _01954_);
  or _34837_ (_02639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _34838_ (_02640_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _34839_ (_02641_, _02640_, _02639_);
  and _34840_ (_02642_, _02641_, _02150_);
  or _34841_ (_02643_, _02642_, _02638_);
  and _34842_ (_02644_, _02643_, _02131_);
  or _34843_ (_02645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _34844_ (_02646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _34845_ (_02647_, _02646_, _02645_);
  and _34846_ (_02648_, _02647_, _01954_);
  or _34847_ (_02649_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _34848_ (_02650_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _34849_ (_02651_, _02650_, _02649_);
  and _34850_ (_02652_, _02651_, _02150_);
  or _34851_ (_02653_, _02652_, _02648_);
  and _34852_ (_02654_, _02653_, _02144_);
  or _34853_ (_02655_, _02654_, _02644_);
  and _34854_ (_02656_, _02655_, _02077_);
  or _34855_ (_02657_, _02656_, _02634_);
  and _34856_ (_02658_, _02657_, _02065_);
  or _34857_ (_02659_, _02658_, _02612_);
  and _34858_ (_02660_, _02659_, _02005_);
  and _34859_ (_02661_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _34860_ (_02662_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _34861_ (_02663_, _02662_, _02661_);
  and _34862_ (_02664_, _02663_, _01954_);
  and _34863_ (_02665_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and _34864_ (_02666_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _34865_ (_02667_, _02666_, _02665_);
  and _34866_ (_02668_, _02667_, _02150_);
  or _34867_ (_02669_, _02668_, _02664_);
  or _34868_ (_02670_, _02669_, _02144_);
  and _34869_ (_02671_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _34870_ (_02672_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _34871_ (_02673_, _02672_, _02671_);
  and _34872_ (_02674_, _02673_, _01954_);
  and _34873_ (_02675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and _34874_ (_02676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _34875_ (_02677_, _02676_, _02675_);
  and _34876_ (_02678_, _02677_, _02150_);
  or _34877_ (_02679_, _02678_, _02674_);
  or _34878_ (_02680_, _02679_, _02131_);
  and _34879_ (_02681_, _02680_, _02157_);
  and _34880_ (_02682_, _02681_, _02670_);
  or _34881_ (_02683_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _34882_ (_02684_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _34883_ (_02685_, _02684_, _02683_);
  and _34884_ (_02686_, _02685_, _01954_);
  or _34885_ (_02687_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _34886_ (_02688_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and _34887_ (_02689_, _02688_, _02687_);
  and _34888_ (_02690_, _02689_, _02150_);
  or _34889_ (_02691_, _02690_, _02686_);
  or _34890_ (_02692_, _02691_, _02144_);
  or _34891_ (_02693_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _34892_ (_02694_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and _34893_ (_02695_, _02694_, _02693_);
  and _34894_ (_02696_, _02695_, _01954_);
  or _34895_ (_02697_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _34896_ (_02698_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _34897_ (_02699_, _02698_, _02697_);
  and _34898_ (_02700_, _02699_, _02150_);
  or _34899_ (_02701_, _02700_, _02696_);
  or _34900_ (_02702_, _02701_, _02131_);
  and _34901_ (_02703_, _02702_, _02077_);
  and _34902_ (_02704_, _02703_, _02692_);
  or _34903_ (_02705_, _02704_, _02682_);
  and _34904_ (_02707_, _02705_, _02065_);
  and _34905_ (_02708_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _34906_ (_02709_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _34907_ (_02710_, _02709_, _02708_);
  and _34908_ (_02711_, _02710_, _01954_);
  and _34909_ (_02712_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _34910_ (_02713_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _34911_ (_02714_, _02713_, _02712_);
  and _34912_ (_02716_, _02714_, _02150_);
  or _34913_ (_02717_, _02716_, _02711_);
  or _34914_ (_02718_, _02717_, _02144_);
  and _34915_ (_02719_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _34916_ (_02720_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _34917_ (_02721_, _02720_, _02719_);
  and _34918_ (_02722_, _02721_, _01954_);
  and _34919_ (_02723_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _34920_ (_02724_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _34921_ (_02725_, _02724_, _02723_);
  and _34922_ (_02726_, _02725_, _02150_);
  or _34923_ (_02727_, _02726_, _02722_);
  or _34924_ (_02728_, _02727_, _02131_);
  and _34925_ (_02729_, _02728_, _02157_);
  and _34926_ (_02730_, _02729_, _02718_);
  or _34927_ (_02731_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _34928_ (_02732_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _34929_ (_02733_, _02732_, _02150_);
  and _34930_ (_02734_, _02733_, _02731_);
  or _34931_ (_02735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _34932_ (_02736_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _34933_ (_02737_, _02736_, _01954_);
  and _34934_ (_02738_, _02737_, _02735_);
  or _34935_ (_02739_, _02738_, _02734_);
  or _34936_ (_02740_, _02739_, _02144_);
  or _34937_ (_02741_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _34938_ (_02742_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _34939_ (_02743_, _02742_, _02150_);
  and _34940_ (_02744_, _02743_, _02741_);
  or _34941_ (_02745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _34942_ (_02746_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _34943_ (_02747_, _02746_, _01954_);
  and _34944_ (_02748_, _02747_, _02745_);
  or _34945_ (_02749_, _02748_, _02744_);
  or _34946_ (_02750_, _02749_, _02131_);
  and _34947_ (_02751_, _02750_, _02077_);
  and _34948_ (_02752_, _02751_, _02740_);
  or _34949_ (_02753_, _02752_, _02730_);
  and _34950_ (_02754_, _02753_, _02194_);
  or _34951_ (_02755_, _02754_, _02707_);
  and _34952_ (_02756_, _02755_, _02143_);
  or _34953_ (_02757_, _02756_, _02660_);
  or _34954_ (_02758_, _02757_, _02054_);
  and _34955_ (_02759_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and _34956_ (_02760_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _34957_ (_02761_, _02760_, _02759_);
  and _34958_ (_02762_, _02761_, _02150_);
  and _34959_ (_02763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _34960_ (_02764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _34961_ (_02765_, _02764_, _02763_);
  and _34962_ (_02766_, _02765_, _01954_);
  or _34963_ (_02767_, _02766_, _02762_);
  or _34964_ (_02768_, _02767_, _02144_);
  and _34965_ (_02769_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _34966_ (_02770_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _34967_ (_02771_, _02770_, _02769_);
  and _34968_ (_02772_, _02771_, _02150_);
  and _34969_ (_02773_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _34970_ (_02774_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _34971_ (_02775_, _02774_, _02773_);
  and _34972_ (_02776_, _02775_, _01954_);
  or _34973_ (_02777_, _02776_, _02772_);
  or _34974_ (_02778_, _02777_, _02131_);
  and _34975_ (_02779_, _02778_, _02157_);
  and _34976_ (_02780_, _02779_, _02768_);
  or _34977_ (_02781_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _34978_ (_02782_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and _34979_ (_02783_, _02782_, _01954_);
  and _34980_ (_02785_, _02783_, _02781_);
  or _34981_ (_02786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _34982_ (_02787_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _34983_ (_02788_, _02787_, _02150_);
  and _34984_ (_02789_, _02788_, _02786_);
  or _34985_ (_02790_, _02789_, _02785_);
  or _34986_ (_02791_, _02790_, _02144_);
  or _34987_ (_02792_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _34988_ (_02793_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and _34989_ (_02794_, _02793_, _01954_);
  and _34990_ (_02795_, _02794_, _02792_);
  or _34991_ (_02796_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _34992_ (_02797_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _34993_ (_02798_, _02797_, _02150_);
  and _34994_ (_02799_, _02798_, _02796_);
  or _34995_ (_02800_, _02799_, _02795_);
  or _34996_ (_02801_, _02800_, _02131_);
  and _34997_ (_02802_, _02801_, _02077_);
  and _34998_ (_02803_, _02802_, _02791_);
  or _34999_ (_02804_, _02803_, _02780_);
  and _35000_ (_02805_, _02804_, _02194_);
  and _35001_ (_02806_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _35002_ (_02807_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _35003_ (_02808_, _02807_, _01954_);
  or _35004_ (_02809_, _02808_, _02806_);
  and _35005_ (_02810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _35006_ (_02811_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _35007_ (_02812_, _02811_, _02150_);
  or _35008_ (_02813_, _02812_, _02810_);
  and _35009_ (_02814_, _02813_, _02809_);
  or _35010_ (_02815_, _02814_, _02144_);
  and _35011_ (_02816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _35012_ (_02817_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _35013_ (_02818_, _02817_, _01954_);
  or _35014_ (_02819_, _02818_, _02816_);
  and _35015_ (_02820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _35016_ (_02821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _35017_ (_02822_, _02821_, _02150_);
  or _35018_ (_02823_, _02822_, _02820_);
  and _35019_ (_02824_, _02823_, _02819_);
  or _35020_ (_02825_, _02824_, _02131_);
  and _35021_ (_02826_, _02825_, _02157_);
  and _35022_ (_02827_, _02826_, _02815_);
  or _35023_ (_02828_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _35024_ (_02829_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _35025_ (_02830_, _02829_, _02828_);
  or _35026_ (_02831_, _02830_, _02150_);
  or _35027_ (_02832_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _35028_ (_02833_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _35029_ (_02834_, _02833_, _02832_);
  or _35030_ (_02835_, _02834_, _01954_);
  and _35031_ (_02836_, _02835_, _02831_);
  or _35032_ (_02837_, _02836_, _02144_);
  or _35033_ (_02838_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _35034_ (_02839_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _35035_ (_02840_, _02839_, _02838_);
  or _35036_ (_02841_, _02840_, _02150_);
  or _35037_ (_02842_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _35038_ (_02843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _35039_ (_02844_, _02843_, _02842_);
  or _35040_ (_02845_, _02844_, _01954_);
  and _35041_ (_02846_, _02845_, _02841_);
  or _35042_ (_02847_, _02846_, _02131_);
  and _35043_ (_02848_, _02847_, _02077_);
  and _35044_ (_02849_, _02848_, _02837_);
  or _35045_ (_02850_, _02849_, _02827_);
  and _35046_ (_02851_, _02850_, _02065_);
  or _35047_ (_02852_, _02851_, _02805_);
  and _35048_ (_02853_, _02852_, _02143_);
  and _35049_ (_02854_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _35050_ (_02855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _35051_ (_02856_, _02855_, _02854_);
  and _35052_ (_02857_, _02856_, _01954_);
  and _35053_ (_02858_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _35054_ (_02859_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _35055_ (_02860_, _02859_, _02858_);
  and _35056_ (_02861_, _02860_, _02150_);
  or _35057_ (_02862_, _02861_, _02857_);
  and _35058_ (_02863_, _02862_, _02131_);
  and _35059_ (_02864_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _35060_ (_02865_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _35061_ (_02866_, _02865_, _02864_);
  and _35062_ (_02867_, _02866_, _01954_);
  and _35063_ (_02868_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _35064_ (_02869_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _35065_ (_02870_, _02869_, _02868_);
  and _35066_ (_02871_, _02870_, _02150_);
  or _35067_ (_02872_, _02871_, _02867_);
  and _35068_ (_02873_, _02872_, _02144_);
  or _35069_ (_02874_, _02873_, _02863_);
  and _35070_ (_02875_, _02874_, _02157_);
  or _35071_ (_02876_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _35072_ (_02877_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _35073_ (_02878_, _02877_, _02876_);
  and _35074_ (_02879_, _02878_, _01954_);
  or _35075_ (_02880_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _35076_ (_02881_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _35077_ (_02882_, _02881_, _02880_);
  and _35078_ (_02883_, _02882_, _02150_);
  or _35079_ (_02884_, _02883_, _02879_);
  and _35080_ (_02885_, _02884_, _02131_);
  or _35081_ (_02886_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _35082_ (_02887_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _35083_ (_02888_, _02887_, _02886_);
  and _35084_ (_02889_, _02888_, _01954_);
  or _35085_ (_02890_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _35086_ (_02891_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _35087_ (_02892_, _02891_, _02890_);
  and _35088_ (_02893_, _02892_, _02150_);
  or _35089_ (_02894_, _02893_, _02889_);
  and _35090_ (_02895_, _02894_, _02144_);
  or _35091_ (_02896_, _02895_, _02885_);
  and _35092_ (_02897_, _02896_, _02077_);
  or _35093_ (_02898_, _02897_, _02875_);
  and _35094_ (_02899_, _02898_, _02065_);
  and _35095_ (_02900_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and _35096_ (_02901_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or _35097_ (_02902_, _02901_, _02900_);
  and _35098_ (_02903_, _02902_, _01954_);
  and _35099_ (_02904_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and _35100_ (_02905_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or _35101_ (_02906_, _02905_, _02904_);
  and _35102_ (_02907_, _02906_, _02150_);
  or _35103_ (_02908_, _02907_, _02903_);
  and _35104_ (_02909_, _02908_, _02131_);
  and _35105_ (_02910_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  and _35106_ (_02911_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or _35107_ (_02912_, _02911_, _02910_);
  and _35108_ (_02913_, _02912_, _01954_);
  and _35109_ (_02914_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and _35110_ (_02915_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or _35111_ (_02916_, _02915_, _02914_);
  and _35112_ (_02917_, _02916_, _02150_);
  or _35113_ (_02918_, _02917_, _02913_);
  and _35114_ (_02919_, _02918_, _02144_);
  or _35115_ (_02920_, _02919_, _02909_);
  and _35116_ (_02921_, _02920_, _02157_);
  or _35117_ (_02922_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _35118_ (_02923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and _35119_ (_02924_, _02923_, _02922_);
  and _35120_ (_02925_, _02924_, _01954_);
  or _35121_ (_02926_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or _35122_ (_02927_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and _35123_ (_02928_, _02927_, _02926_);
  and _35124_ (_02929_, _02928_, _02150_);
  or _35125_ (_02930_, _02929_, _02925_);
  and _35126_ (_02931_, _02930_, _02131_);
  or _35127_ (_02932_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or _35128_ (_02933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  and _35129_ (_02934_, _02933_, _02932_);
  and _35130_ (_02935_, _02934_, _01954_);
  or _35131_ (_02936_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or _35132_ (_02937_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and _35133_ (_02938_, _02937_, _02936_);
  and _35134_ (_02939_, _02938_, _02150_);
  or _35135_ (_02940_, _02939_, _02935_);
  and _35136_ (_02941_, _02940_, _02144_);
  or _35137_ (_02942_, _02941_, _02931_);
  and _35138_ (_02943_, _02942_, _02077_);
  or _35139_ (_02944_, _02943_, _02921_);
  and _35140_ (_02945_, _02944_, _02194_);
  or _35141_ (_02946_, _02945_, _02899_);
  and _35142_ (_02947_, _02946_, _02005_);
  or _35143_ (_02948_, _02947_, _02853_);
  or _35144_ (_02949_, _02948_, _02374_);
  and _35145_ (_02950_, _02949_, _02758_);
  or _35146_ (_02951_, _02950_, _01748_);
  and _35147_ (_02952_, _02951_, _02566_);
  or _35148_ (_02953_, _02952_, _02141_);
  not _35149_ (_02954_, _02141_);
  or _35150_ (_02955_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _35151_ (_02956_, _02955_, _27355_);
  and _35152_ (_02715_, _02956_, _02953_);
  nor _35153_ (_02957_, _02138_, _01623_);
  nor _35154_ (_02958_, _02138_, _01862_);
  nor _35155_ (_02959_, _02958_, _02957_);
  nor _35156_ (_02960_, _02138_, _02084_);
  nor _35157_ (_02961_, _02138_, _02074_);
  nor _35158_ (_02962_, _02961_, _02960_);
  and _35159_ (_02963_, _02962_, _02959_);
  and _35160_ (_02964_, _02137_, _02063_);
  nor _35161_ (_02965_, _02138_, _01959_);
  nor _35162_ (_02966_, _02965_, _02964_);
  nor _35163_ (_02967_, _01650_, _01620_);
  and _35164_ (_02968_, _02967_, _02137_);
  not _35165_ (_02969_, _02968_);
  and _35166_ (_02970_, _02969_, _02966_);
  and _35167_ (_02971_, _02970_, _02137_);
  and _35168_ (_02972_, _02971_, _02963_);
  not _35169_ (_02973_, _02972_);
  and _35170_ (_02974_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _35171_ (_02975_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25182_);
  and _35172_ (_02976_, _02975_, _25168_);
  and _35173_ (_02977_, _02976_, _25574_);
  nor _35174_ (_02978_, _26521_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not _35175_ (_02979_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _35176_ (_02980_, _02976_, _02979_);
  and _35177_ (_02981_, _02980_, _24073_);
  or _35178_ (_02982_, _02981_, _02978_);
  or _35179_ (_02983_, _02982_, _02977_);
  and _35180_ (_02985_, _02983_, _02972_);
  or _35181_ (_03577_, _02985_, _02974_);
  and _35182_ (_02986_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand _35183_ (_02987_, _02975_, _25172_);
  nor _35184_ (_02988_, _02987_, _25514_);
  nor _35185_ (_02989_, _26512_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35186_ (_02990_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _35187_ (_02991_, _02975_, _25177_);
  or _35188_ (_02992_, _02991_, _02990_);
  and _35189_ (_02993_, _02975_, _25174_);
  or _35190_ (_02994_, _02993_, _02992_);
  and _35191_ (_02995_, _02994_, _24023_);
  or _35192_ (_02996_, _02995_, _02989_);
  or _35193_ (_02997_, _02996_, _02988_);
  and _35194_ (_02998_, _02997_, _02972_);
  or _35195_ (_03581_, _02998_, _02986_);
  and _35196_ (_02999_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _35197_ (_03000_, _02975_, _25175_);
  nor _35198_ (_03001_, _03000_, _25514_);
  nor _35199_ (_03002_, _26505_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _35200_ (_03003_, _25175_, _25182_);
  and _35201_ (_03004_, _24059_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35202_ (_03005_, _03004_, _03003_);
  or _35203_ (_03006_, _03005_, _03002_);
  or _35204_ (_03007_, _03006_, _03001_);
  and _35205_ (_03008_, _03007_, _02972_);
  or _35206_ (_03587_, _03008_, _02999_);
  and _35207_ (_03009_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _35208_ (_03010_, _02991_, _25574_);
  nor _35209_ (_03011_, _26497_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _35210_ (_03012_, _25177_, _25182_);
  and _35211_ (_03013_, _24009_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35212_ (_03014_, _03013_, _03012_);
  or _35213_ (_03015_, _03014_, _03011_);
  or _35214_ (_03016_, _03015_, _03010_);
  and _35215_ (_03017_, _03016_, _02972_);
  or _35216_ (_03591_, _03017_, _03009_);
  and _35217_ (_03018_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand _35218_ (_03019_, _02990_, _25168_);
  nor _35219_ (_03020_, _03019_, _25514_);
  nor _35220_ (_03021_, _26489_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _35221_ (_03022_, _25168_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _35222_ (_03023_, _23958_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35223_ (_03024_, _03023_, _03022_);
  or _35224_ (_03025_, _03024_, _03021_);
  or _35225_ (_03026_, _03025_, _03020_);
  and _35226_ (_03027_, _03026_, _02972_);
  or _35227_ (_03595_, _03027_, _03018_);
  and _35228_ (_03028_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand _35229_ (_03029_, _02990_, _25172_);
  nor _35230_ (_03030_, _03029_, _25514_);
  nor _35231_ (_03031_, _26482_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _35232_ (_03032_, _25172_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _35233_ (_03033_, _23995_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35234_ (_03034_, _03033_, _03032_);
  or _35235_ (_03035_, _03034_, _03031_);
  or _35236_ (_03036_, _03035_, _03030_);
  and _35237_ (_03037_, _03036_, _02972_);
  or _35238_ (_03600_, _03037_, _03028_);
  and _35239_ (_03038_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand _35240_ (_03040_, _02990_, _25175_);
  nor _35241_ (_03041_, _03040_, _25514_);
  nor _35242_ (_03042_, _26475_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _35243_ (_03043_, _25175_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _35244_ (_03044_, _24040_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _35245_ (_03045_, _03044_, _03043_);
  or _35246_ (_03046_, _03045_, _03042_);
  or _35247_ (_03047_, _03046_, _03041_);
  and _35248_ (_03048_, _03047_, _02972_);
  or _35249_ (_03605_, _03048_, _03038_);
  and _35250_ (_03050_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _35251_ (_03051_, _02990_, _25177_);
  not _35252_ (_03052_, _03051_);
  nor _35253_ (_03053_, _03052_, _25514_);
  nand _35254_ (_03054_, _26543_, _02979_);
  or _35255_ (_03055_, _23978_, _02979_);
  and _35256_ (_03056_, _03055_, _03052_);
  and _35257_ (_03057_, _03056_, _03054_);
  or _35258_ (_03058_, _03057_, _03053_);
  and _35259_ (_03059_, _03058_, _02972_);
  or _35260_ (_03607_, _03059_, _03050_);
  and _35261_ (_03060_, _02983_, _02137_);
  and _35262_ (_03061_, _02957_, _01862_);
  and _35263_ (_03062_, _03061_, _02962_);
  and _35264_ (_03063_, _03062_, _02970_);
  and _35265_ (_03064_, _03063_, _03060_);
  not _35266_ (_03065_, _03063_);
  and _35267_ (_03066_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _35268_ (_03613_, _03066_, _03064_);
  and _35269_ (_03067_, _02997_, _02137_);
  and _35270_ (_03069_, _03063_, _03067_);
  and _35271_ (_03070_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _35272_ (_03616_, _03070_, _03069_);
  and _35273_ (_03071_, _03007_, _02137_);
  and _35274_ (_03072_, _03063_, _03071_);
  and _35275_ (_03073_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _35276_ (_03619_, _03073_, _03072_);
  and _35277_ (_03074_, _03016_, _02137_);
  and _35278_ (_03075_, _03063_, _03074_);
  and _35279_ (_03076_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _35280_ (_03622_, _03076_, _03075_);
  and _35281_ (_03077_, _03026_, _02137_);
  and _35282_ (_03078_, _03063_, _03077_);
  and _35283_ (_03079_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _35284_ (_03626_, _03079_, _03078_);
  and _35285_ (_03080_, _03036_, _02137_);
  and _35286_ (_03081_, _03063_, _03080_);
  and _35287_ (_03082_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _35288_ (_03629_, _03082_, _03081_);
  and _35289_ (_03083_, _03047_, _02137_);
  and _35290_ (_03085_, _03063_, _03083_);
  and _35291_ (_03086_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _35292_ (_03632_, _03086_, _03085_);
  and _35293_ (_03087_, _03058_, _02137_);
  and _35294_ (_03088_, _03063_, _03087_);
  and _35295_ (_03089_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _35296_ (_03634_, _03089_, _03088_);
  and _35297_ (_03090_, _02958_, _01623_);
  and _35298_ (_03091_, _03090_, _02962_);
  and _35299_ (_03092_, _03091_, _02970_);
  and _35300_ (_03093_, _03092_, _03060_);
  not _35301_ (_03094_, _03092_);
  and _35302_ (_03095_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _35303_ (_03641_, _03095_, _03093_);
  and _35304_ (_03096_, _03092_, _03067_);
  and _35305_ (_03097_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _35306_ (_03644_, _03097_, _03096_);
  and _35307_ (_03098_, _03092_, _03071_);
  and _35308_ (_03099_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _35309_ (_03647_, _03099_, _03098_);
  and _35310_ (_03101_, _03092_, _03074_);
  and _35311_ (_03102_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _35312_ (_03650_, _03102_, _03101_);
  and _35313_ (_03103_, _03092_, _03077_);
  and _35314_ (_03104_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _35315_ (_03653_, _03104_, _03103_);
  and _35316_ (_03105_, _03092_, _03080_);
  and _35317_ (_03106_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _35318_ (_03656_, _03106_, _03105_);
  and _35319_ (_03107_, _03092_, _03083_);
  and _35320_ (_03109_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _35321_ (_03659_, _03109_, _03107_);
  and _35322_ (_03110_, _03092_, _03087_);
  and _35323_ (_03111_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _35324_ (_03662_, _03111_, _03110_);
  and _35325_ (_03112_, _02958_, _02957_);
  and _35326_ (_03113_, _03112_, _02962_);
  and _35327_ (_03114_, _03113_, _02970_);
  and _35328_ (_03115_, _03114_, _03060_);
  not _35329_ (_03116_, _03114_);
  and _35330_ (_03118_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _35331_ (_03667_, _03118_, _03115_);
  and _35332_ (_03119_, _03114_, _03067_);
  and _35333_ (_03120_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _35334_ (_03670_, _03120_, _03119_);
  and _35335_ (_03121_, _03114_, _03071_);
  and _35336_ (_03122_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _35337_ (_03673_, _03122_, _03121_);
  and _35338_ (_03123_, _03114_, _03074_);
  and _35339_ (_03124_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _35340_ (_03676_, _03124_, _03123_);
  and _35341_ (_03126_, _03114_, _03077_);
  and _35342_ (_03127_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _35343_ (_03679_, _03127_, _03126_);
  and _35344_ (_03128_, _03114_, _03080_);
  and _35345_ (_03129_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _35346_ (_03682_, _03129_, _03128_);
  and _35347_ (_03130_, _03114_, _03083_);
  and _35348_ (_03131_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _35349_ (_03685_, _03131_, _03130_);
  and _35350_ (_03133_, _03114_, _03087_);
  and _35351_ (_03134_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _35352_ (_03688_, _03134_, _03133_);
  and _35353_ (_03135_, _02960_, _02074_);
  and _35354_ (_03136_, _03135_, _02959_);
  and _35355_ (_03137_, _03136_, _02970_);
  and _35356_ (_03138_, _03137_, _03060_);
  not _35357_ (_03139_, _03137_);
  and _35358_ (_03140_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _35359_ (_03694_, _03140_, _03138_);
  and _35360_ (_03142_, _03137_, _03067_);
  and _35361_ (_03143_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _35362_ (_03697_, _03143_, _03142_);
  and _35363_ (_03144_, _03137_, _03071_);
  and _35364_ (_03145_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _35365_ (_03700_, _03145_, _03144_);
  and _35366_ (_03146_, _03137_, _03074_);
  and _35367_ (_03147_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _35368_ (_03704_, _03147_, _03146_);
  and _35369_ (_03148_, _03137_, _03077_);
  and _35370_ (_03150_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _35371_ (_03707_, _03150_, _03148_);
  and _35372_ (_03151_, _03137_, _03080_);
  and _35373_ (_03152_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _35374_ (_03710_, _03152_, _03151_);
  and _35375_ (_03153_, _03137_, _03083_);
  and _35376_ (_03154_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _35377_ (_03713_, _03154_, _03153_);
  and _35378_ (_03155_, _03137_, _03087_);
  and _35379_ (_03156_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _35380_ (_03716_, _03156_, _03155_);
  and _35381_ (_03159_, _03135_, _03061_);
  and _35382_ (_03160_, _03159_, _02970_);
  and _35383_ (_03161_, _03160_, _03060_);
  not _35384_ (_03162_, _03160_);
  and _35385_ (_03163_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _35386_ (_03720_, _03163_, _03161_);
  and _35387_ (_03164_, _03160_, _03067_);
  and _35388_ (_03165_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _35389_ (_03723_, _03165_, _03164_);
  and _35390_ (_03167_, _03160_, _03071_);
  and _35391_ (_03168_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _35392_ (_03726_, _03168_, _03167_);
  and _35393_ (_03169_, _03160_, _03074_);
  and _35394_ (_03170_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _35395_ (_03729_, _03170_, _03169_);
  and _35396_ (_03171_, _03160_, _03077_);
  and _35397_ (_03172_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _35398_ (_03733_, _03172_, _03171_);
  and _35399_ (_03173_, _03160_, _03080_);
  and _35400_ (_03174_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _35401_ (_03736_, _03174_, _03173_);
  and _35402_ (_03175_, _03160_, _03083_);
  and _35403_ (_03176_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _35404_ (_03739_, _03176_, _03175_);
  and _35405_ (_03177_, _03160_, _03087_);
  and _35406_ (_03178_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _35407_ (_03741_, _03178_, _03177_);
  and _35408_ (_03179_, _03135_, _03090_);
  and _35409_ (_03180_, _03179_, _02970_);
  and _35410_ (_03181_, _03180_, _03060_);
  not _35411_ (_03182_, _03180_);
  and _35412_ (_03183_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _35413_ (_03745_, _03183_, _03181_);
  and _35414_ (_03184_, _03180_, _03067_);
  and _35415_ (_03185_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _35416_ (_03748_, _03185_, _03184_);
  and _35417_ (_03186_, _03180_, _03071_);
  and _35418_ (_03187_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _35419_ (_03751_, _03187_, _03186_);
  and _35420_ (_03188_, _03180_, _03074_);
  and _35421_ (_03189_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _35422_ (_03754_, _03189_, _03188_);
  and _35423_ (_03190_, _03180_, _03077_);
  and _35424_ (_03191_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _35425_ (_03758_, _03191_, _03190_);
  and _35426_ (_03192_, _03180_, _03080_);
  and _35427_ (_03193_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _35428_ (_03761_, _03193_, _03192_);
  and _35429_ (_03194_, _03180_, _03083_);
  and _35430_ (_03195_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _35431_ (_03764_, _03195_, _03194_);
  and _35432_ (_03196_, _03180_, _03087_);
  and _35433_ (_03197_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _35434_ (_03766_, _03197_, _03196_);
  and _35435_ (_03198_, _03135_, _03112_);
  and _35436_ (_03199_, _03198_, _02970_);
  and _35437_ (_03200_, _03199_, _03060_);
  not _35438_ (_03201_, _03199_);
  and _35439_ (_03202_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _35440_ (_03771_, _03202_, _03200_);
  and _35441_ (_03203_, _03199_, _03067_);
  and _35442_ (_03204_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _35443_ (_03774_, _03204_, _03203_);
  and _35444_ (_03205_, _03199_, _03071_);
  and _35445_ (_03206_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _35446_ (_03777_, _03206_, _03205_);
  and _35447_ (_03207_, _03199_, _03074_);
  and _35448_ (_03208_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _35449_ (_03780_, _03208_, _03207_);
  and _35450_ (_03209_, _03199_, _03077_);
  and _35451_ (_03210_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _35452_ (_03784_, _03210_, _03209_);
  and _35453_ (_03211_, _03199_, _03080_);
  and _35454_ (_03212_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _35455_ (_03787_, _03212_, _03211_);
  and _35456_ (_03213_, _03199_, _03083_);
  and _35457_ (_03214_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _35458_ (_03790_, _03214_, _03213_);
  and _35459_ (_03215_, _03199_, _03087_);
  and _35460_ (_03216_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _35461_ (_03793_, _03216_, _03215_);
  and _35462_ (_03217_, _02961_, _02084_);
  and _35463_ (_03218_, _03217_, _02959_);
  and _35464_ (_03219_, _03218_, _02970_);
  and _35465_ (_03220_, _03219_, _03060_);
  not _35466_ (_03221_, _03219_);
  and _35467_ (_03222_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _35468_ (_03799_, _03222_, _03220_);
  and _35469_ (_03223_, _03219_, _03067_);
  and _35470_ (_03224_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _35471_ (_03802_, _03224_, _03223_);
  and _35472_ (_03225_, _03219_, _03071_);
  and _35473_ (_03226_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _35474_ (_03805_, _03226_, _03225_);
  and _35475_ (_03227_, _03219_, _03074_);
  and _35476_ (_03228_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _35477_ (_03808_, _03228_, _03227_);
  and _35478_ (_03229_, _03219_, _03077_);
  and _35479_ (_03230_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _35480_ (_03812_, _03230_, _03229_);
  and _35481_ (_03231_, _03219_, _03080_);
  and _35482_ (_03232_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _35483_ (_03815_, _03232_, _03231_);
  and _35484_ (_03233_, _03219_, _03083_);
  and _35485_ (_03234_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _35486_ (_03818_, _03234_, _03233_);
  and _35487_ (_03235_, _03219_, _03087_);
  and _35488_ (_03236_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _35489_ (_03820_, _03236_, _03235_);
  and _35490_ (_03237_, _03217_, _03061_);
  and _35491_ (_03238_, _03237_, _02970_);
  and _35492_ (_03239_, _03238_, _03060_);
  not _35493_ (_03240_, _03238_);
  and _35494_ (_03241_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _35495_ (_03824_, _03241_, _03239_);
  and _35496_ (_03242_, _03238_, _03067_);
  and _35497_ (_03243_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _35498_ (_03827_, _03243_, _03242_);
  and _35499_ (_03244_, _03238_, _03071_);
  and _35500_ (_03245_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _35501_ (_03830_, _03245_, _03244_);
  and _35502_ (_03246_, _03238_, _03074_);
  and _35503_ (_03247_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _35504_ (_03833_, _03247_, _03246_);
  and _35505_ (_03248_, _03238_, _03077_);
  and _35506_ (_03249_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _35507_ (_03837_, _03249_, _03248_);
  and _35508_ (_03250_, _03238_, _03080_);
  and _35509_ (_03251_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _35510_ (_03840_, _03251_, _03250_);
  and _35511_ (_03252_, _03238_, _03083_);
  and _35512_ (_03253_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _35513_ (_03843_, _03253_, _03252_);
  and _35514_ (_03254_, _03238_, _03087_);
  and _35515_ (_03255_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _35516_ (_03845_, _03255_, _03254_);
  and _35517_ (_03256_, _03217_, _03090_);
  and _35518_ (_03257_, _03256_, _02970_);
  and _35519_ (_03258_, _03257_, _03060_);
  not _35520_ (_03259_, _03257_);
  and _35521_ (_03260_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _35522_ (_03850_, _03260_, _03258_);
  and _35523_ (_03261_, _03257_, _03067_);
  and _35524_ (_03262_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _35525_ (_03853_, _03262_, _03261_);
  and _35526_ (_03263_, _03257_, _03071_);
  and _35527_ (_03264_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _35528_ (_03856_, _03264_, _03263_);
  and _35529_ (_03265_, _03257_, _03074_);
  and _35530_ (_03266_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _35531_ (_03859_, _03266_, _03265_);
  and _35532_ (_03267_, _03257_, _03077_);
  and _35533_ (_03268_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _35534_ (_03862_, _03268_, _03267_);
  and _35535_ (_03269_, _03257_, _03080_);
  and _35536_ (_03270_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _35537_ (_03865_, _03270_, _03269_);
  and _35538_ (_03271_, _03257_, _03083_);
  and _35539_ (_03272_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _35540_ (_03868_, _03272_, _03271_);
  and _35541_ (_03273_, _03257_, _03087_);
  and _35542_ (_03274_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _35543_ (_03871_, _03274_, _03273_);
  and _35544_ (_03275_, _03217_, _03112_);
  and _35545_ (_03276_, _03275_, _02970_);
  and _35546_ (_03277_, _03276_, _03060_);
  not _35547_ (_03278_, _03276_);
  and _35548_ (_03279_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _35549_ (_03875_, _03279_, _03277_);
  and _35550_ (_03280_, _03276_, _03067_);
  and _35551_ (_03281_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _35552_ (_03878_, _03281_, _03280_);
  and _35553_ (_03282_, _03276_, _03071_);
  and _35554_ (_03283_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _35555_ (_03881_, _03283_, _03282_);
  and _35556_ (_03284_, _03276_, _03074_);
  and _35557_ (_03285_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _35558_ (_03884_, _03285_, _03284_);
  and _35559_ (_03286_, _03276_, _03077_);
  and _35560_ (_03287_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _35561_ (_03887_, _03287_, _03286_);
  and _35562_ (_03288_, _03276_, _03080_);
  and _35563_ (_03289_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _35564_ (_03891_, _03289_, _03288_);
  and _35565_ (_03290_, _03276_, _03083_);
  and _35566_ (_03291_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _35567_ (_03894_, _03291_, _03290_);
  and _35568_ (_03292_, _03276_, _03087_);
  and _35569_ (_03293_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _35570_ (_03896_, _03293_, _03292_);
  and _35571_ (_03294_, _02961_, _02960_);
  and _35572_ (_03295_, _03294_, _02959_);
  and _35573_ (_03296_, _03295_, _02970_);
  and _35574_ (_03297_, _03296_, _03060_);
  not _35575_ (_03298_, _03296_);
  and _35576_ (_03299_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _35577_ (_03901_, _03299_, _03297_);
  and _35578_ (_03300_, _03296_, _03067_);
  and _35579_ (_03301_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _35580_ (_03904_, _03301_, _03300_);
  and _35581_ (_03303_, _03296_, _03071_);
  and _35582_ (_03304_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _35583_ (_03907_, _03304_, _03303_);
  and _35584_ (_03305_, _03296_, _03074_);
  and _35585_ (_03306_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _35586_ (_03910_, _03306_, _03305_);
  and _35587_ (_03307_, _03296_, _03077_);
  and _35588_ (_03308_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _35589_ (_03913_, _03308_, _03307_);
  and _35590_ (_03309_, _03296_, _03080_);
  and _35591_ (_03310_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _35592_ (_03917_, _03310_, _03309_);
  and _35593_ (_03311_, _03296_, _03083_);
  and _35594_ (_03312_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _35595_ (_03920_, _03312_, _03311_);
  and _35596_ (_03313_, _03296_, _03087_);
  and _35597_ (_03314_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _35598_ (_03922_, _03314_, _03313_);
  and _35599_ (_03315_, _03294_, _03061_);
  and _35600_ (_03316_, _03315_, _02970_);
  and _35601_ (_03317_, _03316_, _03060_);
  not _35602_ (_03318_, _03316_);
  and _35603_ (_03319_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _35604_ (_03926_, _03319_, _03317_);
  and _35605_ (_03320_, _03316_, _03067_);
  and _35606_ (_03321_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _35607_ (_03929_, _03321_, _03320_);
  and _35608_ (_03322_, _03316_, _03071_);
  and _35609_ (_03323_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _35610_ (_03932_, _03323_, _03322_);
  and _35611_ (_03324_, _03316_, _03074_);
  and _35612_ (_03325_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _35613_ (_03935_, _03325_, _03324_);
  and _35614_ (_03326_, _03316_, _03077_);
  and _35615_ (_03327_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _35616_ (_03938_, _03327_, _03326_);
  and _35617_ (_03328_, _03316_, _03080_);
  and _35618_ (_03329_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _35619_ (_03942_, _03329_, _03328_);
  and _35620_ (_03330_, _03316_, _03083_);
  and _35621_ (_03331_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _35622_ (_03945_, _03331_, _03330_);
  and _35623_ (_03332_, _03316_, _03087_);
  and _35624_ (_03333_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _35625_ (_03947_, _03333_, _03332_);
  and _35626_ (_03334_, _03294_, _03090_);
  and _35627_ (_03335_, _03334_, _02970_);
  and _35628_ (_03336_, _03335_, _03060_);
  not _35629_ (_03337_, _03335_);
  and _35630_ (_03338_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _35631_ (_03952_, _03338_, _03336_);
  and _35632_ (_03339_, _03335_, _03067_);
  and _35633_ (_03340_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _35634_ (_03955_, _03340_, _03339_);
  and _35635_ (_03341_, _03335_, _03071_);
  and _35636_ (_03342_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _35637_ (_03958_, _03342_, _03341_);
  and _35638_ (_03343_, _03335_, _03074_);
  and _35639_ (_03344_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _35640_ (_03961_, _03344_, _03343_);
  and _35641_ (_03345_, _03335_, _03077_);
  and _35642_ (_03346_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _35643_ (_03964_, _03346_, _03345_);
  and _35644_ (_03347_, _03335_, _03080_);
  and _35645_ (_03348_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _35646_ (_03967_, _03348_, _03347_);
  and _35647_ (_03349_, _03335_, _03083_);
  and _35648_ (_03350_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _35649_ (_03970_, _03350_, _03349_);
  and _35650_ (_03351_, _03335_, _03087_);
  and _35651_ (_03352_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _35652_ (_03973_, _03352_, _03351_);
  and _35653_ (_03353_, _03294_, _03112_);
  and _35654_ (_03354_, _03353_, _02970_);
  and _35655_ (_03355_, _03354_, _03060_);
  not _35656_ (_03356_, _03354_);
  and _35657_ (_03357_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _35658_ (_03977_, _03357_, _03355_);
  and _35659_ (_03358_, _03354_, _03067_);
  and _35660_ (_03359_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _35661_ (_03980_, _03359_, _03358_);
  and _35662_ (_03360_, _03354_, _03071_);
  and _35663_ (_03361_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _35664_ (_03983_, _03361_, _03360_);
  and _35665_ (_03362_, _03354_, _03074_);
  and _35666_ (_03363_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _35667_ (_03987_, _03363_, _03362_);
  and _35668_ (_03364_, _03354_, _03077_);
  and _35669_ (_03365_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _35670_ (_03990_, _03365_, _03364_);
  and _35671_ (_03366_, _03354_, _03080_);
  and _35672_ (_03367_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _35673_ (_03993_, _03367_, _03366_);
  and _35674_ (_03368_, _03354_, _03083_);
  and _35675_ (_03369_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _35676_ (_03997_, _03369_, _03368_);
  and _35677_ (_03370_, _03354_, _03087_);
  and _35678_ (_03371_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _35679_ (_03999_, _03371_, _03370_);
  not _35680_ (_03372_, _02967_);
  and _35681_ (_03373_, _02964_, _25085_);
  and _35682_ (_03374_, _03373_, _03372_);
  and _35683_ (_03375_, _03374_, _02963_);
  and _35684_ (_03376_, _03375_, _03060_);
  not _35685_ (_03377_, _03375_);
  and _35686_ (_03378_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or _35687_ (_04005_, _03378_, _03376_);
  and _35688_ (_03379_, _03375_, _03067_);
  and _35689_ (_03380_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or _35690_ (_04008_, _03380_, _03379_);
  and _35691_ (_03381_, _03375_, _03071_);
  and _35692_ (_03382_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or _35693_ (_04011_, _03382_, _03381_);
  and _35694_ (_03383_, _03375_, _03074_);
  and _35695_ (_03384_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or _35696_ (_04014_, _03384_, _03383_);
  and _35697_ (_03385_, _03375_, _03077_);
  and _35698_ (_03386_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or _35699_ (_04017_, _03386_, _03385_);
  and _35700_ (_03387_, _03375_, _03080_);
  and _35701_ (_03388_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or _35702_ (_04021_, _03388_, _03387_);
  and _35703_ (_03389_, _03375_, _03083_);
  and _35704_ (_03390_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or _35705_ (_04024_, _03390_, _03389_);
  and _35706_ (_03391_, _03375_, _03087_);
  and _35707_ (_03392_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or _35708_ (_04026_, _03392_, _03391_);
  and _35709_ (_03393_, _03374_, _03062_);
  and _35710_ (_03394_, _03393_, _03060_);
  not _35711_ (_03395_, _03393_);
  and _35712_ (_03396_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _35713_ (_04030_, _03396_, _03394_);
  and _35714_ (_03397_, _03393_, _03067_);
  and _35715_ (_03398_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _35716_ (_04033_, _03398_, _03397_);
  and _35717_ (_03399_, _03393_, _03071_);
  and _35718_ (_03400_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _35719_ (_04036_, _03400_, _03399_);
  and _35720_ (_03401_, _03393_, _03074_);
  and _35721_ (_03402_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _35722_ (_04039_, _03402_, _03401_);
  and _35723_ (_03403_, _03393_, _03077_);
  and _35724_ (_03404_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _35725_ (_04042_, _03404_, _03403_);
  and _35726_ (_03405_, _03393_, _03080_);
  and _35727_ (_03406_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _35728_ (_04045_, _03406_, _03405_);
  and _35729_ (_03407_, _03393_, _03083_);
  and _35730_ (_03408_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _35731_ (_04049_, _03408_, _03407_);
  and _35732_ (_03409_, _03393_, _03087_);
  and _35733_ (_03410_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _35734_ (_04051_, _03410_, _03409_);
  and _35735_ (_03411_, _03374_, _03091_);
  and _35736_ (_03412_, _03411_, _03060_);
  not _35737_ (_03413_, _03411_);
  and _35738_ (_03414_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _35739_ (_04055_, _03414_, _03412_);
  and _35740_ (_03415_, _03411_, _03067_);
  and _35741_ (_03416_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _35742_ (_04058_, _03416_, _03415_);
  and _35743_ (_03417_, _03411_, _03071_);
  and _35744_ (_03418_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _35745_ (_04061_, _03418_, _03417_);
  and _35746_ (_03419_, _03411_, _03074_);
  and _35747_ (_03420_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _35748_ (_04064_, _03420_, _03419_);
  and _35749_ (_03421_, _03411_, _03077_);
  and _35750_ (_03422_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _35751_ (_04067_, _03422_, _03421_);
  and _35752_ (_03423_, _03411_, _03080_);
  and _35753_ (_03424_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _35754_ (_04070_, _03424_, _03423_);
  and _35755_ (_03425_, _03411_, _03083_);
  and _35756_ (_03426_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _35757_ (_04073_, _03426_, _03425_);
  and _35758_ (_03427_, _03411_, _03087_);
  and _35759_ (_03428_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _35760_ (_04076_, _03428_, _03427_);
  and _35761_ (_03429_, _03374_, _03113_);
  and _35762_ (_03430_, _03429_, _03060_);
  not _35763_ (_03431_, _03429_);
  and _35764_ (_03432_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or _35765_ (_04079_, _03432_, _03430_);
  and _35766_ (_03433_, _03429_, _03067_);
  and _35767_ (_03434_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or _35768_ (_04082_, _03434_, _03433_);
  and _35769_ (_03435_, _03429_, _03071_);
  and _35770_ (_03436_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or _35771_ (_04085_, _03436_, _03435_);
  and _35772_ (_03437_, _03429_, _03074_);
  and _35773_ (_03438_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or _35774_ (_04088_, _03438_, _03437_);
  and _35775_ (_03439_, _03429_, _03077_);
  and _35776_ (_03440_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or _35777_ (_04091_, _03440_, _03439_);
  and _35778_ (_03441_, _03429_, _03080_);
  and _35779_ (_03442_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or _35780_ (_04094_, _03442_, _03441_);
  and _35781_ (_03444_, _03429_, _03083_);
  and _35782_ (_03445_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or _35783_ (_04097_, _03445_, _03444_);
  and _35784_ (_03446_, _03429_, _03087_);
  and _35785_ (_03447_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or _35786_ (_04100_, _03447_, _03446_);
  and _35787_ (_03448_, _03374_, _03136_);
  and _35788_ (_03449_, _03448_, _03060_);
  not _35789_ (_03450_, _03448_);
  and _35790_ (_03451_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or _35791_ (_04104_, _03451_, _03449_);
  and _35792_ (_03452_, _03448_, _03067_);
  and _35793_ (_03453_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or _35794_ (_04107_, _03453_, _03452_);
  and _35795_ (_03454_, _03448_, _03071_);
  and _35796_ (_03455_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or _35797_ (_04110_, _03455_, _03454_);
  and _35798_ (_03456_, _03448_, _03074_);
  and _35799_ (_03457_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or _35800_ (_04113_, _03457_, _03456_);
  and _35801_ (_03458_, _03448_, _03077_);
  and _35802_ (_03459_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or _35803_ (_04116_, _03459_, _03458_);
  and _35804_ (_03460_, _03448_, _03080_);
  and _35805_ (_03461_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or _35806_ (_04119_, _03461_, _03460_);
  and _35807_ (_03462_, _03448_, _03083_);
  and _35808_ (_03463_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or _35809_ (_04122_, _03463_, _03462_);
  and _35810_ (_03464_, _03448_, _03087_);
  and _35811_ (_03465_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _35812_ (_04124_, _03465_, _03464_);
  and _35813_ (_03466_, _03374_, _03159_);
  and _35814_ (_03467_, _03466_, _03060_);
  not _35815_ (_03468_, _03466_);
  and _35816_ (_03469_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _35817_ (_04129_, _03469_, _03467_);
  and _35818_ (_03470_, _03466_, _03067_);
  and _35819_ (_03471_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _35820_ (_04132_, _03471_, _03470_);
  and _35821_ (_03472_, _03466_, _03071_);
  and _35822_ (_03473_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _35823_ (_04135_, _03473_, _03472_);
  and _35824_ (_03474_, _03466_, _03074_);
  and _35825_ (_03475_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _35826_ (_04138_, _03475_, _03474_);
  and _35827_ (_03476_, _03466_, _03077_);
  and _35828_ (_03477_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _35829_ (_04141_, _03477_, _03476_);
  and _35830_ (_03478_, _03466_, _03080_);
  and _35831_ (_03479_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _35832_ (_04144_, _03479_, _03478_);
  and _35833_ (_03480_, _03466_, _03083_);
  and _35834_ (_03481_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _35835_ (_04147_, _03481_, _03480_);
  and _35836_ (_03482_, _03466_, _03087_);
  and _35837_ (_03483_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _35838_ (_04150_, _03483_, _03482_);
  and _35839_ (_03484_, _03374_, _03179_);
  and _35840_ (_03485_, _03484_, _03060_);
  not _35841_ (_03486_, _03484_);
  and _35842_ (_03487_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _35843_ (_04153_, _03487_, _03485_);
  and _35844_ (_03488_, _03484_, _03067_);
  and _35845_ (_03489_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _35846_ (_04157_, _03489_, _03488_);
  and _35847_ (_03490_, _03484_, _03071_);
  and _35848_ (_03491_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _35849_ (_04160_, _03491_, _03490_);
  and _35850_ (_03492_, _03484_, _03074_);
  and _35851_ (_03493_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _35852_ (_04163_, _03493_, _03492_);
  and _35853_ (_03494_, _03484_, _03077_);
  and _35854_ (_03495_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _35855_ (_04166_, _03495_, _03494_);
  and _35856_ (_03496_, _03484_, _03080_);
  and _35857_ (_03497_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _35858_ (_04169_, _03497_, _03496_);
  and _35859_ (_03498_, _03484_, _03083_);
  and _35860_ (_03499_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _35861_ (_04172_, _03499_, _03498_);
  and _35862_ (_03500_, _03484_, _03087_);
  and _35863_ (_03501_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _35864_ (_04174_, _03501_, _03500_);
  and _35865_ (_03502_, _03374_, _03198_);
  and _35866_ (_03503_, _03502_, _03060_);
  not _35867_ (_03504_, _03502_);
  and _35868_ (_03505_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or _35869_ (_04178_, _03505_, _03503_);
  and _35870_ (_03506_, _03502_, _03067_);
  and _35871_ (_03507_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or _35872_ (_04181_, _03507_, _03506_);
  and _35873_ (_03508_, _03502_, _03071_);
  and _35874_ (_03509_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or _35875_ (_04185_, _03509_, _03508_);
  and _35876_ (_03510_, _03502_, _03074_);
  and _35877_ (_03511_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or _35878_ (_04188_, _03511_, _03510_);
  and _35879_ (_03512_, _03502_, _03077_);
  and _35880_ (_03513_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or _35881_ (_04192_, _03513_, _03512_);
  and _35882_ (_03514_, _03502_, _03080_);
  and _35883_ (_03515_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or _35884_ (_04195_, _03515_, _03514_);
  and _35885_ (_03516_, _03502_, _03083_);
  and _35886_ (_03517_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or _35887_ (_04198_, _03517_, _03516_);
  and _35888_ (_03518_, _03502_, _03087_);
  and _35889_ (_03519_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or _35890_ (_04200_, _03519_, _03518_);
  and _35891_ (_03520_, _03374_, _03218_);
  and _35892_ (_03521_, _03520_, _03060_);
  not _35893_ (_03522_, _03520_);
  and _35894_ (_03523_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _35895_ (_04204_, _03523_, _03521_);
  and _35896_ (_03524_, _03520_, _03067_);
  and _35897_ (_03525_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _35898_ (_04207_, _03525_, _03524_);
  and _35899_ (_03526_, _03520_, _03071_);
  and _35900_ (_03527_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _35901_ (_04210_, _03527_, _03526_);
  and _35902_ (_03528_, _03520_, _03074_);
  and _35903_ (_03529_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _35904_ (_04213_, _03529_, _03528_);
  and _35905_ (_03530_, _03520_, _03077_);
  and _35906_ (_03531_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _35907_ (_04216_, _03531_, _03530_);
  and _35908_ (_03532_, _03520_, _03080_);
  and _35909_ (_03533_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _35910_ (_04219_, _03533_, _03532_);
  and _35911_ (_03534_, _03520_, _03083_);
  and _35912_ (_03535_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _35913_ (_04222_, _03535_, _03534_);
  and _35914_ (_03536_, _03520_, _03087_);
  and _35915_ (_03537_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _35916_ (_04225_, _03537_, _03536_);
  and _35917_ (_03538_, _03374_, _03237_);
  and _35918_ (_03539_, _03538_, _03060_);
  not _35919_ (_03540_, _03538_);
  and _35920_ (_03541_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or _35921_ (_04228_, _03541_, _03539_);
  and _35922_ (_03542_, _03538_, _03067_);
  and _35923_ (_03543_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or _35924_ (_04231_, _03543_, _03542_);
  and _35925_ (_03544_, _03538_, _03071_);
  and _35926_ (_03545_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or _35927_ (_04234_, _03545_, _03544_);
  and _35928_ (_03546_, _03538_, _03074_);
  and _35929_ (_03547_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or _35930_ (_04238_, _03547_, _03546_);
  and _35931_ (_03548_, _03538_, _03077_);
  and _35932_ (_03549_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or _35933_ (_04241_, _03549_, _03548_);
  and _35934_ (_03550_, _03538_, _03080_);
  and _35935_ (_03551_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or _35936_ (_04244_, _03551_, _03550_);
  and _35937_ (_03552_, _03538_, _03083_);
  and _35938_ (_03553_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or _35939_ (_04247_, _03553_, _03552_);
  and _35940_ (_03554_, _03538_, _03087_);
  and _35941_ (_03555_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or _35942_ (_04249_, _03555_, _03554_);
  and _35943_ (_03556_, _03374_, _03256_);
  and _35944_ (_03557_, _03556_, _03060_);
  not _35945_ (_03558_, _03556_);
  and _35946_ (_03559_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or _35947_ (_04253_, _03559_, _03557_);
  and _35948_ (_03560_, _03556_, _03067_);
  and _35949_ (_03561_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or _35950_ (_04256_, _03561_, _03560_);
  and _35951_ (_03562_, _03556_, _03071_);
  and _35952_ (_03563_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or _35953_ (_04259_, _03563_, _03562_);
  and _35954_ (_03564_, _03556_, _03074_);
  and _35955_ (_03565_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or _35956_ (_04262_, _03565_, _03564_);
  and _35957_ (_03566_, _03556_, _03077_);
  and _35958_ (_03567_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or _35959_ (_04266_, _03567_, _03566_);
  and _35960_ (_03568_, _03556_, _03080_);
  and _35961_ (_03569_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or _35962_ (_04269_, _03569_, _03568_);
  and _35963_ (_03570_, _03556_, _03083_);
  and _35964_ (_03571_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or _35965_ (_04272_, _03571_, _03570_);
  and _35966_ (_03572_, _03556_, _03087_);
  and _35967_ (_03573_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or _35968_ (_04274_, _03573_, _03572_);
  and _35969_ (_03574_, _03374_, _03275_);
  and _35970_ (_03575_, _03574_, _03060_);
  not _35971_ (_03576_, _03574_);
  and _35972_ (_03578_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _35973_ (_04278_, _03578_, _03575_);
  and _35974_ (_03579_, _03574_, _03067_);
  and _35975_ (_03580_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _35976_ (_04281_, _03580_, _03579_);
  and _35977_ (_03582_, _03574_, _03071_);
  and _35978_ (_03583_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _35979_ (_04284_, _03583_, _03582_);
  and _35980_ (_03585_, _03574_, _03074_);
  and _35981_ (_03586_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _35982_ (_04287_, _03586_, _03585_);
  and _35983_ (_03588_, _03574_, _03077_);
  and _35984_ (_03589_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _35985_ (_04290_, _03589_, _03588_);
  and _35986_ (_03590_, _03574_, _03080_);
  and _35987_ (_03592_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _35988_ (_04294_, _03592_, _03590_);
  and _35989_ (_03593_, _03574_, _03083_);
  and _35990_ (_03594_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _35991_ (_04297_, _03594_, _03593_);
  and _35992_ (_03596_, _03574_, _03087_);
  and _35993_ (_03597_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _35994_ (_04300_, _03597_, _03596_);
  and _35995_ (_03598_, _03374_, _03295_);
  and _35996_ (_03599_, _03598_, _03060_);
  not _35997_ (_03601_, _03598_);
  and _35998_ (_03602_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _35999_ (_04303_, _03602_, _03599_);
  and _36000_ (_03603_, _03598_, _03067_);
  and _36001_ (_03604_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _36002_ (_04306_, _03604_, _03603_);
  and _36003_ (_03606_, _03598_, _03071_);
  and _36004_ (_03608_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _36005_ (_04309_, _03608_, _03606_);
  and _36006_ (_03609_, _03598_, _03074_);
  and _36007_ (_03610_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _36008_ (_04312_, _03610_, _03609_);
  and _36009_ (_03611_, _03598_, _03077_);
  and _36010_ (_03612_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _36011_ (_04315_, _03612_, _03611_);
  and _36012_ (_03614_, _03598_, _03080_);
  and _36013_ (_03615_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _36014_ (_04319_, _03615_, _03614_);
  and _36015_ (_03617_, _03598_, _03083_);
  and _36016_ (_03618_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _36017_ (_04322_, _03618_, _03617_);
  and _36018_ (_03620_, _03598_, _03087_);
  and _36019_ (_03621_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _36020_ (_04324_, _03621_, _03620_);
  and _36021_ (_03623_, _03374_, _03315_);
  and _36022_ (_03624_, _03623_, _03060_);
  not _36023_ (_03625_, _03623_);
  and _36024_ (_03627_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or _36025_ (_04328_, _03627_, _03624_);
  and _36026_ (_03628_, _03623_, _03067_);
  and _36027_ (_03630_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or _36028_ (_04331_, _03630_, _03628_);
  and _36029_ (_03631_, _03623_, _03071_);
  and _36030_ (_03633_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or _36031_ (_04334_, _03633_, _03631_);
  and _36032_ (_03635_, _03623_, _03074_);
  and _36033_ (_03636_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or _36034_ (_04337_, _03636_, _03635_);
  and _36035_ (_03637_, _03623_, _03077_);
  and _36036_ (_03638_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or _36037_ (_04340_, _03638_, _03637_);
  and _36038_ (_03639_, _03623_, _03080_);
  and _36039_ (_03640_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or _36040_ (_04343_, _03640_, _03639_);
  and _36041_ (_03642_, _03623_, _03083_);
  and _36042_ (_03643_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or _36043_ (_04347_, _03643_, _03642_);
  and _36044_ (_03645_, _03623_, _03087_);
  and _36045_ (_03646_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or _36046_ (_04349_, _03646_, _03645_);
  and _36047_ (_03648_, _03374_, _03334_);
  and _36048_ (_03649_, _03648_, _03060_);
  not _36049_ (_03651_, _03648_);
  and _36050_ (_03652_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or _36051_ (_04353_, _03652_, _03649_);
  and _36052_ (_03654_, _03648_, _03067_);
  and _36053_ (_03655_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or _36054_ (_04356_, _03655_, _03654_);
  and _36055_ (_03657_, _03648_, _03071_);
  and _36056_ (_03658_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or _36057_ (_04359_, _03658_, _03657_);
  and _36058_ (_03660_, _03648_, _03074_);
  and _36059_ (_03661_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or _36060_ (_04362_, _03661_, _03660_);
  and _36061_ (_03663_, _03648_, _03077_);
  and _36062_ (_03664_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or _36063_ (_04365_, _03664_, _03663_);
  and _36064_ (_03665_, _03648_, _03080_);
  and _36065_ (_03666_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or _36066_ (_04368_, _03666_, _03665_);
  and _36067_ (_03668_, _03648_, _03083_);
  and _36068_ (_03669_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or _36069_ (_04371_, _03669_, _03668_);
  and _36070_ (_03671_, _03648_, _03087_);
  and _36071_ (_03672_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or _36072_ (_04374_, _03672_, _03671_);
  and _36073_ (_03674_, _03374_, _03353_);
  and _36074_ (_03675_, _03674_, _03060_);
  not _36075_ (_03677_, _03674_);
  and _36076_ (_03678_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _36077_ (_04377_, _03678_, _03675_);
  and _36078_ (_03680_, _03674_, _03067_);
  and _36079_ (_03681_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _36080_ (_04380_, _03681_, _03680_);
  and _36081_ (_03683_, _03674_, _03071_);
  and _36082_ (_03684_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _36083_ (_04383_, _03684_, _03683_);
  and _36084_ (_03686_, _03674_, _03074_);
  and _36085_ (_03687_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _36086_ (_04386_, _03687_, _03686_);
  and _36087_ (_03689_, _03674_, _03077_);
  and _36088_ (_03690_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _36089_ (_04389_, _03690_, _03689_);
  and _36090_ (_03691_, _03674_, _03080_);
  and _36091_ (_03692_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _36092_ (_04392_, _03692_, _03691_);
  and _36093_ (_03693_, _03674_, _03083_);
  and _36094_ (_03695_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _36095_ (_04395_, _03695_, _03693_);
  and _36096_ (_03696_, _03674_, _03087_);
  and _36097_ (_03698_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _36098_ (_04399_, _03698_, _03696_);
  and _36099_ (_03699_, _02965_, _02064_);
  and _36100_ (_03701_, _03699_, _03372_);
  and _36101_ (_03702_, _03701_, _02963_);
  and _36102_ (_03703_, _03702_, _03060_);
  not _36103_ (_03705_, _03702_);
  and _36104_ (_03706_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _36105_ (_04406_, _03706_, _03703_);
  and _36106_ (_03708_, _03702_, _03067_);
  and _36107_ (_03709_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _36108_ (_04409_, _03709_, _03708_);
  and _36109_ (_03711_, _03702_, _03071_);
  and _36110_ (_03712_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _36111_ (_04412_, _03712_, _03711_);
  and _36112_ (_03714_, _03702_, _03074_);
  and _36113_ (_03715_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _36114_ (_04415_, _03715_, _03714_);
  and _36115_ (_03717_, _03702_, _03077_);
  and _36116_ (_03718_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _36117_ (_04418_, _03718_, _03717_);
  and _36118_ (_03719_, _03702_, _03080_);
  and _36119_ (_03721_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _36120_ (_04421_, _03721_, _03719_);
  and _36121_ (_03722_, _03702_, _03083_);
  and _36122_ (_03724_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _36123_ (_04424_, _03724_, _03722_);
  and _36124_ (_03725_, _03702_, _03087_);
  and _36125_ (_03727_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _36126_ (_04427_, _03727_, _03725_);
  and _36127_ (_03728_, _03701_, _03062_);
  and _36128_ (_03730_, _03728_, _03060_);
  not _36129_ (_03731_, _03728_);
  and _36130_ (_03732_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or _36131_ (_04430_, _03732_, _03730_);
  and _36132_ (_03734_, _03728_, _03067_);
  and _36133_ (_03735_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or _36134_ (_04433_, _03735_, _03734_);
  and _36135_ (_03737_, _03728_, _03071_);
  and _36136_ (_03738_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or _36137_ (_04436_, _03738_, _03737_);
  and _36138_ (_03740_, _03728_, _03074_);
  and _36139_ (_03742_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or _36140_ (_04439_, _03742_, _03740_);
  and _36141_ (_03743_, _03728_, _03077_);
  and _36142_ (_03744_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or _36143_ (_04442_, _03744_, _03743_);
  and _36144_ (_03746_, _03728_, _03080_);
  and _36145_ (_03747_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or _36146_ (_04445_, _03747_, _03746_);
  and _36147_ (_03749_, _03728_, _03083_);
  and _36148_ (_03750_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or _36149_ (_04448_, _03750_, _03749_);
  and _36150_ (_03752_, _03728_, _03087_);
  and _36151_ (_03753_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or _36152_ (_04451_, _03753_, _03752_);
  and _36153_ (_03755_, _03701_, _03091_);
  and _36154_ (_03756_, _03755_, _03060_);
  not _36155_ (_03757_, _03755_);
  and _36156_ (_03759_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or _36157_ (_04455_, _03759_, _03756_);
  and _36158_ (_03760_, _03755_, _03067_);
  and _36159_ (_03762_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or _36160_ (_04458_, _03762_, _03760_);
  and _36161_ (_03763_, _03755_, _03071_);
  and _36162_ (_03765_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or _36163_ (_04461_, _03765_, _03763_);
  and _36164_ (_03767_, _03755_, _03074_);
  and _36165_ (_03768_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or _36166_ (_04464_, _03768_, _03767_);
  and _36167_ (_03769_, _03755_, _03077_);
  and _36168_ (_03770_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or _36169_ (_04467_, _03770_, _03769_);
  and _36170_ (_03772_, _03755_, _03080_);
  and _36171_ (_03773_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or _36172_ (_04470_, _03773_, _03772_);
  and _36173_ (_03775_, _03755_, _03083_);
  and _36174_ (_03776_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or _36175_ (_04473_, _03776_, _03775_);
  and _36176_ (_03778_, _03755_, _03087_);
  and _36177_ (_03779_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or _36178_ (_04475_, _03779_, _03778_);
  and _36179_ (_03781_, _03701_, _03113_);
  and _36180_ (_03783_, _03781_, _03060_);
  not _36181_ (_03785_, _03781_);
  and _36182_ (_03786_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _36183_ (_04480_, _03786_, _03783_);
  and _36184_ (_03788_, _03781_, _03067_);
  and _36185_ (_03789_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _36186_ (_04483_, _03789_, _03788_);
  and _36187_ (_03791_, _03781_, _03071_);
  and _36188_ (_03792_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _36189_ (_04486_, _03792_, _03791_);
  and _36190_ (_03794_, _03781_, _03074_);
  and _36191_ (_03795_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _36192_ (_04489_, _03795_, _03794_);
  and _36193_ (_03796_, _03781_, _03077_);
  and _36194_ (_03797_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _36195_ (_04492_, _03797_, _03796_);
  and _36196_ (_03798_, _03781_, _03080_);
  and _36197_ (_03800_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _36198_ (_04495_, _03800_, _03798_);
  and _36199_ (_03801_, _03781_, _03083_);
  and _36200_ (_03803_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _36201_ (_04498_, _03803_, _03801_);
  and _36202_ (_03804_, _03781_, _03087_);
  and _36203_ (_03806_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _36204_ (_04501_, _03806_, _03804_);
  and _36205_ (_03807_, _03701_, _03136_);
  and _36206_ (_03809_, _03807_, _03060_);
  not _36207_ (_03810_, _03807_);
  and _36208_ (_03811_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _36209_ (_04505_, _03811_, _03809_);
  and _36210_ (_03813_, _03807_, _03067_);
  and _36211_ (_03814_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _36212_ (_04508_, _03814_, _03813_);
  and _36213_ (_03816_, _03807_, _03071_);
  and _36214_ (_03817_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _36215_ (_04511_, _03817_, _03816_);
  and _36216_ (_03819_, _03807_, _03074_);
  and _36217_ (_03821_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _36218_ (_04514_, _03821_, _03819_);
  and _36219_ (_03822_, _03807_, _03077_);
  and _36220_ (_03823_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _36221_ (_04517_, _03823_, _03822_);
  and _36222_ (_03825_, _03807_, _03080_);
  and _36223_ (_03826_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _36224_ (_04520_, _03826_, _03825_);
  and _36225_ (_03828_, _03807_, _03083_);
  and _36226_ (_03829_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _36227_ (_04523_, _03829_, _03828_);
  and _36228_ (_03831_, _03807_, _03087_);
  and _36229_ (_03832_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _36230_ (_04526_, _03832_, _03831_);
  and _36231_ (_03834_, _03701_, _03159_);
  and _36232_ (_03835_, _03834_, _03060_);
  not _36233_ (_03836_, _03834_);
  and _36234_ (_03838_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or _36235_ (_04529_, _03838_, _03835_);
  and _36236_ (_03839_, _03834_, _03067_);
  and _36237_ (_03841_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or _36238_ (_04533_, _03841_, _03839_);
  and _36239_ (_03842_, _03834_, _03071_);
  and _36240_ (_03844_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or _36241_ (_04536_, _03844_, _03842_);
  and _36242_ (_03846_, _03834_, _03074_);
  and _36243_ (_03847_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or _36244_ (_04539_, _03847_, _03846_);
  and _36245_ (_03848_, _03834_, _03077_);
  and _36246_ (_03849_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or _36247_ (_04542_, _03849_, _03848_);
  and _36248_ (_03851_, _03834_, _03080_);
  and _36249_ (_03852_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or _36250_ (_04545_, _03852_, _03851_);
  and _36251_ (_03854_, _03834_, _03083_);
  and _36252_ (_03855_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or _36253_ (_04548_, _03855_, _03854_);
  and _36254_ (_03857_, _03834_, _03087_);
  and _36255_ (_03858_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or _36256_ (_04550_, _03858_, _03857_);
  and _36257_ (_03860_, _03701_, _03179_);
  and _36258_ (_03861_, _03860_, _03060_);
  not _36259_ (_03863_, _03860_);
  and _36260_ (_03864_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or _36261_ (_04554_, _03864_, _03861_);
  and _36262_ (_03866_, _03860_, _03067_);
  and _36263_ (_03867_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or _36264_ (_04557_, _03867_, _03866_);
  and _36265_ (_03869_, _03860_, _03071_);
  and _36266_ (_03870_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or _36267_ (_04561_, _03870_, _03869_);
  and _36268_ (_03872_, _03860_, _03074_);
  and _36269_ (_03873_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or _36270_ (_04565_, _03873_, _03872_);
  and _36271_ (_03874_, _03860_, _03077_);
  and _36272_ (_03876_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or _36273_ (_04568_, _03876_, _03874_);
  and _36274_ (_03877_, _03860_, _03080_);
  and _36275_ (_03879_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or _36276_ (_04571_, _03879_, _03877_);
  and _36277_ (_03880_, _03860_, _03083_);
  and _36278_ (_03882_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or _36279_ (_04574_, _03882_, _03880_);
  and _36280_ (_03883_, _03860_, _03087_);
  and _36281_ (_03885_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or _36282_ (_04576_, _03885_, _03883_);
  and _36283_ (_03886_, _03701_, _03198_);
  and _36284_ (_03888_, _03886_, _03060_);
  not _36285_ (_03889_, _03886_);
  and _36286_ (_03890_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _36287_ (_04580_, _03890_, _03888_);
  and _36288_ (_03892_, _03886_, _03067_);
  and _36289_ (_03893_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _36290_ (_04583_, _03893_, _03892_);
  and _36291_ (_03895_, _03886_, _03071_);
  and _36292_ (_03897_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _36293_ (_04586_, _03897_, _03895_);
  and _36294_ (_03898_, _03886_, _03074_);
  and _36295_ (_03899_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _36296_ (_04589_, _03899_, _03898_);
  and _36297_ (_03900_, _03886_, _03077_);
  and _36298_ (_03902_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _36299_ (_04592_, _03902_, _03900_);
  and _36300_ (_03903_, _03886_, _03080_);
  and _36301_ (_03905_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _36302_ (_04595_, _03905_, _03903_);
  and _36303_ (_03906_, _03886_, _03083_);
  and _36304_ (_03908_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _36305_ (_04598_, _03908_, _03906_);
  and _36306_ (_03909_, _03886_, _03087_);
  and _36307_ (_03911_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _36308_ (_04601_, _03911_, _03909_);
  and _36309_ (_03912_, _03701_, _03218_);
  and _36310_ (_03914_, _03912_, _03060_);
  not _36311_ (_03915_, _03912_);
  and _36312_ (_03916_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or _36313_ (_04605_, _03916_, _03914_);
  and _36314_ (_03918_, _03912_, _03067_);
  and _36315_ (_03919_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or _36316_ (_04608_, _03919_, _03918_);
  and _36317_ (_03921_, _03912_, _03071_);
  and _36318_ (_03923_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or _36319_ (_04611_, _03923_, _03921_);
  and _36320_ (_03924_, _03912_, _03074_);
  and _36321_ (_03925_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or _36322_ (_04614_, _03925_, _03924_);
  and _36323_ (_03927_, _03912_, _03077_);
  and _36324_ (_03928_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or _36325_ (_04618_, _03928_, _03927_);
  and _36326_ (_03930_, _03912_, _03080_);
  and _36327_ (_03931_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or _36328_ (_04621_, _03931_, _03930_);
  and _36329_ (_03933_, _03912_, _03083_);
  and _36330_ (_03934_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or _36331_ (_04624_, _03934_, _03933_);
  and _36332_ (_03936_, _03912_, _03087_);
  and _36333_ (_03937_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or _36334_ (_04626_, _03937_, _03936_);
  and _36335_ (_03939_, _03701_, _03237_);
  and _36336_ (_03940_, _03939_, _03060_);
  not _36337_ (_03941_, _03939_);
  and _36338_ (_03943_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _36339_ (_04630_, _03943_, _03940_);
  and _36340_ (_03944_, _03939_, _03067_);
  and _36341_ (_03946_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _36342_ (_04633_, _03946_, _03944_);
  and _36343_ (_03948_, _03939_, _03071_);
  and _36344_ (_03949_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _36345_ (_04636_, _03949_, _03948_);
  and _36346_ (_03950_, _03939_, _03074_);
  and _36347_ (_03951_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _36348_ (_04639_, _03951_, _03950_);
  and _36349_ (_03953_, _03939_, _03077_);
  and _36350_ (_03954_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _36351_ (_04642_, _03954_, _03953_);
  and _36352_ (_03956_, _03939_, _03080_);
  and _36353_ (_03957_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _36354_ (_04646_, _03957_, _03956_);
  and _36355_ (_03959_, _03939_, _03083_);
  and _36356_ (_03960_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _36357_ (_04649_, _03960_, _03959_);
  and _36358_ (_03962_, _03939_, _03087_);
  and _36359_ (_03963_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _36360_ (_04651_, _03963_, _03962_);
  and _36361_ (_03965_, _03701_, _03256_);
  and _36362_ (_03966_, _03965_, _03060_);
  not _36363_ (_03968_, _03965_);
  and _36364_ (_03969_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _36365_ (_04655_, _03969_, _03966_);
  and _36366_ (_03971_, _03965_, _03067_);
  and _36367_ (_03972_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _36368_ (_04658_, _03972_, _03971_);
  and _36369_ (_03974_, _03965_, _03071_);
  and _36370_ (_03975_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _36371_ (_04661_, _03975_, _03974_);
  and _36372_ (_03976_, _03965_, _03074_);
  and _36373_ (_03978_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _36374_ (_04664_, _03978_, _03976_);
  and _36375_ (_03979_, _03965_, _03077_);
  and _36376_ (_03981_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _36377_ (_04667_, _03981_, _03979_);
  and _36378_ (_03982_, _03965_, _03080_);
  and _36379_ (_03984_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _36380_ (_04670_, _03984_, _03982_);
  and _36381_ (_03986_, _03965_, _03083_);
  and _36382_ (_03988_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _36383_ (_04673_, _03988_, _03986_);
  and _36384_ (_03989_, _03965_, _03087_);
  and _36385_ (_03991_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _36386_ (_04676_, _03991_, _03989_);
  and _36387_ (_03992_, _03701_, _03275_);
  and _36388_ (_03994_, _03992_, _03060_);
  not _36389_ (_03995_, _03992_);
  and _36390_ (_03996_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or _36391_ (_04679_, _03996_, _03994_);
  and _36392_ (_03998_, _03992_, _03067_);
  and _36393_ (_04000_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or _36394_ (_04682_, _04000_, _03998_);
  and _36395_ (_04001_, _03992_, _03071_);
  and _36396_ (_04002_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or _36397_ (_04685_, _04002_, _04001_);
  and _36398_ (_04003_, _03992_, _03074_);
  and _36399_ (_04004_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or _36400_ (_04688_, _04004_, _04003_);
  and _36401_ (_04006_, _03992_, _03077_);
  and _36402_ (_04007_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or _36403_ (_04691_, _04007_, _04006_);
  and _36404_ (_04009_, _03992_, _03080_);
  and _36405_ (_04010_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _36406_ (_04694_, _04010_, _04009_);
  and _36407_ (_04012_, _03992_, _03083_);
  and _36408_ (_04013_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or _36409_ (_04698_, _04013_, _04012_);
  and _36410_ (_04015_, _03992_, _03087_);
  and _36411_ (_04016_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or _36412_ (_04700_, _04016_, _04015_);
  and _36413_ (_04018_, _03701_, _03295_);
  and _36414_ (_04019_, _04018_, _03060_);
  not _36415_ (_04020_, _04018_);
  and _36416_ (_04022_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or _36417_ (_04704_, _04022_, _04019_);
  and _36418_ (_04023_, _04018_, _03067_);
  and _36419_ (_04025_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or _36420_ (_04708_, _04025_, _04023_);
  and _36421_ (_04027_, _04018_, _03071_);
  and _36422_ (_04028_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or _36423_ (_04711_, _04028_, _04027_);
  and _36424_ (_04029_, _04018_, _03074_);
  and _36425_ (_04031_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or _36426_ (_04714_, _04031_, _04029_);
  and _36427_ (_04032_, _04018_, _03077_);
  and _36428_ (_04034_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or _36429_ (_04717_, _04034_, _04032_);
  and _36430_ (_04035_, _04018_, _03080_);
  and _36431_ (_04037_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or _36432_ (_04720_, _04037_, _04035_);
  and _36433_ (_04038_, _04018_, _03083_);
  and _36434_ (_04040_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or _36435_ (_04723_, _04040_, _04038_);
  and _36436_ (_04041_, _04018_, _03087_);
  and _36437_ (_04043_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _36438_ (_04726_, _04043_, _04041_);
  and _36439_ (_04044_, _03701_, _03315_);
  and _36440_ (_04046_, _04044_, _03060_);
  not _36441_ (_04047_, _04044_);
  and _36442_ (_04048_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _36443_ (_04730_, _04048_, _04046_);
  and _36444_ (_04050_, _04044_, _03067_);
  and _36445_ (_04052_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _36446_ (_04733_, _04052_, _04050_);
  and _36447_ (_04053_, _04044_, _03071_);
  and _36448_ (_04054_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _36449_ (_04736_, _04054_, _04053_);
  and _36450_ (_04056_, _04044_, _03074_);
  and _36451_ (_04057_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _36452_ (_04739_, _04057_, _04056_);
  and _36453_ (_04059_, _04044_, _03077_);
  and _36454_ (_04060_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _36455_ (_04742_, _04060_, _04059_);
  and _36456_ (_04062_, _04044_, _03080_);
  and _36457_ (_04063_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _36458_ (_04745_, _04063_, _04062_);
  and _36459_ (_04065_, _04044_, _03083_);
  and _36460_ (_04066_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _36461_ (_04748_, _04066_, _04065_);
  and _36462_ (_04068_, _04044_, _03087_);
  and _36463_ (_04069_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _36464_ (_04750_, _04069_, _04068_);
  and _36465_ (_04071_, _03701_, _03334_);
  and _36466_ (_04072_, _04071_, _03060_);
  not _36467_ (_04074_, _04071_);
  and _36468_ (_04075_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _36469_ (_04754_, _04075_, _04072_);
  and _36470_ (_04077_, _04071_, _03067_);
  and _36471_ (_04078_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _36472_ (_04757_, _04078_, _04077_);
  and _36473_ (_04080_, _04071_, _03071_);
  and _36474_ (_04081_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _36475_ (_04760_, _04081_, _04080_);
  and _36476_ (_04083_, _04071_, _03074_);
  and _36477_ (_04084_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _36478_ (_04763_, _04084_, _04083_);
  and _36479_ (_04086_, _04071_, _03077_);
  and _36480_ (_04087_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _36481_ (_04766_, _04087_, _04086_);
  and _36482_ (_04089_, _04071_, _03080_);
  and _36483_ (_04090_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _36484_ (_04769_, _04090_, _04089_);
  and _36485_ (_04092_, _04071_, _03083_);
  and _36486_ (_04093_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _36487_ (_04772_, _04093_, _04092_);
  and _36488_ (_04095_, _04071_, _03087_);
  and _36489_ (_04096_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _36490_ (_04775_, _04096_, _04095_);
  and _36491_ (_04098_, _03701_, _03353_);
  and _36492_ (_04099_, _04098_, _03060_);
  not _36493_ (_04101_, _04098_);
  and _36494_ (_04102_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or _36495_ (_04779_, _04102_, _04099_);
  and _36496_ (_04103_, _04098_, _03067_);
  and _36497_ (_04105_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or _36498_ (_04782_, _04105_, _04103_);
  and _36499_ (_04106_, _04098_, _03071_);
  and _36500_ (_04108_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or _36501_ (_04785_, _04108_, _04106_);
  and _36502_ (_04109_, _04098_, _03074_);
  and _36503_ (_04111_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or _36504_ (_04788_, _04111_, _04109_);
  and _36505_ (_04112_, _04098_, _03077_);
  and _36506_ (_04114_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or _36507_ (_04791_, _04114_, _04112_);
  and _36508_ (_04115_, _04098_, _03080_);
  and _36509_ (_04117_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _36510_ (_04794_, _04117_, _04115_);
  and _36511_ (_04118_, _04098_, _03083_);
  and _36512_ (_04120_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or _36513_ (_04797_, _04120_, _04118_);
  and _36514_ (_04121_, _04098_, _03087_);
  and _36515_ (_04123_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _36516_ (_04799_, _04123_, _04121_);
  and _36517_ (_04125_, _02965_, _02964_);
  and _36518_ (_04126_, _04125_, _03372_);
  and _36519_ (_04127_, _04126_, _02963_);
  and _36520_ (_04128_, _04127_, _03060_);
  not _36521_ (_04130_, _04127_);
  and _36522_ (_04131_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or _36523_ (_04805_, _04131_, _04128_);
  and _36524_ (_04133_, _04127_, _03067_);
  and _36525_ (_04134_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or _36526_ (_04808_, _04134_, _04133_);
  and _36527_ (_04136_, _04127_, _03071_);
  and _36528_ (_04137_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or _36529_ (_04812_, _04137_, _04136_);
  and _36530_ (_04139_, _04127_, _03074_);
  and _36531_ (_04140_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or _36532_ (_04815_, _04140_, _04139_);
  and _36533_ (_04142_, _04127_, _03077_);
  and _36534_ (_04143_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or _36535_ (_04818_, _04143_, _04142_);
  and _36536_ (_04145_, _04127_, _03080_);
  and _36537_ (_04146_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or _36538_ (_04821_, _04146_, _04145_);
  and _36539_ (_04148_, _04127_, _03083_);
  and _36540_ (_04149_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or _36541_ (_04824_, _04149_, _04148_);
  and _36542_ (_04151_, _04127_, _03087_);
  and _36543_ (_04152_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or _36544_ (_04826_, _04152_, _04151_);
  and _36545_ (_04154_, _04126_, _03062_);
  and _36546_ (_04155_, _04154_, _03060_);
  not _36547_ (_04156_, _04154_);
  and _36548_ (_04158_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _36549_ (_04830_, _04158_, _04155_);
  and _36550_ (_04159_, _04154_, _03067_);
  and _36551_ (_04161_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _36552_ (_04834_, _04161_, _04159_);
  and _36553_ (_04162_, _04154_, _03071_);
  and _36554_ (_04164_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _36555_ (_04837_, _04164_, _04162_);
  and _36556_ (_04165_, _04154_, _03074_);
  and _36557_ (_04167_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _36558_ (_04840_, _04167_, _04165_);
  and _36559_ (_04168_, _04154_, _03077_);
  and _36560_ (_04170_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _36561_ (_04843_, _04170_, _04168_);
  and _36562_ (_04171_, _04154_, _03080_);
  and _36563_ (_04173_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _36564_ (_04846_, _04173_, _04171_);
  and _36565_ (_04175_, _04154_, _03083_);
  and _36566_ (_04176_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _36567_ (_04849_, _04176_, _04175_);
  and _36568_ (_04177_, _04154_, _03087_);
  and _36569_ (_04179_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _36570_ (_04851_, _04179_, _04177_);
  and _36571_ (_04180_, _04126_, _03091_);
  and _36572_ (_04182_, _04180_, _03060_);
  not _36573_ (_04183_, _04180_);
  and _36574_ (_04184_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _36575_ (_04855_, _04184_, _04182_);
  and _36576_ (_04186_, _04180_, _03067_);
  and _36577_ (_04187_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _36578_ (_04858_, _04187_, _04186_);
  and _36579_ (_04189_, _04180_, _03071_);
  and _36580_ (_04191_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _36581_ (_04861_, _04191_, _04189_);
  and _36582_ (_04193_, _04180_, _03074_);
  and _36583_ (_04194_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _36584_ (_04864_, _04194_, _04193_);
  and _36585_ (_04196_, _04180_, _03077_);
  and _36586_ (_04197_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _36587_ (_04867_, _04197_, _04196_);
  and _36588_ (_04199_, _04180_, _03080_);
  and _36589_ (_04201_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _36590_ (_04870_, _04201_, _04199_);
  and _36591_ (_04202_, _04180_, _03083_);
  and _36592_ (_04203_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _36593_ (_04873_, _04203_, _04202_);
  and _36594_ (_04205_, _04180_, _03087_);
  and _36595_ (_04206_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _36596_ (_04876_, _04206_, _04205_);
  and _36597_ (_04208_, _04126_, _03113_);
  and _36598_ (_04209_, _04208_, _03060_);
  not _36599_ (_04211_, _04208_);
  and _36600_ (_04212_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or _36601_ (_04879_, _04212_, _04209_);
  and _36602_ (_04214_, _04208_, _03067_);
  and _36603_ (_04215_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or _36604_ (_04882_, _04215_, _04214_);
  and _36605_ (_04217_, _04208_, _03071_);
  and _36606_ (_04218_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or _36607_ (_04886_, _04218_, _04217_);
  and _36608_ (_04220_, _04208_, _03074_);
  and _36609_ (_04221_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or _36610_ (_04889_, _04221_, _04220_);
  and _36611_ (_04223_, _04208_, _03077_);
  and _36612_ (_04224_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or _36613_ (_04892_, _04224_, _04223_);
  and _36614_ (_04226_, _04208_, _03080_);
  and _36615_ (_04227_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or _36616_ (_04895_, _04227_, _04226_);
  and _36617_ (_04229_, _04208_, _03083_);
  and _36618_ (_04230_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or _36619_ (_04898_, _04230_, _04229_);
  and _36620_ (_04232_, _04208_, _03087_);
  and _36621_ (_04233_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or _36622_ (_04900_, _04233_, _04232_);
  and _36623_ (_04235_, _04126_, _03136_);
  and _36624_ (_04236_, _04235_, _03060_);
  not _36625_ (_04237_, _04235_);
  and _36626_ (_04239_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or _36627_ (_04904_, _04239_, _04236_);
  and _36628_ (_04240_, _04235_, _03067_);
  and _36629_ (_04242_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or _36630_ (_04907_, _04242_, _04240_);
  and _36631_ (_04243_, _04235_, _03071_);
  and _36632_ (_04245_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or _36633_ (_04910_, _04245_, _04243_);
  and _36634_ (_04246_, _04235_, _03074_);
  and _36635_ (_04248_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or _36636_ (_04915_, _04248_, _04246_);
  and _36637_ (_04250_, _04235_, _03077_);
  and _36638_ (_04251_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or _36639_ (_04918_, _04251_, _04250_);
  and _36640_ (_04252_, _04235_, _03080_);
  and _36641_ (_04254_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or _36642_ (_04921_, _04254_, _04252_);
  and _36643_ (_04255_, _04235_, _03083_);
  and _36644_ (_04257_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or _36645_ (_04924_, _04257_, _04255_);
  and _36646_ (_04258_, _04235_, _03087_);
  and _36647_ (_04260_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _36648_ (_04926_, _04260_, _04258_);
  and _36649_ (_04261_, _04126_, _03159_);
  and _36650_ (_04263_, _04261_, _03060_);
  not _36651_ (_04264_, _04261_);
  and _36652_ (_04265_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _36653_ (_04930_, _04265_, _04263_);
  and _36654_ (_04267_, _04261_, _03067_);
  and _36655_ (_04268_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _36656_ (_04933_, _04268_, _04267_);
  and _36657_ (_04270_, _04261_, _03071_);
  and _36658_ (_04271_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _36659_ (_04936_, _04271_, _04270_);
  and _36660_ (_04273_, _04261_, _03074_);
  and _36661_ (_04275_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _36662_ (_04939_, _04275_, _04273_);
  and _36663_ (_04276_, _04261_, _03077_);
  and _36664_ (_04277_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _36665_ (_04942_, _04277_, _04276_);
  and _36666_ (_04279_, _04261_, _03080_);
  and _36667_ (_04280_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _36668_ (_04945_, _04280_, _04279_);
  and _36669_ (_04282_, _04261_, _03083_);
  and _36670_ (_04283_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _36671_ (_04948_, _04283_, _04282_);
  and _36672_ (_04285_, _04261_, _03087_);
  and _36673_ (_04286_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _36674_ (_04951_, _04286_, _04285_);
  and _36675_ (_04288_, _04126_, _03179_);
  and _36676_ (_04289_, _04288_, _03060_);
  not _36677_ (_04291_, _04288_);
  and _36678_ (_04292_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _36679_ (_04954_, _04292_, _04289_);
  and _36680_ (_04295_, _04288_, _03067_);
  and _36681_ (_04296_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _36682_ (_04957_, _04296_, _04295_);
  and _36683_ (_04298_, _04288_, _03071_);
  and _36684_ (_04299_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _36685_ (_04960_, _04299_, _04298_);
  and _36686_ (_04301_, _04288_, _03074_);
  and _36687_ (_04302_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _36688_ (_04963_, _04302_, _04301_);
  and _36689_ (_04304_, _04288_, _03077_);
  and _36690_ (_04305_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _36691_ (_04967_, _04305_, _04304_);
  and _36692_ (_04307_, _04288_, _03080_);
  and _36693_ (_04308_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _36694_ (_04970_, _04308_, _04307_);
  and _36695_ (_04310_, _04288_, _03083_);
  and _36696_ (_04311_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _36697_ (_04973_, _04311_, _04310_);
  and _36698_ (_04313_, _04288_, _03087_);
  and _36699_ (_04314_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _36700_ (_04975_, _04314_, _04313_);
  and _36701_ (_04316_, _04126_, _03198_);
  and _36702_ (_04317_, _04316_, _03060_);
  not _36703_ (_04318_, _04316_);
  and _36704_ (_04320_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or _36705_ (_04979_, _04320_, _04317_);
  and _36706_ (_04321_, _04316_, _03067_);
  and _36707_ (_04323_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or _36708_ (_04982_, _04323_, _04321_);
  and _36709_ (_04325_, _04316_, _03071_);
  and _36710_ (_04326_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or _36711_ (_04985_, _04326_, _04325_);
  and _36712_ (_04327_, _04316_, _03074_);
  and _36713_ (_04329_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or _36714_ (_04988_, _04329_, _04327_);
  and _36715_ (_04330_, _04316_, _03077_);
  and _36716_ (_04332_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or _36717_ (_04991_, _04332_, _04330_);
  and _36718_ (_04333_, _04316_, _03080_);
  and _36719_ (_04335_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or _36720_ (_04995_, _04335_, _04333_);
  and _36721_ (_04336_, _04316_, _03083_);
  and _36722_ (_04338_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or _36723_ (_04998_, _04338_, _04336_);
  and _36724_ (_04339_, _04316_, _03087_);
  and _36725_ (_04341_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or _36726_ (_05000_, _04341_, _04339_);
  and _36727_ (_04342_, _04126_, _03218_);
  and _36728_ (_04344_, _04342_, _03060_);
  not _36729_ (_04345_, _04342_);
  and _36730_ (_04346_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _36731_ (_05004_, _04346_, _04344_);
  and _36732_ (_04348_, _04342_, _03067_);
  and _36733_ (_04350_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _36734_ (_05007_, _04350_, _04348_);
  and _36735_ (_04351_, _04342_, _03071_);
  and _36736_ (_04352_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _36737_ (_05010_, _04352_, _04351_);
  and _36738_ (_04354_, _04342_, _03074_);
  and _36739_ (_04355_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _36740_ (_05013_, _04355_, _04354_);
  and _36741_ (_04357_, _04342_, _03077_);
  and _36742_ (_04358_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _36743_ (_05016_, _04358_, _04357_);
  and _36744_ (_04360_, _04342_, _03080_);
  and _36745_ (_04361_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _36746_ (_05019_, _04361_, _04360_);
  and _36747_ (_04363_, _04342_, _03083_);
  and _36748_ (_04364_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _36749_ (_05023_, _04364_, _04363_);
  and _36750_ (_04366_, _04342_, _03087_);
  and _36751_ (_04367_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _36752_ (_05025_, _04367_, _04366_);
  and _36753_ (_04369_, _04126_, _03237_);
  and _36754_ (_04370_, _04369_, _03060_);
  not _36755_ (_04372_, _04369_);
  and _36756_ (_04373_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or _36757_ (_05029_, _04373_, _04370_);
  and _36758_ (_04375_, _04369_, _03067_);
  and _36759_ (_04376_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or _36760_ (_05032_, _04376_, _04375_);
  and _36761_ (_04378_, _04369_, _03071_);
  and _36762_ (_04379_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or _36763_ (_05035_, _04379_, _04378_);
  and _36764_ (_04381_, _04369_, _03074_);
  and _36765_ (_04382_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or _36766_ (_05038_, _04382_, _04381_);
  and _36767_ (_04384_, _04369_, _03077_);
  and _36768_ (_04385_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or _36769_ (_05041_, _04385_, _04384_);
  and _36770_ (_04387_, _04369_, _03080_);
  and _36771_ (_04388_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or _36772_ (_05044_, _04388_, _04387_);
  and _36773_ (_04390_, _04369_, _03083_);
  and _36774_ (_04391_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or _36775_ (_05047_, _04391_, _04390_);
  and _36776_ (_04393_, _04369_, _03087_);
  and _36777_ (_04394_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or _36778_ (_05050_, _04394_, _04393_);
  and _36779_ (_04396_, _04126_, _03256_);
  and _36780_ (_04398_, _04396_, _03060_);
  not _36781_ (_04400_, _04396_);
  and _36782_ (_04401_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or _36783_ (_05053_, _04401_, _04398_);
  and _36784_ (_04402_, _04396_, _03067_);
  and _36785_ (_04403_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or _36786_ (_05056_, _04403_, _04402_);
  and _36787_ (_04404_, _04396_, _03071_);
  and _36788_ (_04405_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or _36789_ (_05059_, _04405_, _04404_);
  and _36790_ (_04407_, _04396_, _03074_);
  and _36791_ (_04408_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or _36792_ (_05062_, _04408_, _04407_);
  and _36793_ (_04410_, _04396_, _03077_);
  and _36794_ (_04411_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or _36795_ (_05065_, _04411_, _04410_);
  and _36796_ (_04413_, _04396_, _03080_);
  and _36797_ (_04414_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or _36798_ (_05068_, _04414_, _04413_);
  and _36799_ (_04416_, _04396_, _03083_);
  and _36800_ (_04417_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or _36801_ (_05071_, _04417_, _04416_);
  and _36802_ (_04419_, _04396_, _03087_);
  and _36803_ (_04420_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or _36804_ (_05074_, _04420_, _04419_);
  and _36805_ (_04422_, _04126_, _03275_);
  and _36806_ (_04423_, _04422_, _03060_);
  not _36807_ (_04425_, _04422_);
  and _36808_ (_04426_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _36809_ (_05078_, _04426_, _04423_);
  and _36810_ (_04428_, _04422_, _03067_);
  and _36811_ (_04429_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _36812_ (_05081_, _04429_, _04428_);
  and _36813_ (_04431_, _04422_, _03071_);
  and _36814_ (_04432_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _36815_ (_05084_, _04432_, _04431_);
  and _36816_ (_04434_, _04422_, _03074_);
  and _36817_ (_04435_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _36818_ (_05087_, _04435_, _04434_);
  and _36819_ (_04437_, _04422_, _03077_);
  and _36820_ (_04438_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _36821_ (_05090_, _04438_, _04437_);
  and _36822_ (_04440_, _04422_, _03080_);
  and _36823_ (_04441_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _36824_ (_05093_, _04441_, _04440_);
  and _36825_ (_04443_, _04422_, _03083_);
  and _36826_ (_04444_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _36827_ (_05096_, _04444_, _04443_);
  and _36828_ (_04446_, _04422_, _03087_);
  and _36829_ (_04447_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _36830_ (_05098_, _04447_, _04446_);
  and _36831_ (_04449_, _04126_, _03295_);
  and _36832_ (_04450_, _04449_, _03060_);
  not _36833_ (_04452_, _04449_);
  and _36834_ (_04453_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _36835_ (_05103_, _04453_, _04450_);
  and _36836_ (_04454_, _04449_, _03067_);
  and _36837_ (_04456_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _36838_ (_05106_, _04456_, _04454_);
  and _36839_ (_04457_, _04449_, _03071_);
  and _36840_ (_04459_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _36841_ (_05109_, _04459_, _04457_);
  and _36842_ (_04460_, _04449_, _03074_);
  and _36843_ (_04462_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _36844_ (_05112_, _04462_, _04460_);
  and _36845_ (_04463_, _04449_, _03077_);
  and _36846_ (_04465_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _36847_ (_05115_, _04465_, _04463_);
  and _36848_ (_04466_, _04449_, _03080_);
  and _36849_ (_04468_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _36850_ (_05118_, _04468_, _04466_);
  and _36851_ (_04469_, _04449_, _03083_);
  and _36852_ (_04471_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _36853_ (_05121_, _04471_, _04469_);
  and _36854_ (_04472_, _04449_, _03087_);
  and _36855_ (_04474_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _36856_ (_05123_, _04474_, _04472_);
  and _36857_ (_04476_, _04126_, _03315_);
  and _36858_ (_04477_, _04476_, _03060_);
  not _36859_ (_04478_, _04476_);
  and _36860_ (_04479_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or _36861_ (_05127_, _04479_, _04477_);
  and _36862_ (_04481_, _04476_, _03067_);
  and _36863_ (_04482_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or _36864_ (_05130_, _04482_, _04481_);
  and _36865_ (_04484_, _04476_, _03071_);
  and _36866_ (_04485_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or _36867_ (_05133_, _04485_, _04484_);
  and _36868_ (_04487_, _04476_, _03074_);
  and _36869_ (_04488_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or _36870_ (_05136_, _04488_, _04487_);
  and _36871_ (_04490_, _04476_, _03077_);
  and _36872_ (_04491_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or _36873_ (_05139_, _04491_, _04490_);
  and _36874_ (_04493_, _04476_, _03080_);
  and _36875_ (_04494_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or _36876_ (_05142_, _04494_, _04493_);
  and _36877_ (_04496_, _04476_, _03083_);
  and _36878_ (_04497_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or _36879_ (_05145_, _04497_, _04496_);
  and _36880_ (_04500_, _04476_, _03087_);
  and _36881_ (_04502_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or _36882_ (_05148_, _04502_, _04500_);
  and _36883_ (_04503_, _04126_, _03334_);
  and _36884_ (_04504_, _04503_, _03060_);
  not _36885_ (_04506_, _04503_);
  and _36886_ (_04507_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or _36887_ (_05151_, _04507_, _04504_);
  and _36888_ (_04509_, _04503_, _03067_);
  and _36889_ (_04510_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or _36890_ (_05155_, _04510_, _04509_);
  and _36891_ (_04512_, _04503_, _03071_);
  and _36892_ (_04513_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or _36893_ (_05158_, _04513_, _04512_);
  and _36894_ (_04515_, _04503_, _03074_);
  and _36895_ (_04516_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or _36896_ (_05161_, _04516_, _04515_);
  and _36897_ (_04518_, _04503_, _03077_);
  and _36898_ (_04519_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or _36899_ (_05164_, _04519_, _04518_);
  and _36900_ (_04521_, _04503_, _03080_);
  and _36901_ (_04522_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or _36902_ (_05167_, _04522_, _04521_);
  and _36903_ (_04524_, _04503_, _03083_);
  and _36904_ (_04525_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or _36905_ (_05170_, _04525_, _04524_);
  and _36906_ (_04527_, _04503_, _03087_);
  and _36907_ (_04528_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or _36908_ (_05172_, _04528_, _04527_);
  and _36909_ (_04530_, _04126_, _03353_);
  and _36910_ (_04531_, _04530_, _03060_);
  not _36911_ (_04532_, _04530_);
  and _36912_ (_04534_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _36913_ (_05176_, _04534_, _04531_);
  and _36914_ (_04535_, _04530_, _03067_);
  and _36915_ (_04537_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _36916_ (_05179_, _04537_, _04535_);
  and _36917_ (_04538_, _04530_, _03071_);
  and _36918_ (_04540_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _36919_ (_05183_, _04540_, _04538_);
  and _36920_ (_04541_, _04530_, _03074_);
  and _36921_ (_04543_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _36922_ (_05186_, _04543_, _04541_);
  and _36923_ (_04544_, _04530_, _03077_);
  and _36924_ (_04546_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _36925_ (_05189_, _04546_, _04544_);
  and _36926_ (_04547_, _04530_, _03080_);
  and _36927_ (_04549_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _36928_ (_05192_, _04549_, _04547_);
  and _36929_ (_04551_, _04530_, _03083_);
  and _36930_ (_04552_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _36931_ (_05195_, _04552_, _04551_);
  and _36932_ (_04553_, _04530_, _03087_);
  and _36933_ (_04555_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _36934_ (_05197_, _04555_, _04553_);
  and _36935_ (_04556_, _25446_, _25101_);
  and _36936_ (_04558_, _04556_, _02008_);
  and _36937_ (_04559_, _04558_, _02966_);
  and _36938_ (_04560_, _04559_, _02963_);
  and _36939_ (_04562_, _04560_, _03060_);
  not _36940_ (_04563_, _04560_);
  and _36941_ (_04564_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _36942_ (_05203_, _04564_, _04562_);
  and _36943_ (_04566_, _04560_, _03067_);
  and _36944_ (_04567_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _36945_ (_05207_, _04567_, _04566_);
  and _36946_ (_04569_, _04560_, _03071_);
  and _36947_ (_04570_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _36948_ (_05210_, _04570_, _04569_);
  and _36949_ (_04572_, _04560_, _03074_);
  and _36950_ (_04573_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _36951_ (_05213_, _04573_, _04572_);
  and _36952_ (_04575_, _04560_, _03077_);
  and _36953_ (_04577_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _36954_ (_05216_, _04577_, _04575_);
  and _36955_ (_04578_, _04560_, _03080_);
  and _36956_ (_04579_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _36957_ (_05219_, _04579_, _04578_);
  and _36958_ (_04581_, _04560_, _03083_);
  and _36959_ (_04582_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _36960_ (_05222_, _04582_, _04581_);
  and _36961_ (_04584_, _04560_, _03087_);
  and _36962_ (_04585_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _36963_ (_05224_, _04585_, _04584_);
  and _36964_ (_04587_, _04559_, _03062_);
  and _36965_ (_04588_, _04587_, _03060_);
  not _36966_ (_04590_, _04587_);
  and _36967_ (_04591_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or _36968_ (_05228_, _04591_, _04588_);
  and _36969_ (_04593_, _04587_, _03067_);
  and _36970_ (_04594_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or _36971_ (_05231_, _04594_, _04593_);
  and _36972_ (_04596_, _04587_, _03071_);
  and _36973_ (_04597_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _36974_ (_05235_, _04597_, _04596_);
  and _36975_ (_04599_, _04587_, _03074_);
  and _36976_ (_04600_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _36977_ (_05238_, _04600_, _04599_);
  and _36978_ (_04602_, _04587_, _03077_);
  and _36979_ (_04603_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or _36980_ (_05241_, _04603_, _04602_);
  and _36981_ (_04606_, _04587_, _03080_);
  and _36982_ (_04607_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or _36983_ (_05244_, _04607_, _04606_);
  and _36984_ (_04609_, _04587_, _03083_);
  and _36985_ (_04610_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or _36986_ (_05247_, _04610_, _04609_);
  and _36987_ (_04612_, _04587_, _03087_);
  and _36988_ (_04613_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or _36989_ (_05249_, _04613_, _04612_);
  and _36990_ (_04615_, _04559_, _03091_);
  and _36991_ (_04616_, _04615_, _03060_);
  not _36992_ (_04617_, _04615_);
  and _36993_ (_04619_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or _36994_ (_05253_, _04619_, _04616_);
  and _36995_ (_04620_, _04615_, _03067_);
  and _36996_ (_04622_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _36997_ (_05256_, _04622_, _04620_);
  and _36998_ (_04623_, _04615_, _03071_);
  and _36999_ (_04625_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or _37000_ (_05259_, _04625_, _04623_);
  and _37001_ (_04627_, _04615_, _03074_);
  and _37002_ (_04628_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or _37003_ (_05262_, _04628_, _04627_);
  and _37004_ (_04629_, _04615_, _03077_);
  and _37005_ (_04631_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or _37006_ (_05265_, _04631_, _04629_);
  and _37007_ (_04632_, _04615_, _03080_);
  and _37008_ (_04634_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or _37009_ (_05268_, _04634_, _04632_);
  and _37010_ (_04635_, _04615_, _03083_);
  and _37011_ (_04637_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or _37012_ (_05271_, _04637_, _04635_);
  and _37013_ (_04638_, _04615_, _03087_);
  and _37014_ (_04640_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or _37015_ (_05274_, _04640_, _04638_);
  and _37016_ (_04641_, _04559_, _03113_);
  and _37017_ (_04643_, _04641_, _03060_);
  not _37018_ (_04644_, _04641_);
  and _37019_ (_04645_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _37020_ (_05277_, _04645_, _04643_);
  and _37021_ (_04647_, _04641_, _03067_);
  and _37022_ (_04648_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _37023_ (_05280_, _04648_, _04647_);
  and _37024_ (_04650_, _04641_, _03071_);
  and _37025_ (_04652_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _37026_ (_05283_, _04652_, _04650_);
  and _37027_ (_04653_, _04641_, _03074_);
  and _37028_ (_04654_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _37029_ (_05287_, _04654_, _04653_);
  and _37030_ (_04656_, _04641_, _03077_);
  and _37031_ (_04657_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _37032_ (_05290_, _04657_, _04656_);
  and _37033_ (_04659_, _04641_, _03080_);
  and _37034_ (_04660_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _37035_ (_05293_, _04660_, _04659_);
  and _37036_ (_04662_, _04641_, _03083_);
  and _37037_ (_04663_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _37038_ (_05296_, _04663_, _04662_);
  and _37039_ (_04665_, _04641_, _03087_);
  and _37040_ (_04666_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _37041_ (_05298_, _04666_, _04665_);
  and _37042_ (_04668_, _04559_, _03136_);
  and _37043_ (_04669_, _04668_, _03060_);
  not _37044_ (_04671_, _04668_);
  and _37045_ (_04672_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _37046_ (_05302_, _04672_, _04669_);
  and _37047_ (_04674_, _04668_, _03067_);
  and _37048_ (_04675_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _37049_ (_05305_, _04675_, _04674_);
  and _37050_ (_04677_, _04668_, _03071_);
  and _37051_ (_04678_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _37052_ (_05308_, _04678_, _04677_);
  and _37053_ (_04680_, _04668_, _03074_);
  and _37054_ (_04681_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _37055_ (_05311_, _04681_, _04680_);
  and _37056_ (_04683_, _04668_, _03077_);
  and _37057_ (_04684_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _37058_ (_05315_, _04684_, _04683_);
  and _37059_ (_04686_, _04668_, _03080_);
  and _37060_ (_04687_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _37061_ (_05318_, _04687_, _04686_);
  and _37062_ (_04689_, _04668_, _03083_);
  and _37063_ (_04690_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _37064_ (_05321_, _04690_, _04689_);
  and _37065_ (_04692_, _04668_, _03087_);
  and _37066_ (_04693_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _37067_ (_05323_, _04693_, _04692_);
  and _37068_ (_04695_, _04559_, _03159_);
  and _37069_ (_04696_, _04695_, _03060_);
  not _37070_ (_04697_, _04695_);
  and _37071_ (_04699_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or _37072_ (_05327_, _04699_, _04696_);
  and _37073_ (_04701_, _04695_, _03067_);
  and _37074_ (_04702_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _37075_ (_05330_, _04702_, _04701_);
  and _37076_ (_04703_, _04695_, _03071_);
  and _37077_ (_04705_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or _37078_ (_05333_, _04705_, _04703_);
  and _37079_ (_04706_, _04695_, _03074_);
  and _37080_ (_04709_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _37081_ (_05336_, _04709_, _04706_);
  and _37082_ (_04710_, _04695_, _03077_);
  and _37083_ (_04712_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or _37084_ (_05339_, _04712_, _04710_);
  and _37085_ (_04713_, _04695_, _03080_);
  and _37086_ (_04715_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _37087_ (_05342_, _04715_, _04713_);
  and _37088_ (_04716_, _04695_, _03083_);
  and _37089_ (_04718_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or _37090_ (_05345_, _04718_, _04716_);
  and _37091_ (_04719_, _04695_, _03087_);
  and _37092_ (_04721_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _37093_ (_05348_, _04721_, _04719_);
  and _37094_ (_04722_, _04559_, _03179_);
  and _37095_ (_04724_, _04722_, _03060_);
  not _37096_ (_04725_, _04722_);
  and _37097_ (_04727_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or _37098_ (_05351_, _04727_, _04724_);
  and _37099_ (_04728_, _04722_, _03067_);
  and _37100_ (_04729_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or _37101_ (_05354_, _04729_, _04728_);
  and _37102_ (_04731_, _04722_, _03071_);
  and _37103_ (_04732_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _37104_ (_05357_, _04732_, _04731_);
  and _37105_ (_04734_, _04722_, _03074_);
  and _37106_ (_04735_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or _37107_ (_05360_, _04735_, _04734_);
  and _37108_ (_04737_, _04722_, _03077_);
  and _37109_ (_04738_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or _37110_ (_05363_, _04738_, _04737_);
  and _37111_ (_04740_, _04722_, _03080_);
  and _37112_ (_04741_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or _37113_ (_05367_, _04741_, _04740_);
  and _37114_ (_04743_, _04722_, _03083_);
  and _37115_ (_04744_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or _37116_ (_05370_, _04744_, _04743_);
  and _37117_ (_04746_, _04722_, _03087_);
  and _37118_ (_04747_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or _37119_ (_05372_, _04747_, _04746_);
  and _37120_ (_04749_, _04559_, _03198_);
  and _37121_ (_04751_, _04749_, _03060_);
  not _37122_ (_04752_, _04749_);
  and _37123_ (_04753_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _37124_ (_05376_, _04753_, _04751_);
  and _37125_ (_04755_, _04749_, _03067_);
  and _37126_ (_04756_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _37127_ (_05379_, _04756_, _04755_);
  and _37128_ (_04758_, _04749_, _03071_);
  and _37129_ (_04759_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _37130_ (_05382_, _04759_, _04758_);
  and _37131_ (_04761_, _04749_, _03074_);
  and _37132_ (_04762_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _37133_ (_05385_, _04762_, _04761_);
  and _37134_ (_04764_, _04749_, _03077_);
  and _37135_ (_04765_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _37136_ (_05388_, _04765_, _04764_);
  and _37137_ (_04767_, _04749_, _03080_);
  and _37138_ (_04768_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _37139_ (_05391_, _04768_, _04767_);
  and _37140_ (_04770_, _04749_, _03083_);
  and _37141_ (_04771_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _37142_ (_05395_, _04771_, _04770_);
  and _37143_ (_04773_, _04749_, _03087_);
  and _37144_ (_04774_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _37145_ (_05397_, _04774_, _04773_);
  and _37146_ (_04776_, _04559_, _03218_);
  and _37147_ (_04777_, _04776_, _03060_);
  not _37148_ (_04778_, _04776_);
  and _37149_ (_04780_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or _37150_ (_05401_, _04780_, _04777_);
  and _37151_ (_04781_, _04776_, _03067_);
  and _37152_ (_04783_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _37153_ (_05404_, _04783_, _04781_);
  and _37154_ (_04784_, _04776_, _03071_);
  and _37155_ (_04786_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or _37156_ (_05407_, _04786_, _04784_);
  and _37157_ (_04787_, _04776_, _03074_);
  and _37158_ (_04789_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _37159_ (_05410_, _04789_, _04787_);
  and _37160_ (_04790_, _04776_, _03077_);
  and _37161_ (_04792_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or _37162_ (_05413_, _04792_, _04790_);
  and _37163_ (_04793_, _04776_, _03080_);
  and _37164_ (_04795_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _37165_ (_05416_, _04795_, _04793_);
  and _37166_ (_04796_, _04776_, _03083_);
  and _37167_ (_04798_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or _37168_ (_05419_, _04798_, _04796_);
  and _37169_ (_04800_, _04776_, _03087_);
  and _37170_ (_04801_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or _37171_ (_05422_, _04801_, _04800_);
  and _37172_ (_04802_, _04559_, _03237_);
  and _37173_ (_04803_, _04802_, _03060_);
  not _37174_ (_04804_, _04802_);
  and _37175_ (_04806_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _37176_ (_05426_, _04806_, _04803_);
  and _37177_ (_04807_, _04802_, _03067_);
  and _37178_ (_04809_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _37179_ (_05429_, _04809_, _04807_);
  and _37180_ (_04811_, _04802_, _03071_);
  and _37181_ (_04813_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _37182_ (_05432_, _04813_, _04811_);
  and _37183_ (_04814_, _04802_, _03074_);
  and _37184_ (_04816_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _37185_ (_05435_, _04816_, _04814_);
  and _37186_ (_04817_, _04802_, _03077_);
  and _37187_ (_04819_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _37188_ (_05438_, _04819_, _04817_);
  and _37189_ (_04820_, _04802_, _03080_);
  and _37190_ (_04822_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _37191_ (_05441_, _04822_, _04820_);
  and _37192_ (_04823_, _04802_, _03083_);
  and _37193_ (_04825_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _37194_ (_05444_, _04825_, _04823_);
  and _37195_ (_04827_, _04802_, _03087_);
  and _37196_ (_04828_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _37197_ (_05446_, _04828_, _04827_);
  and _37198_ (_04829_, _04559_, _03256_);
  and _37199_ (_04831_, _04829_, _03060_);
  not _37200_ (_04832_, _04829_);
  and _37201_ (_04833_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _37202_ (_05450_, _04833_, _04831_);
  and _37203_ (_04835_, _04829_, _03067_);
  and _37204_ (_04836_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _37205_ (_05453_, _04836_, _04835_);
  and _37206_ (_04838_, _04829_, _03071_);
  and _37207_ (_04839_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _37208_ (_05456_, _04839_, _04838_);
  and _37209_ (_04841_, _04829_, _03074_);
  and _37210_ (_04842_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _37211_ (_05459_, _04842_, _04841_);
  and _37212_ (_04844_, _04829_, _03077_);
  and _37213_ (_04845_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _37214_ (_05462_, _04845_, _04844_);
  and _37215_ (_04847_, _04829_, _03080_);
  and _37216_ (_04848_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _37217_ (_05465_, _04848_, _04847_);
  and _37218_ (_04850_, _04829_, _03083_);
  and _37219_ (_04852_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _37220_ (_05468_, _04852_, _04850_);
  and _37221_ (_04853_, _04829_, _03087_);
  and _37222_ (_04854_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _37223_ (_05471_, _04854_, _04853_);
  and _37224_ (_04856_, _04559_, _03275_);
  and _37225_ (_04857_, _04856_, _03060_);
  not _37226_ (_04859_, _04856_);
  and _37227_ (_04860_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or _37228_ (_05475_, _04860_, _04857_);
  and _37229_ (_04862_, _04856_, _03067_);
  and _37230_ (_04863_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _37231_ (_05478_, _04863_, _04862_);
  and _37232_ (_04865_, _04856_, _03071_);
  and _37233_ (_04866_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _37234_ (_05481_, _04866_, _04865_);
  and _37235_ (_04868_, _04856_, _03074_);
  and _37236_ (_04869_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or _37237_ (_05484_, _04869_, _04868_);
  and _37238_ (_04871_, _04856_, _03077_);
  and _37239_ (_04872_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or _37240_ (_05487_, _04872_, _04871_);
  and _37241_ (_04874_, _04856_, _03080_);
  and _37242_ (_04875_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or _37243_ (_05490_, _04875_, _04874_);
  and _37244_ (_04877_, _04856_, _03083_);
  and _37245_ (_04878_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or _37246_ (_05493_, _04878_, _04877_);
  and _37247_ (_04880_, _04856_, _03087_);
  and _37248_ (_04881_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _37249_ (_05495_, _04881_, _04880_);
  and _37250_ (_04883_, _04559_, _03295_);
  and _37251_ (_04884_, _04883_, _03060_);
  not _37252_ (_04885_, _04883_);
  and _37253_ (_04887_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or _37254_ (_05499_, _04887_, _04884_);
  and _37255_ (_04888_, _04883_, _03067_);
  and _37256_ (_04890_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or _37257_ (_05503_, _04890_, _04888_);
  and _37258_ (_04891_, _04883_, _03071_);
  and _37259_ (_04893_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or _37260_ (_05506_, _04893_, _04891_);
  and _37261_ (_04894_, _04883_, _03074_);
  and _37262_ (_04896_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _37263_ (_05509_, _04896_, _04894_);
  and _37264_ (_04897_, _04883_, _03077_);
  and _37265_ (_04899_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or _37266_ (_05512_, _04899_, _04897_);
  and _37267_ (_04901_, _04883_, _03080_);
  and _37268_ (_04902_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or _37269_ (_05515_, _04902_, _04901_);
  and _37270_ (_04903_, _04883_, _03083_);
  and _37271_ (_04905_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or _37272_ (_05518_, _04905_, _04903_);
  and _37273_ (_04906_, _04883_, _03087_);
  and _37274_ (_04908_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or _37275_ (_05520_, _04908_, _04906_);
  and _37276_ (_04909_, _04559_, _03315_);
  and _37277_ (_04911_, _04909_, _03060_);
  not _37278_ (_04912_, _04909_);
  and _37279_ (_04913_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _37280_ (_05524_, _04913_, _04911_);
  and _37281_ (_04916_, _04909_, _03067_);
  and _37282_ (_04917_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _37283_ (_05527_, _04917_, _04916_);
  and _37284_ (_04919_, _04909_, _03071_);
  and _37285_ (_04920_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _37286_ (_05530_, _04920_, _04919_);
  and _37287_ (_04922_, _04909_, _03074_);
  and _37288_ (_04923_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _37289_ (_05533_, _04923_, _04922_);
  and _37290_ (_04925_, _04909_, _03077_);
  and _37291_ (_04927_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _37292_ (_05536_, _04927_, _04925_);
  and _37293_ (_04928_, _04909_, _03080_);
  and _37294_ (_04929_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _37295_ (_05539_, _04929_, _04928_);
  and _37296_ (_04931_, _04909_, _03083_);
  and _37297_ (_04932_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _37298_ (_05542_, _04932_, _04931_);
  and _37299_ (_04934_, _04909_, _03087_);
  and _37300_ (_04935_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _37301_ (_05545_, _04935_, _04934_);
  and _37302_ (_04937_, _04559_, _03334_);
  and _37303_ (_04938_, _04937_, _03060_);
  not _37304_ (_04940_, _04937_);
  and _37305_ (_04941_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _37306_ (_05548_, _04941_, _04938_);
  and _37307_ (_04943_, _04937_, _03067_);
  and _37308_ (_04944_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _37309_ (_05551_, _04944_, _04943_);
  and _37310_ (_04946_, _04937_, _03071_);
  and _37311_ (_04947_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _37312_ (_05555_, _04947_, _04946_);
  and _37313_ (_04949_, _04937_, _03074_);
  and _37314_ (_04950_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _37315_ (_05558_, _04950_, _04949_);
  and _37316_ (_04952_, _04937_, _03077_);
  and _37317_ (_04953_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _37318_ (_05561_, _04953_, _04952_);
  and _37319_ (_04955_, _04937_, _03080_);
  and _37320_ (_04956_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _37321_ (_05564_, _04956_, _04955_);
  and _37322_ (_04958_, _04937_, _03083_);
  and _37323_ (_04959_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _37324_ (_05567_, _04959_, _04958_);
  and _37325_ (_04961_, _04937_, _03087_);
  and _37326_ (_04962_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _37327_ (_05569_, _04962_, _04961_);
  and _37328_ (_04964_, _04559_, _03353_);
  and _37329_ (_04965_, _04964_, _03060_);
  not _37330_ (_04966_, _04964_);
  and _37331_ (_04968_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or _37332_ (_05573_, _04968_, _04965_);
  and _37333_ (_04969_, _04964_, _03067_);
  and _37334_ (_04971_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or _37335_ (_05576_, _04971_, _04969_);
  and _37336_ (_04972_, _04964_, _03071_);
  and _37337_ (_04974_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _37338_ (_05579_, _04974_, _04972_);
  and _37339_ (_04976_, _04964_, _03074_);
  and _37340_ (_04977_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _37341_ (_05583_, _04977_, _04976_);
  and _37342_ (_04978_, _04964_, _03077_);
  and _37343_ (_04980_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or _37344_ (_05586_, _04980_, _04978_);
  and _37345_ (_04981_, _04964_, _03080_);
  and _37346_ (_04983_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or _37347_ (_05589_, _04983_, _04981_);
  and _37348_ (_04984_, _04964_, _03083_);
  and _37349_ (_04986_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or _37350_ (_05592_, _04986_, _04984_);
  and _37351_ (_04987_, _04964_, _03087_);
  and _37352_ (_04989_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or _37353_ (_05594_, _04989_, _04987_);
  and _37354_ (_04990_, _04558_, _03373_);
  and _37355_ (_04992_, _04990_, _02963_);
  and _37356_ (_04993_, _04992_, _03060_);
  not _37357_ (_04994_, _04992_);
  and _37358_ (_04996_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or _37359_ (_05598_, _04996_, _04993_);
  and _37360_ (_04997_, _04992_, _03067_);
  and _37361_ (_04999_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or _37362_ (_05601_, _04999_, _04997_);
  and _37363_ (_05001_, _04992_, _03071_);
  and _37364_ (_05002_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or _37365_ (_05604_, _05002_, _05001_);
  and _37366_ (_05003_, _04992_, _03074_);
  and _37367_ (_05005_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or _37368_ (_05608_, _05005_, _05003_);
  and _37369_ (_05006_, _04992_, _03077_);
  and _37370_ (_05008_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or _37371_ (_05611_, _05008_, _05006_);
  and _37372_ (_05009_, _04992_, _03080_);
  and _37373_ (_05011_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _37374_ (_05614_, _05011_, _05009_);
  and _37375_ (_05012_, _04992_, _03083_);
  and _37376_ (_05014_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or _37377_ (_05617_, _05014_, _05012_);
  and _37378_ (_05015_, _04992_, _03087_);
  and _37379_ (_05017_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _37380_ (_05619_, _05017_, _05015_);
  and _37381_ (_05018_, _04990_, _03062_);
  and _37382_ (_05020_, _05018_, _03060_);
  not _37383_ (_05021_, _05018_);
  and _37384_ (_05022_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _37385_ (_05623_, _05022_, _05020_);
  and _37386_ (_05024_, _05018_, _03067_);
  and _37387_ (_05026_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _37388_ (_05626_, _05026_, _05024_);
  and _37389_ (_05027_, _05018_, _03071_);
  and _37390_ (_05028_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _37391_ (_05629_, _05028_, _05027_);
  and _37392_ (_05030_, _05018_, _03074_);
  and _37393_ (_05031_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _37394_ (_05632_, _05031_, _05030_);
  and _37395_ (_05033_, _05018_, _03077_);
  and _37396_ (_05034_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _37397_ (_05636_, _05034_, _05033_);
  and _37398_ (_05036_, _05018_, _03080_);
  and _37399_ (_05037_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _37400_ (_05639_, _05037_, _05036_);
  and _37401_ (_05039_, _05018_, _03083_);
  and _37402_ (_05040_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _37403_ (_05642_, _05040_, _05039_);
  and _37404_ (_05042_, _05018_, _03087_);
  and _37405_ (_05043_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _37406_ (_05644_, _05043_, _05042_);
  and _37407_ (_05045_, _04990_, _03091_);
  and _37408_ (_05046_, _05045_, _03060_);
  not _37409_ (_05048_, _05045_);
  and _37410_ (_05049_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _37411_ (_05648_, _05049_, _05046_);
  and _37412_ (_05051_, _05045_, _03067_);
  and _37413_ (_05052_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _37414_ (_05651_, _05052_, _05051_);
  and _37415_ (_05054_, _05045_, _03071_);
  and _37416_ (_05055_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _37417_ (_05654_, _05055_, _05054_);
  and _37418_ (_05057_, _05045_, _03074_);
  and _37419_ (_05058_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _37420_ (_05657_, _05058_, _05057_);
  and _37421_ (_05060_, _05045_, _03077_);
  and _37422_ (_05061_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _37423_ (_05660_, _05061_, _05060_);
  and _37424_ (_05063_, _05045_, _03080_);
  and _37425_ (_05064_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _37426_ (_05663_, _05064_, _05063_);
  and _37427_ (_05066_, _05045_, _03083_);
  and _37428_ (_05067_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _37429_ (_05666_, _05067_, _05066_);
  and _37430_ (_05069_, _05045_, _03087_);
  and _37431_ (_05070_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _37432_ (_05669_, _05070_, _05069_);
  and _37433_ (_05072_, _04990_, _03113_);
  and _37434_ (_05073_, _05072_, _03060_);
  not _37435_ (_05075_, _05072_);
  and _37436_ (_05076_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or _37437_ (_05672_, _05076_, _05073_);
  and _37438_ (_05077_, _05072_, _03067_);
  and _37439_ (_05079_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or _37440_ (_05675_, _05079_, _05077_);
  and _37441_ (_05080_, _05072_, _03071_);
  and _37442_ (_05082_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or _37443_ (_05678_, _05082_, _05080_);
  and _37444_ (_05083_, _05072_, _03074_);
  and _37445_ (_05085_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or _37446_ (_05681_, _05085_, _05083_);
  and _37447_ (_05086_, _05072_, _03077_);
  and _37448_ (_05088_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or _37449_ (_05684_, _05088_, _05086_);
  and _37450_ (_05089_, _05072_, _03080_);
  and _37451_ (_05091_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or _37452_ (_05688_, _05091_, _05089_);
  and _37453_ (_05092_, _05072_, _03083_);
  and _37454_ (_05094_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or _37455_ (_05691_, _05094_, _05092_);
  and _37456_ (_05095_, _05072_, _03087_);
  and _37457_ (_05097_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _37458_ (_05693_, _05097_, _05095_);
  and _37459_ (_05099_, _04990_, _03136_);
  and _37460_ (_05100_, _05099_, _03060_);
  not _37461_ (_05101_, _05099_);
  and _37462_ (_05102_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or _37463_ (_05697_, _05102_, _05100_);
  and _37464_ (_05104_, _05099_, _03067_);
  and _37465_ (_05105_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or _37466_ (_05700_, _05105_, _05104_);
  and _37467_ (_05107_, _05099_, _03071_);
  and _37468_ (_05108_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or _37469_ (_05703_, _05108_, _05107_);
  and _37470_ (_05110_, _05099_, _03074_);
  and _37471_ (_05111_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or _37472_ (_05706_, _05111_, _05110_);
  and _37473_ (_05113_, _05099_, _03077_);
  and _37474_ (_05114_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or _37475_ (_05709_, _05114_, _05113_);
  and _37476_ (_05116_, _05099_, _03080_);
  and _37477_ (_05117_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _37478_ (_05712_, _05117_, _05116_);
  and _37479_ (_05119_, _05099_, _03083_);
  and _37480_ (_05120_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or _37481_ (_05716_, _05120_, _05119_);
  and _37482_ (_05122_, _05099_, _03087_);
  and _37483_ (_05124_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or _37484_ (_05718_, _05124_, _05122_);
  and _37485_ (_05125_, _04990_, _03159_);
  and _37486_ (_05126_, _05125_, _03060_);
  not _37487_ (_05128_, _05125_);
  and _37488_ (_05129_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _37489_ (_05722_, _05129_, _05126_);
  and _37490_ (_05131_, _05125_, _03067_);
  and _37491_ (_05132_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _37492_ (_05725_, _05132_, _05131_);
  and _37493_ (_05134_, _05125_, _03071_);
  and _37494_ (_05135_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _37495_ (_05728_, _05135_, _05134_);
  and _37496_ (_05137_, _05125_, _03074_);
  and _37497_ (_05138_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _37498_ (_05731_, _05138_, _05137_);
  and _37499_ (_05140_, _05125_, _03077_);
  and _37500_ (_05141_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _37501_ (_05734_, _05141_, _05140_);
  and _37502_ (_05143_, _05125_, _03080_);
  and _37503_ (_05144_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _37504_ (_05737_, _05144_, _05143_);
  and _37505_ (_05146_, _05125_, _03083_);
  and _37506_ (_05147_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _37507_ (_05740_, _05147_, _05146_);
  and _37508_ (_05149_, _05125_, _03087_);
  and _37509_ (_05150_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _37510_ (_05743_, _05150_, _05149_);
  and _37511_ (_05152_, _04990_, _03179_);
  and _37512_ (_05153_, _05152_, _03060_);
  not _37513_ (_05154_, _05152_);
  and _37514_ (_05156_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _37515_ (_05746_, _05156_, _05153_);
  and _37516_ (_05157_, _05152_, _03067_);
  and _37517_ (_05159_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _37518_ (_05749_, _05159_, _05157_);
  and _37519_ (_05160_, _05152_, _03071_);
  and _37520_ (_05162_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _37521_ (_05752_, _05162_, _05160_);
  and _37522_ (_05163_, _05152_, _03074_);
  and _37523_ (_05165_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _37524_ (_05755_, _05165_, _05163_);
  and _37525_ (_05166_, _05152_, _03077_);
  and _37526_ (_05168_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _37527_ (_05758_, _05168_, _05166_);
  and _37528_ (_05169_, _05152_, _03080_);
  and _37529_ (_05171_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _37530_ (_05761_, _05171_, _05169_);
  and _37531_ (_05173_, _05152_, _03083_);
  and _37532_ (_05174_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _37533_ (_05764_, _05174_, _05173_);
  and _37534_ (_05175_, _05152_, _03087_);
  and _37535_ (_05177_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _37536_ (_05767_, _05177_, _05175_);
  and _37537_ (_05178_, _04990_, _03198_);
  and _37538_ (_05180_, _05178_, _03060_);
  not _37539_ (_05181_, _05178_);
  and _37540_ (_05182_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or _37541_ (_05771_, _05182_, _05180_);
  and _37542_ (_05184_, _05178_, _03067_);
  and _37543_ (_05185_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or _37544_ (_05774_, _05185_, _05184_);
  and _37545_ (_05187_, _05178_, _03071_);
  and _37546_ (_05188_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or _37547_ (_05777_, _05188_, _05187_);
  and _37548_ (_05190_, _05178_, _03074_);
  and _37549_ (_05191_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or _37550_ (_05780_, _05191_, _05190_);
  and _37551_ (_05193_, _05178_, _03077_);
  and _37552_ (_05194_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or _37553_ (_05783_, _05194_, _05193_);
  and _37554_ (_05196_, _05178_, _03080_);
  and _37555_ (_05198_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _37556_ (_05786_, _05198_, _05196_);
  and _37557_ (_05199_, _05178_, _03083_);
  and _37558_ (_05200_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or _37559_ (_05789_, _05200_, _05199_);
  and _37560_ (_05201_, _05178_, _03087_);
  and _37561_ (_05202_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or _37562_ (_05791_, _05202_, _05201_);
  and _37563_ (_05204_, _04990_, _03218_);
  and _37564_ (_05205_, _05204_, _03060_);
  not _37565_ (_05206_, _05204_);
  and _37566_ (_05208_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _37567_ (_05796_, _05208_, _05205_);
  and _37568_ (_05209_, _05204_, _03067_);
  and _37569_ (_05211_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _37570_ (_05799_, _05211_, _05209_);
  and _37571_ (_05212_, _05204_, _03071_);
  and _37572_ (_05214_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _37573_ (_05802_, _05214_, _05212_);
  and _37574_ (_05215_, _05204_, _03074_);
  and _37575_ (_05217_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _37576_ (_05805_, _05217_, _05215_);
  and _37577_ (_05218_, _05204_, _03077_);
  and _37578_ (_05220_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _37579_ (_05808_, _05220_, _05218_);
  and _37580_ (_05221_, _05204_, _03080_);
  and _37581_ (_05223_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _37582_ (_05811_, _05223_, _05221_);
  and _37583_ (_05225_, _05204_, _03083_);
  and _37584_ (_05226_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _37585_ (_05814_, _05226_, _05225_);
  and _37586_ (_05227_, _05204_, _03087_);
  and _37587_ (_05229_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _37588_ (_05816_, _05229_, _05227_);
  and _37589_ (_05230_, _04990_, _03237_);
  and _37590_ (_05232_, _05230_, _03060_);
  not _37591_ (_05233_, _05230_);
  and _37592_ (_05234_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or _37593_ (_05820_, _05234_, _05232_);
  and _37594_ (_05236_, _05230_, _03067_);
  and _37595_ (_05237_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or _37596_ (_05823_, _05237_, _05236_);
  and _37597_ (_05239_, _05230_, _03071_);
  and _37598_ (_05240_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or _37599_ (_05826_, _05240_, _05239_);
  and _37600_ (_05242_, _05230_, _03074_);
  and _37601_ (_05243_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or _37602_ (_05829_, _05243_, _05242_);
  and _37603_ (_05245_, _05230_, _03077_);
  and _37604_ (_05246_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or _37605_ (_05832_, _05246_, _05245_);
  and _37606_ (_05248_, _05230_, _03080_);
  and _37607_ (_05250_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or _37608_ (_05835_, _05250_, _05248_);
  and _37609_ (_05251_, _05230_, _03083_);
  and _37610_ (_05252_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or _37611_ (_05838_, _05252_, _05251_);
  and _37612_ (_05254_, _05230_, _03087_);
  and _37613_ (_05255_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or _37614_ (_05841_, _05255_, _05254_);
  and _37615_ (_05257_, _04990_, _03256_);
  and _37616_ (_05258_, _05257_, _03060_);
  not _37617_ (_05260_, _05257_);
  and _37618_ (_05261_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or _37619_ (_05844_, _05261_, _05258_);
  and _37620_ (_05263_, _05257_, _03067_);
  and _37621_ (_05264_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or _37622_ (_05848_, _05264_, _05263_);
  and _37623_ (_05266_, _05257_, _03071_);
  and _37624_ (_05267_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or _37625_ (_05851_, _05267_, _05266_);
  and _37626_ (_05269_, _05257_, _03074_);
  and _37627_ (_05270_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or _37628_ (_05854_, _05270_, _05269_);
  and _37629_ (_05272_, _05257_, _03077_);
  and _37630_ (_05273_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or _37631_ (_05857_, _05273_, _05272_);
  and _37632_ (_05275_, _05257_, _03080_);
  and _37633_ (_05276_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or _37634_ (_05860_, _05276_, _05275_);
  and _37635_ (_05278_, _05257_, _03083_);
  and _37636_ (_05279_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or _37637_ (_05863_, _05279_, _05278_);
  and _37638_ (_05281_, _05257_, _03087_);
  and _37639_ (_05282_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or _37640_ (_05866_, _05282_, _05281_);
  and _37641_ (_05284_, _04990_, _03275_);
  and _37642_ (_05285_, _05284_, _03060_);
  not _37643_ (_05286_, _05284_);
  and _37644_ (_05288_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _37645_ (_05869_, _05288_, _05285_);
  and _37646_ (_05289_, _05284_, _03067_);
  and _37647_ (_05291_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _37648_ (_05872_, _05291_, _05289_);
  and _37649_ (_05292_, _05284_, _03071_);
  and _37650_ (_05294_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _37651_ (_05876_, _05294_, _05292_);
  and _37652_ (_05295_, _05284_, _03074_);
  and _37653_ (_05297_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _37654_ (_05879_, _05297_, _05295_);
  and _37655_ (_05299_, _05284_, _03077_);
  and _37656_ (_05300_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _37657_ (_05882_, _05300_, _05299_);
  and _37658_ (_05301_, _05284_, _03080_);
  and _37659_ (_05303_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _37660_ (_05885_, _05303_, _05301_);
  and _37661_ (_05304_, _05284_, _03083_);
  and _37662_ (_05306_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _37663_ (_05888_, _05306_, _05304_);
  and _37664_ (_05307_, _05284_, _03087_);
  and _37665_ (_05309_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _37666_ (_05890_, _05309_, _05307_);
  and _37667_ (_05310_, _04990_, _03295_);
  and _37668_ (_05312_, _05310_, _03060_);
  not _37669_ (_05313_, _05310_);
  and _37670_ (_05314_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _37671_ (_05894_, _05314_, _05312_);
  and _37672_ (_05316_, _05310_, _03067_);
  and _37673_ (_05317_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _37674_ (_05897_, _05317_, _05316_);
  and _37675_ (_05319_, _05310_, _03071_);
  and _37676_ (_05320_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _37677_ (_05900_, _05320_, _05319_);
  and _37678_ (_05322_, _05310_, _03074_);
  and _37679_ (_05324_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _37680_ (_05904_, _05324_, _05322_);
  and _37681_ (_05325_, _05310_, _03077_);
  and _37682_ (_05326_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _37683_ (_05907_, _05326_, _05325_);
  and _37684_ (_05328_, _05310_, _03080_);
  and _37685_ (_05329_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _37686_ (_05910_, _05329_, _05328_);
  and _37687_ (_05331_, _05310_, _03083_);
  and _37688_ (_05332_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _37689_ (_05913_, _05332_, _05331_);
  and _37690_ (_05334_, _05310_, _03087_);
  and _37691_ (_05335_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _37692_ (_05915_, _05335_, _05334_);
  and _37693_ (_05337_, _04990_, _03315_);
  and _37694_ (_05338_, _05337_, _03060_);
  not _37695_ (_05340_, _05337_);
  and _37696_ (_05341_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or _37697_ (_05919_, _05341_, _05338_);
  and _37698_ (_05343_, _05337_, _03067_);
  and _37699_ (_05344_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or _37700_ (_05922_, _05344_, _05343_);
  and _37701_ (_05346_, _05337_, _03071_);
  and _37702_ (_05347_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or _37703_ (_05925_, _05347_, _05346_);
  and _37704_ (_05349_, _05337_, _03074_);
  and _37705_ (_05350_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or _37706_ (_05928_, _05350_, _05349_);
  and _37707_ (_05352_, _05337_, _03077_);
  and _37708_ (_05353_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or _37709_ (_05931_, _05353_, _05352_);
  and _37710_ (_05355_, _05337_, _03080_);
  and _37711_ (_05356_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _37712_ (_05934_, _05356_, _05355_);
  and _37713_ (_05358_, _05337_, _03083_);
  and _37714_ (_05359_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or _37715_ (_05937_, _05359_, _05358_);
  and _37716_ (_05361_, _05337_, _03087_);
  and _37717_ (_05362_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or _37718_ (_05940_, _05362_, _05361_);
  and _37719_ (_05364_, _04990_, _03334_);
  and _37720_ (_05365_, _05364_, _03060_);
  not _37721_ (_05366_, _05364_);
  and _37722_ (_05368_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or _37723_ (_05943_, _05368_, _05365_);
  and _37724_ (_05369_, _05364_, _03067_);
  and _37725_ (_05371_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or _37726_ (_05946_, _05371_, _05369_);
  and _37727_ (_05373_, _05364_, _03071_);
  and _37728_ (_05374_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or _37729_ (_05949_, _05374_, _05373_);
  and _37730_ (_05375_, _05364_, _03074_);
  and _37731_ (_05377_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or _37732_ (_05952_, _05377_, _05375_);
  and _37733_ (_05378_, _05364_, _03077_);
  and _37734_ (_05380_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or _37735_ (_05956_, _05380_, _05378_);
  and _37736_ (_05381_, _05364_, _03080_);
  and _37737_ (_05383_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or _37738_ (_05959_, _05383_, _05381_);
  and _37739_ (_05384_, _05364_, _03083_);
  and _37740_ (_05386_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or _37741_ (_05962_, _05386_, _05384_);
  and _37742_ (_05387_, _05364_, _03087_);
  and _37743_ (_05389_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _37744_ (_05964_, _05389_, _05387_);
  and _37745_ (_05390_, _04990_, _03353_);
  and _37746_ (_05392_, _05390_, _03060_);
  not _37747_ (_05393_, _05390_);
  and _37748_ (_05394_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _37749_ (_05968_, _05394_, _05392_);
  and _37750_ (_05396_, _05390_, _03067_);
  and _37751_ (_05398_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _37752_ (_05971_, _05398_, _05396_);
  and _37753_ (_05399_, _05390_, _03071_);
  and _37754_ (_05400_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _37755_ (_05974_, _05400_, _05399_);
  and _37756_ (_05402_, _05390_, _03074_);
  and _37757_ (_05403_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _37758_ (_05977_, _05403_, _05402_);
  and _37759_ (_05405_, _05390_, _03077_);
  and _37760_ (_05406_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _37761_ (_05980_, _05406_, _05405_);
  and _37762_ (_05408_, _05390_, _03080_);
  and _37763_ (_05409_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _37764_ (_05984_, _05409_, _05408_);
  and _37765_ (_05411_, _05390_, _03083_);
  and _37766_ (_05412_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _37767_ (_05987_, _05412_, _05411_);
  and _37768_ (_05414_, _05390_, _03087_);
  and _37769_ (_05415_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _37770_ (_05989_, _05415_, _05414_);
  and _37771_ (_05417_, _04558_, _03699_);
  and _37772_ (_05418_, _05417_, _02963_);
  and _37773_ (_05420_, _05418_, _03060_);
  not _37774_ (_05421_, _05418_);
  and _37775_ (_05423_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _37776_ (_05993_, _05423_, _05420_);
  and _37777_ (_05424_, _05418_, _03067_);
  and _37778_ (_05425_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _37779_ (_05996_, _05425_, _05424_);
  and _37780_ (_05427_, _05418_, _03071_);
  and _37781_ (_05428_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _37782_ (_05999_, _05428_, _05427_);
  and _37783_ (_05430_, _05418_, _03074_);
  and _37784_ (_05431_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _37785_ (_06002_, _05431_, _05430_);
  and _37786_ (_05433_, _05418_, _03077_);
  and _37787_ (_05434_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _37788_ (_06005_, _05434_, _05433_);
  and _37789_ (_05436_, _05418_, _03080_);
  and _37790_ (_05437_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _37791_ (_06009_, _05437_, _05436_);
  and _37792_ (_05439_, _05418_, _03083_);
  and _37793_ (_05440_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _37794_ (_06012_, _05440_, _05439_);
  and _37795_ (_05442_, _05418_, _03087_);
  and _37796_ (_05443_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _37797_ (_06014_, _05443_, _05442_);
  and _37798_ (_05445_, _05417_, _03062_);
  and _37799_ (_05447_, _05445_, _03060_);
  not _37800_ (_05448_, _05445_);
  and _37801_ (_05449_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or _37802_ (_06018_, _05449_, _05447_);
  and _37803_ (_05451_, _05445_, _03067_);
  and _37804_ (_05452_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or _37805_ (_06021_, _05452_, _05451_);
  and _37806_ (_05454_, _05445_, _03071_);
  and _37807_ (_05455_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or _37808_ (_06024_, _05455_, _05454_);
  and _37809_ (_05457_, _05445_, _03074_);
  and _37810_ (_05458_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or _37811_ (_06027_, _05458_, _05457_);
  and _37812_ (_05460_, _05445_, _03077_);
  and _37813_ (_05461_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or _37814_ (_06030_, _05461_, _05460_);
  and _37815_ (_05463_, _05445_, _03080_);
  and _37816_ (_05464_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or _37817_ (_06033_, _05464_, _05463_);
  and _37818_ (_05466_, _05445_, _03083_);
  and _37819_ (_05467_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or _37820_ (_06037_, _05467_, _05466_);
  and _37821_ (_05469_, _05445_, _03087_);
  and _37822_ (_05470_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _37823_ (_06039_, _05470_, _05469_);
  and _37824_ (_05472_, _05417_, _03091_);
  and _37825_ (_05473_, _05472_, _03060_);
  not _37826_ (_05474_, _05472_);
  and _37827_ (_05476_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or _37828_ (_06043_, _05476_, _05473_);
  and _37829_ (_05477_, _05472_, _03067_);
  and _37830_ (_05479_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or _37831_ (_06046_, _05479_, _05477_);
  and _37832_ (_05480_, _05472_, _03071_);
  and _37833_ (_05482_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or _37834_ (_06049_, _05482_, _05480_);
  and _37835_ (_05483_, _05472_, _03074_);
  and _37836_ (_05485_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or _37837_ (_06052_, _05485_, _05483_);
  and _37838_ (_05486_, _05472_, _03077_);
  and _37839_ (_05488_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or _37840_ (_06055_, _05488_, _05486_);
  and _37841_ (_05489_, _05472_, _03080_);
  and _37842_ (_05491_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or _37843_ (_06058_, _05491_, _05489_);
  and _37844_ (_05492_, _05472_, _03083_);
  and _37845_ (_05494_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or _37846_ (_06061_, _05494_, _05492_);
  and _37847_ (_05496_, _05472_, _03087_);
  and _37848_ (_05497_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or _37849_ (_06064_, _05497_, _05496_);
  and _37850_ (_05498_, _05417_, _03113_);
  and _37851_ (_05500_, _05498_, _03060_);
  not _37852_ (_05501_, _05498_);
  and _37853_ (_05502_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _37854_ (_06067_, _05502_, _05500_);
  and _37855_ (_05504_, _05498_, _03067_);
  and _37856_ (_05505_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _37857_ (_06070_, _05505_, _05504_);
  and _37858_ (_05507_, _05498_, _03071_);
  and _37859_ (_05508_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _37860_ (_06073_, _05508_, _05507_);
  and _37861_ (_05510_, _05498_, _03074_);
  and _37862_ (_05511_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _37863_ (_06076_, _05511_, _05510_);
  and _37864_ (_05513_, _05498_, _03077_);
  and _37865_ (_05514_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _37866_ (_06079_, _05514_, _05513_);
  and _37867_ (_05516_, _05498_, _03080_);
  and _37868_ (_05517_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _37869_ (_06082_, _05517_, _05516_);
  and _37870_ (_05519_, _05498_, _03083_);
  and _37871_ (_05521_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _37872_ (_06085_, _05521_, _05519_);
  and _37873_ (_05522_, _05498_, _03087_);
  and _37874_ (_05523_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _37875_ (_06088_, _05523_, _05522_);
  and _37876_ (_05525_, _05417_, _03136_);
  and _37877_ (_05526_, _05525_, _03060_);
  not _37878_ (_05528_, _05525_);
  and _37879_ (_05529_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _37880_ (_06092_, _05529_, _05526_);
  and _37881_ (_05531_, _05525_, _03067_);
  and _37882_ (_05532_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _37883_ (_06095_, _05532_, _05531_);
  and _37884_ (_05534_, _05525_, _03071_);
  and _37885_ (_05535_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _37886_ (_06098_, _05535_, _05534_);
  and _37887_ (_05537_, _05525_, _03074_);
  and _37888_ (_05538_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _37889_ (_06101_, _05538_, _05537_);
  and _37890_ (_05540_, _05525_, _03077_);
  and _37891_ (_05541_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _37892_ (_06104_, _05541_, _05540_);
  and _37893_ (_05543_, _05525_, _03080_);
  and _37894_ (_05544_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _37895_ (_06107_, _05544_, _05543_);
  and _37896_ (_05546_, _05525_, _03083_);
  and _37897_ (_05547_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _37898_ (_06110_, _05547_, _05546_);
  and _37899_ (_05549_, _05525_, _03087_);
  and _37900_ (_05550_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _37901_ (_06112_, _05550_, _05549_);
  and _37902_ (_05552_, _05417_, _03159_);
  and _37903_ (_05553_, _05552_, _03060_);
  not _37904_ (_05554_, _05552_);
  and _37905_ (_05556_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or _37906_ (_06117_, _05556_, _05553_);
  and _37907_ (_05557_, _05552_, _03067_);
  and _37908_ (_05559_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or _37909_ (_06120_, _05559_, _05557_);
  and _37910_ (_05560_, _05552_, _03071_);
  and _37911_ (_05562_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or _37912_ (_06123_, _05562_, _05560_);
  and _37913_ (_05563_, _05552_, _03074_);
  and _37914_ (_05565_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or _37915_ (_06126_, _05565_, _05563_);
  and _37916_ (_05566_, _05552_, _03077_);
  and _37917_ (_05568_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or _37918_ (_06129_, _05568_, _05566_);
  and _37919_ (_05570_, _05552_, _03080_);
  and _37920_ (_05571_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or _37921_ (_06132_, _05571_, _05570_);
  and _37922_ (_05572_, _05552_, _03083_);
  and _37923_ (_05574_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or _37924_ (_06135_, _05574_, _05572_);
  and _37925_ (_05575_, _05552_, _03087_);
  and _37926_ (_05577_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _37927_ (_06137_, _05577_, _05575_);
  and _37928_ (_05578_, _05417_, _03179_);
  and _37929_ (_05580_, _05578_, _03060_);
  not _37930_ (_05581_, _05578_);
  and _37931_ (_05582_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or _37932_ (_06141_, _05582_, _05580_);
  and _37933_ (_05584_, _05578_, _03067_);
  and _37934_ (_05585_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or _37935_ (_06144_, _05585_, _05584_);
  and _37936_ (_05587_, _05578_, _03071_);
  and _37937_ (_05588_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or _37938_ (_06147_, _05588_, _05587_);
  and _37939_ (_05590_, _05578_, _03074_);
  and _37940_ (_05591_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or _37941_ (_06150_, _05591_, _05590_);
  and _37942_ (_05593_, _05578_, _03077_);
  and _37943_ (_05595_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or _37944_ (_06153_, _05595_, _05593_);
  and _37945_ (_05596_, _05578_, _03080_);
  and _37946_ (_05597_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or _37947_ (_06156_, _05597_, _05596_);
  and _37948_ (_05599_, _05578_, _03083_);
  and _37949_ (_05600_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or _37950_ (_06159_, _05600_, _05599_);
  and _37951_ (_05602_, _05578_, _03087_);
  and _37952_ (_05603_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or _37953_ (_06162_, _05603_, _05602_);
  and _37954_ (_05605_, _05417_, _03198_);
  and _37955_ (_05606_, _05605_, _03060_);
  not _37956_ (_05607_, _05605_);
  and _37957_ (_05609_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _37958_ (_06165_, _05609_, _05606_);
  and _37959_ (_05610_, _05605_, _03067_);
  and _37960_ (_05612_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _37961_ (_06169_, _05612_, _05610_);
  and _37962_ (_05613_, _05605_, _03071_);
  and _37963_ (_05615_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _37964_ (_06172_, _05615_, _05613_);
  and _37965_ (_05616_, _05605_, _03074_);
  and _37966_ (_05618_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _37967_ (_06175_, _05618_, _05616_);
  and _37968_ (_05620_, _05605_, _03077_);
  and _37969_ (_05621_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _37970_ (_06178_, _05621_, _05620_);
  and _37971_ (_05622_, _05605_, _03080_);
  and _37972_ (_05624_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _37973_ (_06181_, _05624_, _05622_);
  and _37974_ (_05625_, _05605_, _03083_);
  and _37975_ (_05627_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _37976_ (_06184_, _05627_, _05625_);
  and _37977_ (_05628_, _05605_, _03087_);
  and _37978_ (_05630_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _37979_ (_06186_, _05630_, _05628_);
  and _37980_ (_05631_, _05417_, _03218_);
  and _37981_ (_05633_, _05631_, _03060_);
  not _37982_ (_05634_, _05631_);
  and _37983_ (_05635_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or _37984_ (_06190_, _05635_, _05633_);
  and _37985_ (_05637_, _05631_, _03067_);
  and _37986_ (_05638_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or _37987_ (_06193_, _05638_, _05637_);
  and _37988_ (_05640_, _05631_, _03071_);
  and _37989_ (_05641_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or _37990_ (_06197_, _05641_, _05640_);
  and _37991_ (_05643_, _05631_, _03074_);
  and _37992_ (_05645_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or _37993_ (_06200_, _05645_, _05643_);
  and _37994_ (_05646_, _05631_, _03077_);
  and _37995_ (_05647_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or _37996_ (_06203_, _05647_, _05646_);
  and _37997_ (_05649_, _05631_, _03080_);
  and _37998_ (_05650_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or _37999_ (_06206_, _05650_, _05649_);
  and _38000_ (_05652_, _05631_, _03083_);
  and _38001_ (_05653_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or _38002_ (_06209_, _05653_, _05652_);
  and _38003_ (_05655_, _05631_, _03087_);
  and _38004_ (_05656_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _38005_ (_06211_, _05656_, _05655_);
  and _38006_ (_05658_, _05417_, _03237_);
  and _38007_ (_05659_, _05658_, _03060_);
  not _38008_ (_05661_, _05658_);
  and _38009_ (_05662_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _38010_ (_06215_, _05662_, _05659_);
  and _38011_ (_05664_, _05658_, _03067_);
  and _38012_ (_05665_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _38013_ (_06218_, _05665_, _05664_);
  and _38014_ (_05667_, _05658_, _03071_);
  and _38015_ (_05668_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _38016_ (_06221_, _05668_, _05667_);
  and _38017_ (_05670_, _05658_, _03074_);
  and _38018_ (_05671_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _38019_ (_06224_, _05671_, _05670_);
  and _38020_ (_05673_, _05658_, _03077_);
  and _38021_ (_05674_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _38022_ (_06227_, _05674_, _05673_);
  and _38023_ (_05676_, _05658_, _03080_);
  and _38024_ (_05677_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _38025_ (_06230_, _05677_, _05676_);
  and _38026_ (_05679_, _05658_, _03083_);
  and _38027_ (_05680_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _38028_ (_06233_, _05680_, _05679_);
  and _38029_ (_05682_, _05658_, _03087_);
  and _38030_ (_05683_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _38031_ (_06236_, _05683_, _05682_);
  and _38032_ (_05685_, _05417_, _03256_);
  and _38033_ (_05686_, _05685_, _03060_);
  not _38034_ (_05687_, _05685_);
  and _38035_ (_05689_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _38036_ (_06239_, _05689_, _05686_);
  and _38037_ (_05690_, _05685_, _03067_);
  and _38038_ (_05692_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _38039_ (_06242_, _05692_, _05690_);
  and _38040_ (_05694_, _05685_, _03071_);
  and _38041_ (_05695_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _38042_ (_06245_, _05695_, _05694_);
  and _38043_ (_05696_, _05685_, _03074_);
  and _38044_ (_05698_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _38045_ (_06249_, _05698_, _05696_);
  and _38046_ (_05699_, _05685_, _03077_);
  and _38047_ (_05701_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _38048_ (_06252_, _05701_, _05699_);
  and _38049_ (_05702_, _05685_, _03080_);
  and _38050_ (_05704_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _38051_ (_06255_, _05704_, _05702_);
  and _38052_ (_05705_, _05685_, _03083_);
  and _38053_ (_05707_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _38054_ (_06258_, _05707_, _05705_);
  and _38055_ (_05708_, _05685_, _03087_);
  and _38056_ (_05710_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _38057_ (_06260_, _05710_, _05708_);
  and _38058_ (_05711_, _05417_, _03275_);
  and _38059_ (_05713_, _05711_, _03060_);
  not _38060_ (_05714_, _05711_);
  and _38061_ (_05715_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or _38062_ (_06264_, _05715_, _05713_);
  and _38063_ (_05717_, _05711_, _03067_);
  and _38064_ (_05719_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or _38065_ (_06267_, _05719_, _05717_);
  and _38066_ (_05720_, _05711_, _03071_);
  and _38067_ (_05721_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or _38068_ (_06270_, _05721_, _05720_);
  and _38069_ (_05723_, _05711_, _03074_);
  and _38070_ (_05724_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or _38071_ (_06273_, _05724_, _05723_);
  and _38072_ (_05726_, _05711_, _03077_);
  and _38073_ (_05727_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or _38074_ (_06277_, _05727_, _05726_);
  and _38075_ (_05729_, _05711_, _03080_);
  and _38076_ (_05730_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or _38077_ (_06280_, _05730_, _05729_);
  and _38078_ (_05732_, _05711_, _03083_);
  and _38079_ (_05733_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or _38080_ (_06283_, _05733_, _05732_);
  and _38081_ (_05735_, _05711_, _03087_);
  and _38082_ (_05736_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or _38083_ (_06286_, _05736_, _05735_);
  and _38084_ (_05738_, _05417_, _03295_);
  and _38085_ (_05739_, _05738_, _03060_);
  not _38086_ (_05741_, _05738_);
  and _38087_ (_05742_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or _38088_ (_06289_, _05742_, _05739_);
  and _38089_ (_05744_, _05738_, _03067_);
  and _38090_ (_05745_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or _38091_ (_06292_, _05745_, _05744_);
  and _38092_ (_05747_, _05738_, _03071_);
  and _38093_ (_05748_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or _38094_ (_06295_, _05748_, _05747_);
  and _38095_ (_05750_, _05738_, _03074_);
  and _38096_ (_05751_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or _38097_ (_06298_, _05751_, _05750_);
  and _38098_ (_05753_, _05738_, _03077_);
  and _38099_ (_05754_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or _38100_ (_06301_, _05754_, _05753_);
  and _38101_ (_05756_, _05738_, _03080_);
  and _38102_ (_05757_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _38103_ (_06305_, _05757_, _05756_);
  and _38104_ (_05759_, _05738_, _03083_);
  and _38105_ (_05760_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or _38106_ (_06308_, _05760_, _05759_);
  and _38107_ (_05762_, _05738_, _03087_);
  and _38108_ (_05763_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _38109_ (_06310_, _05763_, _05762_);
  and _38110_ (_05765_, _05417_, _03315_);
  and _38111_ (_05766_, _05765_, _03060_);
  not _38112_ (_05768_, _05765_);
  and _38113_ (_05769_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _38114_ (_06314_, _05769_, _05766_);
  and _38115_ (_05770_, _05765_, _03067_);
  and _38116_ (_05772_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _38117_ (_06317_, _05772_, _05770_);
  and _38118_ (_05773_, _05765_, _03071_);
  and _38119_ (_05775_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _38120_ (_06320_, _05775_, _05773_);
  and _38121_ (_05776_, _05765_, _03074_);
  and _38122_ (_05778_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _38123_ (_06323_, _05778_, _05776_);
  and _38124_ (_05779_, _05765_, _03077_);
  and _38125_ (_05781_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _38126_ (_06326_, _05781_, _05779_);
  and _38127_ (_05782_, _05765_, _03080_);
  and _38128_ (_05784_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _38129_ (_06329_, _05784_, _05782_);
  and _38130_ (_05785_, _05765_, _03083_);
  and _38131_ (_05787_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _38132_ (_06333_, _05787_, _05785_);
  and _38133_ (_05788_, _05765_, _03087_);
  and _38134_ (_05790_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _38135_ (_06335_, _05790_, _05788_);
  and _38136_ (_05792_, _05417_, _03334_);
  and _38137_ (_05793_, _05792_, _03060_);
  not _38138_ (_05794_, _05792_);
  and _38139_ (_05795_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _38140_ (_06339_, _05795_, _05793_);
  and _38141_ (_05797_, _05792_, _03067_);
  and _38142_ (_05798_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _38143_ (_06342_, _05798_, _05797_);
  and _38144_ (_05800_, _05792_, _03071_);
  and _38145_ (_05801_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _38146_ (_06345_, _05801_, _05800_);
  and _38147_ (_05803_, _05792_, _03074_);
  and _38148_ (_05804_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _38149_ (_06348_, _05804_, _05803_);
  and _38150_ (_05806_, _05792_, _03077_);
  and _38151_ (_05807_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _38152_ (_06351_, _05807_, _05806_);
  and _38153_ (_05809_, _05792_, _03080_);
  and _38154_ (_05810_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _38155_ (_06354_, _05810_, _05809_);
  and _38156_ (_05812_, _05792_, _03083_);
  and _38157_ (_05813_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _38158_ (_06357_, _05813_, _05812_);
  and _38159_ (_05815_, _05792_, _03087_);
  and _38160_ (_05817_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _38161_ (_06360_, _05817_, _05815_);
  and _38162_ (_05818_, _05417_, _03353_);
  and _38163_ (_05819_, _05818_, _03060_);
  not _38164_ (_05821_, _05818_);
  and _38165_ (_05822_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or _38166_ (_06363_, _05822_, _05819_);
  and _38167_ (_05824_, _05818_, _03067_);
  and _38168_ (_05825_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or _38169_ (_06366_, _05825_, _05824_);
  and _38170_ (_05827_, _05818_, _03071_);
  and _38171_ (_05828_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or _38172_ (_06369_, _05828_, _05827_);
  and _38173_ (_05830_, _05818_, _03074_);
  and _38174_ (_05831_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or _38175_ (_06372_, _05831_, _05830_);
  and _38176_ (_05833_, _05818_, _03077_);
  and _38177_ (_05834_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or _38178_ (_06375_, _05834_, _05833_);
  and _38179_ (_05836_, _05818_, _03080_);
  and _38180_ (_05837_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or _38181_ (_06378_, _05837_, _05836_);
  and _38182_ (_05839_, _05818_, _03083_);
  and _38183_ (_05840_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or _38184_ (_06381_, _05840_, _05839_);
  and _38185_ (_05842_, _05818_, _03087_);
  and _38186_ (_05843_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or _38187_ (_06384_, _05843_, _05842_);
  and _38188_ (_05845_, _04558_, _04125_);
  and _38189_ (_05846_, _05845_, _02963_);
  and _38190_ (_05847_, _05846_, _03060_);
  not _38191_ (_05849_, _05846_);
  and _38192_ (_05850_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or _38193_ (_06389_, _05850_, _05847_);
  and _38194_ (_05852_, _05846_, _03067_);
  and _38195_ (_05853_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or _38196_ (_06392_, _05853_, _05852_);
  and _38197_ (_05855_, _05846_, _03071_);
  and _38198_ (_05856_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or _38199_ (_06395_, _05856_, _05855_);
  and _38200_ (_05858_, _05846_, _03074_);
  and _38201_ (_05859_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or _38202_ (_06398_, _05859_, _05858_);
  and _38203_ (_05861_, _05846_, _03077_);
  and _38204_ (_05862_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or _38205_ (_06401_, _05862_, _05861_);
  and _38206_ (_05864_, _05846_, _03080_);
  and _38207_ (_05865_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or _38208_ (_06404_, _05865_, _05864_);
  and _38209_ (_05867_, _05846_, _03083_);
  and _38210_ (_05868_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or _38211_ (_06407_, _05868_, _05867_);
  and _38212_ (_05870_, _05846_, _03087_);
  and _38213_ (_05871_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or _38214_ (_06409_, _05871_, _05870_);
  and _38215_ (_05873_, _05845_, _03062_);
  and _38216_ (_05874_, _05873_, _03060_);
  not _38217_ (_05875_, _05873_);
  and _38218_ (_05877_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _38219_ (_06413_, _05877_, _05874_);
  and _38220_ (_05878_, _05873_, _03067_);
  and _38221_ (_05880_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _38222_ (_06416_, _05880_, _05878_);
  and _38223_ (_05881_, _05873_, _03071_);
  and _38224_ (_05883_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _38225_ (_06419_, _05883_, _05881_);
  and _38226_ (_05884_, _05873_, _03074_);
  and _38227_ (_05886_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _38228_ (_06422_, _05886_, _05884_);
  and _38229_ (_05887_, _05873_, _03077_);
  and _38230_ (_05889_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _38231_ (_06425_, _05889_, _05887_);
  and _38232_ (_05891_, _05873_, _03080_);
  and _38233_ (_05892_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _38234_ (_06428_, _05892_, _05891_);
  and _38235_ (_05893_, _05873_, _03083_);
  and _38236_ (_05895_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _38237_ (_06431_, _05895_, _05893_);
  and _38238_ (_05896_, _05873_, _03087_);
  and _38239_ (_05898_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _38240_ (_06434_, _05898_, _05896_);
  and _38241_ (_05899_, _05845_, _03091_);
  and _38242_ (_05901_, _05899_, _03060_);
  not _38243_ (_05902_, _05899_);
  and _38244_ (_05903_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _38245_ (_06438_, _05903_, _05901_);
  and _38246_ (_05905_, _05899_, _03067_);
  and _38247_ (_05906_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _38248_ (_06441_, _05906_, _05905_);
  and _38249_ (_05908_, _05899_, _03071_);
  and _38250_ (_05909_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _38251_ (_06444_, _05909_, _05908_);
  and _38252_ (_05911_, _05899_, _03074_);
  and _38253_ (_05912_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _38254_ (_06447_, _05912_, _05911_);
  and _38255_ (_05914_, _05899_, _03077_);
  and _38256_ (_05916_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _38257_ (_06450_, _05916_, _05914_);
  and _38258_ (_05917_, _05899_, _03080_);
  and _38259_ (_05918_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _38260_ (_06453_, _05918_, _05917_);
  and _38261_ (_05920_, _05899_, _03083_);
  and _38262_ (_05921_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _38263_ (_06456_, _05921_, _05920_);
  and _38264_ (_05923_, _05899_, _03087_);
  and _38265_ (_05924_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _38266_ (_06458_, _05924_, _05923_);
  and _38267_ (_05926_, _05845_, _03113_);
  and _38268_ (_05927_, _05926_, _03060_);
  not _38269_ (_05929_, _05926_);
  and _38270_ (_05930_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or _38271_ (_06462_, _05930_, _05927_);
  and _38272_ (_05932_, _05926_, _03067_);
  and _38273_ (_05933_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or _38274_ (_06466_, _05933_, _05932_);
  and _38275_ (_05935_, _05926_, _03071_);
  and _38276_ (_05936_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or _38277_ (_06469_, _05936_, _05935_);
  and _38278_ (_05938_, _05926_, _03074_);
  and _38279_ (_05939_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or _38280_ (_06472_, _05939_, _05938_);
  and _38281_ (_05941_, _05926_, _03077_);
  and _38282_ (_05942_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or _38283_ (_06475_, _05942_, _05941_);
  and _38284_ (_05944_, _05926_, _03080_);
  and _38285_ (_05945_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or _38286_ (_06478_, _05945_, _05944_);
  and _38287_ (_05947_, _05926_, _03083_);
  and _38288_ (_05948_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or _38289_ (_06481_, _05948_, _05947_);
  and _38290_ (_05950_, _05926_, _03087_);
  and _38291_ (_05951_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or _38292_ (_06483_, _05951_, _05950_);
  and _38293_ (_05953_, _05845_, _03136_);
  and _38294_ (_05954_, _05953_, _03060_);
  not _38295_ (_05955_, _05953_);
  and _38296_ (_05957_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or _38297_ (_06487_, _05957_, _05954_);
  and _38298_ (_05958_, _05953_, _03067_);
  and _38299_ (_05960_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or _38300_ (_06490_, _05960_, _05958_);
  and _38301_ (_05961_, _05953_, _03071_);
  and _38302_ (_05963_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or _38303_ (_06493_, _05963_, _05961_);
  and _38304_ (_05965_, _05953_, _03074_);
  and _38305_ (_05966_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or _38306_ (_06496_, _05966_, _05965_);
  and _38307_ (_05967_, _05953_, _03077_);
  and _38308_ (_05969_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or _38309_ (_06499_, _05969_, _05967_);
  and _38310_ (_05970_, _05953_, _03080_);
  and _38311_ (_05972_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or _38312_ (_06502_, _05972_, _05970_);
  and _38313_ (_05973_, _05953_, _03083_);
  and _38314_ (_05975_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or _38315_ (_06505_, _05975_, _05973_);
  and _38316_ (_05976_, _05953_, _03087_);
  and _38317_ (_05978_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or _38318_ (_06508_, _05978_, _05976_);
  and _38319_ (_05979_, _05845_, _03159_);
  and _38320_ (_05981_, _05979_, _03060_);
  not _38321_ (_05982_, _05979_);
  and _38322_ (_05983_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _38323_ (_06511_, _05983_, _05981_);
  and _38324_ (_05985_, _05979_, _03067_);
  and _38325_ (_05986_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _38326_ (_06514_, _05986_, _05985_);
  and _38327_ (_05988_, _05979_, _03071_);
  and _38328_ (_05990_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _38329_ (_06518_, _05990_, _05988_);
  and _38330_ (_05991_, _05979_, _03074_);
  and _38331_ (_05992_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _38332_ (_06521_, _05992_, _05991_);
  and _38333_ (_05994_, _05979_, _03077_);
  and _38334_ (_05995_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _38335_ (_06525_, _05995_, _05994_);
  and _38336_ (_05997_, _05979_, _03080_);
  and _38337_ (_05998_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _38338_ (_06528_, _05998_, _05997_);
  and _38339_ (_06000_, _05979_, _03083_);
  and _38340_ (_06001_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _38341_ (_06531_, _06001_, _06000_);
  and _38342_ (_06003_, _05979_, _03087_);
  and _38343_ (_06004_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _38344_ (_06533_, _06004_, _06003_);
  and _38345_ (_06006_, _05845_, _03179_);
  and _38346_ (_06007_, _06006_, _03060_);
  not _38347_ (_06008_, _06006_);
  and _38348_ (_06010_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _38349_ (_06537_, _06010_, _06007_);
  and _38350_ (_06011_, _06006_, _03067_);
  and _38351_ (_06013_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _38352_ (_06540_, _06013_, _06011_);
  and _38353_ (_06015_, _06006_, _03071_);
  and _38354_ (_06016_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _38355_ (_06543_, _06016_, _06015_);
  and _38356_ (_06017_, _06006_, _03074_);
  and _38357_ (_06019_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _38358_ (_06547_, _06019_, _06017_);
  and _38359_ (_06020_, _06006_, _03077_);
  and _38360_ (_06022_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _38361_ (_06550_, _06022_, _06020_);
  and _38362_ (_06023_, _06006_, _03080_);
  and _38363_ (_06025_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _38364_ (_06553_, _06025_, _06023_);
  and _38365_ (_06026_, _06006_, _03083_);
  and _38366_ (_06028_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _38367_ (_06556_, _06028_, _06026_);
  and _38368_ (_06029_, _06006_, _03087_);
  and _38369_ (_06031_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _38370_ (_06558_, _06031_, _06029_);
  and _38371_ (_06032_, _05845_, _03198_);
  and _38372_ (_06034_, _06032_, _03060_);
  not _38373_ (_06035_, _06032_);
  and _38374_ (_06036_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or _38375_ (_06562_, _06036_, _06034_);
  and _38376_ (_06038_, _06032_, _03067_);
  and _38377_ (_06040_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or _38378_ (_06565_, _06040_, _06038_);
  and _38379_ (_06041_, _06032_, _03071_);
  and _38380_ (_06042_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or _38381_ (_06568_, _06042_, _06041_);
  and _38382_ (_06044_, _06032_, _03074_);
  and _38383_ (_06045_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or _38384_ (_06571_, _06045_, _06044_);
  and _38385_ (_06047_, _06032_, _03077_);
  and _38386_ (_06048_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or _38387_ (_06574_, _06048_, _06047_);
  and _38388_ (_06050_, _06032_, _03080_);
  and _38389_ (_06051_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or _38390_ (_06577_, _06051_, _06050_);
  and _38391_ (_06053_, _06032_, _03083_);
  and _38392_ (_06054_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or _38393_ (_06580_, _06054_, _06053_);
  and _38394_ (_06056_, _06032_, _03087_);
  and _38395_ (_06057_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or _38396_ (_06583_, _06057_, _06056_);
  and _38397_ (_06059_, _05845_, _03218_);
  and _38398_ (_06060_, _06059_, _03060_);
  not _38399_ (_06062_, _06059_);
  and _38400_ (_06063_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _38401_ (_06586_, _06063_, _06060_);
  and _38402_ (_06065_, _06059_, _03067_);
  and _38403_ (_06066_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _38404_ (_06589_, _06066_, _06065_);
  and _38405_ (_06068_, _06059_, _03071_);
  and _38406_ (_06069_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _38407_ (_06592_, _06069_, _06068_);
  and _38408_ (_06071_, _06059_, _03074_);
  and _38409_ (_06072_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _38410_ (_06595_, _06072_, _06071_);
  and _38411_ (_06074_, _06059_, _03077_);
  and _38412_ (_06075_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _38413_ (_06599_, _06075_, _06074_);
  and _38414_ (_06077_, _06059_, _03080_);
  and _38415_ (_06078_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _38416_ (_06602_, _06078_, _06077_);
  and _38417_ (_06080_, _06059_, _03083_);
  and _38418_ (_06081_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _38419_ (_06605_, _06081_, _06080_);
  and _38420_ (_06083_, _06059_, _03087_);
  and _38421_ (_06084_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _38422_ (_06607_, _06084_, _06083_);
  and _38423_ (_06086_, _05845_, _03237_);
  and _38424_ (_06087_, _06086_, _03060_);
  not _38425_ (_06089_, _06086_);
  and _38426_ (_06090_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or _38427_ (_06611_, _06090_, _06087_);
  and _38428_ (_06091_, _06086_, _03067_);
  and _38429_ (_06093_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or _38430_ (_06614_, _06093_, _06091_);
  and _38431_ (_06094_, _06086_, _03071_);
  and _38432_ (_06096_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or _38433_ (_06617_, _06096_, _06094_);
  and _38434_ (_06097_, _06086_, _03074_);
  and _38435_ (_06099_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or _38436_ (_06620_, _06099_, _06097_);
  and _38437_ (_06100_, _06086_, _03077_);
  and _38438_ (_06102_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or _38439_ (_06623_, _06102_, _06100_);
  and _38440_ (_06103_, _06086_, _03080_);
  and _38441_ (_06105_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or _38442_ (_06627_, _06105_, _06103_);
  and _38443_ (_06106_, _06086_, _03083_);
  and _38444_ (_06108_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or _38445_ (_06630_, _06108_, _06106_);
  and _38446_ (_06109_, _06086_, _03087_);
  and _38447_ (_06111_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or _38448_ (_06632_, _06111_, _06109_);
  and _38449_ (_06113_, _05845_, _03256_);
  and _38450_ (_06114_, _06113_, _03060_);
  not _38451_ (_06115_, _06113_);
  and _38452_ (_06116_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or _38453_ (_06636_, _06116_, _06114_);
  and _38454_ (_06118_, _06113_, _03067_);
  and _38455_ (_06119_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or _38456_ (_06639_, _06119_, _06118_);
  and _38457_ (_06121_, _06113_, _03071_);
  and _38458_ (_06122_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or _38459_ (_06642_, _06122_, _06121_);
  and _38460_ (_06124_, _06113_, _03074_);
  and _38461_ (_06125_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or _38462_ (_06645_, _06125_, _06124_);
  and _38463_ (_06127_, _06113_, _03077_);
  and _38464_ (_06128_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or _38465_ (_06648_, _06128_, _06127_);
  and _38466_ (_06130_, _06113_, _03080_);
  and _38467_ (_06131_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or _38468_ (_06651_, _06131_, _06130_);
  and _38469_ (_06133_, _06113_, _03083_);
  and _38470_ (_06134_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or _38471_ (_06654_, _06134_, _06133_);
  and _38472_ (_06136_, _06113_, _03087_);
  and _38473_ (_06138_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or _38474_ (_06657_, _06138_, _06136_);
  and _38475_ (_06139_, _05845_, _03275_);
  and _38476_ (_06140_, _06139_, _03060_);
  not _38477_ (_06142_, _06139_);
  and _38478_ (_06143_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _38479_ (_06660_, _06143_, _06140_);
  and _38480_ (_06145_, _06139_, _03067_);
  and _38481_ (_06146_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _38482_ (_06663_, _06146_, _06145_);
  and _38483_ (_06148_, _06139_, _03071_);
  and _38484_ (_06149_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _38485_ (_06666_, _06149_, _06148_);
  and _38486_ (_06151_, _06139_, _03074_);
  and _38487_ (_06152_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _38488_ (_06669_, _06152_, _06151_);
  and _38489_ (_06154_, _06139_, _03077_);
  and _38490_ (_06155_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _38491_ (_06672_, _06155_, _06154_);
  and _38492_ (_06157_, _06139_, _03080_);
  and _38493_ (_06158_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _38494_ (_06675_, _06158_, _06157_);
  and _38495_ (_06160_, _06139_, _03083_);
  and _38496_ (_06161_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _38497_ (_06679_, _06161_, _06160_);
  and _38498_ (_06163_, _06139_, _03087_);
  and _38499_ (_06164_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _38500_ (_06681_, _06164_, _06163_);
  and _38501_ (_06166_, _05845_, _03295_);
  and _38502_ (_06167_, _06166_, _03060_);
  not _38503_ (_06168_, _06166_);
  and _38504_ (_06170_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _38505_ (_06685_, _06170_, _06167_);
  and _38506_ (_06171_, _06166_, _03067_);
  and _38507_ (_06173_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _38508_ (_06688_, _06173_, _06171_);
  and _38509_ (_06174_, _06166_, _03071_);
  and _38510_ (_06176_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _38511_ (_06691_, _06176_, _06174_);
  and _38512_ (_06177_, _06166_, _03074_);
  and _38513_ (_06179_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _38514_ (_06694_, _06179_, _06177_);
  and _38515_ (_06180_, _06166_, _03077_);
  and _38516_ (_06182_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _38517_ (_06697_, _06182_, _06180_);
  and _38518_ (_06183_, _06166_, _03080_);
  and _38519_ (_06185_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _38520_ (_06700_, _06185_, _06183_);
  and _38521_ (_06187_, _06166_, _03083_);
  and _38522_ (_06188_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _38523_ (_06703_, _06188_, _06187_);
  and _38524_ (_06189_, _06166_, _03087_);
  and _38525_ (_06191_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _38526_ (_06706_, _06191_, _06189_);
  and _38527_ (_06192_, _05845_, _03315_);
  and _38528_ (_06194_, _06192_, _03060_);
  not _38529_ (_06195_, _06192_);
  and _38530_ (_06196_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or _38531_ (_06710_, _06196_, _06194_);
  and _38532_ (_06198_, _06192_, _03067_);
  and _38533_ (_06199_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or _38534_ (_06713_, _06199_, _06198_);
  and _38535_ (_06201_, _06192_, _03071_);
  and _38536_ (_06202_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or _38537_ (_06716_, _06202_, _06201_);
  and _38538_ (_06204_, _06192_, _03074_);
  and _38539_ (_06205_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or _38540_ (_06719_, _06205_, _06204_);
  and _38541_ (_06207_, _06192_, _03077_);
  and _38542_ (_06208_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or _38543_ (_06722_, _06208_, _06207_);
  and _38544_ (_06210_, _06192_, _03080_);
  and _38545_ (_06212_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or _38546_ (_06725_, _06212_, _06210_);
  and _38547_ (_06213_, _06192_, _03083_);
  and _38548_ (_06214_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or _38549_ (_06728_, _06214_, _06213_);
  and _38550_ (_06216_, _06192_, _03087_);
  and _38551_ (_06217_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or _38552_ (_06730_, _06217_, _06216_);
  and _38553_ (_06219_, _05845_, _03334_);
  and _38554_ (_06220_, _06219_, _03060_);
  not _38555_ (_06222_, _06219_);
  and _38556_ (_06223_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or _38557_ (_06735_, _06223_, _06220_);
  and _38558_ (_06225_, _06219_, _03067_);
  and _38559_ (_06226_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or _38560_ (_06738_, _06226_, _06225_);
  and _38561_ (_06228_, _06219_, _03071_);
  and _38562_ (_06229_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or _38563_ (_06741_, _06229_, _06228_);
  and _38564_ (_06231_, _06219_, _03074_);
  and _38565_ (_06232_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or _38566_ (_06744_, _06232_, _06231_);
  and _38567_ (_06234_, _06219_, _03077_);
  and _38568_ (_06235_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or _38569_ (_06747_, _06235_, _06234_);
  and _38570_ (_06237_, _06219_, _03080_);
  and _38571_ (_06238_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or _38572_ (_06750_, _06238_, _06237_);
  and _38573_ (_06240_, _06219_, _03083_);
  and _38574_ (_06241_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or _38575_ (_06753_, _06241_, _06240_);
  and _38576_ (_06243_, _06219_, _03087_);
  and _38577_ (_06244_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or _38578_ (_06755_, _06244_, _06243_);
  and _38579_ (_06246_, _05845_, _03353_);
  and _38580_ (_06247_, _06246_, _03060_);
  not _38581_ (_06248_, _06246_);
  and _38582_ (_06250_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _38583_ (_06759_, _06250_, _06247_);
  and _38584_ (_06251_, _06246_, _03067_);
  and _38585_ (_06253_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _38586_ (_06762_, _06253_, _06251_);
  and _38587_ (_06254_, _06246_, _03071_);
  and _38588_ (_06256_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _38589_ (_06765_, _06256_, _06254_);
  and _38590_ (_06257_, _06246_, _03074_);
  and _38591_ (_06259_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _38592_ (_06768_, _06259_, _06257_);
  and _38593_ (_06261_, _06246_, _03077_);
  and _38594_ (_06262_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _38595_ (_06771_, _06262_, _06261_);
  and _38596_ (_06263_, _06246_, _03080_);
  and _38597_ (_06265_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _38598_ (_06774_, _06265_, _06263_);
  and _38599_ (_06266_, _06246_, _03083_);
  and _38600_ (_06268_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _38601_ (_06777_, _06268_, _06266_);
  and _38602_ (_06269_, _06246_, _03087_);
  and _38603_ (_06271_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _38604_ (_06780_, _06271_, _06269_);
  and _38605_ (_06272_, _02137_, _26459_);
  and _38606_ (_06274_, _06272_, _02966_);
  and _38607_ (_06275_, _06274_, _02963_);
  and _38608_ (_06276_, _06275_, _03060_);
  not _38609_ (_06278_, _06275_);
  and _38610_ (_06279_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _38611_ (_06787_, _06279_, _06276_);
  and _38612_ (_06281_, _06275_, _03067_);
  and _38613_ (_06282_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _38614_ (_06790_, _06282_, _06281_);
  and _38615_ (_06284_, _06275_, _03071_);
  and _38616_ (_06285_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _38617_ (_06793_, _06285_, _06284_);
  and _38618_ (_06287_, _06275_, _03074_);
  and _38619_ (_06288_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _38620_ (_06796_, _06288_, _06287_);
  and _38621_ (_06290_, _06275_, _03077_);
  and _38622_ (_06291_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _38623_ (_06799_, _06291_, _06290_);
  and _38624_ (_06293_, _06275_, _03080_);
  and _38625_ (_06294_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _38626_ (_06802_, _06294_, _06293_);
  and _38627_ (_06296_, _06275_, _03083_);
  and _38628_ (_06297_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _38629_ (_06805_, _06297_, _06296_);
  and _38630_ (_06299_, _06275_, _03087_);
  and _38631_ (_06300_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _38632_ (_06808_, _06300_, _06299_);
  and _38633_ (_06302_, _06274_, _03062_);
  and _38634_ (_06303_, _06302_, _03060_);
  not _38635_ (_06304_, _06302_);
  and _38636_ (_06306_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or _38637_ (_06812_, _06306_, _06303_);
  and _38638_ (_06307_, _06302_, _03067_);
  and _38639_ (_06309_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or _38640_ (_06815_, _06309_, _06307_);
  and _38641_ (_06311_, _06302_, _03071_);
  and _38642_ (_06312_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or _38643_ (_06818_, _06312_, _06311_);
  and _38644_ (_06313_, _06302_, _03074_);
  and _38645_ (_06315_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or _38646_ (_06821_, _06315_, _06313_);
  and _38647_ (_06316_, _06302_, _03077_);
  and _38648_ (_06318_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or _38649_ (_06824_, _06318_, _06316_);
  and _38650_ (_06319_, _06302_, _03080_);
  and _38651_ (_06321_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or _38652_ (_06827_, _06321_, _06319_);
  and _38653_ (_06322_, _06302_, _03083_);
  and _38654_ (_06324_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or _38655_ (_06830_, _06324_, _06322_);
  and _38656_ (_06325_, _06302_, _03087_);
  and _38657_ (_06327_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or _38658_ (_06832_, _06327_, _06325_);
  and _38659_ (_06328_, _06274_, _03091_);
  and _38660_ (_06330_, _06328_, _03060_);
  not _38661_ (_06331_, _06328_);
  and _38662_ (_06332_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or _38663_ (_06836_, _06332_, _06330_);
  and _38664_ (_06334_, _06328_, _03067_);
  and _38665_ (_06336_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or _38666_ (_06840_, _06336_, _06334_);
  and _38667_ (_06337_, _06328_, _03071_);
  and _38668_ (_06338_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or _38669_ (_06843_, _06338_, _06337_);
  and _38670_ (_06340_, _06328_, _03074_);
  and _38671_ (_06341_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or _38672_ (_06846_, _06341_, _06340_);
  and _38673_ (_06343_, _06328_, _03077_);
  and _38674_ (_06344_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or _38675_ (_06849_, _06344_, _06343_);
  and _38676_ (_06346_, _06328_, _03080_);
  and _38677_ (_06347_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or _38678_ (_06852_, _06347_, _06346_);
  and _38679_ (_06349_, _06328_, _03083_);
  and _38680_ (_06350_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or _38681_ (_06855_, _06350_, _06349_);
  and _38682_ (_06352_, _06328_, _03087_);
  and _38683_ (_06353_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or _38684_ (_06857_, _06353_, _06352_);
  and _38685_ (_06355_, _06274_, _03113_);
  and _38686_ (_06356_, _06355_, _03060_);
  not _38687_ (_06358_, _06355_);
  and _38688_ (_06359_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _38689_ (_06861_, _06359_, _06356_);
  and _38690_ (_06361_, _06355_, _03067_);
  and _38691_ (_06362_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _38692_ (_06864_, _06362_, _06361_);
  and _38693_ (_06364_, _06355_, _03071_);
  and _38694_ (_06365_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _38695_ (_06867_, _06365_, _06364_);
  and _38696_ (_06367_, _06355_, _03074_);
  and _38697_ (_06368_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _38698_ (_06870_, _06368_, _06367_);
  and _38699_ (_06370_, _06355_, _03077_);
  and _38700_ (_06371_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _38701_ (_06873_, _06371_, _06370_);
  and _38702_ (_06373_, _06355_, _03080_);
  and _38703_ (_06374_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _38704_ (_06876_, _06374_, _06373_);
  and _38705_ (_06376_, _06355_, _03083_);
  and _38706_ (_06377_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _38707_ (_06879_, _06377_, _06376_);
  and _38708_ (_06379_, _06355_, _03087_);
  and _38709_ (_06380_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _38710_ (_06882_, _06380_, _06379_);
  and _38711_ (_06382_, _06274_, _03136_);
  and _38712_ (_06383_, _06382_, _03060_);
  not _38713_ (_06385_, _06382_);
  and _38714_ (_06386_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _38715_ (_06885_, _06386_, _06383_);
  and _38716_ (_06387_, _06382_, _03067_);
  and _38717_ (_06388_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _38718_ (_06888_, _06388_, _06387_);
  and _38719_ (_06390_, _06382_, _03071_);
  and _38720_ (_06391_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _38721_ (_06892_, _06391_, _06390_);
  and _38722_ (_06393_, _06382_, _03074_);
  and _38723_ (_06394_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _38724_ (_06895_, _06394_, _06393_);
  and _38725_ (_06396_, _06382_, _03077_);
  and _38726_ (_06397_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _38727_ (_06898_, _06397_, _06396_);
  and _38728_ (_06399_, _06382_, _03080_);
  and _38729_ (_06400_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _38730_ (_06901_, _06400_, _06399_);
  and _38731_ (_06402_, _06382_, _03083_);
  and _38732_ (_06403_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _38733_ (_06904_, _06403_, _06402_);
  and _38734_ (_06405_, _06382_, _03087_);
  and _38735_ (_06406_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _38736_ (_06906_, _06406_, _06405_);
  and _38737_ (_06408_, _06274_, _03159_);
  and _38738_ (_06410_, _06408_, _03060_);
  not _38739_ (_06411_, _06408_);
  and _38740_ (_06412_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or _38741_ (_06910_, _06412_, _06410_);
  and _38742_ (_06414_, _06408_, _03067_);
  and _38743_ (_06415_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or _38744_ (_06913_, _06415_, _06414_);
  and _38745_ (_06417_, _06408_, _03071_);
  and _38746_ (_06418_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or _38747_ (_06916_, _06418_, _06417_);
  and _38748_ (_06420_, _06408_, _03074_);
  and _38749_ (_06421_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or _38750_ (_06920_, _06421_, _06420_);
  and _38751_ (_06423_, _06408_, _03077_);
  and _38752_ (_06424_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or _38753_ (_06923_, _06424_, _06423_);
  and _38754_ (_06426_, _06408_, _03080_);
  and _38755_ (_06427_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or _38756_ (_06926_, _06427_, _06426_);
  and _38757_ (_06429_, _06408_, _03083_);
  and _38758_ (_06430_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or _38759_ (_06929_, _06430_, _06429_);
  and _38760_ (_06432_, _06408_, _03087_);
  and _38761_ (_06433_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or _38762_ (_06931_, _06433_, _06432_);
  and _38763_ (_06435_, _06274_, _03179_);
  and _38764_ (_06436_, _06435_, _03060_);
  not _38765_ (_06437_, _06435_);
  and _38766_ (_06439_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or _38767_ (_06935_, _06439_, _06436_);
  and _38768_ (_06440_, _06435_, _03067_);
  and _38769_ (_06442_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or _38770_ (_06938_, _06442_, _06440_);
  and _38771_ (_06443_, _06435_, _03071_);
  and _38772_ (_06445_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or _38773_ (_06941_, _06445_, _06443_);
  and _38774_ (_06446_, _06435_, _03074_);
  and _38775_ (_06448_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or _38776_ (_06944_, _06448_, _06446_);
  and _38777_ (_06449_, _06435_, _03077_);
  and _38778_ (_06451_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or _38779_ (_06947_, _06451_, _06449_);
  and _38780_ (_06452_, _06435_, _03080_);
  and _38781_ (_06454_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or _38782_ (_06950_, _06454_, _06452_);
  and _38783_ (_06455_, _06435_, _03083_);
  and _38784_ (_06457_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or _38785_ (_06953_, _06457_, _06455_);
  and _38786_ (_06459_, _06435_, _03087_);
  and _38787_ (_06460_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or _38788_ (_06956_, _06460_, _06459_);
  and _38789_ (_06461_, _06274_, _03198_);
  and _38790_ (_06463_, _06461_, _03060_);
  not _38791_ (_06464_, _06461_);
  and _38792_ (_06465_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _38793_ (_06959_, _06465_, _06463_);
  and _38794_ (_06467_, _06461_, _03067_);
  and _38795_ (_06468_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _38796_ (_06962_, _06468_, _06467_);
  and _38797_ (_06470_, _06461_, _03071_);
  and _38798_ (_06471_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _38799_ (_06965_, _06471_, _06470_);
  and _38800_ (_06473_, _06461_, _03074_);
  and _38801_ (_06474_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _38802_ (_06968_, _06474_, _06473_);
  and _38803_ (_06476_, _06461_, _03077_);
  and _38804_ (_06477_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _38805_ (_06972_, _06477_, _06476_);
  and _38806_ (_06479_, _06461_, _03080_);
  and _38807_ (_06480_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _38808_ (_06975_, _06480_, _06479_);
  and _38809_ (_06482_, _06461_, _03083_);
  and _38810_ (_06484_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _38811_ (_06978_, _06484_, _06482_);
  and _38812_ (_06485_, _06461_, _03087_);
  and _38813_ (_06486_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _38814_ (_06980_, _06486_, _06485_);
  and _38815_ (_06488_, _06274_, _03218_);
  and _38816_ (_06489_, _06488_, _03060_);
  not _38817_ (_06491_, _06488_);
  and _38818_ (_06492_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or _38819_ (_06984_, _06492_, _06489_);
  and _38820_ (_06494_, _06488_, _03067_);
  and _38821_ (_06495_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or _38822_ (_06987_, _06495_, _06494_);
  and _38823_ (_06497_, _06488_, _03071_);
  and _38824_ (_06498_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or _38825_ (_06990_, _06498_, _06497_);
  and _38826_ (_06500_, _06488_, _03074_);
  and _38827_ (_06501_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or _38828_ (_06993_, _06501_, _06500_);
  and _38829_ (_06503_, _06488_, _03077_);
  and _38830_ (_06504_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or _38831_ (_06996_, _06504_, _06503_);
  and _38832_ (_06506_, _06488_, _03080_);
  and _38833_ (_06507_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or _38834_ (_07000_, _06507_, _06506_);
  and _38835_ (_06509_, _06488_, _03083_);
  and _38836_ (_06510_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or _38837_ (_07003_, _06510_, _06509_);
  and _38838_ (_06512_, _06488_, _03087_);
  and _38839_ (_06513_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or _38840_ (_07005_, _06513_, _06512_);
  and _38841_ (_06515_, _06274_, _03237_);
  and _38842_ (_06516_, _06515_, _03060_);
  not _38843_ (_06517_, _06515_);
  and _38844_ (_06519_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _38845_ (_07009_, _06519_, _06516_);
  and _38846_ (_06520_, _06515_, _03067_);
  and _38847_ (_06522_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _38848_ (_07012_, _06522_, _06520_);
  and _38849_ (_06523_, _06515_, _03071_);
  and _38850_ (_06526_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _38851_ (_07015_, _06526_, _06523_);
  and _38852_ (_06527_, _06515_, _03074_);
  and _38853_ (_06529_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _38854_ (_07018_, _06529_, _06527_);
  and _38855_ (_06530_, _06515_, _03077_);
  and _38856_ (_06532_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _38857_ (_07021_, _06532_, _06530_);
  and _38858_ (_06534_, _06515_, _03080_);
  and _38859_ (_06535_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _38860_ (_07024_, _06535_, _06534_);
  and _38861_ (_06536_, _06515_, _03083_);
  and _38862_ (_06538_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _38863_ (_07027_, _06538_, _06536_);
  and _38864_ (_06539_, _06515_, _03087_);
  and _38865_ (_06541_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _38866_ (_07030_, _06541_, _06539_);
  and _38867_ (_06542_, _06274_, _03256_);
  and _38868_ (_06544_, _06542_, _03060_);
  not _38869_ (_06545_, _06542_);
  and _38870_ (_06546_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _38871_ (_07033_, _06546_, _06544_);
  and _38872_ (_06548_, _06542_, _03067_);
  and _38873_ (_06549_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _38874_ (_07036_, _06549_, _06548_);
  and _38875_ (_06551_, _06542_, _03071_);
  and _38876_ (_06552_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _38877_ (_07039_, _06552_, _06551_);
  and _38878_ (_06554_, _06542_, _03074_);
  and _38879_ (_06555_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _38880_ (_07042_, _06555_, _06554_);
  and _38881_ (_06557_, _06542_, _03077_);
  and _38882_ (_06559_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _38883_ (_07045_, _06559_, _06557_);
  and _38884_ (_06560_, _06542_, _03080_);
  and _38885_ (_06561_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _38886_ (_07048_, _06561_, _06560_);
  and _38887_ (_06563_, _06542_, _03083_);
  and _38888_ (_06564_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _38889_ (_07052_, _06564_, _06563_);
  and _38890_ (_06566_, _06542_, _03087_);
  and _38891_ (_06567_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _38892_ (_07054_, _06567_, _06566_);
  and _38893_ (_06569_, _06274_, _03275_);
  and _38894_ (_06570_, _06569_, _03060_);
  not _38895_ (_06572_, _06569_);
  and _38896_ (_06573_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or _38897_ (_07058_, _06573_, _06570_);
  and _38898_ (_06575_, _06569_, _03067_);
  and _38899_ (_06576_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or _38900_ (_07061_, _06576_, _06575_);
  and _38901_ (_06578_, _06569_, _03071_);
  and _38902_ (_06579_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or _38903_ (_07064_, _06579_, _06578_);
  and _38904_ (_06581_, _06569_, _03074_);
  and _38905_ (_06582_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or _38906_ (_07067_, _06582_, _06581_);
  and _38907_ (_06584_, _06569_, _03077_);
  and _38908_ (_06585_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or _38909_ (_07070_, _06585_, _06584_);
  and _38910_ (_06587_, _06569_, _03080_);
  and _38911_ (_06588_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or _38912_ (_07073_, _06588_, _06587_);
  and _38913_ (_06590_, _06569_, _03083_);
  and _38914_ (_06591_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or _38915_ (_07076_, _06591_, _06590_);
  and _38916_ (_06593_, _06569_, _03087_);
  and _38917_ (_06594_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or _38918_ (_07079_, _06594_, _06593_);
  and _38919_ (_06596_, _06274_, _03295_);
  and _38920_ (_06597_, _06596_, _03060_);
  not _38921_ (_06598_, _06596_);
  and _38922_ (_06600_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or _38923_ (_07083_, _06600_, _06597_);
  and _38924_ (_06601_, _06596_, _03067_);
  and _38925_ (_06603_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or _38926_ (_07086_, _06603_, _06601_);
  and _38927_ (_06604_, _06596_, _03071_);
  and _38928_ (_06606_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or _38929_ (_07089_, _06606_, _06604_);
  and _38930_ (_06608_, _06596_, _03074_);
  and _38931_ (_06609_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or _38932_ (_07092_, _06609_, _06608_);
  and _38933_ (_06610_, _06596_, _03077_);
  and _38934_ (_06612_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or _38935_ (_07095_, _06612_, _06610_);
  and _38936_ (_06613_, _06596_, _03080_);
  and _38937_ (_06615_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or _38938_ (_07098_, _06615_, _06613_);
  and _38939_ (_06616_, _06596_, _03083_);
  and _38940_ (_06618_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or _38941_ (_07101_, _06618_, _06616_);
  and _38942_ (_06619_, _06596_, _03087_);
  and _38943_ (_06621_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or _38944_ (_07103_, _06621_, _06619_);
  and _38945_ (_06622_, _06274_, _03315_);
  and _38946_ (_06624_, _06622_, _03060_);
  not _38947_ (_06625_, _06622_);
  and _38948_ (_06626_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _38949_ (_07107_, _06626_, _06624_);
  and _38950_ (_06628_, _06622_, _03067_);
  and _38951_ (_06629_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _38952_ (_07110_, _06629_, _06628_);
  and _38953_ (_06631_, _06622_, _03071_);
  and _38954_ (_06633_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _38955_ (_07113_, _06633_, _06631_);
  and _38956_ (_06634_, _06622_, _03074_);
  and _38957_ (_06635_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _38958_ (_07116_, _06635_, _06634_);
  and _38959_ (_06637_, _06622_, _03077_);
  and _38960_ (_06638_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _38961_ (_07119_, _06638_, _06637_);
  and _38962_ (_06640_, _06622_, _03080_);
  and _38963_ (_06641_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _38964_ (_07122_, _06641_, _06640_);
  and _38965_ (_06643_, _06622_, _03083_);
  and _38966_ (_06644_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _38967_ (_07125_, _06644_, _06643_);
  and _38968_ (_06646_, _06622_, _03087_);
  and _38969_ (_06647_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _38970_ (_07128_, _06647_, _06646_);
  and _38971_ (_06649_, _06274_, _03334_);
  and _38972_ (_06650_, _06649_, _03060_);
  not _38973_ (_06652_, _06649_);
  and _38974_ (_06653_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _38975_ (_07132_, _06653_, _06650_);
  and _38976_ (_06655_, _06649_, _03067_);
  and _38977_ (_06656_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _38978_ (_07135_, _06656_, _06655_);
  and _38979_ (_06658_, _06649_, _03071_);
  and _38980_ (_06659_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _38981_ (_07138_, _06659_, _06658_);
  and _38982_ (_06661_, _06649_, _03074_);
  and _38983_ (_06662_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _38984_ (_07141_, _06662_, _06661_);
  and _38985_ (_06664_, _06649_, _03077_);
  and _38986_ (_06665_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _38987_ (_07144_, _06665_, _06664_);
  and _38988_ (_06667_, _06649_, _03080_);
  and _38989_ (_06668_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _38990_ (_07147_, _06668_, _06667_);
  and _38991_ (_06670_, _06649_, _03083_);
  and _38992_ (_06671_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _38993_ (_07150_, _06671_, _06670_);
  and _38994_ (_06673_, _06649_, _03087_);
  and _38995_ (_06674_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _38996_ (_07153_, _06674_, _06673_);
  and _38997_ (_06676_, _06274_, _03353_);
  and _38998_ (_06677_, _06676_, _03060_);
  not _38999_ (_06678_, _06676_);
  and _39000_ (_06680_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or _39001_ (_07156_, _06680_, _06677_);
  and _39002_ (_06682_, _06676_, _03067_);
  and _39003_ (_06683_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or _39004_ (_07160_, _06683_, _06682_);
  and _39005_ (_06684_, _06676_, _03071_);
  and _39006_ (_06686_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or _39007_ (_07163_, _06686_, _06684_);
  and _39008_ (_06687_, _06676_, _03074_);
  and _39009_ (_06689_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or _39010_ (_07166_, _06689_, _06687_);
  and _39011_ (_06690_, _06676_, _03077_);
  and _39012_ (_06692_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or _39013_ (_07169_, _06692_, _06690_);
  and _39014_ (_06693_, _06676_, _03080_);
  and _39015_ (_06695_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or _39016_ (_07172_, _06695_, _06693_);
  and _39017_ (_06696_, _06676_, _03083_);
  and _39018_ (_06698_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or _39019_ (_07175_, _06698_, _06696_);
  and _39020_ (_06699_, _06676_, _03087_);
  and _39021_ (_06701_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or _39022_ (_07177_, _06701_, _06699_);
  and _39023_ (_06702_, _03373_, _26459_);
  and _39024_ (_06704_, _06702_, _02963_);
  and _39025_ (_06705_, _06704_, _03060_);
  not _39026_ (_06707_, _06704_);
  and _39027_ (_06708_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or _39028_ (_07182_, _06708_, _06705_);
  and _39029_ (_06709_, _06704_, _03067_);
  and _39030_ (_06711_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or _39031_ (_07185_, _06711_, _06709_);
  and _39032_ (_06712_, _06704_, _03071_);
  and _39033_ (_06714_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or _39034_ (_07188_, _06714_, _06712_);
  and _39035_ (_06715_, _06704_, _03074_);
  and _39036_ (_06717_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or _39037_ (_07191_, _06717_, _06715_);
  and _39038_ (_06718_, _06704_, _03077_);
  and _39039_ (_06720_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or _39040_ (_07194_, _06720_, _06718_);
  and _39041_ (_06721_, _06704_, _03080_);
  and _39042_ (_06723_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or _39043_ (_07197_, _06723_, _06721_);
  and _39044_ (_06724_, _06704_, _03083_);
  and _39045_ (_06726_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or _39046_ (_07200_, _06726_, _06724_);
  and _39047_ (_06727_, _06704_, _03087_);
  and _39048_ (_06729_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or _39049_ (_07203_, _06729_, _06727_);
  and _39050_ (_06731_, _06702_, _03062_);
  and _39051_ (_06732_, _06731_, _03060_);
  not _39052_ (_06733_, _06731_);
  and _39053_ (_06734_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _39054_ (_07206_, _06734_, _06732_);
  and _39055_ (_06736_, _06731_, _03067_);
  and _39056_ (_06737_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _39057_ (_07209_, _06737_, _06736_);
  and _39058_ (_06739_, _06731_, _03071_);
  and _39059_ (_06740_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _39060_ (_07213_, _06740_, _06739_);
  and _39061_ (_06742_, _06731_, _03074_);
  and _39062_ (_06743_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _39063_ (_07216_, _06743_, _06742_);
  and _39064_ (_06745_, _06731_, _03077_);
  and _39065_ (_06746_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _39066_ (_07219_, _06746_, _06745_);
  and _39067_ (_06748_, _06731_, _03080_);
  and _39068_ (_06749_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _39069_ (_07222_, _06749_, _06748_);
  and _39070_ (_06751_, _06731_, _03083_);
  and _39071_ (_06752_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _39072_ (_07225_, _06752_, _06751_);
  and _39073_ (_06754_, _06731_, _03087_);
  and _39074_ (_06756_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _39075_ (_07227_, _06756_, _06754_);
  and _39076_ (_06757_, _06702_, _03091_);
  and _39077_ (_06758_, _06757_, _03060_);
  not _39078_ (_06760_, _06757_);
  and _39079_ (_06761_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _39080_ (_07231_, _06761_, _06758_);
  and _39081_ (_06763_, _06757_, _03067_);
  and _39082_ (_06764_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _39083_ (_07234_, _06764_, _06763_);
  and _39084_ (_06766_, _06757_, _03071_);
  and _39085_ (_06767_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _39086_ (_07237_, _06767_, _06766_);
  and _39087_ (_06769_, _06757_, _03074_);
  and _39088_ (_06770_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _39089_ (_07241_, _06770_, _06769_);
  and _39090_ (_06772_, _06757_, _03077_);
  and _39091_ (_06773_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _39092_ (_07244_, _06773_, _06772_);
  and _39093_ (_06775_, _06757_, _03080_);
  and _39094_ (_06776_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _39095_ (_07247_, _06776_, _06775_);
  and _39096_ (_06778_, _06757_, _03083_);
  and _39097_ (_06779_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _39098_ (_07250_, _06779_, _06778_);
  and _39099_ (_06781_, _06757_, _03087_);
  and _39100_ (_06782_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _39101_ (_07252_, _06782_, _06781_);
  and _39102_ (_06783_, _06702_, _03113_);
  and _39103_ (_06784_, _06783_, _03060_);
  not _39104_ (_06785_, _06783_);
  and _39105_ (_06786_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or _39106_ (_07256_, _06786_, _06784_);
  and _39107_ (_06788_, _06783_, _03067_);
  and _39108_ (_06789_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or _39109_ (_07259_, _06789_, _06788_);
  and _39110_ (_06791_, _06783_, _03071_);
  and _39111_ (_06792_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or _39112_ (_07262_, _06792_, _06791_);
  and _39113_ (_06794_, _06783_, _03074_);
  and _39114_ (_06795_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or _39115_ (_07265_, _06795_, _06794_);
  and _39116_ (_06797_, _06783_, _03077_);
  and _39117_ (_06798_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or _39118_ (_07268_, _06798_, _06797_);
  and _39119_ (_06800_, _06783_, _03080_);
  and _39120_ (_06801_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or _39121_ (_07271_, _06801_, _06800_);
  and _39122_ (_06803_, _06783_, _03083_);
  and _39123_ (_06804_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or _39124_ (_07274_, _06804_, _06803_);
  and _39125_ (_06806_, _06783_, _03087_);
  and _39126_ (_06807_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or _39127_ (_07277_, _06807_, _06806_);
  and _39128_ (_06809_, _06702_, _03136_);
  and _39129_ (_06810_, _06809_, _03060_);
  not _39130_ (_06811_, _06809_);
  and _39131_ (_06813_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or _39132_ (_07280_, _06813_, _06810_);
  and _39133_ (_06814_, _06809_, _03067_);
  and _39134_ (_06816_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or _39135_ (_07283_, _06816_, _06814_);
  and _39136_ (_06817_, _06809_, _03071_);
  and _39137_ (_06819_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or _39138_ (_07286_, _06819_, _06817_);
  and _39139_ (_06820_, _06809_, _03074_);
  and _39140_ (_06822_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or _39141_ (_07289_, _06822_, _06820_);
  and _39142_ (_06823_, _06809_, _03077_);
  and _39143_ (_06825_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or _39144_ (_07293_, _06825_, _06823_);
  and _39145_ (_06826_, _06809_, _03080_);
  and _39146_ (_06828_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or _39147_ (_07296_, _06828_, _06826_);
  and _39148_ (_06829_, _06809_, _03083_);
  and _39149_ (_06831_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or _39150_ (_07299_, _06831_, _06829_);
  and _39151_ (_06833_, _06809_, _03087_);
  and _39152_ (_06834_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or _39153_ (_07301_, _06834_, _06833_);
  and _39154_ (_06835_, _06702_, _03159_);
  and _39155_ (_06837_, _06835_, _03060_);
  not _39156_ (_06838_, _06835_);
  and _39157_ (_06839_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _39158_ (_07305_, _06839_, _06837_);
  and _39159_ (_06841_, _06835_, _03067_);
  and _39160_ (_06842_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _39161_ (_07308_, _06842_, _06841_);
  and _39162_ (_06844_, _06835_, _03071_);
  and _39163_ (_06845_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _39164_ (_07311_, _06845_, _06844_);
  and _39165_ (_06847_, _06835_, _03074_);
  and _39166_ (_06848_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _39167_ (_07314_, _06848_, _06847_);
  and _39168_ (_06850_, _06835_, _03077_);
  and _39169_ (_06851_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _39170_ (_07317_, _06851_, _06850_);
  and _39171_ (_06853_, _06835_, _03080_);
  and _39172_ (_06854_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _39173_ (_07321_, _06854_, _06853_);
  and _39174_ (_06856_, _06835_, _03083_);
  and _39175_ (_06858_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _39176_ (_07324_, _06858_, _06856_);
  and _39177_ (_06859_, _06835_, _03087_);
  and _39178_ (_06860_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _39179_ (_07326_, _06860_, _06859_);
  and _39180_ (_06862_, _06702_, _03179_);
  and _39181_ (_06863_, _06862_, _03060_);
  not _39182_ (_06865_, _06862_);
  and _39183_ (_06866_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _39184_ (_07330_, _06866_, _06863_);
  and _39185_ (_06868_, _06862_, _03067_);
  and _39186_ (_06869_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _39187_ (_07333_, _06869_, _06868_);
  and _39188_ (_06871_, _06862_, _03071_);
  and _39189_ (_06872_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _39190_ (_07336_, _06872_, _06871_);
  and _39191_ (_06874_, _06862_, _03074_);
  and _39192_ (_06875_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _39193_ (_07339_, _06875_, _06874_);
  and _39194_ (_06877_, _06862_, _03077_);
  and _39195_ (_06878_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _39196_ (_07342_, _06878_, _06877_);
  and _39197_ (_06880_, _06862_, _03080_);
  and _39198_ (_06881_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _39199_ (_07345_, _06881_, _06880_);
  and _39200_ (_06883_, _06862_, _03083_);
  and _39201_ (_06884_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _39202_ (_07348_, _06884_, _06883_);
  and _39203_ (_06886_, _06862_, _03087_);
  and _39204_ (_06887_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _39205_ (_07351_, _06887_, _06886_);
  and _39206_ (_06889_, _06702_, _03198_);
  and _39207_ (_06890_, _06889_, _03060_);
  not _39208_ (_06891_, _06889_);
  and _39209_ (_06893_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or _39210_ (_07354_, _06893_, _06890_);
  and _39211_ (_06894_, _06889_, _03067_);
  and _39212_ (_06896_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or _39213_ (_07357_, _06896_, _06894_);
  and _39214_ (_06897_, _06889_, _03071_);
  and _39215_ (_06899_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or _39216_ (_07360_, _06899_, _06897_);
  and _39217_ (_06900_, _06889_, _03074_);
  and _39218_ (_06902_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or _39219_ (_07363_, _06902_, _06900_);
  and _39220_ (_06903_, _06889_, _03077_);
  and _39221_ (_06905_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or _39222_ (_07366_, _06905_, _06903_);
  and _39223_ (_06907_, _06889_, _03080_);
  and _39224_ (_06908_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or _39225_ (_07369_, _06908_, _06907_);
  and _39226_ (_06909_, _06889_, _03083_);
  and _39227_ (_06911_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or _39228_ (_07373_, _06911_, _06909_);
  and _39229_ (_06912_, _06889_, _03087_);
  and _39230_ (_06914_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or _39231_ (_07375_, _06914_, _06912_);
  and _39232_ (_06915_, _06702_, _03218_);
  and _39233_ (_06917_, _06915_, _03060_);
  not _39234_ (_06918_, _06915_);
  and _39235_ (_06919_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _39236_ (_07379_, _06919_, _06917_);
  and _39237_ (_06921_, _06915_, _03067_);
  and _39238_ (_06922_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _39239_ (_07382_, _06922_, _06921_);
  and _39240_ (_06924_, _06915_, _03071_);
  and _39241_ (_06925_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _39242_ (_07385_, _06925_, _06924_);
  and _39243_ (_06927_, _06915_, _03074_);
  and _39244_ (_06928_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _39245_ (_07388_, _06928_, _06927_);
  and _39246_ (_06930_, _06915_, _03077_);
  and _39247_ (_06932_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _39248_ (_07391_, _06932_, _06930_);
  and _39249_ (_06933_, _06915_, _03080_);
  and _39250_ (_06934_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _39251_ (_07394_, _06934_, _06933_);
  and _39252_ (_06936_, _06915_, _03083_);
  and _39253_ (_06937_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _39254_ (_07397_, _06937_, _06936_);
  and _39255_ (_06939_, _06915_, _03087_);
  and _39256_ (_06940_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _39257_ (_07400_, _06940_, _06939_);
  and _39258_ (_06942_, _06702_, _03237_);
  and _39259_ (_06943_, _06942_, _03060_);
  not _39260_ (_06945_, _06942_);
  and _39261_ (_06946_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or _39262_ (_07404_, _06946_, _06943_);
  and _39263_ (_06948_, _06942_, _03067_);
  and _39264_ (_06949_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or _39265_ (_07407_, _06949_, _06948_);
  and _39266_ (_06951_, _06942_, _03071_);
  and _39267_ (_06952_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or _39268_ (_07410_, _06952_, _06951_);
  and _39269_ (_06954_, _06942_, _03074_);
  and _39270_ (_06955_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or _39271_ (_07413_, _06955_, _06954_);
  and _39272_ (_06957_, _06942_, _03077_);
  and _39273_ (_06958_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or _39274_ (_07416_, _06958_, _06957_);
  and _39275_ (_06960_, _06942_, _03080_);
  and _39276_ (_06961_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or _39277_ (_07419_, _06961_, _06960_);
  and _39278_ (_06963_, _06942_, _03083_);
  and _39279_ (_06964_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or _39280_ (_07422_, _06964_, _06963_);
  and _39281_ (_06966_, _06942_, _03087_);
  and _39282_ (_06967_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or _39283_ (_07424_, _06967_, _06966_);
  and _39284_ (_06969_, _06702_, _03256_);
  and _39285_ (_06970_, _06969_, _03060_);
  not _39286_ (_06971_, _06969_);
  and _39287_ (_06973_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or _39288_ (_07428_, _06973_, _06970_);
  and _39289_ (_06974_, _06969_, _03067_);
  and _39290_ (_06976_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or _39291_ (_07431_, _06976_, _06974_);
  and _39292_ (_06977_, _06969_, _03071_);
  and _39293_ (_06979_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or _39294_ (_07434_, _06979_, _06977_);
  and _39295_ (_06981_, _06969_, _03074_);
  and _39296_ (_06982_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or _39297_ (_07437_, _06982_, _06981_);
  and _39298_ (_06983_, _06969_, _03077_);
  and _39299_ (_06985_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or _39300_ (_07440_, _06985_, _06983_);
  and _39301_ (_06986_, _06969_, _03080_);
  and _39302_ (_06988_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or _39303_ (_07443_, _06988_, _06986_);
  and _39304_ (_06989_, _06969_, _03083_);
  and _39305_ (_06991_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or _39306_ (_07446_, _06991_, _06989_);
  and _39307_ (_06992_, _06969_, _03087_);
  and _39308_ (_06994_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or _39309_ (_07449_, _06994_, _06992_);
  and _39310_ (_06995_, _06702_, _03275_);
  and _39311_ (_06997_, _06995_, _03060_);
  not _39312_ (_06998_, _06995_);
  and _39313_ (_06999_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _39314_ (_07453_, _06999_, _06997_);
  and _39315_ (_07001_, _06995_, _03067_);
  and _39316_ (_07002_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _39317_ (_07456_, _07002_, _07001_);
  and _39318_ (_07004_, _06995_, _03071_);
  and _39319_ (_07006_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _39320_ (_07459_, _07006_, _07004_);
  and _39321_ (_07007_, _06995_, _03074_);
  and _39322_ (_07008_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _39323_ (_07462_, _07008_, _07007_);
  and _39324_ (_07010_, _06995_, _03077_);
  and _39325_ (_07011_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _39326_ (_07465_, _07011_, _07010_);
  and _39327_ (_07013_, _06995_, _03080_);
  and _39328_ (_07014_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _39329_ (_07468_, _07014_, _07013_);
  and _39330_ (_07016_, _06995_, _03083_);
  and _39331_ (_07017_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _39332_ (_07471_, _07017_, _07016_);
  and _39333_ (_07019_, _06995_, _03087_);
  and _39334_ (_07020_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _39335_ (_07473_, _07020_, _07019_);
  and _39336_ (_07022_, _06702_, _03295_);
  and _39337_ (_07023_, _07022_, _03060_);
  not _39338_ (_07025_, _07022_);
  and _39339_ (_07026_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _39340_ (_07477_, _07026_, _07023_);
  and _39341_ (_07028_, _07022_, _03067_);
  and _39342_ (_07029_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _39343_ (_07481_, _07029_, _07028_);
  and _39344_ (_07031_, _07022_, _03071_);
  and _39345_ (_07032_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _39346_ (_07484_, _07032_, _07031_);
  and _39347_ (_07034_, _07022_, _03074_);
  and _39348_ (_07035_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _39349_ (_07487_, _07035_, _07034_);
  and _39350_ (_07037_, _07022_, _03077_);
  and _39351_ (_07038_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _39352_ (_07490_, _07038_, _07037_);
  and _39353_ (_07040_, _07022_, _03080_);
  and _39354_ (_07041_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _39355_ (_07493_, _07041_, _07040_);
  and _39356_ (_07043_, _07022_, _03083_);
  and _39357_ (_07044_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _39358_ (_07496_, _07044_, _07043_);
  and _39359_ (_07046_, _07022_, _03087_);
  and _39360_ (_07047_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _39361_ (_07498_, _07047_, _07046_);
  and _39362_ (_07049_, _06702_, _03315_);
  and _39363_ (_07050_, _07049_, _03060_);
  not _39364_ (_07051_, _07049_);
  and _39365_ (_07053_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or _39366_ (_07502_, _07053_, _07050_);
  and _39367_ (_07055_, _07049_, _03067_);
  and _39368_ (_07056_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or _39369_ (_07505_, _07056_, _07055_);
  and _39370_ (_07057_, _07049_, _03071_);
  and _39371_ (_07059_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or _39372_ (_07508_, _07059_, _07057_);
  and _39373_ (_07060_, _07049_, _03074_);
  and _39374_ (_07062_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or _39375_ (_07511_, _07062_, _07060_);
  and _39376_ (_07063_, _07049_, _03077_);
  and _39377_ (_07065_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or _39378_ (_07514_, _07065_, _07063_);
  and _39379_ (_07066_, _07049_, _03080_);
  and _39380_ (_07068_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or _39381_ (_07517_, _07068_, _07066_);
  and _39382_ (_07069_, _07049_, _03083_);
  and _39383_ (_07071_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or _39384_ (_07520_, _07071_, _07069_);
  and _39385_ (_07072_, _07049_, _03087_);
  and _39386_ (_07074_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or _39387_ (_07523_, _07074_, _07072_);
  and _39388_ (_07075_, _06702_, _03334_);
  and _39389_ (_07077_, _07075_, _03060_);
  not _39390_ (_07078_, _07075_);
  and _39391_ (_07080_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or _39392_ (_07526_, _07080_, _07077_);
  and _39393_ (_07081_, _07075_, _03067_);
  and _39394_ (_07082_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or _39395_ (_07529_, _07082_, _07081_);
  and _39396_ (_07084_, _07075_, _03071_);
  and _39397_ (_07085_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or _39398_ (_07533_, _07085_, _07084_);
  and _39399_ (_07087_, _07075_, _03074_);
  and _39400_ (_07088_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or _39401_ (_07536_, _07088_, _07087_);
  and _39402_ (_07090_, _07075_, _03077_);
  and _39403_ (_07091_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or _39404_ (_07539_, _07091_, _07090_);
  and _39405_ (_07093_, _07075_, _03080_);
  and _39406_ (_07094_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or _39407_ (_07542_, _07094_, _07093_);
  and _39408_ (_07096_, _07075_, _03083_);
  and _39409_ (_07097_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or _39410_ (_07545_, _07097_, _07096_);
  and _39411_ (_07099_, _07075_, _03087_);
  and _39412_ (_07100_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or _39413_ (_07547_, _07100_, _07099_);
  and _39414_ (_07102_, _06702_, _03353_);
  and _39415_ (_07104_, _07102_, _03060_);
  not _39416_ (_07105_, _07102_);
  and _39417_ (_07106_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _39418_ (_07551_, _07106_, _07104_);
  and _39419_ (_07108_, _07102_, _03067_);
  and _39420_ (_07109_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _39421_ (_07554_, _07109_, _07108_);
  and _39422_ (_07111_, _07102_, _03071_);
  and _39423_ (_07112_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _39424_ (_07557_, _07112_, _07111_);
  and _39425_ (_07114_, _07102_, _03074_);
  and _39426_ (_07115_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _39427_ (_07561_, _07115_, _07114_);
  and _39428_ (_07117_, _07102_, _03077_);
  and _39429_ (_07118_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _39430_ (_07564_, _07118_, _07117_);
  and _39431_ (_07120_, _07102_, _03080_);
  and _39432_ (_07121_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _39433_ (_07567_, _07121_, _07120_);
  and _39434_ (_07123_, _07102_, _03083_);
  and _39435_ (_07124_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _39436_ (_07570_, _07124_, _07123_);
  and _39437_ (_07126_, _07102_, _03087_);
  and _39438_ (_07127_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _39439_ (_07572_, _07127_, _07126_);
  and _39440_ (_07129_, _03699_, _26459_);
  and _39441_ (_07130_, _07129_, _02963_);
  and _39442_ (_07131_, _07130_, _03060_);
  not _39443_ (_07133_, _07130_);
  and _39444_ (_07134_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _39445_ (_07577_, _07134_, _07131_);
  and _39446_ (_07136_, _07130_, _03067_);
  and _39447_ (_07137_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _39448_ (_07580_, _07137_, _07136_);
  and _39449_ (_07139_, _07130_, _03071_);
  and _39450_ (_07140_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _39451_ (_07583_, _07140_, _07139_);
  and _39452_ (_07142_, _07130_, _03074_);
  and _39453_ (_07143_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _39454_ (_07586_, _07143_, _07142_);
  and _39455_ (_07145_, _07130_, _03077_);
  and _39456_ (_07146_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _39457_ (_07589_, _07146_, _07145_);
  and _39458_ (_07148_, _07130_, _03080_);
  and _39459_ (_07149_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _39460_ (_07592_, _07149_, _07148_);
  and _39461_ (_07151_, _07130_, _03083_);
  and _39462_ (_07152_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _39463_ (_07595_, _07152_, _07151_);
  and _39464_ (_07154_, _07130_, _03087_);
  and _39465_ (_07155_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _39466_ (_07598_, _07155_, _07154_);
  and _39467_ (_07157_, _07129_, _03062_);
  and _39468_ (_07158_, _07157_, _03060_);
  not _39469_ (_07159_, _07157_);
  and _39470_ (_07161_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  or _39471_ (_07601_, _07161_, _07158_);
  and _39472_ (_07162_, _07157_, _03067_);
  and _39473_ (_07164_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  or _39474_ (_07604_, _07164_, _07162_);
  and _39475_ (_07165_, _07157_, _03071_);
  and _39476_ (_07167_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  or _39477_ (_07607_, _07167_, _07165_);
  and _39478_ (_07168_, _07157_, _03074_);
  and _39479_ (_07170_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  or _39480_ (_07610_, _07170_, _07168_);
  and _39481_ (_07171_, _07157_, _03077_);
  and _39482_ (_07173_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  or _39483_ (_07614_, _07173_, _07171_);
  and _39484_ (_07174_, _07157_, _03080_);
  and _39485_ (_07176_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  or _39486_ (_07617_, _07176_, _07174_);
  and _39487_ (_07178_, _07157_, _03083_);
  and _39488_ (_07179_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  or _39489_ (_07620_, _07179_, _07178_);
  and _39490_ (_07180_, _07157_, _03087_);
  and _39491_ (_07181_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  or _39492_ (_07622_, _07181_, _07180_);
  and _39493_ (_07183_, _07129_, _03091_);
  and _39494_ (_07184_, _07183_, _03060_);
  not _39495_ (_07186_, _07183_);
  and _39496_ (_07187_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  or _39497_ (_07626_, _07187_, _07184_);
  and _39498_ (_07189_, _07183_, _03067_);
  and _39499_ (_07190_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  or _39500_ (_07629_, _07190_, _07189_);
  and _39501_ (_07192_, _07183_, _03071_);
  and _39502_ (_07193_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  or _39503_ (_07632_, _07193_, _07192_);
  and _39504_ (_07195_, _07183_, _03074_);
  and _39505_ (_07196_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  or _39506_ (_07635_, _07196_, _07195_);
  and _39507_ (_07198_, _07183_, _03077_);
  and _39508_ (_07199_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  or _39509_ (_07638_, _07199_, _07198_);
  and _39510_ (_07201_, _07183_, _03080_);
  and _39511_ (_07202_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  or _39512_ (_07642_, _07202_, _07201_);
  and _39513_ (_07204_, _07183_, _03083_);
  and _39514_ (_07205_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  or _39515_ (_07645_, _07205_, _07204_);
  and _39516_ (_07207_, _07183_, _03087_);
  and _39517_ (_07208_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  or _39518_ (_07647_, _07208_, _07207_);
  and _39519_ (_07210_, _07129_, _03113_);
  and _39520_ (_07211_, _07210_, _03060_);
  not _39521_ (_07212_, _07210_);
  and _39522_ (_07214_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _39523_ (_07651_, _07214_, _07211_);
  and _39524_ (_07215_, _07210_, _03067_);
  and _39525_ (_07217_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _39526_ (_07654_, _07217_, _07215_);
  and _39527_ (_07218_, _07210_, _03071_);
  and _39528_ (_07220_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _39529_ (_07657_, _07220_, _07218_);
  and _39530_ (_07221_, _07210_, _03074_);
  and _39531_ (_07223_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _39532_ (_07660_, _07223_, _07221_);
  and _39533_ (_07224_, _07210_, _03077_);
  and _39534_ (_07226_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _39535_ (_07663_, _07226_, _07224_);
  and _39536_ (_07228_, _07210_, _03080_);
  and _39537_ (_07229_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _39538_ (_07666_, _07229_, _07228_);
  and _39539_ (_07230_, _07210_, _03083_);
  and _39540_ (_07232_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _39541_ (_07669_, _07232_, _07230_);
  and _39542_ (_07233_, _07210_, _03087_);
  and _39543_ (_07235_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _39544_ (_07672_, _07235_, _07233_);
  and _39545_ (_07236_, _07129_, _03136_);
  and _39546_ (_07238_, _07236_, _03060_);
  not _39547_ (_07239_, _07236_);
  and _39548_ (_07240_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _39549_ (_07675_, _07240_, _07238_);
  and _39550_ (_07242_, _07236_, _03067_);
  and _39551_ (_07243_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _39552_ (_07678_, _07243_, _07242_);
  and _39553_ (_07245_, _07236_, _03071_);
  and _39554_ (_07246_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _39555_ (_07681_, _07246_, _07245_);
  and _39556_ (_07248_, _07236_, _03074_);
  and _39557_ (_07249_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _39558_ (_07684_, _07249_, _07248_);
  and _39559_ (_07251_, _07236_, _03077_);
  and _39560_ (_07253_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _39561_ (_07687_, _07253_, _07251_);
  and _39562_ (_07254_, _07236_, _03080_);
  and _39563_ (_07255_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _39564_ (_07690_, _07255_, _07254_);
  and _39565_ (_07257_, _07236_, _03083_);
  and _39566_ (_07258_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _39567_ (_07694_, _07258_, _07257_);
  and _39568_ (_07260_, _07236_, _03087_);
  and _39569_ (_07261_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _39570_ (_07696_, _07261_, _07260_);
  and _39571_ (_07263_, _07129_, _03159_);
  and _39572_ (_07264_, _07263_, _03060_);
  not _39573_ (_07266_, _07263_);
  and _39574_ (_07267_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  or _39575_ (_07700_, _07267_, _07264_);
  and _39576_ (_07269_, _07263_, _03067_);
  and _39577_ (_07270_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  or _39578_ (_07703_, _07270_, _07269_);
  and _39579_ (_07272_, _07263_, _03071_);
  and _39580_ (_07273_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  or _39581_ (_07706_, _07273_, _07272_);
  and _39582_ (_07275_, _07263_, _03074_);
  and _39583_ (_07276_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  or _39584_ (_07709_, _07276_, _07275_);
  and _39585_ (_07278_, _07263_, _03077_);
  and _39586_ (_07279_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  or _39587_ (_07712_, _07279_, _07278_);
  and _39588_ (_07281_, _07263_, _03080_);
  and _39589_ (_07282_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  or _39590_ (_07715_, _07282_, _07281_);
  and _39591_ (_07284_, _07263_, _03083_);
  and _39592_ (_07285_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  or _39593_ (_07718_, _07285_, _07284_);
  and _39594_ (_07287_, _07263_, _03087_);
  and _39595_ (_07288_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  or _39596_ (_07721_, _07288_, _07287_);
  and _39597_ (_07290_, _07129_, _03179_);
  and _39598_ (_07291_, _07290_, _03060_);
  not _39599_ (_07292_, _07290_);
  and _39600_ (_07294_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  or _39601_ (_07725_, _07294_, _07291_);
  and _39602_ (_07295_, _07290_, _03067_);
  and _39603_ (_07297_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  or _39604_ (_07728_, _07297_, _07295_);
  and _39605_ (_07298_, _07290_, _03071_);
  and _39606_ (_07300_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  or _39607_ (_07731_, _07300_, _07298_);
  and _39608_ (_07302_, _07290_, _03074_);
  and _39609_ (_07303_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  or _39610_ (_07734_, _07303_, _07302_);
  and _39611_ (_07304_, _07290_, _03077_);
  and _39612_ (_07306_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  or _39613_ (_07737_, _07306_, _07304_);
  and _39614_ (_07307_, _07290_, _03080_);
  and _39615_ (_07309_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  or _39616_ (_07740_, _07309_, _07307_);
  and _39617_ (_07310_, _07290_, _03083_);
  and _39618_ (_07312_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  or _39619_ (_07743_, _07312_, _07310_);
  and _39620_ (_07313_, _07290_, _03087_);
  and _39621_ (_07315_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  or _39622_ (_07745_, _07315_, _07313_);
  and _39623_ (_07316_, _07129_, _03198_);
  and _39624_ (_07318_, _07316_, _03060_);
  not _39625_ (_07319_, _07316_);
  and _39626_ (_07320_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _39627_ (_07749_, _07320_, _07318_);
  and _39628_ (_07322_, _07316_, _03067_);
  and _39629_ (_07323_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _39630_ (_07752_, _07323_, _07322_);
  and _39631_ (_07325_, _07316_, _03071_);
  and _39632_ (_07327_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _39633_ (_07755_, _07327_, _07325_);
  and _39634_ (_07328_, _07316_, _03074_);
  and _39635_ (_07329_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _39636_ (_07758_, _07329_, _07328_);
  and _39637_ (_07331_, _07316_, _03077_);
  and _39638_ (_07332_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _39639_ (_07761_, _07332_, _07331_);
  and _39640_ (_07334_, _07316_, _03080_);
  and _39641_ (_07335_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _39642_ (_07764_, _07335_, _07334_);
  and _39643_ (_07337_, _07316_, _03083_);
  and _39644_ (_07338_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _39645_ (_07767_, _07338_, _07337_);
  and _39646_ (_07340_, _07316_, _03087_);
  and _39647_ (_07341_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _39648_ (_07770_, _07341_, _07340_);
  and _39649_ (_07343_, _07129_, _03218_);
  and _39650_ (_07344_, _07343_, _03060_);
  not _39651_ (_07346_, _07343_);
  and _39652_ (_07347_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  or _39653_ (_07774_, _07347_, _07344_);
  and _39654_ (_07349_, _07343_, _03067_);
  and _39655_ (_07350_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  or _39656_ (_07777_, _07350_, _07349_);
  and _39657_ (_07352_, _07343_, _03071_);
  and _39658_ (_07353_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  or _39659_ (_07780_, _07353_, _07352_);
  and _39660_ (_07355_, _07343_, _03074_);
  and _39661_ (_07356_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  or _39662_ (_07783_, _07356_, _07355_);
  and _39663_ (_07358_, _07343_, _03077_);
  and _39664_ (_07359_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  or _39665_ (_07786_, _07359_, _07358_);
  and _39666_ (_07361_, _07343_, _03080_);
  and _39667_ (_07362_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  or _39668_ (_07789_, _07362_, _07361_);
  and _39669_ (_07364_, _07343_, _03083_);
  and _39670_ (_07365_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  or _39671_ (_07792_, _07365_, _07364_);
  and _39672_ (_07367_, _07343_, _03087_);
  and _39673_ (_07368_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  or _39674_ (_07794_, _07368_, _07367_);
  and _39675_ (_07370_, _07129_, _03237_);
  and _39676_ (_07371_, _07370_, _03060_);
  not _39677_ (_07372_, _07370_);
  and _39678_ (_07374_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _39679_ (_07798_, _07374_, _07371_);
  and _39680_ (_07376_, _07370_, _03067_);
  and _39681_ (_07377_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _39682_ (_07802_, _07377_, _07376_);
  and _39683_ (_07378_, _07370_, _03071_);
  and _39684_ (_07380_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _39685_ (_07805_, _07380_, _07378_);
  and _39686_ (_07381_, _07370_, _03074_);
  and _39687_ (_07383_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _39688_ (_07808_, _07383_, _07381_);
  and _39689_ (_07384_, _07370_, _03077_);
  and _39690_ (_07386_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _39691_ (_07811_, _07386_, _07384_);
  and _39692_ (_07387_, _07370_, _03080_);
  and _39693_ (_07389_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _39694_ (_07814_, _07389_, _07387_);
  and _39695_ (_07390_, _07370_, _03083_);
  and _39696_ (_07392_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _39697_ (_07817_, _07392_, _07390_);
  and _39698_ (_07393_, _07370_, _03087_);
  and _39699_ (_07395_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _39700_ (_07819_, _07395_, _07393_);
  and _39701_ (_07396_, _07129_, _03256_);
  and _39702_ (_07398_, _07396_, _03060_);
  not _39703_ (_07399_, _07396_);
  and _39704_ (_07401_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _39705_ (_07823_, _07401_, _07398_);
  and _39706_ (_07402_, _07396_, _03067_);
  and _39707_ (_07403_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _39708_ (_07826_, _07403_, _07402_);
  and _39709_ (_07405_, _07396_, _03071_);
  and _39710_ (_07406_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _39711_ (_07829_, _07406_, _07405_);
  and _39712_ (_07408_, _07396_, _03074_);
  and _39713_ (_07409_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _39714_ (_07832_, _07409_, _07408_);
  and _39715_ (_07411_, _07396_, _03077_);
  and _39716_ (_07412_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _39717_ (_07835_, _07412_, _07411_);
  and _39718_ (_07414_, _07396_, _03080_);
  and _39719_ (_07415_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _39720_ (_07838_, _07415_, _07414_);
  and _39721_ (_07417_, _07396_, _03083_);
  and _39722_ (_07418_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _39723_ (_07841_, _07418_, _07417_);
  and _39724_ (_07420_, _07396_, _03087_);
  and _39725_ (_07421_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _39726_ (_07844_, _07421_, _07420_);
  and _39727_ (_07423_, _07129_, _03275_);
  and _39728_ (_07425_, _07423_, _03060_);
  not _39729_ (_07426_, _07423_);
  and _39730_ (_07427_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  or _39731_ (_07847_, _07427_, _07425_);
  and _39732_ (_07429_, _07423_, _03067_);
  and _39733_ (_07430_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  or _39734_ (_07850_, _07430_, _07429_);
  and _39735_ (_07432_, _07423_, _03071_);
  and _39736_ (_07433_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  or _39737_ (_07854_, _07433_, _07432_);
  and _39738_ (_07435_, _07423_, _03074_);
  and _39739_ (_07436_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  or _39740_ (_07857_, _07436_, _07435_);
  and _39741_ (_07438_, _07423_, _03077_);
  and _39742_ (_07439_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  or _39743_ (_07860_, _07439_, _07438_);
  and _39744_ (_07441_, _07423_, _03080_);
  and _39745_ (_07442_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  or _39746_ (_07863_, _07442_, _07441_);
  and _39747_ (_07444_, _07423_, _03083_);
  and _39748_ (_07445_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  or _39749_ (_07866_, _07445_, _07444_);
  and _39750_ (_07447_, _07423_, _03087_);
  and _39751_ (_07448_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  or _39752_ (_07868_, _07448_, _07447_);
  and _39753_ (_07450_, _07129_, _03295_);
  and _39754_ (_07451_, _07450_, _03060_);
  not _39755_ (_07452_, _07450_);
  and _39756_ (_07454_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  or _39757_ (_07872_, _07454_, _07451_);
  and _39758_ (_07455_, _07450_, _03067_);
  and _39759_ (_07457_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  or _39760_ (_07875_, _07457_, _07455_);
  and _39761_ (_07458_, _07450_, _03071_);
  and _39762_ (_07460_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  or _39763_ (_07878_, _07460_, _07458_);
  and _39764_ (_07461_, _07450_, _03074_);
  and _39765_ (_07463_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  or _39766_ (_07882_, _07463_, _07461_);
  and _39767_ (_07464_, _07450_, _03077_);
  and _39768_ (_07466_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  or _39769_ (_07885_, _07466_, _07464_);
  and _39770_ (_07467_, _07450_, _03080_);
  and _39771_ (_07469_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  or _39772_ (_07888_, _07469_, _07467_);
  and _39773_ (_07470_, _07450_, _03083_);
  and _39774_ (_07472_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  or _39775_ (_07891_, _07472_, _07470_);
  and _39776_ (_07474_, _07450_, _03087_);
  and _39777_ (_07475_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or _39778_ (_07893_, _07475_, _07474_);
  and _39779_ (_07476_, _07129_, _03315_);
  and _39780_ (_07478_, _07476_, _03060_);
  not _39781_ (_07479_, _07476_);
  and _39782_ (_07480_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _39783_ (_07897_, _07480_, _07478_);
  and _39784_ (_07482_, _07476_, _03067_);
  and _39785_ (_07483_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _39786_ (_07900_, _07483_, _07482_);
  and _39787_ (_07485_, _07476_, _03071_);
  and _39788_ (_07486_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _39789_ (_07903_, _07486_, _07485_);
  and _39790_ (_07488_, _07476_, _03074_);
  and _39791_ (_07489_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _39792_ (_07906_, _07489_, _07488_);
  and _39793_ (_07491_, _07476_, _03077_);
  and _39794_ (_07492_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _39795_ (_07909_, _07492_, _07491_);
  and _39796_ (_07494_, _07476_, _03080_);
  and _39797_ (_07495_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _39798_ (_07912_, _07495_, _07494_);
  and _39799_ (_07497_, _07476_, _03083_);
  and _39800_ (_07499_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _39801_ (_07915_, _07499_, _07497_);
  and _39802_ (_07500_, _07476_, _03087_);
  and _39803_ (_07501_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _39804_ (_07918_, _07501_, _07500_);
  and _39805_ (_07503_, _07129_, _03334_);
  and _39806_ (_07504_, _07503_, _03060_);
  not _39807_ (_07506_, _07503_);
  and _39808_ (_07507_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _39809_ (_07921_, _07507_, _07504_);
  and _39810_ (_07509_, _07503_, _03067_);
  and _39811_ (_07510_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _39812_ (_07924_, _07510_, _07509_);
  and _39813_ (_07512_, _07503_, _03071_);
  and _39814_ (_07513_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _39815_ (_07927_, _07513_, _07512_);
  and _39816_ (_07515_, _07503_, _03074_);
  and _39817_ (_07516_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _39818_ (_07930_, _07516_, _07515_);
  and _39819_ (_07518_, _07503_, _03077_);
  and _39820_ (_07519_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _39821_ (_07934_, _07519_, _07518_);
  and _39822_ (_07521_, _07503_, _03080_);
  and _39823_ (_07522_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _39824_ (_07937_, _07522_, _07521_);
  and _39825_ (_07524_, _07503_, _03083_);
  and _39826_ (_07525_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _39827_ (_07940_, _07525_, _07524_);
  and _39828_ (_07527_, _07503_, _03087_);
  and _39829_ (_07528_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _39830_ (_07942_, _07528_, _07527_);
  and _39831_ (_07530_, _07129_, _03353_);
  and _39832_ (_07531_, _07530_, _03060_);
  not _39833_ (_07532_, _07530_);
  and _39834_ (_07534_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  or _39835_ (_07946_, _07534_, _07531_);
  and _39836_ (_07535_, _07530_, _03067_);
  and _39837_ (_07537_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  or _39838_ (_07949_, _07537_, _07535_);
  and _39839_ (_07538_, _07530_, _03071_);
  and _39840_ (_07540_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  or _39841_ (_07952_, _07540_, _07538_);
  and _39842_ (_07541_, _07530_, _03074_);
  and _39843_ (_07543_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  or _39844_ (_07955_, _07543_, _07541_);
  and _39845_ (_07544_, _07530_, _03077_);
  and _39846_ (_07546_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  or _39847_ (_07958_, _07546_, _07544_);
  and _39848_ (_07548_, _07530_, _03080_);
  and _39849_ (_07549_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  or _39850_ (_07962_, _07549_, _07548_);
  and _39851_ (_07550_, _07530_, _03083_);
  and _39852_ (_07552_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  or _39853_ (_07965_, _07552_, _07550_);
  and _39854_ (_07553_, _07530_, _03087_);
  and _39855_ (_07555_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  or _39856_ (_07967_, _07555_, _07553_);
  and _39857_ (_07556_, _04125_, _26459_);
  and _39858_ (_07558_, _07556_, _02963_);
  and _39859_ (_07559_, _07558_, _03060_);
  not _39860_ (_07560_, _07558_);
  and _39861_ (_07562_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or _39862_ (_07971_, _07562_, _07559_);
  and _39863_ (_07563_, _07558_, _03067_);
  and _39864_ (_07565_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or _39865_ (_07974_, _07565_, _07563_);
  and _39866_ (_07566_, _07558_, _03071_);
  and _39867_ (_07568_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or _39868_ (_07977_, _07568_, _07566_);
  and _39869_ (_07569_, _07558_, _03074_);
  and _39870_ (_07571_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or _39871_ (_07980_, _07571_, _07569_);
  and _39872_ (_07573_, _07558_, _03077_);
  and _39873_ (_07574_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or _39874_ (_07983_, _07574_, _07573_);
  and _39875_ (_07575_, _07558_, _03080_);
  and _39876_ (_07576_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _39877_ (_07987_, _07576_, _07575_);
  and _39878_ (_07578_, _07558_, _03083_);
  and _39879_ (_07579_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or _39880_ (_07991_, _07579_, _07578_);
  and _39881_ (_07581_, _07558_, _03087_);
  and _39882_ (_07582_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or _39883_ (_07993_, _07582_, _07581_);
  and _39884_ (_07584_, _07556_, _03062_);
  and _39885_ (_07585_, _07584_, _03060_);
  not _39886_ (_07587_, _07584_);
  and _39887_ (_07588_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _39888_ (_07997_, _07588_, _07585_);
  and _39889_ (_07590_, _07584_, _03067_);
  and _39890_ (_07591_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _39891_ (_08000_, _07591_, _07590_);
  and _39892_ (_07593_, _07584_, _03071_);
  and _39893_ (_07594_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _39894_ (_08003_, _07594_, _07593_);
  and _39895_ (_07596_, _07584_, _03074_);
  and _39896_ (_07597_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _39897_ (_08006_, _07597_, _07596_);
  and _39898_ (_07599_, _07584_, _03077_);
  and _39899_ (_07600_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _39900_ (_08009_, _07600_, _07599_);
  and _39901_ (_07602_, _07584_, _03080_);
  and _39902_ (_07603_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _39903_ (_08012_, _07603_, _07602_);
  and _39904_ (_07605_, _07584_, _03083_);
  and _39905_ (_07606_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _39906_ (_08015_, _07606_, _07605_);
  and _39907_ (_07608_, _07584_, _03087_);
  and _39908_ (_07609_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _39909_ (_08018_, _07609_, _07608_);
  and _39910_ (_07611_, _07556_, _03091_);
  and _39911_ (_07612_, _07611_, _03060_);
  not _39912_ (_07613_, _07611_);
  and _39913_ (_07615_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _39914_ (_08021_, _07615_, _07612_);
  and _39915_ (_07616_, _07611_, _03067_);
  and _39916_ (_07618_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _39917_ (_08024_, _07618_, _07616_);
  and _39918_ (_07619_, _07611_, _03071_);
  and _39919_ (_07621_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _39920_ (_08027_, _07621_, _07619_);
  and _39921_ (_07623_, _07611_, _03074_);
  and _39922_ (_07624_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _39923_ (_08030_, _07624_, _07623_);
  and _39924_ (_07625_, _07611_, _03077_);
  and _39925_ (_07627_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _39926_ (_08033_, _07627_, _07625_);
  and _39927_ (_07628_, _07611_, _03080_);
  and _39928_ (_07630_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _39929_ (_08036_, _07630_, _07628_);
  and _39930_ (_07631_, _07611_, _03083_);
  and _39931_ (_07633_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _39932_ (_08039_, _07633_, _07631_);
  and _39933_ (_07634_, _07611_, _03087_);
  and _39934_ (_07636_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _39935_ (_08042_, _07636_, _07634_);
  and _39936_ (_07637_, _07556_, _03113_);
  and _39937_ (_07639_, _07637_, _03060_);
  not _39938_ (_07640_, _07637_);
  and _39939_ (_07641_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or _39940_ (_08046_, _07641_, _07639_);
  and _39941_ (_07643_, _07637_, _03067_);
  and _39942_ (_07644_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or _39943_ (_08049_, _07644_, _07643_);
  and _39944_ (_07646_, _07637_, _03071_);
  and _39945_ (_07648_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or _39946_ (_08052_, _07648_, _07646_);
  and _39947_ (_07649_, _07637_, _03074_);
  and _39948_ (_07650_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or _39949_ (_08055_, _07650_, _07649_);
  and _39950_ (_07652_, _07637_, _03077_);
  and _39951_ (_07653_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or _39952_ (_08058_, _07653_, _07652_);
  and _39953_ (_07655_, _07637_, _03080_);
  and _39954_ (_07656_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or _39955_ (_08061_, _07656_, _07655_);
  and _39956_ (_07658_, _07637_, _03083_);
  and _39957_ (_07659_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or _39958_ (_08064_, _07659_, _07658_);
  and _39959_ (_07661_, _07637_, _03087_);
  and _39960_ (_07662_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _39961_ (_08066_, _07662_, _07661_);
  and _39962_ (_07664_, _07556_, _03136_);
  and _39963_ (_07665_, _07664_, _03060_);
  not _39964_ (_07667_, _07664_);
  and _39965_ (_07668_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or _39966_ (_08071_, _07668_, _07665_);
  and _39967_ (_07670_, _07664_, _03067_);
  and _39968_ (_07671_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or _39969_ (_08074_, _07671_, _07670_);
  and _39970_ (_07673_, _07664_, _03071_);
  and _39971_ (_07674_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or _39972_ (_08077_, _07674_, _07673_);
  and _39973_ (_07676_, _07664_, _03074_);
  and _39974_ (_07677_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or _39975_ (_08080_, _07677_, _07676_);
  and _39976_ (_07679_, _07664_, _03077_);
  and _39977_ (_07680_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or _39978_ (_08083_, _07680_, _07679_);
  and _39979_ (_07682_, _07664_, _03080_);
  and _39980_ (_07683_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or _39981_ (_08086_, _07683_, _07682_);
  and _39982_ (_07685_, _07664_, _03083_);
  and _39983_ (_07686_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or _39984_ (_08089_, _07686_, _07685_);
  and _39985_ (_07688_, _07664_, _03087_);
  and _39986_ (_07689_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or _39987_ (_08091_, _07689_, _07688_);
  and _39988_ (_07691_, _07556_, _03159_);
  and _39989_ (_07692_, _07691_, _03060_);
  not _39990_ (_07693_, _07691_);
  and _39991_ (_07695_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _39992_ (_08095_, _07695_, _07692_);
  and _39993_ (_07697_, _07691_, _03067_);
  and _39994_ (_07698_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _39995_ (_08098_, _07698_, _07697_);
  and _39996_ (_07699_, _07691_, _03071_);
  and _39997_ (_07701_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _39998_ (_08101_, _07701_, _07699_);
  and _39999_ (_07702_, _07691_, _03074_);
  and _40000_ (_07704_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _40001_ (_08104_, _07704_, _07702_);
  and _40002_ (_07705_, _07691_, _03077_);
  and _40003_ (_07707_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _40004_ (_08107_, _07707_, _07705_);
  and _40005_ (_07708_, _07691_, _03080_);
  and _40006_ (_07710_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _40007_ (_08110_, _07710_, _07708_);
  and _40008_ (_07711_, _07691_, _03083_);
  and _40009_ (_07713_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _40010_ (_08113_, _07713_, _07711_);
  and _40011_ (_07714_, _07691_, _03087_);
  and _40012_ (_07716_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _40013_ (_08116_, _07716_, _07714_);
  and _40014_ (_07717_, _07556_, _03179_);
  and _40015_ (_07719_, _07717_, _03060_);
  not _40016_ (_07720_, _07717_);
  and _40017_ (_07722_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _40018_ (_08119_, _07722_, _07719_);
  and _40019_ (_07723_, _07717_, _03067_);
  and _40020_ (_07724_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _40021_ (_08123_, _07724_, _07723_);
  and _40022_ (_07726_, _07717_, _03071_);
  and _40023_ (_07727_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _40024_ (_08126_, _07727_, _07726_);
  and _40025_ (_07729_, _07717_, _03074_);
  and _40026_ (_07730_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _40027_ (_08129_, _07730_, _07729_);
  and _40028_ (_07732_, _07717_, _03077_);
  and _40029_ (_07733_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _40030_ (_08132_, _07733_, _07732_);
  and _40031_ (_07735_, _07717_, _03080_);
  and _40032_ (_07736_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _40033_ (_08135_, _07736_, _07735_);
  and _40034_ (_07738_, _07717_, _03083_);
  and _40035_ (_07739_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _40036_ (_08138_, _07739_, _07738_);
  and _40037_ (_07741_, _07717_, _03087_);
  and _40038_ (_07742_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _40039_ (_08140_, _07742_, _07741_);
  and _40040_ (_07744_, _07556_, _03198_);
  and _40041_ (_07746_, _07744_, _03060_);
  not _40042_ (_07747_, _07744_);
  and _40043_ (_07748_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or _40044_ (_08144_, _07748_, _07746_);
  and _40045_ (_07750_, _07744_, _03067_);
  and _40046_ (_07751_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or _40047_ (_08147_, _07751_, _07750_);
  and _40048_ (_07753_, _07744_, _03071_);
  and _40049_ (_07754_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or _40050_ (_08151_, _07754_, _07753_);
  and _40051_ (_07756_, _07744_, _03074_);
  and _40052_ (_07757_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or _40053_ (_08154_, _07757_, _07756_);
  and _40054_ (_07759_, _07744_, _03077_);
  and _40055_ (_07760_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or _40056_ (_08157_, _07760_, _07759_);
  and _40057_ (_07762_, _07744_, _03080_);
  and _40058_ (_07763_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or _40059_ (_08160_, _07763_, _07762_);
  and _40060_ (_07765_, _07744_, _03083_);
  and _40061_ (_07766_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or _40062_ (_08163_, _07766_, _07765_);
  and _40063_ (_07768_, _07744_, _03087_);
  and _40064_ (_07769_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _40065_ (_08165_, _07769_, _07768_);
  and _40066_ (_07771_, _07556_, _03218_);
  and _40067_ (_07772_, _07771_, _03060_);
  not _40068_ (_07773_, _07771_);
  and _40069_ (_07775_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _40070_ (_08169_, _07775_, _07772_);
  and _40071_ (_07776_, _07771_, _03067_);
  and _40072_ (_07778_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _40073_ (_08172_, _07778_, _07776_);
  and _40074_ (_07779_, _07771_, _03071_);
  and _40075_ (_07781_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _40076_ (_08175_, _07781_, _07779_);
  and _40077_ (_07782_, _07771_, _03074_);
  and _40078_ (_07784_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _40079_ (_08178_, _07784_, _07782_);
  and _40080_ (_07785_, _07771_, _03077_);
  and _40081_ (_07787_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _40082_ (_08181_, _07787_, _07785_);
  and _40083_ (_07788_, _07771_, _03080_);
  and _40084_ (_07790_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _40085_ (_08184_, _07790_, _07788_);
  and _40086_ (_07791_, _07771_, _03083_);
  and _40087_ (_07793_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _40088_ (_08187_, _07793_, _07791_);
  and _40089_ (_07795_, _07771_, _03087_);
  and _40090_ (_07796_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _40091_ (_08190_, _07796_, _07795_);
  and _40092_ (_07797_, _07556_, _03237_);
  and _40093_ (_07799_, _07797_, _03060_);
  not _40094_ (_07800_, _07797_);
  and _40095_ (_07801_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or _40096_ (_08193_, _07801_, _07799_);
  and _40097_ (_07803_, _07797_, _03067_);
  and _40098_ (_07804_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or _40099_ (_08196_, _07804_, _07803_);
  and _40100_ (_07806_, _07797_, _03071_);
  and _40101_ (_07807_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or _40102_ (_08199_, _07807_, _07806_);
  and _40103_ (_07809_, _07797_, _03074_);
  and _40104_ (_07810_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or _40105_ (_08203_, _07810_, _07809_);
  and _40106_ (_07812_, _07797_, _03077_);
  and _40107_ (_07813_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or _40108_ (_08206_, _07813_, _07812_);
  and _40109_ (_07815_, _07797_, _03080_);
  and _40110_ (_07816_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or _40111_ (_08209_, _07816_, _07815_);
  and _40112_ (_07818_, _07797_, _03083_);
  and _40113_ (_07820_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or _40114_ (_08212_, _07820_, _07818_);
  and _40115_ (_07821_, _07797_, _03087_);
  and _40116_ (_07822_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or _40117_ (_08214_, _07822_, _07821_);
  and _40118_ (_07824_, _07556_, _03256_);
  and _40119_ (_07825_, _07824_, _03060_);
  not _40120_ (_07827_, _07824_);
  and _40121_ (_07828_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or _40122_ (_08218_, _07828_, _07825_);
  and _40123_ (_07830_, _07824_, _03067_);
  and _40124_ (_07831_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or _40125_ (_08221_, _07831_, _07830_);
  and _40126_ (_07833_, _07824_, _03071_);
  and _40127_ (_07834_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or _40128_ (_08224_, _07834_, _07833_);
  and _40129_ (_07836_, _07824_, _03074_);
  and _40130_ (_07837_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or _40131_ (_08227_, _07837_, _07836_);
  and _40132_ (_07839_, _07824_, _03077_);
  and _40133_ (_07840_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or _40134_ (_08231_, _07840_, _07839_);
  and _40135_ (_07842_, _07824_, _03080_);
  and _40136_ (_07843_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or _40137_ (_08234_, _07843_, _07842_);
  and _40138_ (_07845_, _07824_, _03083_);
  and _40139_ (_07846_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or _40140_ (_08237_, _07846_, _07845_);
  and _40141_ (_07848_, _07824_, _03087_);
  and _40142_ (_07849_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _40143_ (_08239_, _07849_, _07848_);
  and _40144_ (_07851_, _07556_, _03275_);
  and _40145_ (_07852_, _07851_, _03060_);
  not _40146_ (_07853_, _07851_);
  and _40147_ (_07855_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _40148_ (_08243_, _07855_, _07852_);
  and _40149_ (_07856_, _07851_, _03067_);
  and _40150_ (_07858_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _40151_ (_08246_, _07858_, _07856_);
  and _40152_ (_07859_, _07851_, _03071_);
  and _40153_ (_07861_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _40154_ (_08249_, _07861_, _07859_);
  and _40155_ (_07862_, _07851_, _03074_);
  and _40156_ (_07864_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _40157_ (_08252_, _07864_, _07862_);
  and _40158_ (_07865_, _07851_, _03077_);
  and _40159_ (_07867_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _40160_ (_08255_, _07867_, _07865_);
  and _40161_ (_07869_, _07851_, _03080_);
  and _40162_ (_07870_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _40163_ (_08258_, _07870_, _07869_);
  and _40164_ (_07871_, _07851_, _03083_);
  and _40165_ (_07873_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _40166_ (_08261_, _07873_, _07871_);
  and _40167_ (_07874_, _07851_, _03087_);
  and _40168_ (_07876_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _40169_ (_08264_, _07876_, _07874_);
  and _40170_ (_07877_, _07556_, _03295_);
  and _40171_ (_07879_, _07877_, _03060_);
  not _40172_ (_07880_, _07877_);
  and _40173_ (_07881_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _40174_ (_08267_, _07881_, _07879_);
  and _40175_ (_07883_, _07877_, _03067_);
  and _40176_ (_07884_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _40177_ (_08270_, _07884_, _07883_);
  and _40178_ (_07886_, _07877_, _03071_);
  and _40179_ (_07887_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _40180_ (_08273_, _07887_, _07886_);
  and _40181_ (_07889_, _07877_, _03074_);
  and _40182_ (_07890_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _40183_ (_08276_, _07890_, _07889_);
  and _40184_ (_07892_, _07877_, _03077_);
  and _40185_ (_07894_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _40186_ (_08279_, _07894_, _07892_);
  and _40187_ (_07895_, _07877_, _03080_);
  and _40188_ (_07896_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _40189_ (_08283_, _07896_, _07895_);
  and _40190_ (_07898_, _07877_, _03083_);
  and _40191_ (_07899_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _40192_ (_08286_, _07899_, _07898_);
  and _40193_ (_07901_, _07877_, _03087_);
  and _40194_ (_07902_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _40195_ (_08288_, _07902_, _07901_);
  and _40196_ (_07904_, _07556_, _03315_);
  and _40197_ (_07905_, _07904_, _03060_);
  not _40198_ (_07907_, _07904_);
  and _40199_ (_07908_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or _40200_ (_08292_, _07908_, _07905_);
  and _40201_ (_07910_, _07904_, _03067_);
  and _40202_ (_07911_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or _40203_ (_08295_, _07911_, _07910_);
  and _40204_ (_07913_, _07904_, _03071_);
  and _40205_ (_07914_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or _40206_ (_08298_, _07914_, _07913_);
  and _40207_ (_07916_, _07904_, _03074_);
  and _40208_ (_07917_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or _40209_ (_08301_, _07917_, _07916_);
  and _40210_ (_07919_, _07904_, _03077_);
  and _40211_ (_07920_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or _40212_ (_08304_, _07920_, _07919_);
  and _40213_ (_07922_, _07904_, _03080_);
  and _40214_ (_07923_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _40215_ (_08307_, _07923_, _07922_);
  and _40216_ (_07925_, _07904_, _03083_);
  and _40217_ (_07926_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or _40218_ (_08311_, _07926_, _07925_);
  and _40219_ (_07928_, _07904_, _03087_);
  and _40220_ (_07929_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _40221_ (_08313_, _07929_, _07928_);
  and _40222_ (_07931_, _07556_, _03334_);
  and _40223_ (_07932_, _07931_, _03060_);
  not _40224_ (_07933_, _07931_);
  and _40225_ (_07935_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or _40226_ (_08317_, _07935_, _07932_);
  and _40227_ (_07936_, _07931_, _03067_);
  and _40228_ (_07938_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or _40229_ (_08320_, _07938_, _07936_);
  and _40230_ (_07939_, _07931_, _03071_);
  and _40231_ (_07941_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or _40232_ (_08323_, _07941_, _07939_);
  and _40233_ (_07943_, _07931_, _03074_);
  and _40234_ (_07944_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or _40235_ (_08326_, _07944_, _07943_);
  and _40236_ (_07945_, _07931_, _03077_);
  and _40237_ (_07947_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or _40238_ (_08329_, _07947_, _07945_);
  and _40239_ (_07948_, _07931_, _03080_);
  and _40240_ (_07950_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or _40241_ (_08332_, _07950_, _07948_);
  and _40242_ (_07951_, _07931_, _03083_);
  and _40243_ (_07953_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or _40244_ (_08335_, _07953_, _07951_);
  and _40245_ (_07954_, _07931_, _03087_);
  and _40246_ (_07956_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or _40247_ (_08338_, _07956_, _07954_);
  and _40248_ (_07957_, _07556_, _03353_);
  and _40249_ (_07959_, _07957_, _03060_);
  not _40250_ (_07960_, _07957_);
  and _40251_ (_07961_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _40252_ (_08341_, _07961_, _07959_);
  and _40253_ (_07963_, _07957_, _03067_);
  and _40254_ (_07964_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _40255_ (_08344_, _07964_, _07963_);
  and _40256_ (_07966_, _07957_, _03071_);
  and _40257_ (_07968_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _40258_ (_08347_, _07968_, _07966_);
  and _40259_ (_07969_, _07957_, _03074_);
  and _40260_ (_07970_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _40261_ (_08350_, _07970_, _07969_);
  and _40262_ (_07972_, _07957_, _03077_);
  and _40263_ (_07973_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _40264_ (_08353_, _07973_, _07972_);
  and _40265_ (_07975_, _07957_, _03080_);
  and _40266_ (_07976_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _40267_ (_08356_, _07976_, _07975_);
  and _40268_ (_07978_, _07957_, _03083_);
  and _40269_ (_07979_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _40270_ (_08359_, _07979_, _07978_);
  and _40271_ (_07981_, _07957_, _03087_);
  and _40272_ (_07982_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _40273_ (_08362_, _07982_, _07981_);
  and _40274_ (_07984_, _02137_, _26939_);
  and _40275_ (_07985_, _07984_, _02966_);
  and _40276_ (_07986_, _07985_, _02963_);
  and _40277_ (_07988_, _07986_, _03060_);
  not _40278_ (_07989_, _07986_);
  and _40279_ (_07990_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _40280_ (_08367_, _07990_, _07988_);
  and _40281_ (_07992_, _07986_, _03067_);
  and _40282_ (_07994_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _40283_ (_08370_, _07994_, _07992_);
  and _40284_ (_07995_, _07986_, _03071_);
  and _40285_ (_07996_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _40286_ (_08373_, _07996_, _07995_);
  and _40287_ (_07998_, _07986_, _03074_);
  and _40288_ (_07999_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _40289_ (_08376_, _07999_, _07998_);
  and _40290_ (_08001_, _07986_, _03077_);
  and _40291_ (_08002_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _40292_ (_08379_, _08002_, _08001_);
  and _40293_ (_08004_, _07986_, _03080_);
  and _40294_ (_08005_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _40295_ (_08382_, _08005_, _08004_);
  and _40296_ (_08007_, _07986_, _03083_);
  and _40297_ (_08008_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _40298_ (_08385_, _08008_, _08007_);
  and _40299_ (_08010_, _07986_, _03087_);
  and _40300_ (_08011_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _40301_ (_08388_, _08011_, _08010_);
  and _40302_ (_08013_, _07985_, _03062_);
  and _40303_ (_08014_, _08013_, _03060_);
  not _40304_ (_08016_, _08013_);
  and _40305_ (_08017_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or _40306_ (_08392_, _08017_, _08014_);
  and _40307_ (_08019_, _08013_, _03067_);
  and _40308_ (_08020_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or _40309_ (_08395_, _08020_, _08019_);
  and _40310_ (_08022_, _08013_, _03071_);
  and _40311_ (_08023_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or _40312_ (_08398_, _08023_, _08022_);
  and _40313_ (_08025_, _08013_, _03074_);
  and _40314_ (_08026_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or _40315_ (_08401_, _08026_, _08025_);
  and _40316_ (_08028_, _08013_, _03077_);
  and _40317_ (_08029_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or _40318_ (_08404_, _08029_, _08028_);
  and _40319_ (_08031_, _08013_, _03080_);
  and _40320_ (_08032_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _40321_ (_08407_, _08032_, _08031_);
  and _40322_ (_08034_, _08013_, _03083_);
  and _40323_ (_08035_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or _40324_ (_08410_, _08035_, _08034_);
  and _40325_ (_08037_, _08013_, _03087_);
  and _40326_ (_08038_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or _40327_ (_08412_, _08038_, _08037_);
  and _40328_ (_08040_, _07985_, _03091_);
  and _40329_ (_08041_, _08040_, _03060_);
  not _40330_ (_08043_, _08040_);
  and _40331_ (_08044_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _40332_ (_08417_, _08044_, _08041_);
  and _40333_ (_08045_, _08040_, _03067_);
  and _40334_ (_08047_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or _40335_ (_08420_, _08047_, _08045_);
  and _40336_ (_08048_, _08040_, _03071_);
  and _40337_ (_08050_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or _40338_ (_08423_, _08050_, _08048_);
  and _40339_ (_08051_, _08040_, _03074_);
  and _40340_ (_08053_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or _40341_ (_08426_, _08053_, _08051_);
  and _40342_ (_08054_, _08040_, _03077_);
  and _40343_ (_08056_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or _40344_ (_08429_, _08056_, _08054_);
  and _40345_ (_08057_, _08040_, _03080_);
  and _40346_ (_08059_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or _40347_ (_08432_, _08059_, _08057_);
  and _40348_ (_08060_, _08040_, _03083_);
  and _40349_ (_08062_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or _40350_ (_08435_, _08062_, _08060_);
  and _40351_ (_08063_, _08040_, _03087_);
  and _40352_ (_08065_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or _40353_ (_08437_, _08065_, _08063_);
  and _40354_ (_08067_, _07985_, _03113_);
  and _40355_ (_08068_, _08067_, _03060_);
  not _40356_ (_08069_, _08067_);
  and _40357_ (_08070_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _40358_ (_08441_, _08070_, _08068_);
  and _40359_ (_08072_, _08067_, _03067_);
  and _40360_ (_08073_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _40361_ (_08445_, _08073_, _08072_);
  and _40362_ (_08075_, _08067_, _03071_);
  and _40363_ (_08076_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _40364_ (_08448_, _08076_, _08075_);
  and _40365_ (_08078_, _08067_, _03074_);
  and _40366_ (_08079_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _40367_ (_08451_, _08079_, _08078_);
  and _40368_ (_08081_, _08067_, _03077_);
  and _40369_ (_08082_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _40370_ (_08454_, _08082_, _08081_);
  and _40371_ (_08084_, _08067_, _03080_);
  and _40372_ (_08085_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _40373_ (_08457_, _08085_, _08084_);
  and _40374_ (_08087_, _08067_, _03083_);
  and _40375_ (_08088_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _40376_ (_08460_, _08088_, _08087_);
  and _40377_ (_08090_, _08067_, _03087_);
  and _40378_ (_08092_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _40379_ (_08462_, _08092_, _08090_);
  and _40380_ (_08093_, _07985_, _03136_);
  and _40381_ (_08094_, _08093_, _03060_);
  not _40382_ (_08096_, _08093_);
  and _40383_ (_08097_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _40384_ (_08466_, _08097_, _08094_);
  and _40385_ (_08099_, _08093_, _03067_);
  and _40386_ (_08100_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _40387_ (_08469_, _08100_, _08099_);
  and _40388_ (_08102_, _08093_, _03071_);
  and _40389_ (_08103_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _40390_ (_08472_, _08103_, _08102_);
  and _40391_ (_08105_, _08093_, _03074_);
  and _40392_ (_08106_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _40393_ (_08475_, _08106_, _08105_);
  and _40394_ (_08108_, _08093_, _03077_);
  and _40395_ (_08109_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _40396_ (_08478_, _08109_, _08108_);
  and _40397_ (_08111_, _08093_, _03080_);
  and _40398_ (_08112_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _40399_ (_08481_, _08112_, _08111_);
  and _40400_ (_08114_, _08093_, _03083_);
  and _40401_ (_08115_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _40402_ (_08484_, _08115_, _08114_);
  and _40403_ (_08117_, _08093_, _03087_);
  and _40404_ (_08118_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _40405_ (_08487_, _08118_, _08117_);
  and _40406_ (_08120_, _07985_, _03159_);
  and _40407_ (_08121_, _08120_, _03060_);
  not _40408_ (_08122_, _08120_);
  and _40409_ (_08124_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or _40410_ (_08490_, _08124_, _08121_);
  and _40411_ (_08125_, _08120_, _03067_);
  and _40412_ (_08127_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or _40413_ (_08493_, _08127_, _08125_);
  and _40414_ (_08128_, _08120_, _03071_);
  and _40415_ (_08130_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or _40416_ (_08497_, _08130_, _08128_);
  and _40417_ (_08131_, _08120_, _03074_);
  and _40418_ (_08133_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or _40419_ (_08500_, _08133_, _08131_);
  and _40420_ (_08134_, _08120_, _03077_);
  and _40421_ (_08136_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or _40422_ (_08503_, _08136_, _08134_);
  and _40423_ (_08137_, _08120_, _03080_);
  and _40424_ (_08139_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or _40425_ (_08506_, _08139_, _08137_);
  and _40426_ (_08141_, _08120_, _03083_);
  and _40427_ (_08142_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or _40428_ (_08509_, _08142_, _08141_);
  and _40429_ (_08143_, _08120_, _03087_);
  and _40430_ (_08145_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or _40431_ (_08511_, _08145_, _08143_);
  and _40432_ (_08146_, _07985_, _03179_);
  and _40433_ (_08148_, _08146_, _03060_);
  not _40434_ (_08149_, _08146_);
  and _40435_ (_08150_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _40436_ (_08515_, _08150_, _08148_);
  and _40437_ (_08152_, _08146_, _03067_);
  and _40438_ (_08153_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or _40439_ (_08518_, _08153_, _08152_);
  and _40440_ (_08155_, _08146_, _03071_);
  and _40441_ (_08156_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or _40442_ (_08521_, _08156_, _08155_);
  and _40443_ (_08158_, _08146_, _03074_);
  and _40444_ (_08159_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or _40445_ (_08525_, _08159_, _08158_);
  and _40446_ (_08161_, _08146_, _03077_);
  and _40447_ (_08162_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or _40448_ (_08528_, _08162_, _08161_);
  and _40449_ (_08164_, _08146_, _03080_);
  and _40450_ (_08166_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or _40451_ (_08531_, _08166_, _08164_);
  and _40452_ (_08167_, _08146_, _03083_);
  and _40453_ (_08168_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or _40454_ (_08534_, _08168_, _08167_);
  and _40455_ (_08170_, _08146_, _03087_);
  and _40456_ (_08171_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or _40457_ (_08536_, _08171_, _08170_);
  and _40458_ (_08173_, _07985_, _03198_);
  and _40459_ (_08174_, _08173_, _03060_);
  not _40460_ (_08176_, _08173_);
  and _40461_ (_08177_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _40462_ (_08540_, _08177_, _08174_);
  and _40463_ (_08179_, _08173_, _03067_);
  and _40464_ (_08180_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _40465_ (_08543_, _08180_, _08179_);
  and _40466_ (_08182_, _08173_, _03071_);
  and _40467_ (_08183_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _40468_ (_08546_, _08183_, _08182_);
  and _40469_ (_08185_, _08173_, _03074_);
  and _40470_ (_08186_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _40471_ (_08549_, _08186_, _08185_);
  and _40472_ (_08188_, _08173_, _03077_);
  and _40473_ (_08189_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _40474_ (_08552_, _08189_, _08188_);
  and _40475_ (_08191_, _08173_, _03080_);
  and _40476_ (_08192_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _40477_ (_08555_, _08192_, _08191_);
  and _40478_ (_08194_, _08173_, _03083_);
  and _40479_ (_08195_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _40480_ (_08558_, _08195_, _08194_);
  and _40481_ (_08197_, _08173_, _03087_);
  and _40482_ (_08198_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _40483_ (_08561_, _08198_, _08197_);
  and _40484_ (_08200_, _07985_, _03218_);
  and _40485_ (_08201_, _08200_, _03060_);
  not _40486_ (_08202_, _08200_);
  and _40487_ (_08204_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _40488_ (_08564_, _08204_, _08201_);
  and _40489_ (_08205_, _08200_, _03067_);
  and _40490_ (_08207_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or _40491_ (_08567_, _08207_, _08205_);
  and _40492_ (_08208_, _08200_, _03071_);
  and _40493_ (_08210_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or _40494_ (_08570_, _08210_, _08208_);
  and _40495_ (_08211_, _08200_, _03074_);
  and _40496_ (_08213_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or _40497_ (_08573_, _08213_, _08211_);
  and _40498_ (_08215_, _08200_, _03077_);
  and _40499_ (_08216_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or _40500_ (_08577_, _08216_, _08215_);
  and _40501_ (_08217_, _08200_, _03080_);
  and _40502_ (_08219_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or _40503_ (_08580_, _08219_, _08217_);
  and _40504_ (_08220_, _08200_, _03083_);
  and _40505_ (_08222_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or _40506_ (_08583_, _08222_, _08220_);
  and _40507_ (_08223_, _08200_, _03087_);
  and _40508_ (_08225_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _40509_ (_08585_, _08225_, _08223_);
  and _40510_ (_08226_, _07985_, _03237_);
  and _40511_ (_08228_, _08226_, _03060_);
  not _40512_ (_08229_, _08226_);
  and _40513_ (_08230_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _40514_ (_08589_, _08230_, _08228_);
  and _40515_ (_08232_, _08226_, _03067_);
  and _40516_ (_08233_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _40517_ (_08592_, _08233_, _08232_);
  and _40518_ (_08235_, _08226_, _03071_);
  and _40519_ (_08236_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _40520_ (_08595_, _08236_, _08235_);
  and _40521_ (_08238_, _08226_, _03074_);
  and _40522_ (_08240_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _40523_ (_08598_, _08240_, _08238_);
  and _40524_ (_08241_, _08226_, _03077_);
  and _40525_ (_08242_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _40526_ (_08601_, _08242_, _08241_);
  and _40527_ (_08244_, _08226_, _03080_);
  and _40528_ (_08245_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _40529_ (_08605_, _08245_, _08244_);
  and _40530_ (_08247_, _08226_, _03083_);
  and _40531_ (_08248_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _40532_ (_08608_, _08248_, _08247_);
  and _40533_ (_08250_, _08226_, _03087_);
  and _40534_ (_08251_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _40535_ (_08610_, _08251_, _08250_);
  and _40536_ (_08253_, _07985_, _03256_);
  and _40537_ (_08254_, _08253_, _03060_);
  not _40538_ (_08256_, _08253_);
  and _40539_ (_08257_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _40540_ (_08614_, _08257_, _08254_);
  and _40541_ (_08259_, _08253_, _03067_);
  and _40542_ (_08260_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _40543_ (_08617_, _08260_, _08259_);
  and _40544_ (_08262_, _08253_, _03071_);
  and _40545_ (_08263_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _40546_ (_08620_, _08263_, _08262_);
  and _40547_ (_08265_, _08253_, _03074_);
  and _40548_ (_08266_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _40549_ (_08623_, _08266_, _08265_);
  and _40550_ (_08268_, _08253_, _03077_);
  and _40551_ (_08269_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _40552_ (_08626_, _08269_, _08268_);
  and _40553_ (_08271_, _08253_, _03080_);
  and _40554_ (_08272_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _40555_ (_08629_, _08272_, _08271_);
  and _40556_ (_08274_, _08253_, _03083_);
  and _40557_ (_08275_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _40558_ (_08632_, _08275_, _08274_);
  and _40559_ (_08277_, _08253_, _03087_);
  and _40560_ (_08278_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _40561_ (_08635_, _08278_, _08277_);
  and _40562_ (_08280_, _07985_, _03275_);
  and _40563_ (_08281_, _08280_, _03060_);
  not _40564_ (_08282_, _08280_);
  and _40565_ (_08284_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or _40566_ (_08638_, _08284_, _08281_);
  and _40567_ (_08285_, _08280_, _03067_);
  and _40568_ (_08287_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or _40569_ (_08641_, _08287_, _08285_);
  and _40570_ (_08289_, _08280_, _03071_);
  and _40571_ (_08290_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or _40572_ (_08644_, _08290_, _08289_);
  and _40573_ (_08291_, _08280_, _03074_);
  and _40574_ (_08293_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or _40575_ (_08647_, _08293_, _08291_);
  and _40576_ (_08294_, _08280_, _03077_);
  and _40577_ (_08296_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or _40578_ (_08650_, _08296_, _08294_);
  and _40579_ (_08297_, _08280_, _03080_);
  and _40580_ (_08299_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or _40581_ (_08653_, _08299_, _08297_);
  and _40582_ (_08300_, _08280_, _03083_);
  and _40583_ (_08302_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or _40584_ (_08657_, _08302_, _08300_);
  and _40585_ (_08303_, _08280_, _03087_);
  and _40586_ (_08305_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or _40587_ (_08659_, _08305_, _08303_);
  and _40588_ (_08306_, _07985_, _03295_);
  and _40589_ (_08308_, _08306_, _03060_);
  not _40590_ (_08309_, _08306_);
  and _40591_ (_08310_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _40592_ (_08663_, _08310_, _08308_);
  and _40593_ (_08312_, _08306_, _03067_);
  and _40594_ (_08314_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or _40595_ (_08666_, _08314_, _08312_);
  and _40596_ (_08315_, _08306_, _03071_);
  and _40597_ (_08316_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or _40598_ (_08669_, _08316_, _08315_);
  and _40599_ (_08318_, _08306_, _03074_);
  and _40600_ (_08319_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or _40601_ (_08672_, _08319_, _08318_);
  and _40602_ (_08321_, _08306_, _03077_);
  and _40603_ (_08322_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or _40604_ (_08675_, _08322_, _08321_);
  and _40605_ (_08324_, _08306_, _03080_);
  and _40606_ (_08325_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or _40607_ (_08678_, _08325_, _08324_);
  and _40608_ (_08327_, _08306_, _03083_);
  and _40609_ (_08328_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or _40610_ (_08681_, _08328_, _08327_);
  and _40611_ (_08330_, _08306_, _03087_);
  and _40612_ (_08331_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or _40613_ (_08684_, _08331_, _08330_);
  and _40614_ (_08333_, _07985_, _03315_);
  and _40615_ (_08334_, _08333_, _03060_);
  not _40616_ (_08336_, _08333_);
  and _40617_ (_08337_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _40618_ (_08688_, _08337_, _08334_);
  and _40619_ (_08339_, _08333_, _03067_);
  and _40620_ (_08340_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _40621_ (_08691_, _08340_, _08339_);
  and _40622_ (_08342_, _08333_, _03071_);
  and _40623_ (_08343_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _40624_ (_08694_, _08343_, _08342_);
  and _40625_ (_08345_, _08333_, _03074_);
  and _40626_ (_08346_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _40627_ (_08697_, _08346_, _08345_);
  and _40628_ (_08348_, _08333_, _03077_);
  and _40629_ (_08349_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _40630_ (_08700_, _08349_, _08348_);
  and _40631_ (_08351_, _08333_, _03080_);
  and _40632_ (_08352_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _40633_ (_08703_, _08352_, _08351_);
  and _40634_ (_08354_, _08333_, _03083_);
  and _40635_ (_08355_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _40636_ (_08706_, _08355_, _08354_);
  and _40637_ (_08357_, _08333_, _03087_);
  and _40638_ (_08358_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _40639_ (_08708_, _08358_, _08357_);
  and _40640_ (_08360_, _07985_, _03334_);
  and _40641_ (_08361_, _08360_, _03060_);
  not _40642_ (_08363_, _08360_);
  and _40643_ (_08364_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _40644_ (_08712_, _08364_, _08361_);
  and _40645_ (_08365_, _08360_, _03067_);
  and _40646_ (_08366_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _40647_ (_08715_, _08366_, _08365_);
  and _40648_ (_08368_, _08360_, _03071_);
  and _40649_ (_08369_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _40650_ (_08718_, _08369_, _08368_);
  and _40651_ (_08371_, _08360_, _03074_);
  and _40652_ (_08372_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _40653_ (_08721_, _08372_, _08371_);
  and _40654_ (_08374_, _08360_, _03077_);
  and _40655_ (_08375_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _40656_ (_08724_, _08375_, _08374_);
  and _40657_ (_08377_, _08360_, _03080_);
  and _40658_ (_08378_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _40659_ (_08727_, _08378_, _08377_);
  and _40660_ (_08380_, _08360_, _03083_);
  and _40661_ (_08381_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _40662_ (_08730_, _08381_, _08380_);
  and _40663_ (_08383_, _08360_, _03087_);
  and _40664_ (_08384_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _40665_ (_08733_, _08384_, _08383_);
  and _40666_ (_08386_, _07985_, _03353_);
  and _40667_ (_08387_, _08386_, _03060_);
  not _40668_ (_08389_, _08386_);
  and _40669_ (_08390_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _40670_ (_08737_, _08390_, _08387_);
  and _40671_ (_08391_, _08386_, _03067_);
  and _40672_ (_08393_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or _40673_ (_08740_, _08393_, _08391_);
  and _40674_ (_08394_, _08386_, _03071_);
  and _40675_ (_08396_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or _40676_ (_08743_, _08396_, _08394_);
  and _40677_ (_08397_, _08386_, _03074_);
  and _40678_ (_08399_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or _40679_ (_08746_, _08399_, _08397_);
  and _40680_ (_08400_, _08386_, _03077_);
  and _40681_ (_08402_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or _40682_ (_08749_, _08402_, _08400_);
  and _40683_ (_08403_, _08386_, _03080_);
  and _40684_ (_08405_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or _40685_ (_08752_, _08405_, _08403_);
  and _40686_ (_08406_, _08386_, _03083_);
  and _40687_ (_08408_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or _40688_ (_08755_, _08408_, _08406_);
  and _40689_ (_08409_, _08386_, _03087_);
  and _40690_ (_08411_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or _40691_ (_08757_, _08411_, _08409_);
  and _40692_ (_08413_, _03373_, _26939_);
  and _40693_ (_08414_, _08413_, _02963_);
  and _40694_ (_08415_, _08414_, _03060_);
  not _40695_ (_08416_, _08414_);
  and _40696_ (_08418_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  or _40697_ (_08762_, _08418_, _08415_);
  and _40698_ (_08419_, _08414_, _03067_);
  and _40699_ (_08421_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  or _40700_ (_08765_, _08421_, _08419_);
  and _40701_ (_08422_, _08414_, _03071_);
  and _40702_ (_08424_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or _40703_ (_08768_, _08424_, _08422_);
  and _40704_ (_08425_, _08414_, _03074_);
  and _40705_ (_08427_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or _40706_ (_08771_, _08427_, _08425_);
  and _40707_ (_08428_, _08414_, _03077_);
  and _40708_ (_08430_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or _40709_ (_08774_, _08430_, _08428_);
  and _40710_ (_08431_, _08414_, _03080_);
  and _40711_ (_08433_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or _40712_ (_08777_, _08433_, _08431_);
  and _40713_ (_08434_, _08414_, _03083_);
  and _40714_ (_08436_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or _40715_ (_08780_, _08436_, _08434_);
  and _40716_ (_08438_, _08414_, _03087_);
  and _40717_ (_08439_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  or _40718_ (_08783_, _08439_, _08438_);
  and _40719_ (_08440_, _08413_, _03062_);
  and _40720_ (_08442_, _08440_, _03060_);
  not _40721_ (_08443_, _08440_);
  and _40722_ (_08444_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _40723_ (_08786_, _08444_, _08442_);
  and _40724_ (_08446_, _08440_, _03067_);
  and _40725_ (_08447_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _40726_ (_08790_, _08447_, _08446_);
  and _40727_ (_08449_, _08440_, _03071_);
  and _40728_ (_08450_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _40729_ (_08793_, _08450_, _08449_);
  and _40730_ (_08452_, _08440_, _03074_);
  and _40731_ (_08453_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _40732_ (_08796_, _08453_, _08452_);
  and _40733_ (_08455_, _08440_, _03077_);
  and _40734_ (_08456_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _40735_ (_08799_, _08456_, _08455_);
  and _40736_ (_08458_, _08440_, _03080_);
  and _40737_ (_08459_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _40738_ (_08802_, _08459_, _08458_);
  and _40739_ (_08461_, _08440_, _03083_);
  and _40740_ (_08463_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _40741_ (_08805_, _08463_, _08461_);
  and _40742_ (_08464_, _08440_, _03087_);
  and _40743_ (_08465_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _40744_ (_08807_, _08465_, _08464_);
  and _40745_ (_08467_, _08413_, _03091_);
  and _40746_ (_08468_, _08467_, _03060_);
  not _40747_ (_08470_, _08467_);
  and _40748_ (_08471_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _40749_ (_08811_, _08471_, _08468_);
  and _40750_ (_08473_, _08467_, _03067_);
  and _40751_ (_08474_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _40752_ (_08814_, _08474_, _08473_);
  and _40753_ (_08476_, _08467_, _03071_);
  and _40754_ (_08477_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _40755_ (_08818_, _08477_, _08476_);
  and _40756_ (_08479_, _08467_, _03074_);
  and _40757_ (_08480_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _40758_ (_08821_, _08480_, _08479_);
  and _40759_ (_08482_, _08467_, _03077_);
  and _40760_ (_08483_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _40761_ (_08824_, _08483_, _08482_);
  and _40762_ (_08485_, _08467_, _03080_);
  and _40763_ (_08486_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _40764_ (_08827_, _08486_, _08485_);
  and _40765_ (_08488_, _08467_, _03083_);
  and _40766_ (_08489_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _40767_ (_08830_, _08489_, _08488_);
  and _40768_ (_08491_, _08467_, _03087_);
  and _40769_ (_08492_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _40770_ (_08832_, _08492_, _08491_);
  and _40771_ (_08494_, _08413_, _03113_);
  and _40772_ (_08495_, _08494_, _03060_);
  not _40773_ (_08496_, _08494_);
  and _40774_ (_08498_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  or _40775_ (_08836_, _08498_, _08495_);
  and _40776_ (_08499_, _08494_, _03067_);
  and _40777_ (_08501_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  or _40778_ (_08839_, _08501_, _08499_);
  and _40779_ (_08502_, _08494_, _03071_);
  and _40780_ (_08504_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or _40781_ (_08843_, _08504_, _08502_);
  and _40782_ (_08505_, _08494_, _03074_);
  and _40783_ (_08507_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or _40784_ (_08847_, _08507_, _08505_);
  and _40785_ (_08508_, _08494_, _03077_);
  and _40786_ (_08510_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or _40787_ (_08850_, _08510_, _08508_);
  and _40788_ (_08512_, _08494_, _03080_);
  and _40789_ (_08513_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  or _40790_ (_08854_, _08513_, _08512_);
  and _40791_ (_08514_, _08494_, _03083_);
  and _40792_ (_08516_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or _40793_ (_08857_, _08516_, _08514_);
  and _40794_ (_08517_, _08494_, _03087_);
  and _40795_ (_08519_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or _40796_ (_08859_, _08519_, _08517_);
  and _40797_ (_08520_, _08413_, _03136_);
  and _40798_ (_08522_, _08520_, _03060_);
  not _40799_ (_08523_, _08520_);
  and _40800_ (_08524_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or _40801_ (_08863_, _08524_, _08522_);
  and _40802_ (_08526_, _08520_, _03067_);
  and _40803_ (_08527_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or _40804_ (_08867_, _08527_, _08526_);
  and _40805_ (_08529_, _08520_, _03071_);
  and _40806_ (_08530_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  or _40807_ (_08870_, _08530_, _08529_);
  and _40808_ (_08532_, _08520_, _03074_);
  and _40809_ (_08533_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  or _40810_ (_08873_, _08533_, _08532_);
  and _40811_ (_08535_, _08520_, _03077_);
  and _40812_ (_08537_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  or _40813_ (_08877_, _08537_, _08535_);
  and _40814_ (_08538_, _08520_, _03080_);
  and _40815_ (_08539_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or _40816_ (_08880_, _08539_, _08538_);
  and _40817_ (_08541_, _08520_, _03083_);
  and _40818_ (_08542_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  or _40819_ (_08883_, _08542_, _08541_);
  and _40820_ (_08544_, _08520_, _03087_);
  and _40821_ (_08545_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or _40822_ (_08886_, _08545_, _08544_);
  and _40823_ (_08547_, _08413_, _03159_);
  and _40824_ (_08548_, _08547_, _03060_);
  not _40825_ (_08550_, _08547_);
  and _40826_ (_08551_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _40827_ (_08890_, _08551_, _08548_);
  and _40828_ (_08553_, _08547_, _03067_);
  and _40829_ (_08554_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _40830_ (_08893_, _08554_, _08553_);
  and _40831_ (_08556_, _08547_, _03071_);
  and _40832_ (_08557_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _40833_ (_08896_, _08557_, _08556_);
  and _40834_ (_08559_, _08547_, _03074_);
  and _40835_ (_08560_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _40836_ (_08900_, _08560_, _08559_);
  and _40837_ (_08562_, _08547_, _03077_);
  and _40838_ (_08563_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _40839_ (_08904_, _08563_, _08562_);
  and _40840_ (_08565_, _08547_, _03080_);
  and _40841_ (_08566_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _40842_ (_08907_, _08566_, _08565_);
  and _40843_ (_08568_, _08547_, _03083_);
  and _40844_ (_08569_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _40845_ (_08911_, _08569_, _08568_);
  and _40846_ (_08571_, _08547_, _03087_);
  and _40847_ (_08572_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _40848_ (_08913_, _08572_, _08571_);
  and _40849_ (_08574_, _08413_, _03179_);
  and _40850_ (_08575_, _08574_, _03060_);
  not _40851_ (_08576_, _08574_);
  and _40852_ (_08578_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _40853_ (_08917_, _08578_, _08575_);
  and _40854_ (_08579_, _08574_, _03067_);
  and _40855_ (_08581_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _40856_ (_08920_, _08581_, _08579_);
  and _40857_ (_08582_, _08574_, _03071_);
  and _40858_ (_08584_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _40859_ (_08923_, _08584_, _08582_);
  and _40860_ (_08586_, _08574_, _03074_);
  and _40861_ (_08587_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _40862_ (_08926_, _08587_, _08586_);
  and _40863_ (_08588_, _08574_, _03077_);
  and _40864_ (_08590_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _40865_ (_08929_, _08590_, _08588_);
  and _40866_ (_08591_, _08574_, _03080_);
  and _40867_ (_08593_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _40868_ (_08933_, _08593_, _08591_);
  and _40869_ (_08594_, _08574_, _03083_);
  and _40870_ (_08596_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _40871_ (_08936_, _08596_, _08594_);
  and _40872_ (_08597_, _08574_, _03087_);
  and _40873_ (_08599_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _40874_ (_08938_, _08599_, _08597_);
  and _40875_ (_08600_, _08413_, _03198_);
  and _40876_ (_08602_, _08600_, _03060_);
  not _40877_ (_08603_, _08600_);
  and _40878_ (_08604_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  or _40879_ (_08942_, _08604_, _08602_);
  and _40880_ (_08606_, _08600_, _03067_);
  and _40881_ (_08607_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  or _40882_ (_08945_, _08607_, _08606_);
  and _40883_ (_08609_, _08600_, _03071_);
  and _40884_ (_08611_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or _40885_ (_08948_, _08611_, _08609_);
  and _40886_ (_08612_, _08600_, _03074_);
  and _40887_ (_08613_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or _40888_ (_08951_, _08613_, _08612_);
  and _40889_ (_08615_, _08600_, _03077_);
  and _40890_ (_08616_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or _40891_ (_08954_, _08616_, _08615_);
  and _40892_ (_08618_, _08600_, _03080_);
  and _40893_ (_08619_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  or _40894_ (_08957_, _08619_, _08618_);
  and _40895_ (_08621_, _08600_, _03083_);
  and _40896_ (_08622_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or _40897_ (_08960_, _08622_, _08621_);
  and _40898_ (_08624_, _08600_, _03087_);
  and _40899_ (_08625_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or _40900_ (_08963_, _08625_, _08624_);
  and _40901_ (_08627_, _08413_, _03218_);
  and _40902_ (_08628_, _08627_, _03060_);
  not _40903_ (_08630_, _08627_);
  and _40904_ (_08631_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _40905_ (_08966_, _08631_, _08628_);
  and _40906_ (_08633_, _08627_, _03067_);
  and _40907_ (_08634_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _40908_ (_08969_, _08634_, _08633_);
  and _40909_ (_08636_, _08627_, _03071_);
  and _40910_ (_08637_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _40911_ (_08972_, _08637_, _08636_);
  and _40912_ (_08639_, _08627_, _03074_);
  and _40913_ (_08640_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _40914_ (_08975_, _08640_, _08639_);
  and _40915_ (_08642_, _08627_, _03077_);
  and _40916_ (_08643_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _40917_ (_08978_, _08643_, _08642_);
  and _40918_ (_08645_, _08627_, _03080_);
  and _40919_ (_08646_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _40920_ (_08981_, _08646_, _08645_);
  and _40921_ (_08648_, _08627_, _03083_);
  and _40922_ (_08649_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _40923_ (_08985_, _08649_, _08648_);
  and _40924_ (_08651_, _08627_, _03087_);
  and _40925_ (_08652_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _40926_ (_08987_, _08652_, _08651_);
  and _40927_ (_08654_, _08413_, _03237_);
  and _40928_ (_08655_, _08654_, _03060_);
  not _40929_ (_08656_, _08654_);
  and _40930_ (_08658_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or _40931_ (_08991_, _08658_, _08655_);
  and _40932_ (_08660_, _08654_, _03067_);
  and _40933_ (_08661_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or _40934_ (_08994_, _08661_, _08660_);
  and _40935_ (_08662_, _08654_, _03071_);
  and _40936_ (_08664_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  or _40937_ (_08997_, _08664_, _08662_);
  and _40938_ (_08665_, _08654_, _03074_);
  and _40939_ (_08667_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or _40940_ (_09000_, _08667_, _08665_);
  and _40941_ (_08668_, _08654_, _03077_);
  and _40942_ (_08670_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or _40943_ (_09003_, _08670_, _08668_);
  and _40944_ (_08671_, _08654_, _03080_);
  and _40945_ (_08673_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or _40946_ (_09006_, _08673_, _08671_);
  and _40947_ (_08674_, _08654_, _03083_);
  and _40948_ (_08676_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or _40949_ (_09009_, _08676_, _08674_);
  and _40950_ (_08677_, _08654_, _03087_);
  and _40951_ (_08679_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or _40952_ (_09012_, _08679_, _08677_);
  and _40953_ (_08680_, _08413_, _03256_);
  and _40954_ (_08682_, _08680_, _03060_);
  not _40955_ (_08683_, _08680_);
  and _40956_ (_08685_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  or _40957_ (_09016_, _08685_, _08682_);
  and _40958_ (_08686_, _08680_, _03067_);
  and _40959_ (_08687_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  or _40960_ (_09019_, _08687_, _08686_);
  and _40961_ (_08689_, _08680_, _03071_);
  and _40962_ (_08690_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or _40963_ (_09022_, _08690_, _08689_);
  and _40964_ (_08692_, _08680_, _03074_);
  and _40965_ (_08693_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  or _40966_ (_09025_, _08693_, _08692_);
  and _40967_ (_08695_, _08680_, _03077_);
  and _40968_ (_08696_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  or _40969_ (_09028_, _08696_, _08695_);
  and _40970_ (_08698_, _08680_, _03080_);
  and _40971_ (_08699_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or _40972_ (_09031_, _08699_, _08698_);
  and _40973_ (_08701_, _08680_, _03083_);
  and _40974_ (_08702_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  or _40975_ (_09034_, _08702_, _08701_);
  and _40976_ (_08704_, _08680_, _03087_);
  and _40977_ (_08705_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  or _40978_ (_09036_, _08705_, _08704_);
  and _40979_ (_08707_, _08413_, _03275_);
  and _40980_ (_08709_, _08707_, _03060_);
  not _40981_ (_08710_, _08707_);
  and _40982_ (_08711_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _40983_ (_09040_, _08711_, _08709_);
  and _40984_ (_08713_, _08707_, _03067_);
  and _40985_ (_08714_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _40986_ (_09043_, _08714_, _08713_);
  and _40987_ (_08716_, _08707_, _03071_);
  and _40988_ (_08717_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _40989_ (_09046_, _08717_, _08716_);
  and _40990_ (_08719_, _08707_, _03074_);
  and _40991_ (_08720_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _40992_ (_09049_, _08720_, _08719_);
  and _40993_ (_08722_, _08707_, _03077_);
  and _40994_ (_08723_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _40995_ (_09052_, _08723_, _08722_);
  and _40996_ (_08725_, _08707_, _03080_);
  and _40997_ (_08726_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _40998_ (_09055_, _08726_, _08725_);
  and _40999_ (_08728_, _08707_, _03083_);
  and _41000_ (_08729_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _41001_ (_09058_, _08729_, _08728_);
  and _41002_ (_08731_, _08707_, _03087_);
  and _41003_ (_08732_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _41004_ (_09061_, _08732_, _08731_);
  and _41005_ (_08734_, _08413_, _03295_);
  and _41006_ (_08735_, _08734_, _03060_);
  not _41007_ (_08736_, _08734_);
  and _41008_ (_08738_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _41009_ (_09065_, _08738_, _08735_);
  and _41010_ (_08739_, _08734_, _03067_);
  and _41011_ (_08741_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _41012_ (_09068_, _08741_, _08739_);
  and _41013_ (_08742_, _08734_, _03071_);
  and _41014_ (_08744_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _41015_ (_09071_, _08744_, _08742_);
  and _41016_ (_08745_, _08734_, _03074_);
  and _41017_ (_08747_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _41018_ (_09074_, _08747_, _08745_);
  and _41019_ (_08748_, _08734_, _03077_);
  and _41020_ (_08750_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _41021_ (_09077_, _08750_, _08748_);
  and _41022_ (_08751_, _08734_, _03080_);
  and _41023_ (_08753_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _41024_ (_09080_, _08753_, _08751_);
  and _41025_ (_08754_, _08734_, _03083_);
  and _41026_ (_08756_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _41027_ (_09083_, _08756_, _08754_);
  and _41028_ (_08758_, _08734_, _03087_);
  and _41029_ (_08759_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _41030_ (_09085_, _08759_, _08758_);
  and _41031_ (_08760_, _08413_, _03315_);
  and _41032_ (_08761_, _08760_, _03060_);
  not _41033_ (_08763_, _08760_);
  and _41034_ (_08764_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or _41035_ (_09089_, _08764_, _08761_);
  and _41036_ (_08766_, _08760_, _03067_);
  and _41037_ (_08767_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or _41038_ (_09093_, _08767_, _08766_);
  and _41039_ (_08769_, _08760_, _03071_);
  and _41040_ (_08770_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or _41041_ (_09096_, _08770_, _08769_);
  and _41042_ (_08772_, _08760_, _03074_);
  and _41043_ (_08773_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or _41044_ (_09099_, _08773_, _08772_);
  and _41045_ (_08775_, _08760_, _03077_);
  and _41046_ (_08776_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  or _41047_ (_09102_, _08776_, _08775_);
  and _41048_ (_08778_, _08760_, _03080_);
  and _41049_ (_08779_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or _41050_ (_09105_, _08779_, _08778_);
  and _41051_ (_08781_, _08760_, _03083_);
  and _41052_ (_08782_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or _41053_ (_09108_, _08782_, _08781_);
  and _41054_ (_08784_, _08760_, _03087_);
  and _41055_ (_08785_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  or _41056_ (_09110_, _08785_, _08784_);
  and _41057_ (_08787_, _08413_, _03334_);
  and _41058_ (_08788_, _08787_, _03060_);
  not _41059_ (_08789_, _08787_);
  and _41060_ (_08791_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  or _41061_ (_09114_, _08791_, _08788_);
  and _41062_ (_08792_, _08787_, _03067_);
  and _41063_ (_08794_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  or _41064_ (_09117_, _08794_, _08792_);
  and _41065_ (_08795_, _08787_, _03071_);
  and _41066_ (_08797_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  or _41067_ (_09120_, _08797_, _08795_);
  and _41068_ (_08798_, _08787_, _03074_);
  and _41069_ (_08800_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  or _41070_ (_09123_, _08800_, _08798_);
  and _41071_ (_08801_, _08787_, _03077_);
  and _41072_ (_08803_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or _41073_ (_09126_, _08803_, _08801_);
  and _41074_ (_08804_, _08787_, _03080_);
  and _41075_ (_08806_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  or _41076_ (_09129_, _08806_, _08804_);
  and _41077_ (_08808_, _08787_, _03083_);
  and _41078_ (_08809_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  or _41079_ (_09132_, _08809_, _08808_);
  and _41080_ (_08810_, _08787_, _03087_);
  and _41081_ (_08812_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or _41082_ (_09135_, _08812_, _08810_);
  and _41083_ (_08813_, _08413_, _03353_);
  and _41084_ (_08815_, _08813_, _03060_);
  not _41085_ (_08816_, _08813_);
  and _41086_ (_08817_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _41087_ (_09138_, _08817_, _08815_);
  and _41088_ (_08819_, _08813_, _03067_);
  and _41089_ (_08820_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _41090_ (_09141_, _08820_, _08819_);
  and _41091_ (_08822_, _08813_, _03071_);
  and _41092_ (_08823_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _41093_ (_09145_, _08823_, _08822_);
  and _41094_ (_08825_, _08813_, _03074_);
  and _41095_ (_08826_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _41096_ (_09148_, _08826_, _08825_);
  and _41097_ (_08828_, _08813_, _03077_);
  and _41098_ (_08829_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _41099_ (_09151_, _08829_, _08828_);
  and _41100_ (_08831_, _08813_, _03080_);
  and _41101_ (_08833_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _41102_ (_09154_, _08833_, _08831_);
  and _41103_ (_08834_, _08813_, _03083_);
  and _41104_ (_08835_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _41105_ (_09157_, _08835_, _08834_);
  and _41106_ (_08837_, _08813_, _03087_);
  and _41107_ (_08838_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _41108_ (_09159_, _08838_, _08837_);
  and _41109_ (_08840_, _03699_, _26939_);
  and _41110_ (_08842_, _08840_, _02963_);
  and _41111_ (_08844_, _08842_, _03060_);
  not _41112_ (_08845_, _08842_);
  and _41113_ (_08846_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _41114_ (_09164_, _08846_, _08844_);
  and _41115_ (_08848_, _08842_, _03067_);
  and _41116_ (_08849_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _41117_ (_09167_, _08849_, _08848_);
  and _41118_ (_08851_, _08842_, _03071_);
  and _41119_ (_08852_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _41120_ (_09170_, _08852_, _08851_);
  and _41121_ (_08855_, _08842_, _03074_);
  and _41122_ (_08856_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _41123_ (_09173_, _08856_, _08855_);
  and _41124_ (_08858_, _08842_, _03077_);
  and _41125_ (_08860_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _41126_ (_09176_, _08860_, _08858_);
  and _41127_ (_08861_, _08842_, _03080_);
  and _41128_ (_08862_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _41129_ (_09179_, _08862_, _08861_);
  and _41130_ (_08865_, _08842_, _03083_);
  and _41131_ (_08866_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _41132_ (_09182_, _08866_, _08865_);
  and _41133_ (_08868_, _08842_, _03087_);
  and _41134_ (_08869_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _41135_ (_09185_, _08869_, _08868_);
  and _41136_ (_08871_, _08840_, _03062_);
  and _41137_ (_08872_, _08871_, _03060_);
  not _41138_ (_08874_, _08871_);
  and _41139_ (_08875_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or _41140_ (_09188_, _08875_, _08872_);
  and _41141_ (_08878_, _08871_, _03067_);
  and _41142_ (_08879_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or _41143_ (_09191_, _08879_, _08878_);
  and _41144_ (_08881_, _08871_, _03071_);
  and _41145_ (_08882_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or _41146_ (_09194_, _08882_, _08881_);
  and _41147_ (_08884_, _08871_, _03074_);
  and _41148_ (_08885_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or _41149_ (_09198_, _08885_, _08884_);
  and _41150_ (_08888_, _08871_, _03077_);
  and _41151_ (_08889_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or _41152_ (_09201_, _08889_, _08888_);
  and _41153_ (_08891_, _08871_, _03080_);
  and _41154_ (_08892_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or _41155_ (_09204_, _08892_, _08891_);
  and _41156_ (_08894_, _08871_, _03083_);
  and _41157_ (_08895_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or _41158_ (_09207_, _08895_, _08894_);
  and _41159_ (_08897_, _08871_, _03087_);
  and _41160_ (_08899_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or _41161_ (_09209_, _08899_, _08897_);
  and _41162_ (_08901_, _08840_, _03091_);
  and _41163_ (_08902_, _08901_, _03060_);
  not _41164_ (_08903_, _08901_);
  and _41165_ (_08905_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or _41166_ (_09213_, _08905_, _08902_);
  and _41167_ (_08906_, _08901_, _03067_);
  and _41168_ (_08908_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or _41169_ (_09216_, _08908_, _08906_);
  and _41170_ (_08910_, _08901_, _03071_);
  and _41171_ (_08912_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or _41172_ (_09219_, _08912_, _08910_);
  and _41173_ (_08914_, _08901_, _03074_);
  and _41174_ (_08915_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or _41175_ (_09222_, _08915_, _08914_);
  and _41176_ (_08916_, _08901_, _03077_);
  and _41177_ (_08918_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or _41178_ (_09226_, _08918_, _08916_);
  and _41179_ (_08919_, _08901_, _03080_);
  and _41180_ (_08921_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or _41181_ (_09229_, _08921_, _08919_);
  and _41182_ (_08922_, _08901_, _03083_);
  and _41183_ (_08924_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or _41184_ (_09232_, _08924_, _08922_);
  and _41185_ (_08925_, _08901_, _03087_);
  and _41186_ (_08927_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _41187_ (_09234_, _08927_, _08925_);
  and _41188_ (_08928_, _08840_, _03113_);
  and _41189_ (_08930_, _08928_, _03060_);
  not _41190_ (_08931_, _08928_);
  and _41191_ (_08932_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _41192_ (_09238_, _08932_, _08930_);
  and _41193_ (_08934_, _08928_, _03067_);
  and _41194_ (_08935_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _41195_ (_09241_, _08935_, _08934_);
  and _41196_ (_08937_, _08928_, _03071_);
  and _41197_ (_08939_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _41198_ (_09244_, _08939_, _08937_);
  and _41199_ (_08940_, _08928_, _03074_);
  and _41200_ (_08941_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _41201_ (_09247_, _08941_, _08940_);
  and _41202_ (_08943_, _08928_, _03077_);
  and _41203_ (_08944_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _41204_ (_09250_, _08944_, _08943_);
  and _41205_ (_08946_, _08928_, _03080_);
  and _41206_ (_08947_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _41207_ (_09253_, _08947_, _08946_);
  and _41208_ (_08949_, _08928_, _03083_);
  and _41209_ (_08950_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _41210_ (_09256_, _08950_, _08949_);
  and _41211_ (_08952_, _08928_, _03087_);
  and _41212_ (_08953_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _41213_ (_09259_, _08953_, _08952_);
  and _41214_ (_08955_, _08840_, _03136_);
  and _41215_ (_08956_, _08955_, _03060_);
  not _41216_ (_08958_, _08955_);
  and _41217_ (_08959_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _41218_ (_09262_, _08959_, _08956_);
  and _41219_ (_08961_, _08955_, _03067_);
  and _41220_ (_08962_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _41221_ (_09265_, _08962_, _08961_);
  and _41222_ (_08964_, _08955_, _03071_);
  and _41223_ (_08965_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _41224_ (_09268_, _08965_, _08964_);
  and _41225_ (_08967_, _08955_, _03074_);
  and _41226_ (_08968_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _41227_ (_09271_, _08968_, _08967_);
  and _41228_ (_08970_, _08955_, _03077_);
  and _41229_ (_08971_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _41230_ (_09274_, _08971_, _08970_);
  and _41231_ (_08973_, _08955_, _03080_);
  and _41232_ (_08974_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _41233_ (_09278_, _08974_, _08973_);
  and _41234_ (_08976_, _08955_, _03083_);
  and _41235_ (_08977_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _41236_ (_09281_, _08977_, _08976_);
  and _41237_ (_08979_, _08955_, _03087_);
  and _41238_ (_08980_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _41239_ (_09284_, _08980_, _08979_);
  and _41240_ (_08982_, _08840_, _03159_);
  and _41241_ (_08983_, _08982_, _03060_);
  not _41242_ (_08984_, _08982_);
  and _41243_ (_08986_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or _41244_ (_09287_, _08986_, _08983_);
  and _41245_ (_08988_, _08982_, _03067_);
  and _41246_ (_08989_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or _41247_ (_09290_, _08989_, _08988_);
  and _41248_ (_08990_, _08982_, _03071_);
  and _41249_ (_08992_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or _41250_ (_09293_, _08992_, _08990_);
  and _41251_ (_08993_, _08982_, _03074_);
  and _41252_ (_08995_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or _41253_ (_09296_, _08995_, _08993_);
  and _41254_ (_08996_, _08982_, _03077_);
  and _41255_ (_08998_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or _41256_ (_09299_, _08998_, _08996_);
  and _41257_ (_08999_, _08982_, _03080_);
  and _41258_ (_09001_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or _41259_ (_09302_, _09001_, _08999_);
  and _41260_ (_09002_, _08982_, _03083_);
  and _41261_ (_09004_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or _41262_ (_09306_, _09004_, _09002_);
  and _41263_ (_09005_, _08982_, _03087_);
  and _41264_ (_09007_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or _41265_ (_09308_, _09007_, _09005_);
  and _41266_ (_09008_, _08840_, _03179_);
  and _41267_ (_09010_, _09008_, _03060_);
  not _41268_ (_09011_, _09008_);
  and _41269_ (_09013_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or _41270_ (_09312_, _09013_, _09010_);
  and _41271_ (_09014_, _09008_, _03067_);
  and _41272_ (_09015_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or _41273_ (_09315_, _09015_, _09014_);
  and _41274_ (_09017_, _09008_, _03071_);
  and _41275_ (_09018_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or _41276_ (_09318_, _09018_, _09017_);
  and _41277_ (_09020_, _09008_, _03074_);
  and _41278_ (_09021_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or _41279_ (_09321_, _09021_, _09020_);
  and _41280_ (_09023_, _09008_, _03077_);
  and _41281_ (_09024_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or _41282_ (_09324_, _09024_, _09023_);
  and _41283_ (_09026_, _09008_, _03080_);
  and _41284_ (_09027_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _41285_ (_09327_, _09027_, _09026_);
  and _41286_ (_09029_, _09008_, _03083_);
  and _41287_ (_09030_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or _41288_ (_09330_, _09030_, _09029_);
  and _41289_ (_09032_, _09008_, _03087_);
  and _41290_ (_09033_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or _41291_ (_09333_, _09033_, _09032_);
  and _41292_ (_09035_, _08840_, _03198_);
  and _41293_ (_09037_, _09035_, _03060_);
  not _41294_ (_09038_, _09035_);
  and _41295_ (_09039_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _41296_ (_09337_, _09039_, _09037_);
  and _41297_ (_09041_, _09035_, _03067_);
  and _41298_ (_09042_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _41299_ (_09340_, _09042_, _09041_);
  and _41300_ (_09044_, _09035_, _03071_);
  and _41301_ (_09045_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _41302_ (_09343_, _09045_, _09044_);
  and _41303_ (_09047_, _09035_, _03074_);
  and _41304_ (_09048_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _41305_ (_09346_, _09048_, _09047_);
  and _41306_ (_09050_, _09035_, _03077_);
  and _41307_ (_09051_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _41308_ (_09349_, _09051_, _09050_);
  and _41309_ (_09053_, _09035_, _03080_);
  and _41310_ (_09054_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _41311_ (_09352_, _09054_, _09053_);
  and _41312_ (_09056_, _09035_, _03083_);
  and _41313_ (_09057_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _41314_ (_09355_, _09057_, _09056_);
  and _41315_ (_09059_, _09035_, _03087_);
  and _41316_ (_09060_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _41317_ (_09357_, _09060_, _09059_);
  and _41318_ (_09062_, _08840_, _03218_);
  and _41319_ (_09063_, _09062_, _03060_);
  not _41320_ (_09064_, _09062_);
  and _41321_ (_09066_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or _41322_ (_09361_, _09066_, _09063_);
  and _41323_ (_09067_, _09062_, _03067_);
  and _41324_ (_09069_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or _41325_ (_09364_, _09069_, _09067_);
  and _41326_ (_09070_, _09062_, _03071_);
  and _41327_ (_09072_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or _41328_ (_09367_, _09072_, _09070_);
  and _41329_ (_09073_, _09062_, _03074_);
  and _41330_ (_09075_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or _41331_ (_09370_, _09075_, _09073_);
  and _41332_ (_09076_, _09062_, _03077_);
  and _41333_ (_09078_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or _41334_ (_09373_, _09078_, _09076_);
  and _41335_ (_09079_, _09062_, _03080_);
  and _41336_ (_09081_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or _41337_ (_09376_, _09081_, _09079_);
  and _41338_ (_09082_, _09062_, _03083_);
  and _41339_ (_09084_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or _41340_ (_09379_, _09084_, _09082_);
  and _41341_ (_09086_, _09062_, _03087_);
  and _41342_ (_09087_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _41343_ (_09382_, _09087_, _09086_);
  and _41344_ (_09088_, _08840_, _03237_);
  and _41345_ (_09090_, _09088_, _03060_);
  not _41346_ (_09091_, _09088_);
  and _41347_ (_09092_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _41348_ (_09386_, _09092_, _09090_);
  and _41349_ (_09094_, _09088_, _03067_);
  and _41350_ (_09095_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _41351_ (_09389_, _09095_, _09094_);
  and _41352_ (_09097_, _09088_, _03071_);
  and _41353_ (_09098_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _41354_ (_09392_, _09098_, _09097_);
  and _41355_ (_09100_, _09088_, _03074_);
  and _41356_ (_09101_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _41357_ (_09395_, _09101_, _09100_);
  and _41358_ (_09103_, _09088_, _03077_);
  and _41359_ (_09104_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _41360_ (_09398_, _09104_, _09103_);
  and _41361_ (_09106_, _09088_, _03080_);
  and _41362_ (_09107_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _41363_ (_09401_, _09107_, _09106_);
  and _41364_ (_09109_, _09088_, _03083_);
  and _41365_ (_09111_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _41366_ (_09404_, _09111_, _09109_);
  and _41367_ (_09112_, _09088_, _03087_);
  and _41368_ (_09113_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _41369_ (_09406_, _09113_, _09112_);
  and _41370_ (_09115_, _08840_, _03256_);
  and _41371_ (_09116_, _09115_, _03060_);
  not _41372_ (_09118_, _09115_);
  and _41373_ (_09119_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _41374_ (_09410_, _09119_, _09116_);
  and _41375_ (_09121_, _09115_, _03067_);
  and _41376_ (_09122_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _41377_ (_09414_, _09122_, _09121_);
  and _41378_ (_09124_, _09115_, _03071_);
  and _41379_ (_09125_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _41380_ (_09417_, _09125_, _09124_);
  and _41381_ (_09127_, _09115_, _03074_);
  and _41382_ (_09128_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _41383_ (_09420_, _09128_, _09127_);
  and _41384_ (_09130_, _09115_, _03077_);
  and _41385_ (_09131_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _41386_ (_09423_, _09131_, _09130_);
  and _41387_ (_09133_, _09115_, _03080_);
  and _41388_ (_09134_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _41389_ (_09426_, _09134_, _09133_);
  and _41390_ (_09136_, _09115_, _03083_);
  and _41391_ (_09137_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _41392_ (_09429_, _09137_, _09136_);
  and _41393_ (_09139_, _09115_, _03087_);
  and _41394_ (_09140_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _41395_ (_09431_, _09140_, _09139_);
  and _41396_ (_09142_, _08840_, _03275_);
  and _41397_ (_09143_, _09142_, _03060_);
  not _41398_ (_09144_, _09142_);
  and _41399_ (_09146_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or _41400_ (_09435_, _09146_, _09143_);
  and _41401_ (_09147_, _09142_, _03067_);
  and _41402_ (_09149_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or _41403_ (_09438_, _09149_, _09147_);
  and _41404_ (_09150_, _09142_, _03071_);
  and _41405_ (_09152_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or _41406_ (_09441_, _09152_, _09150_);
  and _41407_ (_09153_, _09142_, _03074_);
  and _41408_ (_09155_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or _41409_ (_09444_, _09155_, _09153_);
  and _41410_ (_09156_, _09142_, _03077_);
  and _41411_ (_09158_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or _41412_ (_09447_, _09158_, _09156_);
  and _41413_ (_09160_, _09142_, _03080_);
  and _41414_ (_09161_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or _41415_ (_09450_, _09161_, _09160_);
  and _41416_ (_09162_, _09142_, _03083_);
  and _41417_ (_09163_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or _41418_ (_09453_, _09163_, _09162_);
  and _41419_ (_09165_, _09142_, _03087_);
  and _41420_ (_09166_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or _41421_ (_09456_, _09166_, _09165_);
  and _41422_ (_09168_, _08840_, _03295_);
  and _41423_ (_09169_, _09168_, _03060_);
  not _41424_ (_09171_, _09168_);
  and _41425_ (_09172_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or _41426_ (_09459_, _09172_, _09169_);
  and _41427_ (_09174_, _09168_, _03067_);
  and _41428_ (_09175_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or _41429_ (_09462_, _09175_, _09174_);
  and _41430_ (_09177_, _09168_, _03071_);
  and _41431_ (_09178_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or _41432_ (_09466_, _09178_, _09177_);
  and _41433_ (_09180_, _09168_, _03074_);
  and _41434_ (_09181_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or _41435_ (_09469_, _09181_, _09180_);
  and _41436_ (_09183_, _09168_, _03077_);
  and _41437_ (_09184_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or _41438_ (_09472_, _09184_, _09183_);
  and _41439_ (_09186_, _09168_, _03080_);
  and _41440_ (_09187_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _41441_ (_09476_, _09187_, _09186_);
  and _41442_ (_09189_, _09168_, _03083_);
  and _41443_ (_09190_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or _41444_ (_09479_, _09190_, _09189_);
  and _41445_ (_09192_, _09168_, _03087_);
  and _41446_ (_09193_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _41447_ (_09481_, _09193_, _09192_);
  and _41448_ (_09195_, _08840_, _03315_);
  and _41449_ (_09196_, _09195_, _03060_);
  not _41450_ (_09197_, _09195_);
  and _41451_ (_09199_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _41452_ (_09485_, _09199_, _09196_);
  and _41453_ (_09200_, _09195_, _03067_);
  and _41454_ (_09202_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _41455_ (_09488_, _09202_, _09200_);
  and _41456_ (_09203_, _09195_, _03071_);
  and _41457_ (_09205_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _41458_ (_09491_, _09205_, _09203_);
  and _41459_ (_09206_, _09195_, _03074_);
  and _41460_ (_09208_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _41461_ (_09495_, _09208_, _09206_);
  and _41462_ (_09210_, _09195_, _03077_);
  and _41463_ (_09211_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _41464_ (_09499_, _09211_, _09210_);
  and _41465_ (_09212_, _09195_, _03080_);
  and _41466_ (_09214_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _41467_ (_09502_, _09214_, _09212_);
  and _41468_ (_09215_, _09195_, _03083_);
  and _41469_ (_09217_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _41470_ (_09505_, _09217_, _09215_);
  and _41471_ (_09218_, _09195_, _03087_);
  and _41472_ (_09220_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _41473_ (_09507_, _09220_, _09218_);
  and _41474_ (_09221_, _08840_, _03334_);
  and _41475_ (_09223_, _09221_, _03060_);
  not _41476_ (_09224_, _09221_);
  and _41477_ (_09225_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _41478_ (_09511_, _09225_, _09223_);
  and _41479_ (_09227_, _09221_, _03067_);
  and _41480_ (_09228_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _41481_ (_09514_, _09228_, _09227_);
  and _41482_ (_09230_, _09221_, _03071_);
  and _41483_ (_09231_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _41484_ (_09517_, _09231_, _09230_);
  and _41485_ (_09233_, _09221_, _03074_);
  and _41486_ (_09235_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _41487_ (_09520_, _09235_, _09233_);
  and _41488_ (_09236_, _09221_, _03077_);
  and _41489_ (_09237_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _41490_ (_09523_, _09237_, _09236_);
  and _41491_ (_09239_, _09221_, _03080_);
  and _41492_ (_09240_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _41493_ (_09526_, _09240_, _09239_);
  and _41494_ (_09242_, _09221_, _03083_);
  and _41495_ (_09243_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _41496_ (_09529_, _09243_, _09242_);
  and _41497_ (_09245_, _09221_, _03087_);
  and _41498_ (_09246_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _41499_ (_09532_, _09246_, _09245_);
  and _41500_ (_09248_, _08840_, _03353_);
  and _41501_ (_09249_, _09248_, _03060_);
  not _41502_ (_09251_, _09248_);
  and _41503_ (_09252_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or _41504_ (_09535_, _09252_, _09249_);
  and _41505_ (_09254_, _09248_, _03067_);
  and _41506_ (_09255_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or _41507_ (_09538_, _09255_, _09254_);
  and _41508_ (_09257_, _09248_, _03071_);
  and _41509_ (_09258_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or _41510_ (_09541_, _09258_, _09257_);
  and _41511_ (_09260_, _09248_, _03074_);
  and _41512_ (_09261_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or _41513_ (_09544_, _09261_, _09260_);
  and _41514_ (_09263_, _09248_, _03077_);
  and _41515_ (_09264_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or _41516_ (_09548_, _09264_, _09263_);
  and _41517_ (_09266_, _09248_, _03080_);
  and _41518_ (_09267_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _41519_ (_09551_, _09267_, _09266_);
  and _41520_ (_09269_, _09248_, _03083_);
  and _41521_ (_09270_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or _41522_ (_09554_, _09270_, _09269_);
  and _41523_ (_09272_, _09248_, _03087_);
  and _41524_ (_09273_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or _41525_ (_09556_, _09273_, _09272_);
  and _41526_ (_09275_, _04125_, _26939_);
  and _41527_ (_09276_, _09275_, _02963_);
  not _41528_ (_09277_, _09276_);
  and _41529_ (_09279_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _41530_ (_09280_, _09276_, _03060_);
  or _41531_ (_09561_, _09280_, _09279_);
  and _41532_ (_09282_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _41533_ (_09283_, _09276_, _03067_);
  or _41534_ (_09564_, _09283_, _09282_);
  and _41535_ (_09285_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _41536_ (_09286_, _09276_, _03071_);
  or _41537_ (_09567_, _09286_, _09285_);
  and _41538_ (_09288_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _41539_ (_09289_, _09276_, _03074_);
  or _41540_ (_09570_, _09289_, _09288_);
  and _41541_ (_09291_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _41542_ (_09292_, _09276_, _03077_);
  or _41543_ (_09573_, _09292_, _09291_);
  and _41544_ (_09294_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _41545_ (_09295_, _09276_, _03080_);
  or _41546_ (_09576_, _09295_, _09294_);
  and _41547_ (_09297_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _41548_ (_09298_, _09276_, _03083_);
  or _41549_ (_09579_, _09298_, _09297_);
  and _41550_ (_09300_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _41551_ (_09301_, _09276_, _03087_);
  or _41552_ (_09582_, _09301_, _09300_);
  and _41553_ (_09303_, _09275_, _03062_);
  not _41554_ (_09304_, _09303_);
  and _41555_ (_09305_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and _41556_ (_09307_, _09303_, _03060_);
  or _41557_ (_09585_, _09307_, _09305_);
  and _41558_ (_09309_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and _41559_ (_09310_, _09303_, _03067_);
  or _41560_ (_09588_, _09310_, _09309_);
  and _41561_ (_09311_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and _41562_ (_09313_, _09303_, _03071_);
  or _41563_ (_09591_, _09313_, _09311_);
  and _41564_ (_09314_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and _41565_ (_09316_, _09303_, _03074_);
  or _41566_ (_09594_, _09316_, _09314_);
  and _41567_ (_09317_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  and _41568_ (_09319_, _09303_, _03077_);
  or _41569_ (_09597_, _09319_, _09317_);
  and _41570_ (_09320_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and _41571_ (_09322_, _09303_, _03080_);
  or _41572_ (_09601_, _09322_, _09320_);
  and _41573_ (_09323_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  and _41574_ (_09325_, _09303_, _03083_);
  or _41575_ (_09604_, _09325_, _09323_);
  and _41576_ (_09326_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  and _41577_ (_09328_, _09303_, _03087_);
  or _41578_ (_09606_, _09328_, _09326_);
  and _41579_ (_09329_, _09275_, _03091_);
  not _41580_ (_09331_, _09329_);
  and _41581_ (_09332_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and _41582_ (_09334_, _09329_, _03060_);
  or _41583_ (_09610_, _09334_, _09332_);
  and _41584_ (_09335_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and _41585_ (_09336_, _09329_, _03067_);
  or _41586_ (_09613_, _09336_, _09335_);
  and _41587_ (_09338_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and _41588_ (_09339_, _09329_, _03071_);
  or _41589_ (_09616_, _09339_, _09338_);
  and _41590_ (_09341_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and _41591_ (_09342_, _09329_, _03074_);
  or _41592_ (_09619_, _09342_, _09341_);
  and _41593_ (_09344_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and _41594_ (_09345_, _09329_, _03077_);
  or _41595_ (_09622_, _09345_, _09344_);
  and _41596_ (_09347_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and _41597_ (_09348_, _09329_, _03080_);
  or _41598_ (_09625_, _09348_, _09347_);
  and _41599_ (_09350_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and _41600_ (_09351_, _09329_, _03083_);
  or _41601_ (_09629_, _09351_, _09350_);
  and _41602_ (_09353_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and _41603_ (_09354_, _09329_, _03087_);
  or _41604_ (_09631_, _09354_, _09353_);
  and _41605_ (_09356_, _09275_, _03113_);
  not _41606_ (_09358_, _09356_);
  and _41607_ (_09359_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _41608_ (_09360_, _09356_, _03060_);
  or _41609_ (_09635_, _09360_, _09359_);
  and _41610_ (_09362_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _41611_ (_09363_, _09356_, _03067_);
  or _41612_ (_09638_, _09363_, _09362_);
  and _41613_ (_09365_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _41614_ (_09366_, _09356_, _03071_);
  or _41615_ (_09641_, _09366_, _09365_);
  and _41616_ (_09368_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _41617_ (_09369_, _09356_, _03074_);
  or _41618_ (_09644_, _09369_, _09368_);
  and _41619_ (_09371_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _41620_ (_09372_, _09356_, _03077_);
  or _41621_ (_09647_, _09372_, _09371_);
  and _41622_ (_09374_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _41623_ (_09375_, _09356_, _03080_);
  or _41624_ (_09650_, _09375_, _09374_);
  and _41625_ (_09377_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _41626_ (_09378_, _09356_, _03083_);
  or _41627_ (_09653_, _09378_, _09377_);
  and _41628_ (_09380_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _41629_ (_09381_, _09356_, _03087_);
  or _41630_ (_09656_, _09381_, _09380_);
  and _41631_ (_09383_, _09275_, _03136_);
  not _41632_ (_09384_, _09383_);
  and _41633_ (_09385_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _41634_ (_09387_, _09383_, _03060_);
  or _41635_ (_09659_, _09387_, _09385_);
  and _41636_ (_09388_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _41637_ (_09390_, _09383_, _03067_);
  or _41638_ (_09662_, _09390_, _09388_);
  and _41639_ (_09391_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _41640_ (_09393_, _09383_, _03071_);
  or _41641_ (_09665_, _09393_, _09391_);
  and _41642_ (_09394_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _41643_ (_09396_, _09383_, _03074_);
  or _41644_ (_09668_, _09396_, _09394_);
  and _41645_ (_09397_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _41646_ (_09399_, _09383_, _03077_);
  or _41647_ (_09671_, _09399_, _09397_);
  and _41648_ (_09400_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _41649_ (_09402_, _09383_, _03080_);
  or _41650_ (_09674_, _09402_, _09400_);
  and _41651_ (_09403_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _41652_ (_09405_, _09383_, _03083_);
  or _41653_ (_09677_, _09405_, _09403_);
  and _41654_ (_09407_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _41655_ (_09408_, _09383_, _03087_);
  or _41656_ (_09680_, _09408_, _09407_);
  and _41657_ (_09409_, _09275_, _03159_);
  not _41658_ (_09411_, _09409_);
  and _41659_ (_09412_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and _41660_ (_09413_, _09409_, _03060_);
  or _41661_ (_09684_, _09413_, _09412_);
  and _41662_ (_09415_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and _41663_ (_09416_, _09409_, _03067_);
  or _41664_ (_09687_, _09416_, _09415_);
  and _41665_ (_09418_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  and _41666_ (_09419_, _09409_, _03071_);
  or _41667_ (_09690_, _09419_, _09418_);
  and _41668_ (_09421_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and _41669_ (_09422_, _09409_, _03074_);
  or _41670_ (_09693_, _09422_, _09421_);
  and _41671_ (_09424_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and _41672_ (_09425_, _09409_, _03077_);
  or _41673_ (_09696_, _09425_, _09424_);
  and _41674_ (_09427_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and _41675_ (_09428_, _09409_, _03080_);
  or _41676_ (_09699_, _09428_, _09427_);
  and _41677_ (_09430_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and _41678_ (_09432_, _09409_, _03083_);
  or _41679_ (_09702_, _09432_, _09430_);
  and _41680_ (_09433_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and _41681_ (_09434_, _09409_, _03087_);
  or _41682_ (_09704_, _09434_, _09433_);
  and _41683_ (_09436_, _09275_, _03179_);
  not _41684_ (_09437_, _09436_);
  and _41685_ (_09439_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and _41686_ (_09440_, _09436_, _03060_);
  or _41687_ (_09709_, _09440_, _09439_);
  and _41688_ (_09442_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  and _41689_ (_09443_, _09436_, _03067_);
  or _41690_ (_09713_, _09443_, _09442_);
  and _41691_ (_09445_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and _41692_ (_09446_, _09436_, _03071_);
  or _41693_ (_09717_, _09446_, _09445_);
  and _41694_ (_09448_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  and _41695_ (_09449_, _09436_, _03074_);
  or _41696_ (_09721_, _09449_, _09448_);
  and _41697_ (_09451_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  and _41698_ (_09452_, _09436_, _03077_);
  or _41699_ (_09725_, _09452_, _09451_);
  and _41700_ (_09454_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  and _41701_ (_09455_, _09436_, _03080_);
  or _41702_ (_09729_, _09455_, _09454_);
  and _41703_ (_09457_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  and _41704_ (_09458_, _09436_, _03083_);
  or _41705_ (_09733_, _09458_, _09457_);
  and _41706_ (_09460_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  and _41707_ (_09461_, _09436_, _03087_);
  or _41708_ (_09736_, _09461_, _09460_);
  and _41709_ (_09463_, _09275_, _03198_);
  not _41710_ (_09464_, _09463_);
  and _41711_ (_09465_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _41712_ (_09467_, _09463_, _03060_);
  or _41713_ (_09741_, _09467_, _09465_);
  and _41714_ (_09468_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _41715_ (_09470_, _09463_, _03067_);
  or _41716_ (_09745_, _09470_, _09468_);
  and _41717_ (_09471_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _41718_ (_09473_, _09463_, _03071_);
  or _41719_ (_09749_, _09473_, _09471_);
  and _41720_ (_09475_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _41721_ (_09477_, _09463_, _03074_);
  or _41722_ (_09753_, _09477_, _09475_);
  and _41723_ (_09478_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _41724_ (_09480_, _09463_, _03077_);
  or _41725_ (_09757_, _09480_, _09478_);
  and _41726_ (_09482_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _41727_ (_09483_, _09463_, _03080_);
  or _41728_ (_09761_, _09483_, _09482_);
  and _41729_ (_09484_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _41730_ (_09486_, _09463_, _03083_);
  or _41731_ (_09765_, _09486_, _09484_);
  and _41732_ (_09487_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _41733_ (_09489_, _09463_, _03087_);
  or _41734_ (_09768_, _09489_, _09487_);
  and _41735_ (_09490_, _09275_, _03218_);
  not _41736_ (_09492_, _09490_);
  and _41737_ (_09493_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and _41738_ (_09494_, _09490_, _03060_);
  or _41739_ (_09773_, _09494_, _09493_);
  and _41740_ (_09497_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and _41741_ (_09498_, _09490_, _03067_);
  or _41742_ (_09777_, _09498_, _09497_);
  and _41743_ (_09500_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and _41744_ (_09501_, _09490_, _03071_);
  or _41745_ (_09781_, _09501_, _09500_);
  and _41746_ (_09503_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and _41747_ (_09504_, _09490_, _03074_);
  or _41748_ (_09785_, _09504_, _09503_);
  and _41749_ (_09506_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and _41750_ (_09508_, _09490_, _03077_);
  or _41751_ (_09789_, _09508_, _09506_);
  and _41752_ (_09509_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  and _41753_ (_09510_, _09490_, _03080_);
  or _41754_ (_09793_, _09510_, _09509_);
  and _41755_ (_09512_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and _41756_ (_09513_, _09490_, _03083_);
  or _41757_ (_09797_, _09513_, _09512_);
  and _41758_ (_09515_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and _41759_ (_09516_, _09490_, _03087_);
  or _41760_ (_09800_, _09516_, _09515_);
  and _41761_ (_09518_, _09275_, _03237_);
  not _41762_ (_09519_, _09518_);
  and _41763_ (_09521_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _41764_ (_09522_, _09518_, _03060_);
  or _41765_ (_09805_, _09522_, _09521_);
  and _41766_ (_09524_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _41767_ (_09525_, _09518_, _03067_);
  or _41768_ (_09809_, _09525_, _09524_);
  and _41769_ (_09527_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _41770_ (_09528_, _09518_, _03071_);
  or _41771_ (_09813_, _09528_, _09527_);
  and _41772_ (_09530_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _41773_ (_09531_, _09518_, _03074_);
  or _41774_ (_09817_, _09531_, _09530_);
  and _41775_ (_09533_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _41776_ (_09534_, _09518_, _03077_);
  or _41777_ (_09821_, _09534_, _09533_);
  and _41778_ (_09536_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _41779_ (_09537_, _09518_, _03080_);
  or _41780_ (_09825_, _09537_, _09536_);
  and _41781_ (_09539_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _41782_ (_09540_, _09518_, _03083_);
  or _41783_ (_09829_, _09540_, _09539_);
  and _41784_ (_09542_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _41785_ (_09543_, _09518_, _03087_);
  or _41786_ (_09832_, _09543_, _09542_);
  and _41787_ (_09545_, _09275_, _03256_);
  not _41788_ (_09546_, _09545_);
  and _41789_ (_09547_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _41790_ (_09549_, _09545_, _03060_);
  or _41791_ (_09837_, _09549_, _09547_);
  and _41792_ (_09550_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _41793_ (_09552_, _09545_, _03067_);
  or _41794_ (_09841_, _09552_, _09550_);
  and _41795_ (_09553_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _41796_ (_09555_, _09545_, _03071_);
  or _41797_ (_09845_, _09555_, _09553_);
  and _41798_ (_09557_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _41799_ (_09558_, _09545_, _03074_);
  or _41800_ (_09849_, _09558_, _09557_);
  and _41801_ (_09559_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _41802_ (_09560_, _09545_, _03077_);
  or _41803_ (_09853_, _09560_, _09559_);
  and _41804_ (_09562_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _41805_ (_09563_, _09545_, _03080_);
  or _41806_ (_09857_, _09563_, _09562_);
  and _41807_ (_09565_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _41808_ (_09566_, _09545_, _03083_);
  or _41809_ (_09861_, _09566_, _09565_);
  and _41810_ (_09568_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _41811_ (_09569_, _09545_, _03087_);
  or _41812_ (_09864_, _09569_, _09568_);
  and _41813_ (_09571_, _09275_, _03275_);
  not _41814_ (_09572_, _09571_);
  and _41815_ (_09574_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  and _41816_ (_09575_, _09571_, _03060_);
  or _41817_ (_09869_, _09575_, _09574_);
  and _41818_ (_09577_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and _41819_ (_09578_, _09571_, _03067_);
  or _41820_ (_09873_, _09578_, _09577_);
  and _41821_ (_09580_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and _41822_ (_09581_, _09571_, _03071_);
  or _41823_ (_09877_, _09581_, _09580_);
  and _41824_ (_09583_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and _41825_ (_09584_, _09571_, _03074_);
  or _41826_ (_09881_, _09584_, _09583_);
  and _41827_ (_09586_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and _41828_ (_09587_, _09571_, _03077_);
  or _41829_ (_09885_, _09587_, _09586_);
  and _41830_ (_09589_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and _41831_ (_09590_, _09571_, _03080_);
  or _41832_ (_09889_, _09590_, _09589_);
  and _41833_ (_09592_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  and _41834_ (_09593_, _09571_, _03083_);
  or _41835_ (_09893_, _09593_, _09592_);
  and _41836_ (_09595_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and _41837_ (_09596_, _09571_, _03087_);
  or _41838_ (_09896_, _09596_, _09595_);
  and _41839_ (_09598_, _09275_, _03295_);
  not _41840_ (_09599_, _09598_);
  and _41841_ (_09600_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and _41842_ (_09602_, _09598_, _03060_);
  or _41843_ (_09901_, _09602_, _09600_);
  and _41844_ (_09603_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and _41845_ (_09605_, _09598_, _03067_);
  or _41846_ (_09905_, _09605_, _09603_);
  and _41847_ (_09607_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and _41848_ (_09608_, _09598_, _03071_);
  or _41849_ (_09909_, _09608_, _09607_);
  and _41850_ (_09609_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  and _41851_ (_09611_, _09598_, _03074_);
  or _41852_ (_09913_, _09611_, _09609_);
  and _41853_ (_09612_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  and _41854_ (_09614_, _09598_, _03077_);
  or _41855_ (_09917_, _09614_, _09612_);
  and _41856_ (_09615_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and _41857_ (_09617_, _09598_, _03080_);
  or _41858_ (_09921_, _09617_, _09615_);
  and _41859_ (_09618_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and _41860_ (_09620_, _09598_, _03083_);
  or _41861_ (_09925_, _09620_, _09618_);
  and _41862_ (_09621_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and _41863_ (_09623_, _09598_, _03087_);
  or _41864_ (_09928_, _09623_, _09621_);
  and _41865_ (_09624_, _09275_, _03315_);
  not _41866_ (_09626_, _09624_);
  and _41867_ (_09627_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _41868_ (_09628_, _09624_, _03060_);
  or _41869_ (_09933_, _09628_, _09627_);
  and _41870_ (_09630_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _41871_ (_09632_, _09624_, _03067_);
  or _41872_ (_09937_, _09632_, _09630_);
  and _41873_ (_09633_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _41874_ (_09634_, _09624_, _03071_);
  or _41875_ (_09941_, _09634_, _09633_);
  and _41876_ (_09636_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _41877_ (_09637_, _09624_, _03074_);
  or _41878_ (_09945_, _09637_, _09636_);
  and _41879_ (_09639_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _41880_ (_09640_, _09624_, _03077_);
  or _41881_ (_09949_, _09640_, _09639_);
  and _41882_ (_09642_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _41883_ (_09643_, _09624_, _03080_);
  or _41884_ (_09953_, _09643_, _09642_);
  and _41885_ (_09645_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _41886_ (_09646_, _09624_, _03083_);
  or _41887_ (_09957_, _09646_, _09645_);
  and _41888_ (_09648_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _41889_ (_09649_, _09624_, _03087_);
  or _41890_ (_09960_, _09649_, _09648_);
  and _41891_ (_09651_, _09275_, _03334_);
  not _41892_ (_09652_, _09651_);
  and _41893_ (_09654_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _41894_ (_09655_, _09651_, _03060_);
  or _41895_ (_09965_, _09655_, _09654_);
  and _41896_ (_09657_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _41897_ (_09658_, _09651_, _03067_);
  or _41898_ (_09969_, _09658_, _09657_);
  and _41899_ (_09660_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _41900_ (_09661_, _09651_, _03071_);
  or _41901_ (_09973_, _09661_, _09660_);
  and _41902_ (_09663_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _41903_ (_09664_, _09651_, _03074_);
  or _41904_ (_09977_, _09664_, _09663_);
  and _41905_ (_09666_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _41906_ (_09667_, _09651_, _03077_);
  or _41907_ (_09981_, _09667_, _09666_);
  and _41908_ (_09669_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _41909_ (_09670_, _09651_, _03080_);
  or _41910_ (_09985_, _09670_, _09669_);
  and _41911_ (_09672_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _41912_ (_09673_, _09651_, _03083_);
  or _41913_ (_09989_, _09673_, _09672_);
  and _41914_ (_09675_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _41915_ (_09676_, _09651_, _03087_);
  or _41916_ (_09992_, _09676_, _09675_);
  and _41917_ (_09678_, _09275_, _03353_);
  not _41918_ (_09679_, _09678_);
  and _41919_ (_09681_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  and _41920_ (_09682_, _09678_, _03060_);
  or _41921_ (_09997_, _09682_, _09681_);
  and _41922_ (_09683_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  and _41923_ (_09685_, _09678_, _03067_);
  or _41924_ (_10001_, _09685_, _09683_);
  and _41925_ (_09686_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  and _41926_ (_09688_, _09678_, _03071_);
  or _41927_ (_10005_, _09688_, _09686_);
  and _41928_ (_09689_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  and _41929_ (_09691_, _09678_, _03074_);
  or _41930_ (_10009_, _09691_, _09689_);
  and _41931_ (_09692_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  and _41932_ (_09694_, _09678_, _03077_);
  or _41933_ (_10013_, _09694_, _09692_);
  and _41934_ (_09695_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  and _41935_ (_09697_, _09678_, _03080_);
  or _41936_ (_10017_, _09697_, _09695_);
  and _41937_ (_09698_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  and _41938_ (_09700_, _09678_, _03083_);
  or _41939_ (_10021_, _09700_, _09698_);
  and _41940_ (_09701_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  and _41941_ (_09703_, _09678_, _03087_);
  or _41942_ (_10024_, _09703_, _09701_);
  and _41943_ (_09705_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _41944_ (_09706_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _41945_ (_09707_, _09706_, _09705_);
  and _41946_ (_09708_, _09707_, _01954_);
  and _41947_ (_09710_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and _41948_ (_09711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _41949_ (_09712_, _09711_, _09710_);
  and _41950_ (_09714_, _09712_, _02150_);
  or _41951_ (_09715_, _09714_, _09708_);
  or _41952_ (_09716_, _09715_, _02144_);
  and _41953_ (_09718_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _41954_ (_09719_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _41955_ (_09720_, _09719_, _09718_);
  and _41956_ (_09722_, _09720_, _01954_);
  and _41957_ (_09723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _41958_ (_09724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _41959_ (_09726_, _09724_, _09723_);
  and _41960_ (_09727_, _09726_, _02150_);
  or _41961_ (_09728_, _09727_, _09722_);
  or _41962_ (_09730_, _09728_, _02131_);
  and _41963_ (_09731_, _09730_, _02157_);
  and _41964_ (_09732_, _09731_, _09716_);
  or _41965_ (_09734_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _41966_ (_09735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and _41967_ (_09737_, _09735_, _09734_);
  and _41968_ (_09738_, _09737_, _01954_);
  or _41969_ (_09739_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _41970_ (_09740_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _41971_ (_09742_, _09740_, _09739_);
  and _41972_ (_09743_, _09742_, _02150_);
  or _41973_ (_09744_, _09743_, _09738_);
  or _41974_ (_09746_, _09744_, _02144_);
  or _41975_ (_09747_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _41976_ (_09748_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _41977_ (_09750_, _09748_, _09747_);
  and _41978_ (_09751_, _09750_, _01954_);
  or _41979_ (_09752_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _41980_ (_09754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and _41981_ (_09755_, _09754_, _09752_);
  and _41982_ (_09756_, _09755_, _02150_);
  or _41983_ (_09758_, _09756_, _09751_);
  or _41984_ (_09759_, _09758_, _02131_);
  and _41985_ (_09760_, _09759_, _02077_);
  and _41986_ (_09762_, _09760_, _09746_);
  or _41987_ (_09763_, _09762_, _09732_);
  and _41988_ (_09764_, _09763_, _02065_);
  and _41989_ (_09766_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _41990_ (_09767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _41991_ (_09769_, _09767_, _09766_);
  and _41992_ (_09770_, _09769_, _01954_);
  and _41993_ (_09771_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and _41994_ (_09772_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _41995_ (_09774_, _09772_, _09771_);
  and _41996_ (_09775_, _09774_, _02150_);
  or _41997_ (_09776_, _09775_, _09770_);
  or _41998_ (_09778_, _09776_, _02144_);
  and _41999_ (_09779_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _42000_ (_09780_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _42001_ (_09782_, _09780_, _09779_);
  and _42002_ (_09783_, _09782_, _01954_);
  and _42003_ (_09784_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and _42004_ (_09786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _42005_ (_09787_, _09786_, _09784_);
  and _42006_ (_09788_, _09787_, _02150_);
  or _42007_ (_09790_, _09788_, _09783_);
  or _42008_ (_09791_, _09790_, _02131_);
  and _42009_ (_09792_, _09791_, _02157_);
  and _42010_ (_09794_, _09792_, _09778_);
  or _42011_ (_09795_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _42012_ (_09796_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and _42013_ (_09798_, _09796_, _02150_);
  and _42014_ (_09799_, _09798_, _09795_);
  or _42015_ (_09801_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _42016_ (_09802_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _42017_ (_09803_, _09802_, _01954_);
  and _42018_ (_09804_, _09803_, _09801_);
  or _42019_ (_09806_, _09804_, _09799_);
  or _42020_ (_09807_, _09806_, _02144_);
  or _42021_ (_09808_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _42022_ (_09810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _42023_ (_09811_, _09810_, _02150_);
  and _42024_ (_09812_, _09811_, _09808_);
  or _42025_ (_09814_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _42026_ (_09815_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _42027_ (_09816_, _09815_, _01954_);
  and _42028_ (_09818_, _09816_, _09814_);
  or _42029_ (_09819_, _09818_, _09812_);
  or _42030_ (_09820_, _09819_, _02131_);
  and _42031_ (_09822_, _09820_, _02077_);
  and _42032_ (_09823_, _09822_, _09807_);
  or _42033_ (_09824_, _09823_, _09794_);
  and _42034_ (_09826_, _09824_, _02194_);
  or _42035_ (_09827_, _09826_, _09764_);
  and _42036_ (_09828_, _09827_, _02143_);
  and _42037_ (_09830_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _42038_ (_09831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _42039_ (_09833_, _09831_, _09830_);
  and _42040_ (_09834_, _09833_, _01954_);
  and _42041_ (_09835_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _42042_ (_09836_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _42043_ (_09838_, _09836_, _09835_);
  and _42044_ (_09839_, _09838_, _02150_);
  or _42045_ (_09840_, _09839_, _09834_);
  and _42046_ (_09842_, _09840_, _02131_);
  and _42047_ (_09843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _42048_ (_09844_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _42049_ (_09846_, _09844_, _09843_);
  and _42050_ (_09847_, _09846_, _01954_);
  and _42051_ (_09848_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _42052_ (_09850_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _42053_ (_09851_, _09850_, _09848_);
  and _42054_ (_09852_, _09851_, _02150_);
  or _42055_ (_09854_, _09852_, _09847_);
  and _42056_ (_09855_, _09854_, _02144_);
  or _42057_ (_09856_, _09855_, _09842_);
  and _42058_ (_09858_, _09856_, _02157_);
  or _42059_ (_09859_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _42060_ (_09860_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _42061_ (_09862_, _09860_, _02150_);
  and _42062_ (_09863_, _09862_, _09859_);
  or _42063_ (_09865_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _42064_ (_09866_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _42065_ (_09867_, _09866_, _01954_);
  and _42066_ (_09868_, _09867_, _09865_);
  or _42067_ (_09870_, _09868_, _09863_);
  and _42068_ (_09871_, _09870_, _02131_);
  or _42069_ (_09872_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _42070_ (_09874_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _42071_ (_09875_, _09874_, _02150_);
  and _42072_ (_09876_, _09875_, _09872_);
  or _42073_ (_09878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _42074_ (_09879_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _42075_ (_09880_, _09879_, _01954_);
  and _42076_ (_09882_, _09880_, _09878_);
  or _42077_ (_09883_, _09882_, _09876_);
  and _42078_ (_09884_, _09883_, _02144_);
  or _42079_ (_09886_, _09884_, _09871_);
  and _42080_ (_09887_, _09886_, _02077_);
  or _42081_ (_09888_, _09887_, _09858_);
  and _42082_ (_09890_, _09888_, _02194_);
  and _42083_ (_09891_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _42084_ (_09892_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _42085_ (_09894_, _09892_, _09891_);
  and _42086_ (_09895_, _09894_, _01954_);
  and _42087_ (_09897_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and _42088_ (_09898_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _42089_ (_09899_, _09898_, _09897_);
  and _42090_ (_09900_, _09899_, _02150_);
  or _42091_ (_09902_, _09900_, _09895_);
  and _42092_ (_09903_, _09902_, _02131_);
  and _42093_ (_09904_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _42094_ (_09906_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _42095_ (_09907_, _09906_, _09904_);
  and _42096_ (_09908_, _09907_, _01954_);
  and _42097_ (_09910_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _42098_ (_09911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _42099_ (_09912_, _09911_, _09910_);
  and _42100_ (_09914_, _09912_, _02150_);
  or _42101_ (_09915_, _09914_, _09908_);
  and _42102_ (_09916_, _09915_, _02144_);
  or _42103_ (_09918_, _09916_, _09903_);
  and _42104_ (_09919_, _09918_, _02157_);
  or _42105_ (_09920_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _42106_ (_09922_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _42107_ (_09923_, _09922_, _09920_);
  and _42108_ (_09924_, _09923_, _01954_);
  or _42109_ (_09926_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _42110_ (_09927_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _42111_ (_09929_, _09927_, _09926_);
  and _42112_ (_09930_, _09929_, _02150_);
  or _42113_ (_09931_, _09930_, _09924_);
  and _42114_ (_09932_, _09931_, _02131_);
  or _42115_ (_09934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _42116_ (_09935_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _42117_ (_09936_, _09935_, _09934_);
  and _42118_ (_09938_, _09936_, _01954_);
  or _42119_ (_09939_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _42120_ (_09940_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _42121_ (_09942_, _09940_, _09939_);
  and _42122_ (_09943_, _09942_, _02150_);
  or _42123_ (_09944_, _09943_, _09938_);
  and _42124_ (_09946_, _09944_, _02144_);
  or _42125_ (_09947_, _09946_, _09932_);
  and _42126_ (_09948_, _09947_, _02077_);
  or _42127_ (_09950_, _09948_, _09919_);
  and _42128_ (_09951_, _09950_, _02065_);
  or _42129_ (_09952_, _09951_, _09890_);
  and _42130_ (_09954_, _09952_, _02005_);
  or _42131_ (_09955_, _09954_, _09828_);
  or _42132_ (_09956_, _09955_, _02054_);
  and _42133_ (_09958_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _42134_ (_09959_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _42135_ (_09961_, _09959_, _09958_);
  and _42136_ (_09962_, _09961_, _01954_);
  and _42137_ (_09963_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _42138_ (_09964_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _42139_ (_09966_, _09964_, _09963_);
  and _42140_ (_09967_, _09966_, _02150_);
  or _42141_ (_09968_, _09967_, _09962_);
  or _42142_ (_09970_, _09968_, _02144_);
  and _42143_ (_09971_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _42144_ (_09972_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _42145_ (_09974_, _09972_, _09971_);
  and _42146_ (_09975_, _09974_, _01954_);
  and _42147_ (_09976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _42148_ (_09978_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _42149_ (_09979_, _09978_, _09976_);
  and _42150_ (_09980_, _09979_, _02150_);
  or _42151_ (_09982_, _09980_, _09975_);
  or _42152_ (_09983_, _09982_, _02131_);
  and _42153_ (_09984_, _09983_, _02157_);
  and _42154_ (_09986_, _09984_, _09970_);
  or _42155_ (_09987_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _42156_ (_09988_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and _42157_ (_09990_, _09988_, _02150_);
  and _42158_ (_09991_, _09990_, _09987_);
  or _42159_ (_09993_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _42160_ (_09994_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _42161_ (_09995_, _09994_, _01954_);
  and _42162_ (_09996_, _09995_, _09993_);
  or _42163_ (_09998_, _09996_, _09991_);
  or _42164_ (_09999_, _09998_, _02144_);
  or _42165_ (_10000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _42166_ (_10002_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _42167_ (_10003_, _10002_, _02150_);
  and _42168_ (_10004_, _10003_, _10000_);
  or _42169_ (_10006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _42170_ (_10007_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _42171_ (_10008_, _10007_, _01954_);
  and _42172_ (_10010_, _10008_, _10006_);
  or _42173_ (_10011_, _10010_, _10004_);
  or _42174_ (_10012_, _10011_, _02131_);
  and _42175_ (_10014_, _10012_, _02077_);
  and _42176_ (_10015_, _10014_, _09999_);
  or _42177_ (_10016_, _10015_, _09986_);
  and _42178_ (_10018_, _10016_, _02194_);
  and _42179_ (_10019_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _42180_ (_10020_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _42181_ (_10022_, _10020_, _10019_);
  and _42182_ (_10023_, _10022_, _01954_);
  and _42183_ (_10025_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _42184_ (_10026_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _42185_ (_10027_, _10026_, _10025_);
  and _42186_ (_10028_, _10027_, _02150_);
  or _42187_ (_10029_, _10028_, _10023_);
  or _42188_ (_10030_, _10029_, _02144_);
  and _42189_ (_10031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _42190_ (_10032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _42191_ (_10033_, _10032_, _10031_);
  and _42192_ (_10035_, _10033_, _01954_);
  and _42193_ (_10036_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _42194_ (_10037_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _42195_ (_10039_, _10037_, _10036_);
  and _42196_ (_10040_, _10039_, _02150_);
  or _42197_ (_10041_, _10040_, _10035_);
  or _42198_ (_10043_, _10041_, _02131_);
  and _42199_ (_10044_, _10043_, _02157_);
  and _42200_ (_10045_, _10044_, _10030_);
  or _42201_ (_10047_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _42202_ (_10048_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _42203_ (_10049_, _10048_, _10047_);
  and _42204_ (_10051_, _10049_, _01954_);
  or _42205_ (_10052_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _42206_ (_10053_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _42207_ (_10055_, _10053_, _10052_);
  and _42208_ (_10056_, _10055_, _02150_);
  or _42209_ (_10057_, _10056_, _10051_);
  or _42210_ (_10059_, _10057_, _02144_);
  or _42211_ (_10060_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _42212_ (_10061_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _42213_ (_10062_, _10061_, _10060_);
  and _42214_ (_10063_, _10062_, _01954_);
  or _42215_ (_10064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _42216_ (_10065_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _42217_ (_10066_, _10065_, _10064_);
  and _42218_ (_10067_, _10066_, _02150_);
  or _42219_ (_10068_, _10067_, _10063_);
  or _42220_ (_10069_, _10068_, _02131_);
  and _42221_ (_10070_, _10069_, _02077_);
  and _42222_ (_10071_, _10070_, _10059_);
  or _42223_ (_10072_, _10071_, _10045_);
  and _42224_ (_10073_, _10072_, _02065_);
  or _42225_ (_10074_, _10073_, _10018_);
  and _42226_ (_10075_, _10074_, _02143_);
  or _42227_ (_10076_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _42228_ (_10077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _42229_ (_10078_, _10077_, _10076_);
  and _42230_ (_10079_, _10078_, _01954_);
  or _42231_ (_10080_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _42232_ (_10081_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _42233_ (_10082_, _10081_, _10080_);
  and _42234_ (_10083_, _10082_, _02150_);
  or _42235_ (_10084_, _10083_, _10079_);
  and _42236_ (_10085_, _10084_, _02144_);
  or _42237_ (_10086_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _42238_ (_10087_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _42239_ (_10088_, _10087_, _10086_);
  and _42240_ (_10089_, _10088_, _01954_);
  or _42241_ (_10090_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _42242_ (_10091_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _42243_ (_10092_, _10091_, _10090_);
  and _42244_ (_10093_, _10092_, _02150_);
  or _42245_ (_10094_, _10093_, _10089_);
  and _42246_ (_10095_, _10094_, _02131_);
  or _42247_ (_10096_, _10095_, _10085_);
  and _42248_ (_10097_, _10096_, _02077_);
  and _42249_ (_10098_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _42250_ (_10099_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _42251_ (_10100_, _10099_, _10098_);
  and _42252_ (_10101_, _10100_, _01954_);
  and _42253_ (_10102_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _42254_ (_10103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _42255_ (_10104_, _10103_, _10102_);
  and _42256_ (_10105_, _10104_, _02150_);
  or _42257_ (_10106_, _10105_, _10101_);
  and _42258_ (_10107_, _10106_, _02144_);
  and _42259_ (_10108_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _42260_ (_10109_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _42261_ (_10110_, _10109_, _10108_);
  and _42262_ (_10111_, _10110_, _01954_);
  and _42263_ (_10112_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _42264_ (_10113_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _42265_ (_10114_, _10113_, _10112_);
  and _42266_ (_10115_, _10114_, _02150_);
  or _42267_ (_10116_, _10115_, _10111_);
  and _42268_ (_10117_, _10116_, _02131_);
  or _42269_ (_10118_, _10117_, _10107_);
  and _42270_ (_10119_, _10118_, _02157_);
  or _42271_ (_10120_, _10119_, _10097_);
  and _42272_ (_10121_, _10120_, _02065_);
  or _42273_ (_10122_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _42274_ (_10123_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _42275_ (_10124_, _10123_, _02150_);
  and _42276_ (_10125_, _10124_, _10122_);
  or _42277_ (_10126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _42278_ (_10127_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _42279_ (_10128_, _10127_, _01954_);
  and _42280_ (_10129_, _10128_, _10126_);
  or _42281_ (_10130_, _10129_, _10125_);
  and _42282_ (_10131_, _10130_, _02144_);
  or _42283_ (_10132_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _42284_ (_10133_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _42285_ (_10134_, _10133_, _02150_);
  and _42286_ (_10135_, _10134_, _10132_);
  or _42287_ (_10136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _42288_ (_10137_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _42289_ (_10138_, _10137_, _01954_);
  and _42290_ (_10139_, _10138_, _10136_);
  or _42291_ (_10140_, _10139_, _10135_);
  and _42292_ (_10141_, _10140_, _02131_);
  or _42293_ (_10142_, _10141_, _10131_);
  and _42294_ (_10143_, _10142_, _02077_);
  and _42295_ (_10144_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _42296_ (_10145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _42297_ (_10146_, _10145_, _10144_);
  and _42298_ (_10147_, _10146_, _01954_);
  and _42299_ (_10148_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _42300_ (_10149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _42301_ (_10150_, _10149_, _10148_);
  and _42302_ (_10151_, _10150_, _02150_);
  or _42303_ (_10152_, _10151_, _10147_);
  and _42304_ (_10153_, _10152_, _02144_);
  and _42305_ (_10154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _42306_ (_10155_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _42307_ (_10156_, _10155_, _10154_);
  and _42308_ (_10157_, _10156_, _01954_);
  and _42309_ (_10158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _42310_ (_10159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _42311_ (_10160_, _10159_, _10158_);
  and _42312_ (_10161_, _10160_, _02150_);
  or _42313_ (_10162_, _10161_, _10157_);
  and _42314_ (_10163_, _10162_, _02131_);
  or _42315_ (_10164_, _10163_, _10153_);
  and _42316_ (_10165_, _10164_, _02157_);
  or _42317_ (_10166_, _10165_, _10143_);
  and _42318_ (_10167_, _10166_, _02194_);
  or _42319_ (_10168_, _10167_, _10121_);
  and _42320_ (_10169_, _10168_, _02005_);
  or _42321_ (_10170_, _10169_, _10075_);
  or _42322_ (_10171_, _10170_, _02374_);
  and _42323_ (_10172_, _10171_, _09956_);
  or _42324_ (_10173_, _10172_, _02142_);
  and _42325_ (_10174_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _42326_ (_10175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _42327_ (_10176_, _10175_, _10174_);
  and _42328_ (_10177_, _10176_, _01954_);
  and _42329_ (_10178_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _42330_ (_10179_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _42331_ (_10180_, _10179_, _10178_);
  and _42332_ (_10181_, _10180_, _02150_);
  or _42333_ (_10182_, _10181_, _10177_);
  and _42334_ (_10183_, _10182_, _02131_);
  and _42335_ (_10184_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _42336_ (_10185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _42337_ (_10186_, _10185_, _10184_);
  and _42338_ (_10187_, _10186_, _01954_);
  and _42339_ (_10188_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _42340_ (_10189_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _42341_ (_10190_, _10189_, _10188_);
  and _42342_ (_10191_, _10190_, _02150_);
  or _42343_ (_10192_, _10191_, _10187_);
  and _42344_ (_10193_, _10192_, _02144_);
  or _42345_ (_10194_, _10193_, _10183_);
  and _42346_ (_10195_, _10194_, _02157_);
  or _42347_ (_10196_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _42348_ (_10197_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _42349_ (_10198_, _10197_, _02150_);
  and _42350_ (_10199_, _10198_, _10196_);
  or _42351_ (_10200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _42352_ (_10201_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _42353_ (_10202_, _10201_, _01954_);
  and _42354_ (_10203_, _10202_, _10200_);
  or _42355_ (_10204_, _10203_, _10199_);
  and _42356_ (_10205_, _10204_, _02131_);
  or _42357_ (_10206_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _42358_ (_10207_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _42359_ (_10208_, _10207_, _02150_);
  and _42360_ (_10209_, _10208_, _10206_);
  or _42361_ (_10210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _42362_ (_10211_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _42363_ (_10212_, _10211_, _01954_);
  and _42364_ (_10213_, _10212_, _10210_);
  or _42365_ (_10214_, _10213_, _10209_);
  and _42366_ (_10215_, _10214_, _02144_);
  or _42367_ (_10216_, _10215_, _10205_);
  and _42368_ (_10217_, _10216_, _02077_);
  or _42369_ (_10218_, _10217_, _10195_);
  and _42370_ (_10219_, _10218_, _02194_);
  and _42371_ (_10220_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _42372_ (_10221_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _42373_ (_10222_, _10221_, _10220_);
  and _42374_ (_10223_, _10222_, _01954_);
  and _42375_ (_10224_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _42376_ (_10225_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _42377_ (_10226_, _10225_, _10224_);
  and _42378_ (_10227_, _10226_, _02150_);
  or _42379_ (_10228_, _10227_, _10223_);
  and _42380_ (_10229_, _10228_, _02131_);
  and _42381_ (_10230_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _42382_ (_10231_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _42383_ (_10232_, _10231_, _10230_);
  and _42384_ (_10233_, _10232_, _01954_);
  and _42385_ (_10234_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _42386_ (_10235_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _42387_ (_10236_, _10235_, _10234_);
  and _42388_ (_10237_, _10236_, _02150_);
  or _42389_ (_10238_, _10237_, _10233_);
  and _42390_ (_10239_, _10238_, _02144_);
  or _42391_ (_10240_, _10239_, _10229_);
  and _42392_ (_10241_, _10240_, _02157_);
  or _42393_ (_10242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _42394_ (_10243_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _42395_ (_10244_, _10243_, _10242_);
  and _42396_ (_10245_, _10244_, _01954_);
  or _42397_ (_10246_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _42398_ (_10247_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _42399_ (_10248_, _10247_, _10246_);
  and _42400_ (_10249_, _10248_, _02150_);
  or _42401_ (_10250_, _10249_, _10245_);
  and _42402_ (_10251_, _10250_, _02131_);
  or _42403_ (_10252_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _42404_ (_10253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _42405_ (_10254_, _10253_, _10252_);
  and _42406_ (_10255_, _10254_, _01954_);
  or _42407_ (_10256_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _42408_ (_10257_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _42409_ (_10258_, _10257_, _10256_);
  and _42410_ (_10259_, _10258_, _02150_);
  or _42411_ (_10260_, _10259_, _10255_);
  and _42412_ (_10261_, _10260_, _02144_);
  or _42413_ (_10262_, _10261_, _10251_);
  and _42414_ (_10263_, _10262_, _02077_);
  or _42415_ (_10264_, _10263_, _10241_);
  and _42416_ (_10265_, _10264_, _02065_);
  or _42417_ (_10266_, _10265_, _10219_);
  and _42418_ (_10267_, _10266_, _02005_);
  and _42419_ (_10268_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and _42420_ (_10269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _42421_ (_10270_, _10269_, _10268_);
  and _42422_ (_10271_, _10270_, _01954_);
  and _42423_ (_10272_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _42424_ (_10273_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _42425_ (_10274_, _10273_, _10272_);
  and _42426_ (_10275_, _10274_, _02150_);
  or _42427_ (_10276_, _10275_, _10271_);
  or _42428_ (_10277_, _10276_, _02144_);
  and _42429_ (_10278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _42430_ (_10279_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _42431_ (_10280_, _10279_, _10278_);
  and _42432_ (_10281_, _10280_, _01954_);
  and _42433_ (_10282_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _42434_ (_10283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _42435_ (_10284_, _10283_, _10282_);
  and _42436_ (_10285_, _10284_, _02150_);
  or _42437_ (_10286_, _10285_, _10281_);
  or _42438_ (_10287_, _10286_, _02131_);
  and _42439_ (_10288_, _10287_, _02157_);
  and _42440_ (_10289_, _10288_, _10277_);
  or _42441_ (_10290_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _42442_ (_10291_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _42443_ (_10292_, _10291_, _10290_);
  and _42444_ (_10293_, _10292_, _01954_);
  or _42445_ (_10294_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _42446_ (_10295_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _42447_ (_10296_, _10295_, _10294_);
  and _42448_ (_10297_, _10296_, _02150_);
  or _42449_ (_10298_, _10297_, _10293_);
  or _42450_ (_10299_, _10298_, _02144_);
  or _42451_ (_10300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _42452_ (_10301_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and _42453_ (_10302_, _10301_, _10300_);
  and _42454_ (_10303_, _10302_, _01954_);
  or _42455_ (_10304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _42456_ (_10305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _42457_ (_10306_, _10305_, _10304_);
  and _42458_ (_10307_, _10306_, _02150_);
  or _42459_ (_10308_, _10307_, _10303_);
  or _42460_ (_10309_, _10308_, _02131_);
  and _42461_ (_10310_, _10309_, _02077_);
  and _42462_ (_10311_, _10310_, _10299_);
  or _42463_ (_10312_, _10311_, _10289_);
  and _42464_ (_10313_, _10312_, _02065_);
  and _42465_ (_10314_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _42466_ (_10315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _42467_ (_10316_, _10315_, _10314_);
  and _42468_ (_10317_, _10316_, _01954_);
  and _42469_ (_10318_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _42470_ (_10319_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _42471_ (_10320_, _10319_, _10318_);
  and _42472_ (_10321_, _10320_, _02150_);
  or _42473_ (_10322_, _10321_, _10317_);
  or _42474_ (_10323_, _10322_, _02144_);
  and _42475_ (_10324_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _42476_ (_10325_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _42477_ (_10326_, _10325_, _10324_);
  and _42478_ (_10327_, _10326_, _01954_);
  and _42479_ (_10328_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _42480_ (_10329_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _42481_ (_10330_, _10329_, _10328_);
  and _42482_ (_10331_, _10330_, _02150_);
  or _42483_ (_10332_, _10331_, _10327_);
  or _42484_ (_10333_, _10332_, _02131_);
  and _42485_ (_10334_, _10333_, _02157_);
  and _42486_ (_10335_, _10334_, _10323_);
  or _42487_ (_10336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _42488_ (_10337_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _42489_ (_10338_, _10337_, _02150_);
  and _42490_ (_10339_, _10338_, _10336_);
  or _42491_ (_10340_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _42492_ (_10341_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _42493_ (_10342_, _10341_, _01954_);
  and _42494_ (_10343_, _10342_, _10340_);
  or _42495_ (_10344_, _10343_, _10339_);
  or _42496_ (_10345_, _10344_, _02144_);
  or _42497_ (_10346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _42498_ (_10347_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _42499_ (_10348_, _10347_, _02150_);
  and _42500_ (_10349_, _10348_, _10346_);
  or _42501_ (_10350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _42502_ (_10351_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _42503_ (_10352_, _10351_, _01954_);
  and _42504_ (_10353_, _10352_, _10350_);
  or _42505_ (_10354_, _10353_, _10349_);
  or _42506_ (_10355_, _10354_, _02131_);
  and _42507_ (_10356_, _10355_, _02077_);
  and _42508_ (_10357_, _10356_, _10345_);
  or _42509_ (_10358_, _10357_, _10335_);
  and _42510_ (_10359_, _10358_, _02194_);
  or _42511_ (_10360_, _10359_, _10313_);
  and _42512_ (_10361_, _10360_, _02143_);
  or _42513_ (_10362_, _10361_, _10267_);
  or _42514_ (_10363_, _10362_, _02054_);
  and _42515_ (_10364_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _42516_ (_10365_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _42517_ (_10366_, _10365_, _10364_);
  and _42518_ (_10367_, _10366_, _02150_);
  and _42519_ (_10368_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _42520_ (_10369_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _42521_ (_10370_, _10369_, _10368_);
  and _42522_ (_10371_, _10370_, _01954_);
  or _42523_ (_10372_, _10371_, _10367_);
  or _42524_ (_10373_, _10372_, _02144_);
  and _42525_ (_10374_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _42526_ (_10375_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _42527_ (_10376_, _10375_, _10374_);
  and _42528_ (_10377_, _10376_, _02150_);
  and _42529_ (_10378_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and _42530_ (_10379_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _42531_ (_10380_, _10379_, _10378_);
  and _42532_ (_10381_, _10380_, _01954_);
  or _42533_ (_10382_, _10381_, _10377_);
  or _42534_ (_10383_, _10382_, _02131_);
  and _42535_ (_10384_, _10383_, _02157_);
  and _42536_ (_10385_, _10384_, _10373_);
  or _42537_ (_10386_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _42538_ (_10387_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _42539_ (_10388_, _10387_, _01954_);
  and _42540_ (_10389_, _10388_, _10386_);
  or _42541_ (_10390_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _42542_ (_10391_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _42543_ (_10392_, _10391_, _02150_);
  and _42544_ (_10393_, _10392_, _10390_);
  or _42545_ (_10394_, _10393_, _10389_);
  or _42546_ (_10395_, _10394_, _02144_);
  or _42547_ (_10396_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _42548_ (_10397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _42549_ (_10398_, _10397_, _01954_);
  and _42550_ (_10399_, _10398_, _10396_);
  or _42551_ (_10400_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _42552_ (_10401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and _42553_ (_10402_, _10401_, _02150_);
  and _42554_ (_10403_, _10402_, _10400_);
  or _42555_ (_10404_, _10403_, _10399_);
  or _42556_ (_10405_, _10404_, _02131_);
  and _42557_ (_10406_, _10405_, _02077_);
  and _42558_ (_10407_, _10406_, _10395_);
  or _42559_ (_10408_, _10407_, _10385_);
  and _42560_ (_10409_, _10408_, _02194_);
  and _42561_ (_10410_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _42562_ (_10411_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _42563_ (_10412_, _10411_, _01954_);
  or _42564_ (_10413_, _10412_, _10410_);
  and _42565_ (_10414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _42566_ (_10415_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _42567_ (_10416_, _10415_, _02150_);
  or _42568_ (_10417_, _10416_, _10414_);
  and _42569_ (_10418_, _10417_, _10413_);
  or _42570_ (_10419_, _10418_, _02144_);
  and _42571_ (_10420_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _42572_ (_10421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _42573_ (_10422_, _10421_, _01954_);
  or _42574_ (_10423_, _10422_, _10420_);
  and _42575_ (_10424_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _42576_ (_10425_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _42577_ (_10426_, _10425_, _02150_);
  or _42578_ (_10427_, _10426_, _10424_);
  and _42579_ (_10428_, _10427_, _10423_);
  or _42580_ (_10429_, _10428_, _02131_);
  and _42581_ (_10430_, _10429_, _02157_);
  and _42582_ (_10431_, _10430_, _10419_);
  or _42583_ (_10432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _42584_ (_10433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _42585_ (_10434_, _10433_, _10432_);
  or _42586_ (_10435_, _10434_, _02150_);
  or _42587_ (_10436_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _42588_ (_10437_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _42589_ (_10438_, _10437_, _10436_);
  or _42590_ (_10439_, _10438_, _01954_);
  and _42591_ (_10440_, _10439_, _10435_);
  or _42592_ (_10441_, _10440_, _02144_);
  or _42593_ (_10442_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _42594_ (_10443_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _42595_ (_10444_, _10443_, _10442_);
  or _42596_ (_10445_, _10444_, _02150_);
  or _42597_ (_10446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _42598_ (_10447_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _42599_ (_10448_, _10447_, _10446_);
  or _42600_ (_10449_, _10448_, _01954_);
  and _42601_ (_10450_, _10449_, _10445_);
  or _42602_ (_10451_, _10450_, _02131_);
  and _42603_ (_10452_, _10451_, _02077_);
  and _42604_ (_10453_, _10452_, _10441_);
  or _42605_ (_10454_, _10453_, _10431_);
  and _42606_ (_10455_, _10454_, _02065_);
  or _42607_ (_10456_, _10455_, _10409_);
  and _42608_ (_10457_, _10456_, _02143_);
  and _42609_ (_10458_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _42610_ (_10459_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _42611_ (_10460_, _10459_, _10458_);
  and _42612_ (_10461_, _10460_, _01954_);
  and _42613_ (_10462_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _42614_ (_10463_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _42615_ (_10464_, _10463_, _10462_);
  and _42616_ (_10465_, _10464_, _02150_);
  or _42617_ (_10466_, _10465_, _10461_);
  and _42618_ (_10467_, _10466_, _02131_);
  and _42619_ (_10468_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _42620_ (_10469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _42621_ (_10470_, _10469_, _10468_);
  and _42622_ (_10471_, _10470_, _01954_);
  and _42623_ (_10472_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _42624_ (_10473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _42625_ (_10474_, _10473_, _10472_);
  and _42626_ (_10475_, _10474_, _02150_);
  or _42627_ (_10476_, _10475_, _10471_);
  and _42628_ (_10477_, _10476_, _02144_);
  or _42629_ (_10478_, _10477_, _10467_);
  and _42630_ (_10479_, _10478_, _02157_);
  or _42631_ (_10480_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _42632_ (_10481_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _42633_ (_10482_, _10481_, _10480_);
  and _42634_ (_10483_, _10482_, _01954_);
  or _42635_ (_10484_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _42636_ (_10485_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _42637_ (_10486_, _10485_, _10484_);
  and _42638_ (_10487_, _10486_, _02150_);
  or _42639_ (_10488_, _10487_, _10483_);
  and _42640_ (_10489_, _10488_, _02131_);
  or _42641_ (_10490_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _42642_ (_10491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _42643_ (_10492_, _10491_, _10490_);
  and _42644_ (_10493_, _10492_, _01954_);
  or _42645_ (_10494_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _42646_ (_10495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _42647_ (_10496_, _10495_, _10494_);
  and _42648_ (_10497_, _10496_, _02150_);
  or _42649_ (_10498_, _10497_, _10493_);
  and _42650_ (_10499_, _10498_, _02144_);
  or _42651_ (_10500_, _10499_, _10489_);
  and _42652_ (_10501_, _10500_, _02077_);
  or _42653_ (_10502_, _10501_, _10479_);
  and _42654_ (_10503_, _10502_, _02065_);
  and _42655_ (_10504_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and _42656_ (_10505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or _42657_ (_10506_, _10505_, _10504_);
  and _42658_ (_10507_, _10506_, _01954_);
  and _42659_ (_10508_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and _42660_ (_10509_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _42661_ (_10510_, _10509_, _10508_);
  and _42662_ (_10511_, _10510_, _02150_);
  or _42663_ (_10512_, _10511_, _10507_);
  and _42664_ (_10513_, _10512_, _02131_);
  and _42665_ (_10514_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and _42666_ (_10515_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or _42667_ (_10516_, _10515_, _10514_);
  and _42668_ (_10517_, _10516_, _01954_);
  and _42669_ (_10518_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and _42670_ (_10519_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _42671_ (_10520_, _10519_, _10518_);
  and _42672_ (_10521_, _10520_, _02150_);
  or _42673_ (_10522_, _10521_, _10517_);
  and _42674_ (_10523_, _10522_, _02144_);
  or _42675_ (_10524_, _10523_, _10513_);
  and _42676_ (_10525_, _10524_, _02157_);
  or _42677_ (_10526_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _42678_ (_10527_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and _42679_ (_10528_, _10527_, _10526_);
  and _42680_ (_10529_, _10528_, _01954_);
  or _42681_ (_10530_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or _42682_ (_10531_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and _42683_ (_10532_, _10531_, _10530_);
  and _42684_ (_10533_, _10532_, _02150_);
  or _42685_ (_10534_, _10533_, _10529_);
  and _42686_ (_10535_, _10534_, _02131_);
  or _42687_ (_10536_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _42688_ (_10537_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and _42689_ (_10538_, _10537_, _10536_);
  and _42690_ (_10539_, _10538_, _01954_);
  or _42691_ (_10540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _42692_ (_10541_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and _42693_ (_10542_, _10541_, _10540_);
  and _42694_ (_10543_, _10542_, _02150_);
  or _42695_ (_10544_, _10543_, _10539_);
  and _42696_ (_10545_, _10544_, _02144_);
  or _42697_ (_10546_, _10545_, _10535_);
  and _42698_ (_10547_, _10546_, _02077_);
  or _42699_ (_10548_, _10547_, _10525_);
  and _42700_ (_10549_, _10548_, _02194_);
  or _42701_ (_10550_, _10549_, _10503_);
  and _42702_ (_10551_, _10550_, _02005_);
  or _42703_ (_10552_, _10551_, _10457_);
  or _42704_ (_10553_, _10552_, _02374_);
  and _42705_ (_10554_, _10553_, _10363_);
  or _42706_ (_10555_, _10554_, _01748_);
  and _42707_ (_10556_, _10555_, _10173_);
  or _42708_ (_10557_, _10556_, _02141_);
  or _42709_ (_10558_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _42710_ (_10559_, _10558_, _27355_);
  and _42711_ (_15236_, _10559_, _10557_);
  and _42712_ (_10560_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _42713_ (_10561_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _42714_ (_10562_, _10561_, _10560_);
  and _42715_ (_10563_, _10562_, _01954_);
  and _42716_ (_10564_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _42717_ (_10565_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _42718_ (_10566_, _10565_, _10564_);
  and _42719_ (_10567_, _10566_, _02150_);
  or _42720_ (_10568_, _10567_, _10563_);
  or _42721_ (_10569_, _10568_, _02144_);
  and _42722_ (_10570_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _42723_ (_10571_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _42724_ (_10572_, _10571_, _10570_);
  and _42725_ (_10573_, _10572_, _01954_);
  and _42726_ (_10574_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and _42727_ (_10575_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _42728_ (_10576_, _10575_, _10574_);
  and _42729_ (_10577_, _10576_, _02150_);
  or _42730_ (_10578_, _10577_, _10573_);
  or _42731_ (_10579_, _10578_, _02131_);
  and _42732_ (_10580_, _10579_, _02157_);
  and _42733_ (_10581_, _10580_, _10569_);
  or _42734_ (_10582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _42735_ (_10583_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _42736_ (_10584_, _10583_, _10582_);
  and _42737_ (_10585_, _10584_, _01954_);
  or _42738_ (_10586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _42739_ (_10587_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _42740_ (_10588_, _10587_, _10586_);
  and _42741_ (_10589_, _10588_, _02150_);
  or _42742_ (_10590_, _10589_, _10585_);
  or _42743_ (_10591_, _10590_, _02144_);
  or _42744_ (_10592_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _42745_ (_10593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and _42746_ (_10594_, _10593_, _10592_);
  and _42747_ (_10595_, _10594_, _01954_);
  or _42748_ (_10596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _42749_ (_10597_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _42750_ (_10598_, _10597_, _10596_);
  and _42751_ (_10599_, _10598_, _02150_);
  or _42752_ (_10600_, _10599_, _10595_);
  or _42753_ (_10601_, _10600_, _02131_);
  and _42754_ (_10602_, _10601_, _02077_);
  and _42755_ (_10603_, _10602_, _10591_);
  or _42756_ (_10604_, _10603_, _10581_);
  or _42757_ (_10605_, _10604_, _02194_);
  and _42758_ (_10606_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _42759_ (_10607_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _42760_ (_10608_, _10607_, _10606_);
  and _42761_ (_10609_, _10608_, _01954_);
  and _42762_ (_10610_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _42763_ (_10611_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _42764_ (_10612_, _10611_, _10610_);
  and _42765_ (_10613_, _10612_, _02150_);
  or _42766_ (_10614_, _10613_, _10609_);
  or _42767_ (_10615_, _10614_, _02144_);
  and _42768_ (_10616_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and _42769_ (_10617_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _42770_ (_10618_, _10617_, _10616_);
  and _42771_ (_10619_, _10618_, _01954_);
  and _42772_ (_10620_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _42773_ (_10621_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _42774_ (_10622_, _10621_, _10620_);
  and _42775_ (_10623_, _10622_, _02150_);
  or _42776_ (_10624_, _10623_, _10619_);
  or _42777_ (_10625_, _10624_, _02131_);
  and _42778_ (_10626_, _10625_, _02157_);
  and _42779_ (_10627_, _10626_, _10615_);
  or _42780_ (_10628_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _42781_ (_10629_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and _42782_ (_10630_, _10629_, _02150_);
  and _42783_ (_10631_, _10630_, _10628_);
  or _42784_ (_10632_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _42785_ (_10633_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _42786_ (_10634_, _10633_, _01954_);
  and _42787_ (_10635_, _10634_, _10632_);
  or _42788_ (_10636_, _10635_, _10631_);
  or _42789_ (_10637_, _10636_, _02144_);
  or _42790_ (_10638_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _42791_ (_10639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and _42792_ (_10640_, _10639_, _02150_);
  and _42793_ (_10641_, _10640_, _10638_);
  or _42794_ (_10642_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _42795_ (_10643_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _42796_ (_10644_, _10643_, _01954_);
  and _42797_ (_10645_, _10644_, _10642_);
  or _42798_ (_10646_, _10645_, _10641_);
  or _42799_ (_10647_, _10646_, _02131_);
  and _42800_ (_10648_, _10647_, _02077_);
  and _42801_ (_10649_, _10648_, _10637_);
  or _42802_ (_10650_, _10649_, _10627_);
  or _42803_ (_10651_, _10650_, _02065_);
  and _42804_ (_10652_, _10651_, _02143_);
  and _42805_ (_10653_, _10652_, _10605_);
  and _42806_ (_10654_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _42807_ (_10655_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or _42808_ (_10656_, _10655_, _10654_);
  and _42809_ (_10657_, _10656_, _01954_);
  and _42810_ (_10658_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _42811_ (_10659_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _42812_ (_10660_, _10659_, _10658_);
  and _42813_ (_10661_, _10660_, _02150_);
  or _42814_ (_10662_, _10661_, _10657_);
  and _42815_ (_10663_, _10662_, _02131_);
  and _42816_ (_10664_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _42817_ (_10665_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _42818_ (_10666_, _10665_, _10664_);
  and _42819_ (_10667_, _10666_, _01954_);
  and _42820_ (_10668_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _42821_ (_10669_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _42822_ (_10670_, _10669_, _10668_);
  and _42823_ (_10671_, _10670_, _02150_);
  or _42824_ (_10672_, _10671_, _10667_);
  and _42825_ (_10673_, _10672_, _02144_);
  or _42826_ (_10674_, _10673_, _02077_);
  or _42827_ (_10675_, _10674_, _10663_);
  or _42828_ (_10676_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _42829_ (_10677_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _42830_ (_10678_, _10677_, _02150_);
  and _42831_ (_10679_, _10678_, _10676_);
  or _42832_ (_10680_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _42833_ (_10681_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _42834_ (_10682_, _10681_, _01954_);
  and _42835_ (_10683_, _10682_, _10680_);
  or _42836_ (_10684_, _10683_, _10679_);
  and _42837_ (_10685_, _10684_, _02131_);
  or _42838_ (_10686_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _42839_ (_10687_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _42840_ (_10688_, _10687_, _02150_);
  and _42841_ (_10689_, _10688_, _10686_);
  or _42842_ (_10690_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _42843_ (_10691_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and _42844_ (_10692_, _10691_, _01954_);
  and _42845_ (_10693_, _10692_, _10690_);
  or _42846_ (_10694_, _10693_, _10689_);
  and _42847_ (_10695_, _10694_, _02144_);
  or _42848_ (_10696_, _10695_, _02157_);
  or _42849_ (_10697_, _10696_, _10685_);
  and _42850_ (_10698_, _10697_, _10675_);
  or _42851_ (_10699_, _10698_, _02065_);
  and _42852_ (_10700_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and _42853_ (_10701_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _42854_ (_10702_, _10701_, _10700_);
  and _42855_ (_10703_, _10702_, _01954_);
  and _42856_ (_10704_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _42857_ (_10705_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _42858_ (_10706_, _10705_, _10704_);
  and _42859_ (_10707_, _10706_, _02150_);
  or _42860_ (_10708_, _10707_, _10703_);
  and _42861_ (_10709_, _10708_, _02131_);
  and _42862_ (_10710_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _42863_ (_10711_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _42864_ (_10712_, _10711_, _10710_);
  and _42865_ (_10713_, _10712_, _01954_);
  and _42866_ (_10714_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _42867_ (_10715_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _42868_ (_10716_, _10715_, _10714_);
  and _42869_ (_10717_, _10716_, _02150_);
  or _42870_ (_10719_, _10717_, _10713_);
  and _42871_ (_10720_, _10719_, _02144_);
  or _42872_ (_10721_, _10720_, _02077_);
  or _42873_ (_10722_, _10721_, _10709_);
  or _42874_ (_10723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _42875_ (_10724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and _42876_ (_10725_, _10724_, _10723_);
  and _42877_ (_10726_, _10725_, _01954_);
  or _42878_ (_10727_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _42879_ (_10728_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _42880_ (_10730_, _10728_, _10727_);
  and _42881_ (_10731_, _10730_, _02150_);
  or _42882_ (_10732_, _10731_, _10726_);
  and _42883_ (_10733_, _10732_, _02131_);
  or _42884_ (_10734_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _42885_ (_10735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _42886_ (_10736_, _10735_, _10734_);
  and _42887_ (_10737_, _10736_, _01954_);
  or _42888_ (_10738_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _42889_ (_10739_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _42890_ (_10741_, _10739_, _10738_);
  and _42891_ (_10742_, _10741_, _02150_);
  or _42892_ (_10743_, _10742_, _10737_);
  and _42893_ (_10744_, _10743_, _02144_);
  or _42894_ (_10745_, _10744_, _02157_);
  or _42895_ (_10746_, _10745_, _10733_);
  and _42896_ (_10747_, _10746_, _10722_);
  or _42897_ (_10748_, _10747_, _02194_);
  and _42898_ (_10749_, _10748_, _02005_);
  and _42899_ (_10750_, _10749_, _10699_);
  or _42900_ (_10752_, _10750_, _10653_);
  or _42901_ (_10753_, _10752_, _02054_);
  and _42902_ (_10754_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and _42903_ (_10755_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or _42904_ (_10756_, _10755_, _10754_);
  and _42905_ (_10757_, _10756_, _01954_);
  and _42906_ (_10758_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and _42907_ (_10759_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _42908_ (_10760_, _10759_, _10758_);
  and _42909_ (_10761_, _10760_, _02150_);
  or _42910_ (_10763_, _10761_, _10757_);
  and _42911_ (_10764_, _10763_, _02131_);
  and _42912_ (_10765_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and _42913_ (_10766_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _42914_ (_10767_, _10766_, _10765_);
  and _42915_ (_10768_, _10767_, _01954_);
  and _42916_ (_10769_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and _42917_ (_10770_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or _42918_ (_10771_, _10770_, _10769_);
  and _42919_ (_10772_, _10771_, _02150_);
  or _42920_ (_10774_, _10772_, _10768_);
  and _42921_ (_10775_, _10774_, _02144_);
  or _42922_ (_10776_, _10775_, _02077_);
  or _42923_ (_10777_, _10776_, _10764_);
  or _42924_ (_10778_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _42925_ (_10779_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and _42926_ (_10780_, _10779_, _10778_);
  and _42927_ (_10781_, _10780_, _01954_);
  or _42928_ (_10782_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _42929_ (_10783_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and _42930_ (_10785_, _10783_, _10782_);
  and _42931_ (_10786_, _10785_, _02150_);
  or _42932_ (_10787_, _10786_, _10781_);
  and _42933_ (_10788_, _10787_, _02131_);
  or _42934_ (_10789_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or _42935_ (_10790_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and _42936_ (_10791_, _10790_, _10789_);
  and _42937_ (_10792_, _10791_, _01954_);
  or _42938_ (_10793_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or _42939_ (_10794_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and _42940_ (_10795_, _10794_, _10793_);
  and _42941_ (_10796_, _10795_, _02150_);
  or _42942_ (_10797_, _10796_, _10792_);
  and _42943_ (_10798_, _10797_, _02144_);
  or _42944_ (_10799_, _10798_, _02157_);
  or _42945_ (_10800_, _10799_, _10788_);
  and _42946_ (_10801_, _10800_, _10777_);
  or _42947_ (_10802_, _10801_, _02065_);
  and _42948_ (_10803_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _42949_ (_10804_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _42950_ (_10805_, _10804_, _10803_);
  and _42951_ (_10806_, _10805_, _01954_);
  and _42952_ (_10807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and _42953_ (_10808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _42954_ (_10809_, _10808_, _10807_);
  and _42955_ (_10810_, _10809_, _02150_);
  or _42956_ (_10811_, _10810_, _10806_);
  and _42957_ (_10812_, _10811_, _02131_);
  and _42958_ (_10813_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _42959_ (_10814_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _42960_ (_10815_, _10814_, _10813_);
  and _42961_ (_10816_, _10815_, _01954_);
  and _42962_ (_10817_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and _42963_ (_10818_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _42964_ (_10819_, _10818_, _10817_);
  and _42965_ (_10820_, _10819_, _02150_);
  or _42966_ (_10821_, _10820_, _10816_);
  and _42967_ (_10822_, _10821_, _02144_);
  or _42968_ (_10823_, _10822_, _02077_);
  or _42969_ (_10824_, _10823_, _10812_);
  or _42970_ (_10825_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _42971_ (_10826_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _42972_ (_10827_, _10826_, _10825_);
  and _42973_ (_10828_, _10827_, _01954_);
  or _42974_ (_10829_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _42975_ (_10830_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and _42976_ (_10831_, _10830_, _10829_);
  and _42977_ (_10832_, _10831_, _02150_);
  or _42978_ (_10833_, _10832_, _10828_);
  and _42979_ (_10834_, _10833_, _02131_);
  or _42980_ (_10835_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _42981_ (_10836_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _42982_ (_10837_, _10836_, _10835_);
  and _42983_ (_10838_, _10837_, _01954_);
  or _42984_ (_10839_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _42985_ (_10840_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and _42986_ (_10841_, _10840_, _10839_);
  and _42987_ (_10842_, _10841_, _02150_);
  or _42988_ (_10843_, _10842_, _10838_);
  and _42989_ (_10844_, _10843_, _02144_);
  or _42990_ (_10845_, _10844_, _02157_);
  or _42991_ (_10846_, _10845_, _10834_);
  and _42992_ (_10847_, _10846_, _10824_);
  or _42993_ (_10848_, _10847_, _02194_);
  and _42994_ (_10849_, _10848_, _02005_);
  and _42995_ (_10850_, _10849_, _10802_);
  and _42996_ (_10851_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _42997_ (_10852_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _42998_ (_10853_, _10852_, _10851_);
  and _42999_ (_10854_, _10853_, _02150_);
  and _43000_ (_10855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and _43001_ (_10856_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _43002_ (_10857_, _10856_, _10855_);
  and _43003_ (_10858_, _10857_, _01954_);
  or _43004_ (_10859_, _10858_, _10854_);
  or _43005_ (_10860_, _10859_, _02144_);
  and _43006_ (_10861_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _43007_ (_10862_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _43008_ (_10863_, _10862_, _10861_);
  and _43009_ (_10864_, _10863_, _02150_);
  and _43010_ (_10865_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and _43011_ (_10866_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _43012_ (_10867_, _10866_, _10865_);
  and _43013_ (_10868_, _10867_, _01954_);
  or _43014_ (_10869_, _10868_, _10864_);
  or _43015_ (_10870_, _10869_, _02131_);
  and _43016_ (_10871_, _10870_, _02157_);
  and _43017_ (_10872_, _10871_, _10860_);
  or _43018_ (_10873_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _43019_ (_10874_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _43020_ (_10875_, _10874_, _01954_);
  and _43021_ (_10876_, _10875_, _10873_);
  or _43022_ (_10877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _43023_ (_10878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _43024_ (_10879_, _10878_, _02150_);
  and _43025_ (_10880_, _10879_, _10877_);
  or _43026_ (_10881_, _10880_, _10876_);
  or _43027_ (_10882_, _10881_, _02144_);
  or _43028_ (_10883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _43029_ (_10884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and _43030_ (_10885_, _10884_, _01954_);
  and _43031_ (_10886_, _10885_, _10883_);
  or _43032_ (_10887_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _43033_ (_10888_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _43034_ (_10889_, _10888_, _02150_);
  and _43035_ (_10890_, _10889_, _10887_);
  or _43036_ (_10891_, _10890_, _10886_);
  or _43037_ (_10892_, _10891_, _02131_);
  and _43038_ (_10893_, _10892_, _02077_);
  and _43039_ (_10894_, _10893_, _10882_);
  or _43040_ (_10895_, _10894_, _10872_);
  and _43041_ (_10896_, _10895_, _02194_);
  and _43042_ (_10897_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _43043_ (_10898_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _43044_ (_10899_, _10898_, _01954_);
  or _43045_ (_10900_, _10899_, _10897_);
  and _43046_ (_10901_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _43047_ (_10902_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _43048_ (_10903_, _10902_, _02150_);
  or _43049_ (_10904_, _10903_, _10901_);
  and _43050_ (_10905_, _10904_, _10900_);
  or _43051_ (_10906_, _10905_, _02144_);
  and _43052_ (_10907_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _43053_ (_10908_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _43054_ (_10909_, _10908_, _01954_);
  or _43055_ (_10910_, _10909_, _10907_);
  and _43056_ (_10911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _43057_ (_10912_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _43058_ (_10913_, _10912_, _02150_);
  or _43059_ (_10914_, _10913_, _10911_);
  and _43060_ (_10915_, _10914_, _10910_);
  or _43061_ (_10916_, _10915_, _02131_);
  and _43062_ (_10917_, _10916_, _02157_);
  and _43063_ (_10918_, _10917_, _10906_);
  or _43064_ (_10919_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _43065_ (_10920_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _43066_ (_10921_, _10920_, _10919_);
  or _43067_ (_10922_, _10921_, _02150_);
  or _43068_ (_10923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _43069_ (_10924_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _43070_ (_10925_, _10924_, _10923_);
  or _43071_ (_10926_, _10925_, _01954_);
  and _43072_ (_10927_, _10926_, _10922_);
  or _43073_ (_10928_, _10927_, _02144_);
  or _43074_ (_10929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _43075_ (_10930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _43076_ (_10931_, _10930_, _10929_);
  or _43077_ (_10932_, _10931_, _02150_);
  or _43078_ (_10933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _43079_ (_10934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _43080_ (_10935_, _10934_, _10933_);
  or _43081_ (_10936_, _10935_, _01954_);
  and _43082_ (_10937_, _10936_, _10932_);
  or _43083_ (_10938_, _10937_, _02131_);
  and _43084_ (_10939_, _10938_, _02077_);
  and _43085_ (_10940_, _10939_, _10928_);
  or _43086_ (_10941_, _10940_, _10918_);
  and _43087_ (_10942_, _10941_, _02065_);
  or _43088_ (_10943_, _10942_, _10896_);
  and _43089_ (_10944_, _10943_, _02143_);
  or _43090_ (_10945_, _10944_, _10850_);
  or _43091_ (_10946_, _10945_, _02374_);
  and _43092_ (_10947_, _10946_, _10753_);
  or _43093_ (_10948_, _10947_, _02142_);
  and _43094_ (_10949_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _43095_ (_10950_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _43096_ (_10951_, _10950_, _10949_);
  and _43097_ (_10952_, _10951_, _01954_);
  and _43098_ (_10953_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and _43099_ (_10954_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _43100_ (_10955_, _10954_, _10953_);
  and _43101_ (_10956_, _10955_, _02150_);
  or _43102_ (_10957_, _10956_, _10952_);
  or _43103_ (_10958_, _10957_, _02144_);
  and _43104_ (_10959_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _43105_ (_10960_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _43106_ (_10961_, _10960_, _10959_);
  and _43107_ (_10962_, _10961_, _01954_);
  and _43108_ (_10963_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and _43109_ (_10964_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _43110_ (_10965_, _10964_, _10963_);
  and _43111_ (_10966_, _10965_, _02150_);
  or _43112_ (_10967_, _10966_, _10962_);
  or _43113_ (_10968_, _10967_, _02131_);
  and _43114_ (_10969_, _10968_, _02157_);
  and _43115_ (_10970_, _10969_, _10958_);
  or _43116_ (_10971_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _43117_ (_10972_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _43118_ (_10973_, _10972_, _10971_);
  and _43119_ (_10974_, _10973_, _01954_);
  or _43120_ (_10975_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _43121_ (_10976_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and _43122_ (_10977_, _10976_, _10975_);
  and _43123_ (_10978_, _10977_, _02150_);
  or _43124_ (_10979_, _10978_, _10974_);
  or _43125_ (_10980_, _10979_, _02144_);
  or _43126_ (_10981_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _43127_ (_10982_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _43128_ (_10983_, _10982_, _10981_);
  and _43129_ (_10984_, _10983_, _01954_);
  or _43130_ (_10985_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _43131_ (_10986_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and _43132_ (_10987_, _10986_, _10985_);
  and _43133_ (_10988_, _10987_, _02150_);
  or _43134_ (_10989_, _10988_, _10984_);
  or _43135_ (_10990_, _10989_, _02131_);
  and _43136_ (_10991_, _10990_, _02077_);
  and _43137_ (_10992_, _10991_, _10980_);
  or _43138_ (_10993_, _10992_, _10970_);
  and _43139_ (_10994_, _10993_, _02065_);
  and _43140_ (_10995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _43141_ (_10996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _43142_ (_10997_, _10996_, _10995_);
  and _43143_ (_10998_, _10997_, _01954_);
  and _43144_ (_10999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _43145_ (_11000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _43146_ (_11001_, _11000_, _10999_);
  and _43147_ (_11002_, _11001_, _02150_);
  or _43148_ (_11003_, _11002_, _10998_);
  or _43149_ (_11004_, _11003_, _02144_);
  and _43150_ (_11005_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _43151_ (_11006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _43152_ (_11007_, _11006_, _11005_);
  and _43153_ (_11008_, _11007_, _01954_);
  and _43154_ (_11009_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _43155_ (_11010_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _43156_ (_11011_, _11010_, _11009_);
  and _43157_ (_11012_, _11011_, _02150_);
  or _43158_ (_11013_, _11012_, _11008_);
  or _43159_ (_11014_, _11013_, _02131_);
  and _43160_ (_11015_, _11014_, _02157_);
  and _43161_ (_11016_, _11015_, _11004_);
  or _43162_ (_11017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _43163_ (_11018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _43164_ (_11019_, _11018_, _02150_);
  and _43165_ (_11020_, _11019_, _11017_);
  or _43166_ (_11021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _43167_ (_11022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _43168_ (_11023_, _11022_, _01954_);
  and _43169_ (_11024_, _11023_, _11021_);
  or _43170_ (_11025_, _11024_, _11020_);
  or _43171_ (_11026_, _11025_, _02144_);
  or _43172_ (_11027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _43173_ (_11028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _43174_ (_11029_, _11028_, _02150_);
  and _43175_ (_11030_, _11029_, _11027_);
  or _43176_ (_11031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _43177_ (_11032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _43178_ (_11033_, _11032_, _01954_);
  and _43179_ (_11034_, _11033_, _11031_);
  or _43180_ (_11035_, _11034_, _11030_);
  or _43181_ (_11036_, _11035_, _02131_);
  and _43182_ (_11037_, _11036_, _02077_);
  and _43183_ (_11038_, _11037_, _11026_);
  or _43184_ (_11039_, _11038_, _11016_);
  and _43185_ (_11040_, _11039_, _02194_);
  or _43186_ (_11041_, _11040_, _10994_);
  and _43187_ (_11042_, _11041_, _02143_);
  and _43188_ (_11043_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _43189_ (_11044_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _43190_ (_11045_, _11044_, _11043_);
  and _43191_ (_11046_, _11045_, _01954_);
  and _43192_ (_11047_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _43193_ (_11048_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _43194_ (_11049_, _11048_, _11047_);
  and _43195_ (_11050_, _11049_, _02150_);
  or _43196_ (_11051_, _11050_, _11046_);
  and _43197_ (_11052_, _11051_, _02131_);
  and _43198_ (_11053_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _43199_ (_11054_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _43200_ (_11055_, _11054_, _11053_);
  and _43201_ (_11056_, _11055_, _01954_);
  and _43202_ (_11057_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _43203_ (_11058_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _43204_ (_11059_, _11058_, _11057_);
  and _43205_ (_11060_, _11059_, _02150_);
  or _43206_ (_11061_, _11060_, _11056_);
  and _43207_ (_11062_, _11061_, _02144_);
  or _43208_ (_11063_, _11062_, _11052_);
  and _43209_ (_11064_, _11063_, _02157_);
  or _43210_ (_11065_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _43211_ (_11066_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _43212_ (_11067_, _11066_, _02150_);
  and _43213_ (_11068_, _11067_, _11065_);
  or _43214_ (_11069_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _43215_ (_11070_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _43216_ (_11071_, _11070_, _01954_);
  and _43217_ (_11072_, _11071_, _11069_);
  or _43218_ (_11073_, _11072_, _11068_);
  and _43219_ (_11074_, _11073_, _02131_);
  or _43220_ (_11075_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _43221_ (_11076_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _43222_ (_11077_, _11076_, _02150_);
  and _43223_ (_11078_, _11077_, _11075_);
  or _43224_ (_11079_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _43225_ (_11080_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _43226_ (_11081_, _11080_, _01954_);
  and _43227_ (_11082_, _11081_, _11079_);
  or _43228_ (_11083_, _11082_, _11078_);
  and _43229_ (_11084_, _11083_, _02144_);
  or _43230_ (_11085_, _11084_, _11074_);
  and _43231_ (_11086_, _11085_, _02077_);
  or _43232_ (_11087_, _11086_, _11064_);
  and _43233_ (_11088_, _11087_, _02194_);
  and _43234_ (_11089_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _43235_ (_11090_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _43236_ (_11091_, _11090_, _11089_);
  and _43237_ (_11092_, _11091_, _01954_);
  and _43238_ (_11093_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _43239_ (_11094_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _43240_ (_11095_, _11094_, _11093_);
  and _43241_ (_11096_, _11095_, _02150_);
  or _43242_ (_11097_, _11096_, _11092_);
  and _43243_ (_11098_, _11097_, _02131_);
  and _43244_ (_11099_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _43245_ (_11100_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _43246_ (_11101_, _11100_, _11099_);
  and _43247_ (_11102_, _11101_, _01954_);
  and _43248_ (_11103_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _43249_ (_11104_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _43250_ (_11105_, _11104_, _11103_);
  and _43251_ (_11106_, _11105_, _02150_);
  or _43252_ (_11107_, _11106_, _11102_);
  and _43253_ (_11108_, _11107_, _02144_);
  or _43254_ (_11109_, _11108_, _11098_);
  and _43255_ (_11110_, _11109_, _02157_);
  or _43256_ (_11111_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _43257_ (_11112_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _43258_ (_11113_, _11112_, _11111_);
  and _43259_ (_11114_, _11113_, _01954_);
  or _43260_ (_11115_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _43261_ (_11116_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _43262_ (_11117_, _11116_, _11115_);
  and _43263_ (_11118_, _11117_, _02150_);
  or _43264_ (_11119_, _11118_, _11114_);
  and _43265_ (_11120_, _11119_, _02131_);
  or _43266_ (_11121_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _43267_ (_11122_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _43268_ (_11123_, _11122_, _11121_);
  and _43269_ (_11124_, _11123_, _01954_);
  or _43270_ (_11125_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _43271_ (_11126_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _43272_ (_11127_, _11126_, _11125_);
  and _43273_ (_11128_, _11127_, _02150_);
  or _43274_ (_11129_, _11128_, _11124_);
  and _43275_ (_11130_, _11129_, _02144_);
  or _43276_ (_11131_, _11130_, _11120_);
  and _43277_ (_11132_, _11131_, _02077_);
  or _43278_ (_11133_, _11132_, _11110_);
  and _43279_ (_11134_, _11133_, _02065_);
  or _43280_ (_11135_, _11134_, _11088_);
  and _43281_ (_11136_, _11135_, _02005_);
  or _43282_ (_11137_, _11136_, _11042_);
  or _43283_ (_11138_, _11137_, _02054_);
  and _43284_ (_11139_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _43285_ (_11140_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _43286_ (_11141_, _11140_, _11139_);
  and _43287_ (_11142_, _11141_, _01954_);
  and _43288_ (_11143_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _43289_ (_11144_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _43290_ (_11145_, _11144_, _11143_);
  and _43291_ (_11146_, _11145_, _02150_);
  or _43292_ (_11147_, _11146_, _11142_);
  or _43293_ (_11148_, _11147_, _02144_);
  and _43294_ (_11149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _43295_ (_11150_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _43296_ (_11151_, _11150_, _11149_);
  and _43297_ (_11152_, _11151_, _01954_);
  and _43298_ (_11153_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and _43299_ (_11154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _43300_ (_11155_, _11154_, _11153_);
  and _43301_ (_11156_, _11155_, _02150_);
  or _43302_ (_11157_, _11156_, _11152_);
  or _43303_ (_11158_, _11157_, _02131_);
  and _43304_ (_11159_, _11158_, _02157_);
  and _43305_ (_11160_, _11159_, _11148_);
  or _43306_ (_11161_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _43307_ (_11162_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _43308_ (_11163_, _11162_, _02150_);
  and _43309_ (_11164_, _11163_, _11161_);
  or _43310_ (_11165_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _43311_ (_11166_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _43312_ (_11167_, _11166_, _01954_);
  and _43313_ (_11168_, _11167_, _11165_);
  or _43314_ (_11169_, _11168_, _11164_);
  or _43315_ (_11170_, _11169_, _02144_);
  or _43316_ (_11171_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _43317_ (_11172_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _43318_ (_11173_, _11172_, _02150_);
  and _43319_ (_11174_, _11173_, _11171_);
  or _43320_ (_11175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _43321_ (_11176_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _43322_ (_11177_, _11176_, _01954_);
  and _43323_ (_11178_, _11177_, _11175_);
  or _43324_ (_11179_, _11178_, _11174_);
  or _43325_ (_11180_, _11179_, _02131_);
  and _43326_ (_11181_, _11180_, _02077_);
  and _43327_ (_11182_, _11181_, _11170_);
  or _43328_ (_11183_, _11182_, _11160_);
  and _43329_ (_11184_, _11183_, _02194_);
  and _43330_ (_11185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _43331_ (_11186_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _43332_ (_11187_, _11186_, _11185_);
  and _43333_ (_11188_, _11187_, _01954_);
  and _43334_ (_11189_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _43335_ (_11190_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _43336_ (_11191_, _11190_, _11189_);
  and _43337_ (_11192_, _11191_, _02150_);
  or _43338_ (_11193_, _11192_, _11188_);
  or _43339_ (_11194_, _11193_, _02144_);
  and _43340_ (_11195_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _43341_ (_11196_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _43342_ (_11197_, _11196_, _11195_);
  and _43343_ (_11198_, _11197_, _01954_);
  and _43344_ (_11199_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _43345_ (_11200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _43346_ (_11201_, _11200_, _11199_);
  and _43347_ (_11202_, _11201_, _02150_);
  or _43348_ (_11203_, _11202_, _11198_);
  or _43349_ (_11204_, _11203_, _02131_);
  and _43350_ (_11205_, _11204_, _02157_);
  and _43351_ (_11206_, _11205_, _11194_);
  or _43352_ (_11207_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _43353_ (_11208_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _43354_ (_11209_, _11208_, _11207_);
  and _43355_ (_11210_, _11209_, _01954_);
  or _43356_ (_11211_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _43357_ (_11212_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _43358_ (_11213_, _11212_, _11211_);
  and _43359_ (_11214_, _11213_, _02150_);
  or _43360_ (_11215_, _11214_, _11210_);
  or _43361_ (_11216_, _11215_, _02144_);
  or _43362_ (_11217_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _43363_ (_11218_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _43364_ (_11219_, _11218_, _11217_);
  and _43365_ (_11220_, _11219_, _01954_);
  or _43366_ (_11221_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _43367_ (_11222_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _43368_ (_11223_, _11222_, _11221_);
  and _43369_ (_11224_, _11223_, _02150_);
  or _43370_ (_11225_, _11224_, _11220_);
  or _43371_ (_11226_, _11225_, _02131_);
  and _43372_ (_11227_, _11226_, _02077_);
  and _43373_ (_11228_, _11227_, _11216_);
  or _43374_ (_11229_, _11228_, _11206_);
  and _43375_ (_11230_, _11229_, _02065_);
  or _43376_ (_11231_, _11230_, _11184_);
  and _43377_ (_11232_, _11231_, _02143_);
  or _43378_ (_11233_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _43379_ (_11234_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _43380_ (_11235_, _11234_, _11233_);
  and _43381_ (_11236_, _11235_, _01954_);
  or _43382_ (_11237_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _43383_ (_11238_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _43384_ (_11239_, _11238_, _11237_);
  and _43385_ (_11240_, _11239_, _02150_);
  or _43386_ (_11241_, _11240_, _11236_);
  and _43387_ (_11242_, _11241_, _02144_);
  or _43388_ (_11243_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _43389_ (_11244_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _43390_ (_11245_, _11244_, _11243_);
  and _43391_ (_11246_, _11245_, _01954_);
  or _43392_ (_11247_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _43393_ (_11248_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _43394_ (_11249_, _11248_, _11247_);
  and _43395_ (_11250_, _11249_, _02150_);
  or _43396_ (_11251_, _11250_, _11246_);
  and _43397_ (_11252_, _11251_, _02131_);
  or _43398_ (_11253_, _11252_, _11242_);
  and _43399_ (_11254_, _11253_, _02077_);
  and _43400_ (_11255_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _43401_ (_11256_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _43402_ (_11257_, _11256_, _11255_);
  and _43403_ (_11258_, _11257_, _01954_);
  and _43404_ (_11259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _43405_ (_11260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _43406_ (_11261_, _11260_, _11259_);
  and _43407_ (_11262_, _11261_, _02150_);
  or _43408_ (_11263_, _11262_, _11258_);
  and _43409_ (_11264_, _11263_, _02144_);
  and _43410_ (_11265_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _43411_ (_11266_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _43412_ (_11267_, _11266_, _11265_);
  and _43413_ (_11268_, _11267_, _01954_);
  and _43414_ (_11269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _43415_ (_11270_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _43416_ (_11271_, _11270_, _11269_);
  and _43417_ (_11272_, _11271_, _02150_);
  or _43418_ (_11273_, _11272_, _11268_);
  and _43419_ (_11274_, _11273_, _02131_);
  or _43420_ (_11275_, _11274_, _11264_);
  and _43421_ (_11276_, _11275_, _02157_);
  or _43422_ (_11277_, _11276_, _11254_);
  and _43423_ (_11278_, _11277_, _02065_);
  or _43424_ (_11279_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _43425_ (_11280_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _43426_ (_11281_, _11280_, _02150_);
  and _43427_ (_11282_, _11281_, _11279_);
  or _43428_ (_11283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _43429_ (_11284_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _43430_ (_11285_, _11284_, _01954_);
  and _43431_ (_11286_, _11285_, _11283_);
  or _43432_ (_11287_, _11286_, _11282_);
  and _43433_ (_11288_, _11287_, _02144_);
  or _43434_ (_11289_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _43435_ (_11290_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _43436_ (_11291_, _11290_, _02150_);
  and _43437_ (_11292_, _11291_, _11289_);
  or _43438_ (_11293_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _43439_ (_11294_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _43440_ (_11295_, _11294_, _01954_);
  and _43441_ (_11296_, _11295_, _11293_);
  or _43442_ (_11297_, _11296_, _11292_);
  and _43443_ (_11298_, _11297_, _02131_);
  or _43444_ (_11299_, _11298_, _11288_);
  and _43445_ (_11300_, _11299_, _02077_);
  and _43446_ (_11301_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _43447_ (_11302_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _43448_ (_11303_, _11302_, _11301_);
  and _43449_ (_11304_, _11303_, _01954_);
  and _43450_ (_11305_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _43451_ (_11306_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _43452_ (_11307_, _11306_, _11305_);
  and _43453_ (_11308_, _11307_, _02150_);
  or _43454_ (_11309_, _11308_, _11304_);
  and _43455_ (_11310_, _11309_, _02144_);
  and _43456_ (_11311_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _43457_ (_11312_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _43458_ (_11313_, _11312_, _11311_);
  and _43459_ (_11314_, _11313_, _01954_);
  and _43460_ (_11315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _43461_ (_11316_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _43462_ (_11317_, _11316_, _11315_);
  and _43463_ (_11318_, _11317_, _02150_);
  or _43464_ (_11319_, _11318_, _11314_);
  and _43465_ (_11320_, _11319_, _02131_);
  or _43466_ (_11321_, _11320_, _11310_);
  and _43467_ (_11322_, _11321_, _02157_);
  or _43468_ (_11323_, _11322_, _11300_);
  and _43469_ (_11324_, _11323_, _02194_);
  or _43470_ (_11325_, _11324_, _11278_);
  and _43471_ (_11326_, _11325_, _02005_);
  or _43472_ (_11327_, _11326_, _11232_);
  or _43473_ (_11328_, _11327_, _02374_);
  and _43474_ (_11329_, _11328_, _11138_);
  or _43475_ (_11330_, _11329_, _01748_);
  and _43476_ (_11331_, _11330_, _10948_);
  or _43477_ (_11332_, _11331_, _02141_);
  or _43478_ (_11333_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _43479_ (_11334_, _11333_, _27355_);
  and _43480_ (_15238_, _11334_, _11332_);
  and _43481_ (_11335_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _43482_ (_11336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _43483_ (_11337_, _11336_, _11335_);
  and _43484_ (_11338_, _11337_, _01954_);
  and _43485_ (_11339_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _43486_ (_11340_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _43487_ (_11341_, _11340_, _11339_);
  and _43488_ (_11342_, _11341_, _02150_);
  or _43489_ (_11343_, _11342_, _11338_);
  or _43490_ (_11344_, _11343_, _02144_);
  and _43491_ (_11345_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _43492_ (_11346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _43493_ (_11347_, _11346_, _11345_);
  and _43494_ (_11348_, _11347_, _01954_);
  and _43495_ (_11349_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _43496_ (_11350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _43497_ (_11351_, _11350_, _11349_);
  and _43498_ (_11352_, _11351_, _02150_);
  or _43499_ (_11353_, _11352_, _11348_);
  or _43500_ (_11354_, _11353_, _02131_);
  and _43501_ (_11355_, _11354_, _02157_);
  and _43502_ (_11356_, _11355_, _11344_);
  or _43503_ (_11357_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _43504_ (_11358_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _43505_ (_11359_, _11358_, _11357_);
  and _43506_ (_11360_, _11359_, _01954_);
  or _43507_ (_11361_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _43508_ (_11362_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _43509_ (_11363_, _11362_, _11361_);
  and _43510_ (_11364_, _11363_, _02150_);
  or _43511_ (_11365_, _11364_, _11360_);
  or _43512_ (_11366_, _11365_, _02144_);
  or _43513_ (_11367_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _43514_ (_11368_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _43515_ (_11369_, _11368_, _11367_);
  and _43516_ (_11370_, _11369_, _01954_);
  or _43517_ (_11371_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _43518_ (_11372_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _43519_ (_11373_, _11372_, _11371_);
  and _43520_ (_11374_, _11373_, _02150_);
  or _43521_ (_11375_, _11374_, _11370_);
  or _43522_ (_11376_, _11375_, _02131_);
  and _43523_ (_11377_, _11376_, _02077_);
  and _43524_ (_11378_, _11377_, _11366_);
  or _43525_ (_11379_, _11378_, _11356_);
  and _43526_ (_11380_, _11379_, _02065_);
  and _43527_ (_11381_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _43528_ (_11382_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _43529_ (_11383_, _11382_, _11381_);
  and _43530_ (_11384_, _11383_, _01954_);
  and _43531_ (_11385_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _43532_ (_11386_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _43533_ (_11387_, _11386_, _11385_);
  and _43534_ (_11388_, _11387_, _02150_);
  or _43535_ (_11389_, _11388_, _11384_);
  or _43536_ (_11390_, _11389_, _02144_);
  and _43537_ (_11391_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _43538_ (_11392_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _43539_ (_11393_, _11392_, _11391_);
  and _43540_ (_11394_, _11393_, _01954_);
  and _43541_ (_11395_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _43542_ (_11396_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _43543_ (_11397_, _11396_, _11395_);
  and _43544_ (_11398_, _11397_, _02150_);
  or _43545_ (_11399_, _11398_, _11394_);
  or _43546_ (_11400_, _11399_, _02131_);
  and _43547_ (_11401_, _11400_, _02157_);
  and _43548_ (_11402_, _11401_, _11390_);
  or _43549_ (_11403_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _43550_ (_11404_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and _43551_ (_11405_, _11404_, _02150_);
  and _43552_ (_11406_, _11405_, _11403_);
  or _43553_ (_11407_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _43554_ (_11408_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and _43555_ (_11409_, _11408_, _01954_);
  and _43556_ (_11410_, _11409_, _11407_);
  or _43557_ (_11411_, _11410_, _11406_);
  or _43558_ (_11412_, _11411_, _02144_);
  or _43559_ (_11413_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _43560_ (_11414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _43561_ (_11415_, _11414_, _02150_);
  and _43562_ (_11416_, _11415_, _11413_);
  or _43563_ (_11417_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _43564_ (_11418_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _43565_ (_11419_, _11418_, _01954_);
  and _43566_ (_11420_, _11419_, _11417_);
  or _43567_ (_11421_, _11420_, _11416_);
  or _43568_ (_11422_, _11421_, _02131_);
  and _43569_ (_11423_, _11422_, _02077_);
  and _43570_ (_11424_, _11423_, _11412_);
  or _43571_ (_11425_, _11424_, _11402_);
  and _43572_ (_11426_, _11425_, _02194_);
  or _43573_ (_11427_, _11426_, _11380_);
  and _43574_ (_11428_, _11427_, _02143_);
  and _43575_ (_11429_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _43576_ (_11430_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _43577_ (_11431_, _11430_, _11429_);
  and _43578_ (_11432_, _11431_, _01954_);
  and _43579_ (_11433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _43580_ (_11434_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _43581_ (_11435_, _11434_, _11433_);
  and _43582_ (_11436_, _11435_, _02150_);
  or _43583_ (_11437_, _11436_, _11432_);
  and _43584_ (_11438_, _11437_, _02131_);
  and _43585_ (_11439_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _43586_ (_11440_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _43587_ (_11441_, _11440_, _11439_);
  and _43588_ (_11442_, _11441_, _01954_);
  and _43589_ (_11443_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _43590_ (_11444_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _43591_ (_11445_, _11444_, _11443_);
  and _43592_ (_11446_, _11445_, _02150_);
  or _43593_ (_11447_, _11446_, _11442_);
  and _43594_ (_11448_, _11447_, _02144_);
  or _43595_ (_11449_, _11448_, _11438_);
  and _43596_ (_11450_, _11449_, _02157_);
  or _43597_ (_11451_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _43598_ (_11452_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _43599_ (_11453_, _11452_, _02150_);
  and _43600_ (_11454_, _11453_, _11451_);
  or _43601_ (_11455_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _43602_ (_11456_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _43603_ (_11457_, _11456_, _01954_);
  and _43604_ (_11458_, _11457_, _11455_);
  or _43605_ (_11459_, _11458_, _11454_);
  and _43606_ (_11460_, _11459_, _02131_);
  or _43607_ (_11461_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _43608_ (_11462_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _43609_ (_11463_, _11462_, _02150_);
  and _43610_ (_11464_, _11463_, _11461_);
  or _43611_ (_11465_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _43612_ (_11466_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _43613_ (_11467_, _11466_, _01954_);
  and _43614_ (_11468_, _11467_, _11465_);
  or _43615_ (_11469_, _11468_, _11464_);
  and _43616_ (_11470_, _11469_, _02144_);
  or _43617_ (_11471_, _11470_, _11460_);
  and _43618_ (_11472_, _11471_, _02077_);
  or _43619_ (_11473_, _11472_, _11450_);
  and _43620_ (_11474_, _11473_, _02194_);
  and _43621_ (_11475_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _43622_ (_11476_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _43623_ (_11477_, _11476_, _11475_);
  and _43624_ (_11478_, _11477_, _01954_);
  and _43625_ (_11479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and _43626_ (_11480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _43627_ (_11481_, _11480_, _11479_);
  and _43628_ (_11482_, _11481_, _02150_);
  or _43629_ (_11483_, _11482_, _11478_);
  and _43630_ (_11484_, _11483_, _02131_);
  and _43631_ (_11485_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _43632_ (_11486_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _43633_ (_11487_, _11486_, _11485_);
  and _43634_ (_11488_, _11487_, _01954_);
  and _43635_ (_11489_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _43636_ (_11490_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _43637_ (_11491_, _11490_, _11489_);
  and _43638_ (_11492_, _11491_, _02150_);
  or _43639_ (_11493_, _11492_, _11488_);
  and _43640_ (_11494_, _11493_, _02144_);
  or _43641_ (_11495_, _11494_, _11484_);
  and _43642_ (_11496_, _11495_, _02157_);
  or _43643_ (_11497_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _43644_ (_11498_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _43645_ (_11499_, _11498_, _11497_);
  and _43646_ (_11500_, _11499_, _01954_);
  or _43647_ (_11501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _43648_ (_11502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _43649_ (_11503_, _11502_, _11501_);
  and _43650_ (_11504_, _11503_, _02150_);
  or _43651_ (_11505_, _11504_, _11500_);
  and _43652_ (_11506_, _11505_, _02131_);
  or _43653_ (_11507_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _43654_ (_11508_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _43655_ (_11509_, _11508_, _11507_);
  and _43656_ (_11510_, _11509_, _01954_);
  or _43657_ (_11511_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _43658_ (_11512_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _43659_ (_11513_, _11512_, _11511_);
  and _43660_ (_11514_, _11513_, _02150_);
  or _43661_ (_11515_, _11514_, _11510_);
  and _43662_ (_11516_, _11515_, _02144_);
  or _43663_ (_11517_, _11516_, _11506_);
  and _43664_ (_11518_, _11517_, _02077_);
  or _43665_ (_11519_, _11518_, _11496_);
  and _43666_ (_11520_, _11519_, _02065_);
  or _43667_ (_11521_, _11520_, _11474_);
  and _43668_ (_11522_, _11521_, _02005_);
  or _43669_ (_11523_, _11522_, _11428_);
  or _43670_ (_11524_, _11523_, _02054_);
  and _43671_ (_11525_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _43672_ (_11526_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _43673_ (_11527_, _11526_, _11525_);
  and _43674_ (_11528_, _11527_, _01954_);
  and _43675_ (_11529_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _43676_ (_11530_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _43677_ (_11531_, _11530_, _11529_);
  and _43678_ (_11532_, _11531_, _02150_);
  or _43679_ (_11533_, _11532_, _11528_);
  or _43680_ (_11534_, _11533_, _02144_);
  and _43681_ (_11535_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _43682_ (_11536_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _43683_ (_11537_, _11536_, _11535_);
  and _43684_ (_11538_, _11537_, _01954_);
  and _43685_ (_11539_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _43686_ (_11540_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _43687_ (_11541_, _11540_, _11539_);
  and _43688_ (_11542_, _11541_, _02150_);
  or _43689_ (_11543_, _11542_, _11538_);
  or _43690_ (_11544_, _11543_, _02131_);
  and _43691_ (_11545_, _11544_, _02157_);
  and _43692_ (_11546_, _11545_, _11534_);
  or _43693_ (_11547_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _43694_ (_11548_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _43695_ (_11549_, _11548_, _02150_);
  and _43696_ (_11550_, _11549_, _11547_);
  or _43697_ (_11551_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _43698_ (_11552_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _43699_ (_11553_, _11552_, _01954_);
  and _43700_ (_11554_, _11553_, _11551_);
  or _43701_ (_11555_, _11554_, _11550_);
  or _43702_ (_11556_, _11555_, _02144_);
  or _43703_ (_11557_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _43704_ (_11558_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _43705_ (_11559_, _11558_, _02150_);
  and _43706_ (_11560_, _11559_, _11557_);
  or _43707_ (_11561_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _43708_ (_11562_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and _43709_ (_11563_, _11562_, _01954_);
  and _43710_ (_11564_, _11563_, _11561_);
  or _43711_ (_11565_, _11564_, _11560_);
  or _43712_ (_11566_, _11565_, _02131_);
  and _43713_ (_11567_, _11566_, _02077_);
  and _43714_ (_11568_, _11567_, _11556_);
  or _43715_ (_11569_, _11568_, _11546_);
  and _43716_ (_11570_, _11569_, _02194_);
  and _43717_ (_11571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _43718_ (_11572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _43719_ (_11573_, _11572_, _11571_);
  and _43720_ (_11574_, _11573_, _01954_);
  and _43721_ (_11575_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _43722_ (_11576_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _43723_ (_11577_, _11576_, _11575_);
  and _43724_ (_11578_, _11577_, _02150_);
  or _43725_ (_11579_, _11578_, _11574_);
  or _43726_ (_11580_, _11579_, _02144_);
  and _43727_ (_11581_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _43728_ (_11582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _43729_ (_11583_, _11582_, _11581_);
  and _43730_ (_11584_, _11583_, _01954_);
  and _43731_ (_11585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _43732_ (_11586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _43733_ (_11587_, _11586_, _11585_);
  and _43734_ (_11588_, _11587_, _02150_);
  or _43735_ (_11589_, _11588_, _11584_);
  or _43736_ (_11590_, _11589_, _02131_);
  and _43737_ (_11591_, _11590_, _02157_);
  and _43738_ (_11592_, _11591_, _11580_);
  or _43739_ (_11593_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _43740_ (_11594_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _43741_ (_11595_, _11594_, _11593_);
  and _43742_ (_11596_, _11595_, _01954_);
  or _43743_ (_11597_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _43744_ (_11598_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _43745_ (_11599_, _11598_, _11597_);
  and _43746_ (_11600_, _11599_, _02150_);
  or _43747_ (_11601_, _11600_, _11596_);
  or _43748_ (_11602_, _11601_, _02144_);
  or _43749_ (_11603_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _43750_ (_11604_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _43751_ (_11605_, _11604_, _11603_);
  and _43752_ (_11606_, _11605_, _01954_);
  or _43753_ (_11607_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _43754_ (_11608_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _43755_ (_11609_, _11608_, _11607_);
  and _43756_ (_11610_, _11609_, _02150_);
  or _43757_ (_11611_, _11610_, _11606_);
  or _43758_ (_11612_, _11611_, _02131_);
  and _43759_ (_11613_, _11612_, _02077_);
  and _43760_ (_11614_, _11613_, _11602_);
  or _43761_ (_11615_, _11614_, _11592_);
  and _43762_ (_11616_, _11615_, _02065_);
  or _43763_ (_11617_, _11616_, _11570_);
  and _43764_ (_11618_, _11617_, _02143_);
  or _43765_ (_11619_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _43766_ (_11620_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _43767_ (_11621_, _11620_, _11619_);
  and _43768_ (_11622_, _11621_, _01954_);
  or _43769_ (_11623_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _43770_ (_11624_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and _43771_ (_11625_, _11624_, _11623_);
  and _43772_ (_11626_, _11625_, _02150_);
  or _43773_ (_11627_, _11626_, _11622_);
  and _43774_ (_11628_, _11627_, _02144_);
  or _43775_ (_11629_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _43776_ (_11630_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _43777_ (_11631_, _11630_, _11629_);
  and _43778_ (_11632_, _11631_, _01954_);
  or _43779_ (_11633_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _43780_ (_11634_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _43781_ (_11635_, _11634_, _11633_);
  and _43782_ (_11636_, _11635_, _02150_);
  or _43783_ (_11637_, _11636_, _11632_);
  and _43784_ (_11638_, _11637_, _02131_);
  or _43785_ (_11639_, _11638_, _11628_);
  and _43786_ (_11640_, _11639_, _02077_);
  and _43787_ (_11641_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _43788_ (_11642_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _43789_ (_11643_, _11642_, _11641_);
  and _43790_ (_11644_, _11643_, _01954_);
  and _43791_ (_11645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _43792_ (_11646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _43793_ (_11647_, _11646_, _11645_);
  and _43794_ (_11648_, _11647_, _02150_);
  or _43795_ (_11649_, _11648_, _11644_);
  and _43796_ (_11650_, _11649_, _02144_);
  and _43797_ (_11651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _43798_ (_11652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _43799_ (_11653_, _11652_, _11651_);
  and _43800_ (_11654_, _11653_, _01954_);
  and _43801_ (_11655_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _43802_ (_11656_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _43803_ (_11657_, _11656_, _11655_);
  and _43804_ (_11658_, _11657_, _02150_);
  or _43805_ (_11659_, _11658_, _11654_);
  and _43806_ (_11660_, _11659_, _02131_);
  or _43807_ (_11661_, _11660_, _11650_);
  and _43808_ (_11662_, _11661_, _02157_);
  or _43809_ (_11663_, _11662_, _11640_);
  and _43810_ (_11664_, _11663_, _02065_);
  or _43811_ (_11665_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _43812_ (_11666_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and _43813_ (_11667_, _11666_, _02150_);
  and _43814_ (_11668_, _11667_, _11665_);
  or _43815_ (_11669_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _43816_ (_11670_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _43817_ (_11671_, _11670_, _01954_);
  and _43818_ (_11672_, _11671_, _11669_);
  or _43819_ (_11673_, _11672_, _11668_);
  and _43820_ (_11674_, _11673_, _02144_);
  or _43821_ (_11675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _43822_ (_11676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and _43823_ (_11677_, _11676_, _02150_);
  and _43824_ (_11678_, _11677_, _11675_);
  or _43825_ (_11679_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _43826_ (_11680_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _43827_ (_11681_, _11680_, _01954_);
  and _43828_ (_11682_, _11681_, _11679_);
  or _43829_ (_11683_, _11682_, _11678_);
  and _43830_ (_11684_, _11683_, _02131_);
  or _43831_ (_11685_, _11684_, _11674_);
  and _43832_ (_11686_, _11685_, _02077_);
  and _43833_ (_11687_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _43834_ (_11688_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _43835_ (_11689_, _11688_, _11687_);
  and _43836_ (_11690_, _11689_, _01954_);
  and _43837_ (_11691_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and _43838_ (_11692_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _43839_ (_11693_, _11692_, _11691_);
  and _43840_ (_11694_, _11693_, _02150_);
  or _43841_ (_11695_, _11694_, _11690_);
  and _43842_ (_11696_, _11695_, _02144_);
  and _43843_ (_11697_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and _43844_ (_11698_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _43845_ (_11699_, _11698_, _11697_);
  and _43846_ (_11700_, _11699_, _01954_);
  and _43847_ (_11701_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _43848_ (_11702_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _43849_ (_11703_, _11702_, _11701_);
  and _43850_ (_11704_, _11703_, _02150_);
  or _43851_ (_11705_, _11704_, _11700_);
  and _43852_ (_11706_, _11705_, _02131_);
  or _43853_ (_11707_, _11706_, _11696_);
  and _43854_ (_11708_, _11707_, _02157_);
  or _43855_ (_11709_, _11708_, _11686_);
  and _43856_ (_11710_, _11709_, _02194_);
  or _43857_ (_11711_, _11710_, _11664_);
  and _43858_ (_11712_, _11711_, _02005_);
  or _43859_ (_11713_, _11712_, _11618_);
  or _43860_ (_11714_, _11713_, _02374_);
  and _43861_ (_11715_, _11714_, _11524_);
  or _43862_ (_11716_, _11715_, _02142_);
  and _43863_ (_11717_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _43864_ (_11718_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _43865_ (_11719_, _11718_, _11717_);
  and _43866_ (_11720_, _11719_, _01954_);
  and _43867_ (_11721_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and _43868_ (_11722_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _43869_ (_11723_, _11722_, _11721_);
  and _43870_ (_11724_, _11723_, _02150_);
  or _43871_ (_11725_, _11724_, _11720_);
  or _43872_ (_11726_, _11725_, _02144_);
  and _43873_ (_11727_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _43874_ (_11728_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _43875_ (_11729_, _11728_, _11727_);
  and _43876_ (_11730_, _11729_, _01954_);
  and _43877_ (_11731_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and _43878_ (_11732_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _43879_ (_11733_, _11732_, _11731_);
  and _43880_ (_11734_, _11733_, _02150_);
  or _43881_ (_11735_, _11734_, _11730_);
  or _43882_ (_11736_, _11735_, _02131_);
  and _43883_ (_11737_, _11736_, _02157_);
  and _43884_ (_11738_, _11737_, _11726_);
  or _43885_ (_11739_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _43886_ (_11740_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _43887_ (_11741_, _11740_, _11739_);
  and _43888_ (_11742_, _11741_, _01954_);
  or _43889_ (_11743_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _43890_ (_11744_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and _43891_ (_11745_, _11744_, _11743_);
  and _43892_ (_11746_, _11745_, _02150_);
  or _43893_ (_11747_, _11746_, _11742_);
  or _43894_ (_11748_, _11747_, _02144_);
  or _43895_ (_11749_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _43896_ (_11750_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _43897_ (_11751_, _11750_, _11749_);
  and _43898_ (_11752_, _11751_, _01954_);
  or _43899_ (_11753_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _43900_ (_11754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _43901_ (_11755_, _11754_, _11753_);
  and _43902_ (_11756_, _11755_, _02150_);
  or _43903_ (_11757_, _11756_, _11752_);
  or _43904_ (_11758_, _11757_, _02131_);
  and _43905_ (_11759_, _11758_, _02077_);
  and _43906_ (_11760_, _11759_, _11748_);
  or _43907_ (_11761_, _11760_, _11738_);
  and _43908_ (_11762_, _11761_, _02065_);
  and _43909_ (_11763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _43910_ (_11764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _43911_ (_11765_, _11764_, _11763_);
  and _43912_ (_11766_, _11765_, _01954_);
  and _43913_ (_11767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _43914_ (_11768_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _43915_ (_11769_, _11768_, _11767_);
  and _43916_ (_11770_, _11769_, _02150_);
  or _43917_ (_11771_, _11770_, _11766_);
  or _43918_ (_11772_, _11771_, _02144_);
  and _43919_ (_11773_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _43920_ (_11774_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _43921_ (_11775_, _11774_, _11773_);
  and _43922_ (_11776_, _11775_, _01954_);
  and _43923_ (_11777_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _43924_ (_11778_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _43925_ (_11779_, _11778_, _11777_);
  and _43926_ (_11780_, _11779_, _02150_);
  or _43927_ (_11781_, _11780_, _11776_);
  or _43928_ (_11782_, _11781_, _02131_);
  and _43929_ (_11783_, _11782_, _02157_);
  and _43930_ (_11784_, _11783_, _11772_);
  or _43931_ (_11785_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _43932_ (_11786_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _43933_ (_11787_, _11786_, _02150_);
  and _43934_ (_11788_, _11787_, _11785_);
  or _43935_ (_11789_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _43936_ (_11790_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _43937_ (_11791_, _11790_, _01954_);
  and _43938_ (_11792_, _11791_, _11789_);
  or _43939_ (_11793_, _11792_, _11788_);
  or _43940_ (_11794_, _11793_, _02144_);
  or _43941_ (_11795_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _43942_ (_11796_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _43943_ (_11797_, _11796_, _02150_);
  and _43944_ (_11798_, _11797_, _11795_);
  or _43945_ (_11799_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _43946_ (_11800_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _43947_ (_11801_, _11800_, _01954_);
  and _43948_ (_11802_, _11801_, _11799_);
  or _43949_ (_11803_, _11802_, _11798_);
  or _43950_ (_11804_, _11803_, _02131_);
  and _43951_ (_11805_, _11804_, _02077_);
  and _43952_ (_11806_, _11805_, _11794_);
  or _43953_ (_11807_, _11806_, _11784_);
  and _43954_ (_11808_, _11807_, _02194_);
  or _43955_ (_11809_, _11808_, _11762_);
  and _43956_ (_11810_, _11809_, _02143_);
  and _43957_ (_11811_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _43958_ (_11812_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _43959_ (_11813_, _11812_, _11811_);
  and _43960_ (_11814_, _11813_, _01954_);
  and _43961_ (_11815_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _43962_ (_11816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _43963_ (_11817_, _11816_, _11815_);
  and _43964_ (_11818_, _11817_, _02150_);
  or _43965_ (_11819_, _11818_, _11814_);
  and _43966_ (_11820_, _11819_, _02131_);
  and _43967_ (_11821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _43968_ (_11822_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _43969_ (_11823_, _11822_, _11821_);
  and _43970_ (_11824_, _11823_, _01954_);
  and _43971_ (_11825_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _43972_ (_11826_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _43973_ (_11827_, _11826_, _11825_);
  and _43974_ (_11828_, _11827_, _02150_);
  or _43975_ (_11829_, _11828_, _11824_);
  and _43976_ (_11830_, _11829_, _02144_);
  or _43977_ (_11831_, _11830_, _11820_);
  and _43978_ (_11832_, _11831_, _02157_);
  or _43979_ (_11833_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _43980_ (_11834_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _43981_ (_11835_, _11834_, _02150_);
  and _43982_ (_11836_, _11835_, _11833_);
  or _43983_ (_11837_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _43984_ (_11838_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _43985_ (_11839_, _11838_, _01954_);
  and _43986_ (_11840_, _11839_, _11837_);
  or _43987_ (_11841_, _11840_, _11836_);
  and _43988_ (_11842_, _11841_, _02131_);
  or _43989_ (_11843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _43990_ (_11844_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _43991_ (_11845_, _11844_, _02150_);
  and _43992_ (_11846_, _11845_, _11843_);
  or _43993_ (_11847_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _43994_ (_11848_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _43995_ (_11849_, _11848_, _01954_);
  and _43996_ (_11850_, _11849_, _11847_);
  or _43997_ (_11851_, _11850_, _11846_);
  and _43998_ (_11852_, _11851_, _02144_);
  or _43999_ (_11853_, _11852_, _11842_);
  and _44000_ (_11854_, _11853_, _02077_);
  or _44001_ (_11855_, _11854_, _11832_);
  and _44002_ (_11856_, _11855_, _02194_);
  and _44003_ (_11857_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _44004_ (_11858_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _44005_ (_11859_, _11858_, _11857_);
  and _44006_ (_11860_, _11859_, _01954_);
  and _44007_ (_11861_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _44008_ (_11862_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _44009_ (_11863_, _11862_, _11861_);
  and _44010_ (_11864_, _11863_, _02150_);
  or _44011_ (_11865_, _11864_, _11860_);
  and _44012_ (_11866_, _11865_, _02131_);
  and _44013_ (_11867_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _44014_ (_11868_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _44015_ (_11869_, _11868_, _11867_);
  and _44016_ (_11870_, _11869_, _01954_);
  and _44017_ (_11871_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _44018_ (_11872_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _44019_ (_11873_, _11872_, _11871_);
  and _44020_ (_11874_, _11873_, _02150_);
  or _44021_ (_11875_, _11874_, _11870_);
  and _44022_ (_11876_, _11875_, _02144_);
  or _44023_ (_11877_, _11876_, _11866_);
  and _44024_ (_11878_, _11877_, _02157_);
  or _44025_ (_11879_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _44026_ (_11880_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _44027_ (_11881_, _11880_, _11879_);
  and _44028_ (_11882_, _11881_, _01954_);
  or _44029_ (_11883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _44030_ (_11884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _44031_ (_11885_, _11884_, _11883_);
  and _44032_ (_11886_, _11885_, _02150_);
  or _44033_ (_11887_, _11886_, _11882_);
  and _44034_ (_11888_, _11887_, _02131_);
  or _44035_ (_11889_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _44036_ (_11890_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _44037_ (_11891_, _11890_, _11889_);
  and _44038_ (_11892_, _11891_, _01954_);
  or _44039_ (_11893_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _44040_ (_11894_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _44041_ (_11895_, _11894_, _11893_);
  and _44042_ (_11896_, _11895_, _02150_);
  or _44043_ (_11897_, _11896_, _11892_);
  and _44044_ (_11898_, _11897_, _02144_);
  or _44045_ (_11899_, _11898_, _11888_);
  and _44046_ (_11900_, _11899_, _02077_);
  or _44047_ (_11901_, _11900_, _11878_);
  and _44048_ (_11902_, _11901_, _02065_);
  or _44049_ (_11903_, _11902_, _11856_);
  and _44050_ (_11904_, _11903_, _02005_);
  or _44051_ (_11905_, _11904_, _11810_);
  or _44052_ (_11906_, _11905_, _02054_);
  and _44053_ (_11907_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _44054_ (_11908_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _44055_ (_11909_, _11908_, _11907_);
  and _44056_ (_11910_, _11909_, _01954_);
  and _44057_ (_11911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and _44058_ (_11912_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _44059_ (_11913_, _11912_, _11911_);
  and _44060_ (_11914_, _11913_, _02150_);
  or _44061_ (_11915_, _11914_, _11910_);
  or _44062_ (_11916_, _11915_, _02144_);
  and _44063_ (_11917_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _44064_ (_11918_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _44065_ (_11919_, _11918_, _11917_);
  and _44066_ (_11920_, _11919_, _01954_);
  and _44067_ (_11921_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _44068_ (_11922_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _44069_ (_11923_, _11922_, _11921_);
  and _44070_ (_11924_, _11923_, _02150_);
  or _44071_ (_11925_, _11924_, _11920_);
  or _44072_ (_11926_, _11925_, _02131_);
  and _44073_ (_11927_, _11926_, _02157_);
  and _44074_ (_11928_, _11927_, _11916_);
  or _44075_ (_11929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _44076_ (_11930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and _44077_ (_11931_, _11930_, _02150_);
  and _44078_ (_11932_, _11931_, _11929_);
  or _44079_ (_11933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _44080_ (_11934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _44081_ (_11935_, _11934_, _01954_);
  and _44082_ (_11936_, _11935_, _11933_);
  or _44083_ (_11937_, _11936_, _11932_);
  or _44084_ (_11938_, _11937_, _02144_);
  or _44085_ (_11939_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _44086_ (_11940_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _44087_ (_11941_, _11940_, _02150_);
  and _44088_ (_11942_, _11941_, _11939_);
  or _44089_ (_11943_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _44090_ (_11944_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _44091_ (_11945_, _11944_, _01954_);
  and _44092_ (_11946_, _11945_, _11943_);
  or _44093_ (_11947_, _11946_, _11942_);
  or _44094_ (_11948_, _11947_, _02131_);
  and _44095_ (_11949_, _11948_, _02077_);
  and _44096_ (_11950_, _11949_, _11938_);
  or _44097_ (_11951_, _11950_, _11928_);
  and _44098_ (_11952_, _11951_, _02194_);
  and _44099_ (_11953_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _44100_ (_11954_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _44101_ (_11955_, _11954_, _11953_);
  and _44102_ (_11956_, _11955_, _01954_);
  and _44103_ (_11957_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _44104_ (_11958_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _44105_ (_11959_, _11958_, _11957_);
  and _44106_ (_11960_, _11959_, _02150_);
  or _44107_ (_11961_, _11960_, _11956_);
  or _44108_ (_11962_, _11961_, _02144_);
  and _44109_ (_11963_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _44110_ (_11964_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _44111_ (_11965_, _11964_, _11963_);
  and _44112_ (_11966_, _11965_, _01954_);
  and _44113_ (_11967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _44114_ (_11968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _44115_ (_11969_, _11968_, _11967_);
  and _44116_ (_11970_, _11969_, _02150_);
  or _44117_ (_11971_, _11970_, _11966_);
  or _44118_ (_11972_, _11971_, _02131_);
  and _44119_ (_11973_, _11972_, _02157_);
  and _44120_ (_11974_, _11973_, _11962_);
  or _44121_ (_11975_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _44122_ (_11976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _44123_ (_11977_, _11976_, _11975_);
  and _44124_ (_11978_, _11977_, _01954_);
  or _44125_ (_11979_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _44126_ (_11980_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _44127_ (_11981_, _11980_, _11979_);
  and _44128_ (_11982_, _11981_, _02150_);
  or _44129_ (_11983_, _11982_, _11978_);
  or _44130_ (_11984_, _11983_, _02144_);
  or _44131_ (_11985_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _44132_ (_11986_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _44133_ (_11987_, _11986_, _11985_);
  and _44134_ (_11988_, _11987_, _01954_);
  or _44135_ (_11989_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _44136_ (_11990_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _44137_ (_11991_, _11990_, _11989_);
  and _44138_ (_11992_, _11991_, _02150_);
  or _44139_ (_11993_, _11992_, _11988_);
  or _44140_ (_11994_, _11993_, _02131_);
  and _44141_ (_11995_, _11994_, _02077_);
  and _44142_ (_11996_, _11995_, _11984_);
  or _44143_ (_11997_, _11996_, _11974_);
  and _44144_ (_11998_, _11997_, _02065_);
  or _44145_ (_11999_, _11998_, _11952_);
  and _44146_ (_12000_, _11999_, _02143_);
  or _44147_ (_12001_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _44148_ (_12002_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _44149_ (_12003_, _12002_, _12001_);
  and _44150_ (_12004_, _12003_, _01954_);
  or _44151_ (_12005_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _44152_ (_12006_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _44153_ (_12007_, _12006_, _12005_);
  and _44154_ (_12008_, _12007_, _02150_);
  or _44155_ (_12009_, _12008_, _12004_);
  and _44156_ (_12010_, _12009_, _02144_);
  or _44157_ (_12011_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _44158_ (_12012_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _44159_ (_12013_, _12012_, _12011_);
  and _44160_ (_12014_, _12013_, _01954_);
  or _44161_ (_12015_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _44162_ (_12016_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _44163_ (_12017_, _12016_, _12015_);
  and _44164_ (_12018_, _12017_, _02150_);
  or _44165_ (_12019_, _12018_, _12014_);
  and _44166_ (_12020_, _12019_, _02131_);
  or _44167_ (_12021_, _12020_, _12010_);
  and _44168_ (_12022_, _12021_, _02077_);
  and _44169_ (_12023_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _44170_ (_12024_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _44171_ (_12025_, _12024_, _12023_);
  and _44172_ (_12026_, _12025_, _01954_);
  and _44173_ (_12027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _44174_ (_12028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _44175_ (_12029_, _12028_, _12027_);
  and _44176_ (_12030_, _12029_, _02150_);
  or _44177_ (_12031_, _12030_, _12026_);
  and _44178_ (_12032_, _12031_, _02144_);
  and _44179_ (_12033_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _44180_ (_12034_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _44181_ (_12035_, _12034_, _12033_);
  and _44182_ (_12036_, _12035_, _01954_);
  and _44183_ (_12037_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _44184_ (_12038_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _44185_ (_12039_, _12038_, _12037_);
  and _44186_ (_12040_, _12039_, _02150_);
  or _44187_ (_12041_, _12040_, _12036_);
  and _44188_ (_12042_, _12041_, _02131_);
  or _44189_ (_12043_, _12042_, _12032_);
  and _44190_ (_12044_, _12043_, _02157_);
  or _44191_ (_12045_, _12044_, _12022_);
  and _44192_ (_12046_, _12045_, _02065_);
  or _44193_ (_12047_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _44194_ (_12048_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _44195_ (_12049_, _12048_, _02150_);
  and _44196_ (_12050_, _12049_, _12047_);
  or _44197_ (_12051_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _44198_ (_12052_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _44199_ (_12053_, _12052_, _01954_);
  and _44200_ (_12054_, _12053_, _12051_);
  or _44201_ (_12055_, _12054_, _12050_);
  and _44202_ (_12056_, _12055_, _02144_);
  or _44203_ (_12057_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _44204_ (_12058_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _44205_ (_12059_, _12058_, _02150_);
  and _44206_ (_12060_, _12059_, _12057_);
  or _44207_ (_12061_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _44208_ (_12062_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _44209_ (_12063_, _12062_, _01954_);
  and _44210_ (_12064_, _12063_, _12061_);
  or _44211_ (_12065_, _12064_, _12060_);
  and _44212_ (_12066_, _12065_, _02131_);
  or _44213_ (_12067_, _12066_, _12056_);
  and _44214_ (_12068_, _12067_, _02077_);
  and _44215_ (_12069_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _44216_ (_12070_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _44217_ (_12071_, _12070_, _12069_);
  and _44218_ (_12072_, _12071_, _01954_);
  and _44219_ (_12073_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _44220_ (_12074_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _44221_ (_12075_, _12074_, _12073_);
  and _44222_ (_12076_, _12075_, _02150_);
  or _44223_ (_12077_, _12076_, _12072_);
  and _44224_ (_12078_, _12077_, _02144_);
  and _44225_ (_12079_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _44226_ (_12080_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _44227_ (_12081_, _12080_, _12079_);
  and _44228_ (_12082_, _12081_, _01954_);
  and _44229_ (_12083_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _44230_ (_12084_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _44231_ (_12085_, _12084_, _12083_);
  and _44232_ (_12086_, _12085_, _02150_);
  or _44233_ (_12087_, _12086_, _12082_);
  and _44234_ (_12088_, _12087_, _02131_);
  or _44235_ (_12089_, _12088_, _12078_);
  and _44236_ (_12090_, _12089_, _02157_);
  or _44237_ (_12091_, _12090_, _12068_);
  and _44238_ (_12092_, _12091_, _02194_);
  or _44239_ (_12093_, _12092_, _12046_);
  and _44240_ (_12094_, _12093_, _02005_);
  or _44241_ (_12095_, _12094_, _12000_);
  or _44242_ (_12096_, _12095_, _02374_);
  and _44243_ (_12097_, _12096_, _11906_);
  or _44244_ (_12098_, _12097_, _01748_);
  and _44245_ (_12099_, _12098_, _11716_);
  or _44246_ (_12100_, _12099_, _02141_);
  or _44247_ (_12101_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _44248_ (_12102_, _12101_, _27355_);
  and _44249_ (_15240_, _12102_, _12100_);
  and _44250_ (_12103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _44251_ (_12104_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _44252_ (_12105_, _12104_, _12103_);
  and _44253_ (_12106_, _12105_, _01954_);
  and _44254_ (_12107_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _44255_ (_12108_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _44256_ (_12109_, _12108_, _12107_);
  and _44257_ (_12110_, _12109_, _02150_);
  or _44258_ (_12111_, _12110_, _12106_);
  or _44259_ (_12112_, _12111_, _02144_);
  and _44260_ (_12113_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _44261_ (_12114_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _44262_ (_12115_, _12114_, _12113_);
  and _44263_ (_12116_, _12115_, _01954_);
  and _44264_ (_12117_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and _44265_ (_12118_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _44266_ (_12119_, _12118_, _12117_);
  and _44267_ (_12120_, _12119_, _02150_);
  or _44268_ (_12121_, _12120_, _12116_);
  or _44269_ (_12122_, _12121_, _02131_);
  and _44270_ (_12123_, _12122_, _02157_);
  and _44271_ (_12124_, _12123_, _12112_);
  or _44272_ (_12125_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _44273_ (_12126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and _44274_ (_12127_, _12126_, _12125_);
  and _44275_ (_12128_, _12127_, _01954_);
  or _44276_ (_12129_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _44277_ (_12130_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _44278_ (_12131_, _12130_, _12129_);
  and _44279_ (_12132_, _12131_, _02150_);
  or _44280_ (_12133_, _12132_, _12128_);
  or _44281_ (_12134_, _12133_, _02144_);
  or _44282_ (_12135_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _44283_ (_12136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _44284_ (_12137_, _12136_, _12135_);
  and _44285_ (_12138_, _12137_, _01954_);
  or _44286_ (_12139_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _44287_ (_12140_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _44288_ (_12141_, _12140_, _12139_);
  and _44289_ (_12142_, _12141_, _02150_);
  or _44290_ (_12143_, _12142_, _12138_);
  or _44291_ (_12144_, _12143_, _02131_);
  and _44292_ (_12145_, _12144_, _02077_);
  and _44293_ (_12146_, _12145_, _12134_);
  or _44294_ (_12147_, _12146_, _12124_);
  and _44295_ (_12148_, _12147_, _02065_);
  and _44296_ (_12149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _44297_ (_12150_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _44298_ (_12151_, _12150_, _12149_);
  and _44299_ (_12152_, _12151_, _01954_);
  and _44300_ (_12153_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _44301_ (_12154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _44302_ (_12155_, _12154_, _12153_);
  and _44303_ (_12156_, _12155_, _02150_);
  or _44304_ (_12157_, _12156_, _12152_);
  or _44305_ (_12158_, _12157_, _02144_);
  and _44306_ (_12159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and _44307_ (_12160_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _44308_ (_12161_, _12160_, _12159_);
  and _44309_ (_12162_, _12161_, _01954_);
  and _44310_ (_12163_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _44311_ (_12164_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _44312_ (_12165_, _12164_, _12163_);
  and _44313_ (_12166_, _12165_, _02150_);
  or _44314_ (_12167_, _12166_, _12162_);
  or _44315_ (_12168_, _12167_, _02131_);
  and _44316_ (_12169_, _12168_, _02157_);
  and _44317_ (_12170_, _12169_, _12158_);
  or _44318_ (_12171_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _44319_ (_12172_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _44320_ (_12173_, _12172_, _02150_);
  and _44321_ (_12174_, _12173_, _12171_);
  or _44322_ (_12175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _44323_ (_12176_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _44324_ (_12177_, _12176_, _01954_);
  and _44325_ (_12178_, _12177_, _12175_);
  or _44326_ (_12179_, _12178_, _12174_);
  or _44327_ (_12180_, _12179_, _02144_);
  or _44328_ (_12181_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _44329_ (_12182_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and _44330_ (_12183_, _12182_, _02150_);
  and _44331_ (_12184_, _12183_, _12181_);
  or _44332_ (_12185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _44333_ (_12186_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _44334_ (_12187_, _12186_, _01954_);
  and _44335_ (_12188_, _12187_, _12185_);
  or _44336_ (_12189_, _12188_, _12184_);
  or _44337_ (_12190_, _12189_, _02131_);
  and _44338_ (_12191_, _12190_, _02077_);
  and _44339_ (_12192_, _12191_, _12180_);
  or _44340_ (_12193_, _12192_, _12170_);
  and _44341_ (_12194_, _12193_, _02194_);
  or _44342_ (_12195_, _12194_, _12148_);
  and _44343_ (_12196_, _12195_, _02143_);
  and _44344_ (_12197_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _44345_ (_12198_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _44346_ (_12199_, _12198_, _12197_);
  and _44347_ (_12200_, _12199_, _01954_);
  and _44348_ (_12201_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _44349_ (_12202_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _44350_ (_12203_, _12202_, _12201_);
  and _44351_ (_12204_, _12203_, _02150_);
  or _44352_ (_12205_, _12204_, _12200_);
  and _44353_ (_12206_, _12205_, _02131_);
  and _44354_ (_12207_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _44355_ (_12208_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _44356_ (_12209_, _12208_, _12207_);
  and _44357_ (_12210_, _12209_, _01954_);
  and _44358_ (_12211_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _44359_ (_12212_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _44360_ (_12213_, _12212_, _12211_);
  and _44361_ (_12214_, _12213_, _02150_);
  or _44362_ (_12215_, _12214_, _12210_);
  and _44363_ (_12216_, _12215_, _02144_);
  or _44364_ (_12217_, _12216_, _12206_);
  and _44365_ (_12218_, _12217_, _02157_);
  or _44366_ (_12219_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _44367_ (_12220_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _44368_ (_12221_, _12220_, _02150_);
  and _44369_ (_12222_, _12221_, _12219_);
  or _44370_ (_12223_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _44371_ (_12224_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _44372_ (_12225_, _12224_, _01954_);
  and _44373_ (_12226_, _12225_, _12223_);
  or _44374_ (_12227_, _12226_, _12222_);
  and _44375_ (_12228_, _12227_, _02131_);
  or _44376_ (_12229_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _44377_ (_12230_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _44378_ (_12231_, _12230_, _02150_);
  and _44379_ (_12232_, _12231_, _12229_);
  or _44380_ (_12233_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _44381_ (_12234_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _44382_ (_12235_, _12234_, _01954_);
  and _44383_ (_12236_, _12235_, _12233_);
  or _44384_ (_12237_, _12236_, _12232_);
  and _44385_ (_12238_, _12237_, _02144_);
  or _44386_ (_12239_, _12238_, _12228_);
  and _44387_ (_12240_, _12239_, _02077_);
  or _44388_ (_12241_, _12240_, _12218_);
  and _44389_ (_12242_, _12241_, _02194_);
  and _44390_ (_12243_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _44391_ (_12244_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _44392_ (_12245_, _12244_, _12243_);
  and _44393_ (_12246_, _12245_, _01954_);
  and _44394_ (_12247_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _44395_ (_12248_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _44396_ (_12249_, _12248_, _12247_);
  and _44397_ (_12250_, _12249_, _02150_);
  or _44398_ (_12251_, _12250_, _12246_);
  and _44399_ (_12252_, _12251_, _02131_);
  and _44400_ (_12253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _44401_ (_12254_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _44402_ (_12255_, _12254_, _12253_);
  and _44403_ (_12256_, _12255_, _01954_);
  and _44404_ (_12257_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and _44405_ (_12258_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _44406_ (_12259_, _12258_, _12257_);
  and _44407_ (_12260_, _12259_, _02150_);
  or _44408_ (_12261_, _12260_, _12256_);
  and _44409_ (_12262_, _12261_, _02144_);
  or _44410_ (_12263_, _12262_, _12252_);
  and _44411_ (_12264_, _12263_, _02157_);
  or _44412_ (_12265_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _44413_ (_12266_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and _44414_ (_12267_, _12266_, _12265_);
  and _44415_ (_12268_, _12267_, _01954_);
  or _44416_ (_12269_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _44417_ (_12270_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _44418_ (_12271_, _12270_, _12269_);
  and _44419_ (_12272_, _12271_, _02150_);
  or _44420_ (_12273_, _12272_, _12268_);
  and _44421_ (_12274_, _12273_, _02131_);
  or _44422_ (_12275_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _44423_ (_12276_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _44424_ (_12277_, _12276_, _12275_);
  and _44425_ (_12278_, _12277_, _01954_);
  or _44426_ (_12279_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _44427_ (_12280_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _44428_ (_12281_, _12280_, _12279_);
  and _44429_ (_12282_, _12281_, _02150_);
  or _44430_ (_12283_, _12282_, _12278_);
  and _44431_ (_12284_, _12283_, _02144_);
  or _44432_ (_12285_, _12284_, _12274_);
  and _44433_ (_12286_, _12285_, _02077_);
  or _44434_ (_12287_, _12286_, _12264_);
  and _44435_ (_12288_, _12287_, _02065_);
  or _44436_ (_12289_, _12288_, _12242_);
  and _44437_ (_12290_, _12289_, _02005_);
  or _44438_ (_12291_, _12290_, _12196_);
  or _44439_ (_12292_, _12291_, _02054_);
  and _44440_ (_12293_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _44441_ (_12294_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _44442_ (_12295_, _12294_, _12293_);
  and _44443_ (_12296_, _12295_, _01954_);
  and _44444_ (_12297_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and _44445_ (_12298_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _44446_ (_12299_, _12298_, _12297_);
  and _44447_ (_12300_, _12299_, _02150_);
  or _44448_ (_12301_, _12300_, _12296_);
  or _44449_ (_12302_, _12301_, _02144_);
  and _44450_ (_12303_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _44451_ (_12304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _44452_ (_12305_, _12304_, _12303_);
  and _44453_ (_12306_, _12305_, _01954_);
  and _44454_ (_12307_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _44455_ (_12308_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _44456_ (_12309_, _12308_, _12307_);
  and _44457_ (_12310_, _12309_, _02150_);
  or _44458_ (_12311_, _12310_, _12306_);
  or _44459_ (_12312_, _12311_, _02131_);
  and _44460_ (_12313_, _12312_, _02157_);
  and _44461_ (_12314_, _12313_, _12302_);
  or _44462_ (_12315_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _44463_ (_12316_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and _44464_ (_12317_, _12316_, _02150_);
  and _44465_ (_12318_, _12317_, _12315_);
  or _44466_ (_12319_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _44467_ (_12320_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _44468_ (_12321_, _12320_, _01954_);
  and _44469_ (_12322_, _12321_, _12319_);
  or _44470_ (_12323_, _12322_, _12318_);
  or _44471_ (_12324_, _12323_, _02144_);
  or _44472_ (_12325_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _44473_ (_12326_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and _44474_ (_12327_, _12326_, _02150_);
  and _44475_ (_12328_, _12327_, _12325_);
  or _44476_ (_12329_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _44477_ (_12330_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _44478_ (_12331_, _12330_, _01954_);
  and _44479_ (_12332_, _12331_, _12329_);
  or _44480_ (_12333_, _12332_, _12328_);
  or _44481_ (_12334_, _12333_, _02131_);
  and _44482_ (_12335_, _12334_, _02077_);
  and _44483_ (_12336_, _12335_, _12324_);
  or _44484_ (_12337_, _12336_, _12314_);
  and _44485_ (_12338_, _12337_, _02194_);
  and _44486_ (_12339_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _44487_ (_12340_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _44488_ (_12341_, _12340_, _12339_);
  and _44489_ (_12342_, _12341_, _01954_);
  and _44490_ (_12343_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _44491_ (_12344_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _44492_ (_12345_, _12344_, _12343_);
  and _44493_ (_12346_, _12345_, _02150_);
  or _44494_ (_12347_, _12346_, _12342_);
  or _44495_ (_12348_, _12347_, _02144_);
  and _44496_ (_12349_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _44497_ (_12350_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _44498_ (_12351_, _12350_, _12349_);
  and _44499_ (_12352_, _12351_, _01954_);
  and _44500_ (_12353_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _44501_ (_12354_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _44502_ (_12355_, _12354_, _12353_);
  and _44503_ (_12356_, _12355_, _02150_);
  or _44504_ (_12357_, _12356_, _12352_);
  or _44505_ (_12358_, _12357_, _02131_);
  and _44506_ (_12359_, _12358_, _02157_);
  and _44507_ (_12360_, _12359_, _12348_);
  or _44508_ (_12361_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _44509_ (_12362_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _44510_ (_12363_, _12362_, _12361_);
  and _44511_ (_12364_, _12363_, _01954_);
  or _44512_ (_12365_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _44513_ (_12366_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _44514_ (_12367_, _12366_, _12365_);
  and _44515_ (_12368_, _12367_, _02150_);
  or _44516_ (_12369_, _12368_, _12364_);
  or _44517_ (_12370_, _12369_, _02144_);
  or _44518_ (_12371_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _44519_ (_12372_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _44520_ (_12373_, _12372_, _12371_);
  and _44521_ (_12374_, _12373_, _01954_);
  or _44522_ (_12375_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _44523_ (_12376_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _44524_ (_12377_, _12376_, _12375_);
  and _44525_ (_12378_, _12377_, _02150_);
  or _44526_ (_12379_, _12378_, _12374_);
  or _44527_ (_12380_, _12379_, _02131_);
  and _44528_ (_12381_, _12380_, _02077_);
  and _44529_ (_12382_, _12381_, _12370_);
  or _44530_ (_12383_, _12382_, _12360_);
  and _44531_ (_12384_, _12383_, _02065_);
  or _44532_ (_12385_, _12384_, _12338_);
  and _44533_ (_12386_, _12385_, _02143_);
  or _44534_ (_12387_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _44535_ (_12388_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _44536_ (_12389_, _12388_, _12387_);
  and _44537_ (_12390_, _12389_, _01954_);
  or _44538_ (_12391_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _44539_ (_12392_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and _44540_ (_12393_, _12392_, _12391_);
  and _44541_ (_12394_, _12393_, _02150_);
  or _44542_ (_12395_, _12394_, _12390_);
  and _44543_ (_12396_, _12395_, _02144_);
  or _44544_ (_12397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _44545_ (_12398_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _44546_ (_12399_, _12398_, _12397_);
  and _44547_ (_12400_, _12399_, _01954_);
  or _44548_ (_12401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _44549_ (_12402_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _44550_ (_12403_, _12402_, _12401_);
  and _44551_ (_12404_, _12403_, _02150_);
  or _44552_ (_12405_, _12404_, _12400_);
  and _44553_ (_12406_, _12405_, _02131_);
  or _44554_ (_12407_, _12406_, _12396_);
  and _44555_ (_12408_, _12407_, _02077_);
  and _44556_ (_12409_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and _44557_ (_12410_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _44558_ (_12411_, _12410_, _12409_);
  and _44559_ (_12412_, _12411_, _01954_);
  and _44560_ (_12413_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _44561_ (_12414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _44562_ (_12415_, _12414_, _12413_);
  and _44563_ (_12416_, _12415_, _02150_);
  or _44564_ (_12417_, _12416_, _12412_);
  and _44565_ (_12418_, _12417_, _02144_);
  and _44566_ (_12419_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _44567_ (_12420_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _44568_ (_12421_, _12420_, _12419_);
  and _44569_ (_12422_, _12421_, _01954_);
  and _44570_ (_12423_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _44571_ (_12424_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _44572_ (_12425_, _12424_, _12423_);
  and _44573_ (_12426_, _12425_, _02150_);
  or _44574_ (_12427_, _12426_, _12422_);
  and _44575_ (_12428_, _12427_, _02131_);
  or _44576_ (_12429_, _12428_, _12418_);
  and _44577_ (_12430_, _12429_, _02157_);
  or _44578_ (_12431_, _12430_, _12408_);
  and _44579_ (_12432_, _12431_, _02065_);
  or _44580_ (_12433_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _44581_ (_12434_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and _44582_ (_12435_, _12434_, _02150_);
  and _44583_ (_12436_, _12435_, _12433_);
  or _44584_ (_12437_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _44585_ (_12438_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and _44586_ (_12439_, _12438_, _01954_);
  and _44587_ (_12440_, _12439_, _12437_);
  or _44588_ (_12441_, _12440_, _12436_);
  and _44589_ (_12442_, _12441_, _02144_);
  or _44590_ (_12443_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _44591_ (_12444_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _44592_ (_12445_, _12444_, _02150_);
  and _44593_ (_12446_, _12445_, _12443_);
  or _44594_ (_12447_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _44595_ (_12448_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and _44596_ (_12449_, _12448_, _01954_);
  and _44597_ (_12450_, _12449_, _12447_);
  or _44598_ (_12451_, _12450_, _12446_);
  and _44599_ (_12452_, _12451_, _02131_);
  or _44600_ (_12453_, _12452_, _12442_);
  and _44601_ (_12454_, _12453_, _02077_);
  and _44602_ (_12455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and _44603_ (_12456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _44604_ (_12457_, _12456_, _12455_);
  and _44605_ (_12458_, _12457_, _01954_);
  and _44606_ (_12459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _44607_ (_12460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _44608_ (_12461_, _12460_, _12459_);
  and _44609_ (_12462_, _12461_, _02150_);
  or _44610_ (_12463_, _12462_, _12458_);
  and _44611_ (_12464_, _12463_, _02144_);
  and _44612_ (_12465_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and _44613_ (_12466_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _44614_ (_12467_, _12466_, _12465_);
  and _44615_ (_12468_, _12467_, _01954_);
  and _44616_ (_12469_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _44617_ (_12470_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _44618_ (_12471_, _12470_, _12469_);
  and _44619_ (_12472_, _12471_, _02150_);
  or _44620_ (_12473_, _12472_, _12468_);
  and _44621_ (_12474_, _12473_, _02131_);
  or _44622_ (_12475_, _12474_, _12464_);
  and _44623_ (_12476_, _12475_, _02157_);
  or _44624_ (_12477_, _12476_, _12454_);
  and _44625_ (_12478_, _12477_, _02194_);
  or _44626_ (_12479_, _12478_, _12432_);
  and _44627_ (_12480_, _12479_, _02005_);
  or _44628_ (_12481_, _12480_, _12386_);
  or _44629_ (_12482_, _12481_, _02374_);
  and _44630_ (_12483_, _12482_, _12292_);
  or _44631_ (_12484_, _12483_, _02142_);
  and _44632_ (_12485_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _44633_ (_12486_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _44634_ (_12487_, _12486_, _12485_);
  and _44635_ (_12488_, _12487_, _01954_);
  and _44636_ (_12489_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _44637_ (_12490_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _44638_ (_12491_, _12490_, _12489_);
  and _44639_ (_12492_, _12491_, _02150_);
  or _44640_ (_12493_, _12492_, _12488_);
  or _44641_ (_12494_, _12493_, _02144_);
  and _44642_ (_12495_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _44643_ (_12496_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _44644_ (_12497_, _12496_, _12495_);
  and _44645_ (_12498_, _12497_, _01954_);
  and _44646_ (_12499_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _44647_ (_12500_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _44648_ (_12501_, _12500_, _12499_);
  and _44649_ (_12502_, _12501_, _02150_);
  or _44650_ (_12503_, _12502_, _12498_);
  or _44651_ (_12504_, _12503_, _02131_);
  and _44652_ (_12505_, _12504_, _02157_);
  and _44653_ (_12506_, _12505_, _12494_);
  or _44654_ (_12507_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _44655_ (_12508_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and _44656_ (_12509_, _12508_, _12507_);
  and _44657_ (_12510_, _12509_, _01954_);
  or _44658_ (_12511_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _44659_ (_12512_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _44660_ (_12513_, _12512_, _12511_);
  and _44661_ (_12514_, _12513_, _02150_);
  or _44662_ (_12515_, _12514_, _12510_);
  or _44663_ (_12516_, _12515_, _02144_);
  or _44664_ (_12517_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _44665_ (_12518_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _44666_ (_12519_, _12518_, _12517_);
  and _44667_ (_12520_, _12519_, _01954_);
  or _44668_ (_12521_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _44669_ (_12522_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _44670_ (_12523_, _12522_, _12521_);
  and _44671_ (_12524_, _12523_, _02150_);
  or _44672_ (_12525_, _12524_, _12520_);
  or _44673_ (_12526_, _12525_, _02131_);
  and _44674_ (_12527_, _12526_, _02077_);
  and _44675_ (_12528_, _12527_, _12516_);
  or _44676_ (_12529_, _12528_, _12506_);
  and _44677_ (_12530_, _12529_, _02065_);
  and _44678_ (_12531_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _44679_ (_12532_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _44680_ (_12533_, _12532_, _12531_);
  and _44681_ (_12534_, _12533_, _01954_);
  and _44682_ (_12535_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _44683_ (_12536_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _44684_ (_12537_, _12536_, _12535_);
  and _44685_ (_12538_, _12537_, _02150_);
  or _44686_ (_12539_, _12538_, _12534_);
  or _44687_ (_12540_, _12539_, _02144_);
  and _44688_ (_12541_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _44689_ (_12542_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _44690_ (_12543_, _12542_, _12541_);
  and _44691_ (_12544_, _12543_, _01954_);
  and _44692_ (_12545_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _44693_ (_12546_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _44694_ (_12547_, _12546_, _12545_);
  and _44695_ (_12548_, _12547_, _02150_);
  or _44696_ (_12549_, _12548_, _12544_);
  or _44697_ (_12550_, _12549_, _02131_);
  and _44698_ (_12551_, _12550_, _02157_);
  and _44699_ (_12552_, _12551_, _12540_);
  or _44700_ (_12553_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _44701_ (_12554_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _44702_ (_12555_, _12554_, _02150_);
  and _44703_ (_12556_, _12555_, _12553_);
  or _44704_ (_12557_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _44705_ (_12558_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _44706_ (_12559_, _12558_, _01954_);
  and _44707_ (_12560_, _12559_, _12557_);
  or _44708_ (_12561_, _12560_, _12556_);
  or _44709_ (_12562_, _12561_, _02144_);
  or _44710_ (_12563_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _44711_ (_12564_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _44712_ (_12565_, _12564_, _02150_);
  and _44713_ (_12566_, _12565_, _12563_);
  or _44714_ (_12567_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _44715_ (_12568_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _44716_ (_12569_, _12568_, _01954_);
  and _44717_ (_12570_, _12569_, _12567_);
  or _44718_ (_12571_, _12570_, _12566_);
  or _44719_ (_12572_, _12571_, _02131_);
  and _44720_ (_12573_, _12572_, _02077_);
  and _44721_ (_12574_, _12573_, _12562_);
  or _44722_ (_12575_, _12574_, _12552_);
  and _44723_ (_12576_, _12575_, _02194_);
  or _44724_ (_12577_, _12576_, _12530_);
  and _44725_ (_12578_, _12577_, _02143_);
  and _44726_ (_12579_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _44727_ (_12580_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _44728_ (_12581_, _12580_, _12579_);
  and _44729_ (_12582_, _12581_, _01954_);
  and _44730_ (_12583_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _44731_ (_12584_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _44732_ (_12585_, _12584_, _12583_);
  and _44733_ (_12586_, _12585_, _02150_);
  or _44734_ (_12587_, _12586_, _12582_);
  and _44735_ (_12588_, _12587_, _02131_);
  and _44736_ (_12589_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _44737_ (_12590_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _44738_ (_12591_, _12590_, _12589_);
  and _44739_ (_12592_, _12591_, _01954_);
  and _44740_ (_12593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _44741_ (_12594_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _44742_ (_12595_, _12594_, _12593_);
  and _44743_ (_12596_, _12595_, _02150_);
  or _44744_ (_12597_, _12596_, _12592_);
  and _44745_ (_12598_, _12597_, _02144_);
  or _44746_ (_12599_, _12598_, _12588_);
  and _44747_ (_12600_, _12599_, _02157_);
  or _44748_ (_12601_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _44749_ (_12602_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _44750_ (_12603_, _12602_, _02150_);
  and _44751_ (_12604_, _12603_, _12601_);
  or _44752_ (_12605_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _44753_ (_12606_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _44754_ (_12607_, _12606_, _01954_);
  and _44755_ (_12608_, _12607_, _12605_);
  or _44756_ (_12609_, _12608_, _12604_);
  and _44757_ (_12610_, _12609_, _02131_);
  or _44758_ (_12611_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _44759_ (_12612_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _44760_ (_12613_, _12612_, _02150_);
  and _44761_ (_12614_, _12613_, _12611_);
  or _44762_ (_12615_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _44763_ (_12616_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _44764_ (_12617_, _12616_, _01954_);
  and _44765_ (_12618_, _12617_, _12615_);
  or _44766_ (_12619_, _12618_, _12614_);
  and _44767_ (_12620_, _12619_, _02144_);
  or _44768_ (_12621_, _12620_, _12610_);
  and _44769_ (_12622_, _12621_, _02077_);
  or _44770_ (_12623_, _12622_, _12600_);
  and _44771_ (_12624_, _12623_, _02194_);
  and _44772_ (_12625_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _44773_ (_12626_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _44774_ (_12627_, _12626_, _12625_);
  and _44775_ (_12628_, _12627_, _01954_);
  and _44776_ (_12629_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _44777_ (_12630_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _44778_ (_12631_, _12630_, _12629_);
  and _44779_ (_12632_, _12631_, _02150_);
  or _44780_ (_12633_, _12632_, _12628_);
  and _44781_ (_12634_, _12633_, _02131_);
  and _44782_ (_12635_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _44783_ (_12636_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _44784_ (_12637_, _12636_, _12635_);
  and _44785_ (_12638_, _12637_, _01954_);
  and _44786_ (_12639_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _44787_ (_12640_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _44788_ (_12641_, _12640_, _12639_);
  and _44789_ (_12642_, _12641_, _02150_);
  or _44790_ (_12643_, _12642_, _12638_);
  and _44791_ (_12644_, _12643_, _02144_);
  or _44792_ (_12645_, _12644_, _12634_);
  and _44793_ (_12646_, _12645_, _02157_);
  or _44794_ (_12647_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _44795_ (_12648_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _44796_ (_12649_, _12648_, _12647_);
  and _44797_ (_12650_, _12649_, _01954_);
  or _44798_ (_12651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _44799_ (_12652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _44800_ (_12653_, _12652_, _12651_);
  and _44801_ (_12654_, _12653_, _02150_);
  or _44802_ (_12655_, _12654_, _12650_);
  and _44803_ (_12656_, _12655_, _02131_);
  or _44804_ (_12657_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _44805_ (_12658_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _44806_ (_12659_, _12658_, _12657_);
  and _44807_ (_12660_, _12659_, _01954_);
  or _44808_ (_12661_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _44809_ (_12662_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _44810_ (_12663_, _12662_, _12661_);
  and _44811_ (_12664_, _12663_, _02150_);
  or _44812_ (_12665_, _12664_, _12660_);
  and _44813_ (_12666_, _12665_, _02144_);
  or _44814_ (_12667_, _12666_, _12656_);
  and _44815_ (_12668_, _12667_, _02077_);
  or _44816_ (_12669_, _12668_, _12646_);
  and _44817_ (_12670_, _12669_, _02065_);
  or _44818_ (_12671_, _12670_, _12624_);
  and _44819_ (_12672_, _12671_, _02005_);
  or _44820_ (_12673_, _12672_, _12578_);
  or _44821_ (_12674_, _12673_, _02054_);
  and _44822_ (_12675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _44823_ (_12676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _44824_ (_12677_, _12676_, _12675_);
  and _44825_ (_12678_, _12677_, _01954_);
  and _44826_ (_12679_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _44827_ (_12680_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _44828_ (_12681_, _12680_, _12679_);
  and _44829_ (_12682_, _12681_, _02150_);
  or _44830_ (_12683_, _12682_, _12678_);
  or _44831_ (_12684_, _12683_, _02144_);
  and _44832_ (_12685_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _44833_ (_12686_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _44834_ (_12687_, _12686_, _12685_);
  and _44835_ (_12688_, _12687_, _01954_);
  and _44836_ (_12689_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _44837_ (_12690_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _44838_ (_12691_, _12690_, _12689_);
  and _44839_ (_12692_, _12691_, _02150_);
  or _44840_ (_12693_, _12692_, _12688_);
  or _44841_ (_12694_, _12693_, _02131_);
  and _44842_ (_12695_, _12694_, _02157_);
  and _44843_ (_12696_, _12695_, _12684_);
  or _44844_ (_12697_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _44845_ (_12698_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and _44846_ (_12699_, _12698_, _02150_);
  and _44847_ (_12700_, _12699_, _12697_);
  or _44848_ (_12701_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _44849_ (_12702_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and _44850_ (_12703_, _12702_, _01954_);
  and _44851_ (_12704_, _12703_, _12701_);
  or _44852_ (_12705_, _12704_, _12700_);
  or _44853_ (_12706_, _12705_, _02144_);
  or _44854_ (_12707_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _44855_ (_12708_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _44856_ (_12709_, _12708_, _02150_);
  and _44857_ (_12710_, _12709_, _12707_);
  or _44858_ (_12711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _44859_ (_12712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _44860_ (_12713_, _12712_, _01954_);
  and _44861_ (_12714_, _12713_, _12711_);
  or _44862_ (_12715_, _12714_, _12710_);
  or _44863_ (_12716_, _12715_, _02131_);
  and _44864_ (_12717_, _12716_, _02077_);
  and _44865_ (_12718_, _12717_, _12706_);
  or _44866_ (_12719_, _12718_, _12696_);
  and _44867_ (_12720_, _12719_, _02194_);
  and _44868_ (_12721_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _44869_ (_12722_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _44870_ (_12723_, _12722_, _12721_);
  and _44871_ (_12724_, _12723_, _01954_);
  and _44872_ (_12725_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _44873_ (_12726_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _44874_ (_12727_, _12726_, _12725_);
  and _44875_ (_12728_, _12727_, _02150_);
  or _44876_ (_12729_, _12728_, _12724_);
  or _44877_ (_12730_, _12729_, _02144_);
  and _44878_ (_12731_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _44879_ (_12732_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _44880_ (_12733_, _12732_, _12731_);
  and _44881_ (_12734_, _12733_, _01954_);
  and _44882_ (_12735_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _44883_ (_12736_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _44884_ (_12737_, _12736_, _12735_);
  and _44885_ (_12738_, _12737_, _02150_);
  or _44886_ (_12739_, _12738_, _12734_);
  or _44887_ (_12740_, _12739_, _02131_);
  and _44888_ (_12741_, _12740_, _02157_);
  and _44889_ (_12742_, _12741_, _12730_);
  or _44890_ (_12744_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _44891_ (_12745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _44892_ (_12746_, _12745_, _12744_);
  and _44893_ (_12747_, _12746_, _01954_);
  or _44894_ (_12748_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _44895_ (_12749_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _44896_ (_12750_, _12749_, _12748_);
  and _44897_ (_12751_, _12750_, _02150_);
  or _44898_ (_12752_, _12751_, _12747_);
  or _44899_ (_12753_, _12752_, _02144_);
  or _44900_ (_12754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _44901_ (_12755_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _44902_ (_12756_, _12755_, _12754_);
  and _44903_ (_12757_, _12756_, _01954_);
  or _44904_ (_12758_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _44905_ (_12759_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _44906_ (_12760_, _12759_, _12758_);
  and _44907_ (_12761_, _12760_, _02150_);
  or _44908_ (_12762_, _12761_, _12757_);
  or _44909_ (_12763_, _12762_, _02131_);
  and _44910_ (_12765_, _12763_, _02077_);
  and _44911_ (_12766_, _12765_, _12753_);
  or _44912_ (_12767_, _12766_, _12742_);
  and _44913_ (_12768_, _12767_, _02065_);
  or _44914_ (_12769_, _12768_, _12720_);
  and _44915_ (_12770_, _12769_, _02143_);
  or _44916_ (_12771_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _44917_ (_12772_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _44918_ (_12773_, _12772_, _12771_);
  and _44919_ (_12774_, _12773_, _01954_);
  or _44920_ (_12775_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _44921_ (_12776_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _44922_ (_12777_, _12776_, _12775_);
  and _44923_ (_12778_, _12777_, _02150_);
  or _44924_ (_12779_, _12778_, _12774_);
  and _44925_ (_12780_, _12779_, _02144_);
  or _44926_ (_12781_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _44927_ (_12782_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _44928_ (_12783_, _12782_, _12781_);
  and _44929_ (_12784_, _12783_, _01954_);
  or _44930_ (_12785_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _44931_ (_12786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _44932_ (_12787_, _12786_, _12785_);
  and _44933_ (_12788_, _12787_, _02150_);
  or _44934_ (_12789_, _12788_, _12784_);
  and _44935_ (_12790_, _12789_, _02131_);
  or _44936_ (_12791_, _12790_, _12780_);
  and _44937_ (_12792_, _12791_, _02077_);
  and _44938_ (_12793_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _44939_ (_12794_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _44940_ (_12795_, _12794_, _12793_);
  and _44941_ (_12796_, _12795_, _01954_);
  and _44942_ (_12797_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _44943_ (_12798_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _44944_ (_12799_, _12798_, _12797_);
  and _44945_ (_12800_, _12799_, _02150_);
  or _44946_ (_12801_, _12800_, _12796_);
  and _44947_ (_12802_, _12801_, _02144_);
  and _44948_ (_12803_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _44949_ (_12804_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _44950_ (_12805_, _12804_, _12803_);
  and _44951_ (_12806_, _12805_, _01954_);
  and _44952_ (_12807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _44953_ (_12808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _44954_ (_12809_, _12808_, _12807_);
  and _44955_ (_12810_, _12809_, _02150_);
  or _44956_ (_12811_, _12810_, _12806_);
  and _44957_ (_12812_, _12811_, _02131_);
  or _44958_ (_12813_, _12812_, _12802_);
  and _44959_ (_12814_, _12813_, _02157_);
  or _44960_ (_12815_, _12814_, _12792_);
  and _44961_ (_12816_, _12815_, _02065_);
  or _44962_ (_12817_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _44963_ (_12818_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _44964_ (_12819_, _12818_, _02150_);
  and _44965_ (_12820_, _12819_, _12817_);
  or _44966_ (_12821_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _44967_ (_12822_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _44968_ (_12823_, _12822_, _01954_);
  and _44969_ (_12824_, _12823_, _12821_);
  or _44970_ (_12825_, _12824_, _12820_);
  and _44971_ (_12826_, _12825_, _02144_);
  or _44972_ (_12827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _44973_ (_12828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _44974_ (_12829_, _12828_, _02150_);
  and _44975_ (_12830_, _12829_, _12827_);
  or _44976_ (_12831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _44977_ (_12832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _44978_ (_12833_, _12832_, _01954_);
  and _44979_ (_12834_, _12833_, _12831_);
  or _44980_ (_12835_, _12834_, _12830_);
  and _44981_ (_12836_, _12835_, _02131_);
  or _44982_ (_12837_, _12836_, _12826_);
  and _44983_ (_12838_, _12837_, _02077_);
  and _44984_ (_12839_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _44985_ (_12840_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _44986_ (_12841_, _12840_, _12839_);
  and _44987_ (_12842_, _12841_, _01954_);
  and _44988_ (_12843_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _44989_ (_12844_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _44990_ (_12845_, _12844_, _12843_);
  and _44991_ (_12846_, _12845_, _02150_);
  or _44992_ (_12847_, _12846_, _12842_);
  and _44993_ (_12848_, _12847_, _02144_);
  and _44994_ (_12849_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _44995_ (_12850_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _44996_ (_12851_, _12850_, _12849_);
  and _44997_ (_12852_, _12851_, _01954_);
  and _44998_ (_12853_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _44999_ (_12854_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _45000_ (_12855_, _12854_, _12853_);
  and _45001_ (_12856_, _12855_, _02150_);
  or _45002_ (_12857_, _12856_, _12852_);
  and _45003_ (_12858_, _12857_, _02131_);
  or _45004_ (_12859_, _12858_, _12848_);
  and _45005_ (_12860_, _12859_, _02157_);
  or _45006_ (_12861_, _12860_, _12838_);
  and _45007_ (_12862_, _12861_, _02194_);
  or _45008_ (_12863_, _12862_, _12816_);
  and _45009_ (_12864_, _12863_, _02005_);
  or _45010_ (_12865_, _12864_, _12770_);
  or _45011_ (_12866_, _12865_, _02374_);
  and _45012_ (_12867_, _12866_, _12674_);
  or _45013_ (_12868_, _12867_, _01748_);
  and _45014_ (_12869_, _12868_, _12484_);
  or _45015_ (_12870_, _12869_, _02141_);
  or _45016_ (_12871_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _45017_ (_12872_, _12871_, _27355_);
  and _45018_ (_15242_, _12872_, _12870_);
  and _45019_ (_12873_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _45020_ (_12874_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _45021_ (_12875_, _12874_, _12873_);
  and _45022_ (_12876_, _12875_, _01954_);
  and _45023_ (_12877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _45024_ (_12878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _45025_ (_12879_, _12878_, _12877_);
  and _45026_ (_12880_, _12879_, _02150_);
  or _45027_ (_12881_, _12880_, _12876_);
  or _45028_ (_12882_, _12881_, _02144_);
  and _45029_ (_12883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _45030_ (_12884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _45031_ (_12885_, _12884_, _12883_);
  and _45032_ (_12886_, _12885_, _01954_);
  and _45033_ (_12887_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and _45034_ (_12888_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _45035_ (_12889_, _12888_, _12887_);
  and _45036_ (_12890_, _12889_, _02150_);
  or _45037_ (_12891_, _12890_, _12886_);
  or _45038_ (_12892_, _12891_, _02131_);
  and _45039_ (_12893_, _12892_, _02157_);
  and _45040_ (_12894_, _12893_, _12882_);
  or _45041_ (_12895_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _45042_ (_12896_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _45043_ (_12897_, _12896_, _12895_);
  and _45044_ (_12898_, _12897_, _01954_);
  or _45045_ (_12899_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _45046_ (_12900_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and _45047_ (_12901_, _12900_, _12899_);
  and _45048_ (_12902_, _12901_, _02150_);
  or _45049_ (_12903_, _12902_, _12898_);
  or _45050_ (_12904_, _12903_, _02144_);
  or _45051_ (_12905_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _45052_ (_12906_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _45053_ (_12907_, _12906_, _12905_);
  and _45054_ (_12908_, _12907_, _01954_);
  or _45055_ (_12909_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _45056_ (_12910_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _45057_ (_12911_, _12910_, _12909_);
  and _45058_ (_12912_, _12911_, _02150_);
  or _45059_ (_12913_, _12912_, _12908_);
  or _45060_ (_12914_, _12913_, _02131_);
  and _45061_ (_12915_, _12914_, _02077_);
  and _45062_ (_12916_, _12915_, _12904_);
  or _45063_ (_12917_, _12916_, _12894_);
  and _45064_ (_12918_, _12917_, _02065_);
  and _45065_ (_12919_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _45066_ (_12920_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _45067_ (_12921_, _12920_, _12919_);
  and _45068_ (_12922_, _12921_, _01954_);
  and _45069_ (_12923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and _45070_ (_12924_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _45071_ (_12925_, _12924_, _12923_);
  and _45072_ (_12926_, _12925_, _02150_);
  or _45073_ (_12927_, _12926_, _12922_);
  or _45074_ (_12928_, _12927_, _02144_);
  and _45075_ (_12929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _45076_ (_12930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _45077_ (_12931_, _12930_, _12929_);
  and _45078_ (_12932_, _12931_, _01954_);
  and _45079_ (_12933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _45080_ (_12934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _45081_ (_12935_, _12934_, _12933_);
  and _45082_ (_12936_, _12935_, _02150_);
  or _45083_ (_12937_, _12936_, _12932_);
  or _45084_ (_12938_, _12937_, _02131_);
  and _45085_ (_12939_, _12938_, _02157_);
  and _45086_ (_12940_, _12939_, _12928_);
  or _45087_ (_12941_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _45088_ (_12942_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _45089_ (_12943_, _12942_, _02150_);
  and _45090_ (_12944_, _12943_, _12941_);
  or _45091_ (_12945_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _45092_ (_12946_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _45093_ (_12947_, _12946_, _01954_);
  and _45094_ (_12948_, _12947_, _12945_);
  or _45095_ (_12949_, _12948_, _12944_);
  or _45096_ (_12950_, _12949_, _02144_);
  or _45097_ (_12951_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _45098_ (_12952_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _45099_ (_12953_, _12952_, _02150_);
  and _45100_ (_12954_, _12953_, _12951_);
  or _45101_ (_12955_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _45102_ (_12956_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and _45103_ (_12957_, _12956_, _01954_);
  and _45104_ (_12958_, _12957_, _12955_);
  or _45105_ (_12959_, _12958_, _12954_);
  or _45106_ (_12960_, _12959_, _02131_);
  and _45107_ (_12961_, _12960_, _02077_);
  and _45108_ (_12962_, _12961_, _12950_);
  or _45109_ (_12963_, _12962_, _12940_);
  and _45110_ (_12964_, _12963_, _02194_);
  or _45111_ (_12965_, _12964_, _12918_);
  and _45112_ (_12966_, _12965_, _02143_);
  and _45113_ (_12967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _45114_ (_12968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _45115_ (_12969_, _12968_, _12967_);
  and _45116_ (_12970_, _12969_, _01954_);
  and _45117_ (_12971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _45118_ (_12972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _45119_ (_12973_, _12972_, _12971_);
  and _45120_ (_12974_, _12973_, _02150_);
  or _45121_ (_12975_, _12974_, _12970_);
  and _45122_ (_12976_, _12975_, _02131_);
  and _45123_ (_12977_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _45124_ (_12978_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _45125_ (_12979_, _12978_, _12977_);
  and _45126_ (_12980_, _12979_, _01954_);
  and _45127_ (_12981_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _45128_ (_12982_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _45129_ (_12983_, _12982_, _12981_);
  and _45130_ (_12984_, _12983_, _02150_);
  or _45131_ (_12985_, _12984_, _12980_);
  and _45132_ (_12986_, _12985_, _02144_);
  or _45133_ (_12987_, _12986_, _12976_);
  and _45134_ (_12988_, _12987_, _02157_);
  or _45135_ (_12989_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _45136_ (_12990_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _45137_ (_12991_, _12990_, _02150_);
  and _45138_ (_12992_, _12991_, _12989_);
  or _45139_ (_12993_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _45140_ (_12994_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _45141_ (_12995_, _12994_, _01954_);
  and _45142_ (_12996_, _12995_, _12993_);
  or _45143_ (_12997_, _12996_, _12992_);
  and _45144_ (_12998_, _12997_, _02131_);
  or _45145_ (_12999_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _45146_ (_13000_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _45147_ (_13001_, _13000_, _02150_);
  and _45148_ (_13002_, _13001_, _12999_);
  or _45149_ (_13003_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _45150_ (_13004_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _45151_ (_13005_, _13004_, _01954_);
  and _45152_ (_13006_, _13005_, _13003_);
  or _45153_ (_13007_, _13006_, _13002_);
  and _45154_ (_13008_, _13007_, _02144_);
  or _45155_ (_13009_, _13008_, _12998_);
  and _45156_ (_13010_, _13009_, _02077_);
  or _45157_ (_13011_, _13010_, _12988_);
  and _45158_ (_13012_, _13011_, _02194_);
  and _45159_ (_13013_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _45160_ (_13014_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _45161_ (_13015_, _13014_, _13013_);
  and _45162_ (_13016_, _13015_, _01954_);
  and _45163_ (_13017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _45164_ (_13018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _45165_ (_13019_, _13018_, _13017_);
  and _45166_ (_13020_, _13019_, _02150_);
  or _45167_ (_13021_, _13020_, _13016_);
  and _45168_ (_13022_, _13021_, _02131_);
  and _45169_ (_13023_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _45170_ (_13024_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _45171_ (_13025_, _13024_, _13023_);
  and _45172_ (_13026_, _13025_, _01954_);
  and _45173_ (_13027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _45174_ (_13028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _45175_ (_13029_, _13028_, _13027_);
  and _45176_ (_13030_, _13029_, _02150_);
  or _45177_ (_13031_, _13030_, _13026_);
  and _45178_ (_13032_, _13031_, _02144_);
  or _45179_ (_13033_, _13032_, _13022_);
  and _45180_ (_13034_, _13033_, _02157_);
  or _45181_ (_13035_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _45182_ (_13036_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _45183_ (_13037_, _13036_, _13035_);
  and _45184_ (_13038_, _13037_, _01954_);
  or _45185_ (_13039_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _45186_ (_13040_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _45187_ (_13041_, _13040_, _13039_);
  and _45188_ (_13042_, _13041_, _02150_);
  or _45189_ (_13043_, _13042_, _13038_);
  and _45190_ (_13044_, _13043_, _02131_);
  or _45191_ (_13045_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _45192_ (_13046_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _45193_ (_13047_, _13046_, _13045_);
  and _45194_ (_13048_, _13047_, _01954_);
  or _45195_ (_13049_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _45196_ (_13050_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _45197_ (_13051_, _13050_, _13049_);
  and _45198_ (_13052_, _13051_, _02150_);
  or _45199_ (_13053_, _13052_, _13048_);
  and _45200_ (_13054_, _13053_, _02144_);
  or _45201_ (_13055_, _13054_, _13044_);
  and _45202_ (_13056_, _13055_, _02077_);
  or _45203_ (_13057_, _13056_, _13034_);
  and _45204_ (_13058_, _13057_, _02065_);
  or _45205_ (_13059_, _13058_, _13012_);
  and _45206_ (_13060_, _13059_, _02005_);
  or _45207_ (_13061_, _13060_, _12966_);
  or _45208_ (_13062_, _13061_, _02054_);
  and _45209_ (_13063_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and _45210_ (_13064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _45211_ (_13065_, _13064_, _13063_);
  and _45212_ (_13066_, _13065_, _01954_);
  and _45213_ (_13067_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _45214_ (_13068_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _45215_ (_13069_, _13068_, _13067_);
  and _45216_ (_13070_, _13069_, _02150_);
  or _45217_ (_13071_, _13070_, _13066_);
  or _45218_ (_13072_, _13071_, _02144_);
  and _45219_ (_13073_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _45220_ (_13074_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _45221_ (_13075_, _13074_, _13073_);
  and _45222_ (_13076_, _13075_, _01954_);
  and _45223_ (_13077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _45224_ (_13078_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _45225_ (_13079_, _13078_, _13077_);
  and _45226_ (_13080_, _13079_, _02150_);
  or _45227_ (_13081_, _13080_, _13076_);
  or _45228_ (_13082_, _13081_, _02131_);
  and _45229_ (_13083_, _13082_, _02157_);
  and _45230_ (_13084_, _13083_, _13072_);
  or _45231_ (_13085_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _45232_ (_13086_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _45233_ (_13087_, _13086_, _02150_);
  and _45234_ (_13088_, _13087_, _13085_);
  or _45235_ (_13089_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _45236_ (_13090_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _45237_ (_13091_, _13090_, _01954_);
  and _45238_ (_13092_, _13091_, _13089_);
  or _45239_ (_13093_, _13092_, _13088_);
  or _45240_ (_13094_, _13093_, _02144_);
  or _45241_ (_13095_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _45242_ (_13096_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _45243_ (_13097_, _13096_, _02150_);
  and _45244_ (_13098_, _13097_, _13095_);
  or _45245_ (_13099_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _45246_ (_13100_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and _45247_ (_13101_, _13100_, _01954_);
  and _45248_ (_13102_, _13101_, _13099_);
  or _45249_ (_13103_, _13102_, _13098_);
  or _45250_ (_13104_, _13103_, _02131_);
  and _45251_ (_13105_, _13104_, _02077_);
  and _45252_ (_13106_, _13105_, _13094_);
  or _45253_ (_13107_, _13106_, _13084_);
  and _45254_ (_13108_, _13107_, _02194_);
  and _45255_ (_13109_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _45256_ (_13110_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _45257_ (_13111_, _13110_, _13109_);
  and _45258_ (_13112_, _13111_, _01954_);
  and _45259_ (_13113_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _45260_ (_13114_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _45261_ (_13115_, _13114_, _13113_);
  and _45262_ (_13116_, _13115_, _02150_);
  or _45263_ (_13117_, _13116_, _13112_);
  or _45264_ (_13118_, _13117_, _02144_);
  and _45265_ (_13119_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _45266_ (_13120_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _45267_ (_13121_, _13120_, _13119_);
  and _45268_ (_13122_, _13121_, _01954_);
  and _45269_ (_13123_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _45270_ (_13124_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _45271_ (_13125_, _13124_, _13123_);
  and _45272_ (_13126_, _13125_, _02150_);
  or _45273_ (_13127_, _13126_, _13122_);
  or _45274_ (_13128_, _13127_, _02131_);
  and _45275_ (_13129_, _13128_, _02157_);
  and _45276_ (_13130_, _13129_, _13118_);
  or _45277_ (_13131_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _45278_ (_13132_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _45279_ (_13133_, _13132_, _13131_);
  and _45280_ (_13134_, _13133_, _01954_);
  or _45281_ (_13135_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _45282_ (_13136_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _45283_ (_13137_, _13136_, _13135_);
  and _45284_ (_13138_, _13137_, _02150_);
  or _45285_ (_13139_, _13138_, _13134_);
  or _45286_ (_13140_, _13139_, _02144_);
  or _45287_ (_13141_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _45288_ (_13142_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _45289_ (_13143_, _13142_, _13141_);
  and _45290_ (_13144_, _13143_, _01954_);
  or _45291_ (_13145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _45292_ (_13146_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _45293_ (_13147_, _13146_, _13145_);
  and _45294_ (_13148_, _13147_, _02150_);
  or _45295_ (_13149_, _13148_, _13144_);
  or _45296_ (_13150_, _13149_, _02131_);
  and _45297_ (_13151_, _13150_, _02077_);
  and _45298_ (_13152_, _13151_, _13140_);
  or _45299_ (_13153_, _13152_, _13130_);
  and _45300_ (_13154_, _13153_, _02065_);
  or _45301_ (_13155_, _13154_, _13108_);
  and _45302_ (_13156_, _13155_, _02143_);
  or _45303_ (_13157_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _45304_ (_13158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and _45305_ (_13159_, _13158_, _13157_);
  and _45306_ (_13160_, _13159_, _01954_);
  or _45307_ (_13161_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _45308_ (_13162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _45309_ (_13163_, _13162_, _13161_);
  and _45310_ (_13164_, _13163_, _02150_);
  or _45311_ (_13165_, _13164_, _13160_);
  and _45312_ (_13166_, _13165_, _02144_);
  or _45313_ (_13167_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _45314_ (_13168_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _45315_ (_13169_, _13168_, _13167_);
  and _45316_ (_13170_, _13169_, _01954_);
  or _45317_ (_13171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _45318_ (_13172_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and _45319_ (_13173_, _13172_, _13171_);
  and _45320_ (_13174_, _13173_, _02150_);
  or _45321_ (_13175_, _13174_, _13170_);
  and _45322_ (_13176_, _13175_, _02131_);
  or _45323_ (_13177_, _13176_, _13166_);
  and _45324_ (_13178_, _13177_, _02077_);
  and _45325_ (_13179_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _45326_ (_13180_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _45327_ (_13181_, _13180_, _13179_);
  and _45328_ (_13182_, _13181_, _01954_);
  and _45329_ (_13183_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _45330_ (_13184_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _45331_ (_13185_, _13184_, _13183_);
  and _45332_ (_13186_, _13185_, _02150_);
  or _45333_ (_13187_, _13186_, _13182_);
  and _45334_ (_13188_, _13187_, _02144_);
  and _45335_ (_13189_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _45336_ (_13190_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _45337_ (_13191_, _13190_, _13189_);
  and _45338_ (_13192_, _13191_, _01954_);
  and _45339_ (_13193_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _45340_ (_13194_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _45341_ (_13195_, _13194_, _13193_);
  and _45342_ (_13196_, _13195_, _02150_);
  or _45343_ (_13197_, _13196_, _13192_);
  and _45344_ (_13198_, _13197_, _02131_);
  or _45345_ (_13199_, _13198_, _13188_);
  and _45346_ (_13200_, _13199_, _02157_);
  or _45347_ (_13201_, _13200_, _13178_);
  and _45348_ (_13202_, _13201_, _02065_);
  or _45349_ (_13203_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _45350_ (_13204_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _45351_ (_13205_, _13204_, _02150_);
  and _45352_ (_13206_, _13205_, _13203_);
  or _45353_ (_13207_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _45354_ (_13208_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _45355_ (_13209_, _13208_, _01954_);
  and _45356_ (_13210_, _13209_, _13207_);
  or _45357_ (_13211_, _13210_, _13206_);
  and _45358_ (_13212_, _13211_, _02144_);
  or _45359_ (_13213_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _45360_ (_13214_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _45361_ (_13215_, _13214_, _02150_);
  and _45362_ (_13216_, _13215_, _13213_);
  or _45363_ (_13217_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _45364_ (_13218_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and _45365_ (_13219_, _13218_, _01954_);
  and _45366_ (_13220_, _13219_, _13217_);
  or _45367_ (_13221_, _13220_, _13216_);
  and _45368_ (_13222_, _13221_, _02131_);
  or _45369_ (_13223_, _13222_, _13212_);
  and _45370_ (_13224_, _13223_, _02077_);
  and _45371_ (_13225_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _45372_ (_13226_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _45373_ (_13227_, _13226_, _13225_);
  and _45374_ (_13228_, _13227_, _01954_);
  and _45375_ (_13229_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _45376_ (_13230_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _45377_ (_13231_, _13230_, _13229_);
  and _45378_ (_13232_, _13231_, _02150_);
  or _45379_ (_13233_, _13232_, _13228_);
  and _45380_ (_13234_, _13233_, _02144_);
  and _45381_ (_13235_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _45382_ (_13236_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _45383_ (_13237_, _13236_, _13235_);
  and _45384_ (_13238_, _13237_, _01954_);
  and _45385_ (_13239_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _45386_ (_13240_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _45387_ (_13241_, _13240_, _13239_);
  and _45388_ (_13242_, _13241_, _02150_);
  or _45389_ (_13243_, _13242_, _13238_);
  and _45390_ (_13244_, _13243_, _02131_);
  or _45391_ (_13245_, _13244_, _13234_);
  and _45392_ (_13246_, _13245_, _02157_);
  or _45393_ (_13247_, _13246_, _13224_);
  and _45394_ (_13248_, _13247_, _02194_);
  or _45395_ (_13249_, _13248_, _13202_);
  and _45396_ (_13250_, _13249_, _02005_);
  or _45397_ (_13251_, _13250_, _13156_);
  or _45398_ (_13252_, _13251_, _02374_);
  and _45399_ (_13253_, _13252_, _13062_);
  or _45400_ (_13254_, _13253_, _02142_);
  and _45401_ (_13255_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _45402_ (_13256_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _45403_ (_13257_, _13256_, _13255_);
  and _45404_ (_13258_, _13257_, _01954_);
  and _45405_ (_13259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _45406_ (_13260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _45407_ (_13261_, _13260_, _13259_);
  and _45408_ (_13262_, _13261_, _02150_);
  or _45409_ (_13263_, _13262_, _13258_);
  or _45410_ (_13264_, _13263_, _02144_);
  and _45411_ (_13265_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _45412_ (_13266_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _45413_ (_13267_, _13266_, _13265_);
  and _45414_ (_13268_, _13267_, _01954_);
  and _45415_ (_13269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _45416_ (_13270_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _45417_ (_13271_, _13270_, _13269_);
  and _45418_ (_13272_, _13271_, _02150_);
  or _45419_ (_13273_, _13272_, _13268_);
  or _45420_ (_13274_, _13273_, _02131_);
  and _45421_ (_13275_, _13274_, _02157_);
  and _45422_ (_13276_, _13275_, _13264_);
  or _45423_ (_13277_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _45424_ (_13278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _45425_ (_13279_, _13278_, _13277_);
  and _45426_ (_13280_, _13279_, _01954_);
  or _45427_ (_13281_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _45428_ (_13282_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and _45429_ (_13283_, _13282_, _13281_);
  and _45430_ (_13284_, _13283_, _02150_);
  or _45431_ (_13285_, _13284_, _13280_);
  or _45432_ (_13286_, _13285_, _02144_);
  or _45433_ (_13287_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _45434_ (_13288_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and _45435_ (_13289_, _13288_, _13287_);
  and _45436_ (_13290_, _13289_, _01954_);
  or _45437_ (_13291_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _45438_ (_13292_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _45439_ (_13293_, _13292_, _13291_);
  and _45440_ (_13294_, _13293_, _02150_);
  or _45441_ (_13295_, _13294_, _13290_);
  or _45442_ (_13296_, _13295_, _02131_);
  and _45443_ (_13297_, _13296_, _02077_);
  and _45444_ (_13298_, _13297_, _13286_);
  or _45445_ (_13299_, _13298_, _13276_);
  and _45446_ (_13300_, _13299_, _02065_);
  and _45447_ (_13301_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _45448_ (_13302_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _45449_ (_13303_, _13302_, _13301_);
  and _45450_ (_13304_, _13303_, _01954_);
  and _45451_ (_13305_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _45452_ (_13306_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _45453_ (_13307_, _13306_, _13305_);
  and _45454_ (_13308_, _13307_, _02150_);
  or _45455_ (_13309_, _13308_, _13304_);
  or _45456_ (_13310_, _13309_, _02144_);
  and _45457_ (_13311_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _45458_ (_13312_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _45459_ (_13313_, _13312_, _13311_);
  and _45460_ (_13314_, _13313_, _01954_);
  and _45461_ (_13315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _45462_ (_13316_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _45463_ (_13317_, _13316_, _13315_);
  and _45464_ (_13318_, _13317_, _02150_);
  or _45465_ (_13319_, _13318_, _13314_);
  or _45466_ (_13320_, _13319_, _02131_);
  and _45467_ (_13321_, _13320_, _02157_);
  and _45468_ (_13322_, _13321_, _13310_);
  or _45469_ (_13323_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _45470_ (_13324_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _45471_ (_13325_, _13324_, _02150_);
  and _45472_ (_13326_, _13325_, _13323_);
  or _45473_ (_13327_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _45474_ (_13328_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _45475_ (_13329_, _13328_, _01954_);
  and _45476_ (_13330_, _13329_, _13327_);
  or _45477_ (_13331_, _13330_, _13326_);
  or _45478_ (_13332_, _13331_, _02144_);
  or _45479_ (_13333_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _45480_ (_13334_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _45481_ (_13335_, _13334_, _02150_);
  and _45482_ (_13336_, _13335_, _13333_);
  or _45483_ (_13337_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _45484_ (_13338_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _45485_ (_13339_, _13338_, _01954_);
  and _45486_ (_13340_, _13339_, _13337_);
  or _45487_ (_13341_, _13340_, _13336_);
  or _45488_ (_13342_, _13341_, _02131_);
  and _45489_ (_13343_, _13342_, _02077_);
  and _45490_ (_13344_, _13343_, _13332_);
  or _45491_ (_13345_, _13344_, _13322_);
  and _45492_ (_13346_, _13345_, _02194_);
  or _45493_ (_13347_, _13346_, _13300_);
  and _45494_ (_13348_, _13347_, _02143_);
  and _45495_ (_13349_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _45496_ (_13350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _45497_ (_13351_, _13350_, _13349_);
  and _45498_ (_13352_, _13351_, _01954_);
  and _45499_ (_13353_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _45500_ (_13354_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _45501_ (_13355_, _13354_, _13353_);
  and _45502_ (_13356_, _13355_, _02150_);
  or _45503_ (_13357_, _13356_, _13352_);
  and _45504_ (_13358_, _13357_, _02131_);
  and _45505_ (_13359_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _45506_ (_13360_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _45507_ (_13361_, _13360_, _13359_);
  and _45508_ (_13362_, _13361_, _01954_);
  and _45509_ (_13363_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _45510_ (_13364_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _45511_ (_13365_, _13364_, _13363_);
  and _45512_ (_13366_, _13365_, _02150_);
  or _45513_ (_13367_, _13366_, _13362_);
  and _45514_ (_13368_, _13367_, _02144_);
  or _45515_ (_13369_, _13368_, _13358_);
  and _45516_ (_13370_, _13369_, _02157_);
  or _45517_ (_13371_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _45518_ (_13372_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _45519_ (_13373_, _13372_, _02150_);
  and _45520_ (_13374_, _13373_, _13371_);
  or _45521_ (_13375_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _45522_ (_13376_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _45523_ (_13377_, _13376_, _01954_);
  and _45524_ (_13378_, _13377_, _13375_);
  or _45525_ (_13379_, _13378_, _13374_);
  and _45526_ (_13380_, _13379_, _02131_);
  or _45527_ (_13381_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _45528_ (_13382_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _45529_ (_13383_, _13382_, _02150_);
  and _45530_ (_13384_, _13383_, _13381_);
  or _45531_ (_13385_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _45532_ (_13386_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _45533_ (_13387_, _13386_, _01954_);
  and _45534_ (_13388_, _13387_, _13385_);
  or _45535_ (_13389_, _13388_, _13384_);
  and _45536_ (_13390_, _13389_, _02144_);
  or _45537_ (_13391_, _13390_, _13380_);
  and _45538_ (_13392_, _13391_, _02077_);
  or _45539_ (_13393_, _13392_, _13370_);
  and _45540_ (_13394_, _13393_, _02194_);
  and _45541_ (_13395_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _45542_ (_13396_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _45543_ (_13397_, _13396_, _13395_);
  and _45544_ (_13398_, _13397_, _01954_);
  and _45545_ (_13399_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _45546_ (_13400_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _45547_ (_13401_, _13400_, _13399_);
  and _45548_ (_13402_, _13401_, _02150_);
  or _45549_ (_13403_, _13402_, _13398_);
  and _45550_ (_13404_, _13403_, _02131_);
  and _45551_ (_13405_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _45552_ (_13406_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _45553_ (_13407_, _13406_, _13405_);
  and _45554_ (_13408_, _13407_, _01954_);
  and _45555_ (_13409_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _45556_ (_13410_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _45557_ (_13411_, _13410_, _13409_);
  and _45558_ (_13412_, _13411_, _02150_);
  or _45559_ (_13413_, _13412_, _13408_);
  and _45560_ (_13414_, _13413_, _02144_);
  or _45561_ (_13415_, _13414_, _13404_);
  and _45562_ (_13416_, _13415_, _02157_);
  or _45563_ (_13417_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _45564_ (_13418_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _45565_ (_13419_, _13418_, _13417_);
  and _45566_ (_13420_, _13419_, _01954_);
  or _45567_ (_13421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _45568_ (_13422_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _45569_ (_13423_, _13422_, _13421_);
  and _45570_ (_13424_, _13423_, _02150_);
  or _45571_ (_13425_, _13424_, _13420_);
  and _45572_ (_13426_, _13425_, _02131_);
  or _45573_ (_13427_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _45574_ (_13428_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _45575_ (_13429_, _13428_, _13427_);
  and _45576_ (_13430_, _13429_, _01954_);
  or _45577_ (_13431_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _45578_ (_13432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _45579_ (_13433_, _13432_, _13431_);
  and _45580_ (_13434_, _13433_, _02150_);
  or _45581_ (_13435_, _13434_, _13430_);
  and _45582_ (_13436_, _13435_, _02144_);
  or _45583_ (_13437_, _13436_, _13426_);
  and _45584_ (_13438_, _13437_, _02077_);
  or _45585_ (_13439_, _13438_, _13416_);
  and _45586_ (_13440_, _13439_, _02065_);
  or _45587_ (_13441_, _13440_, _13394_);
  and _45588_ (_13442_, _13441_, _02005_);
  or _45589_ (_13443_, _13442_, _13348_);
  or _45590_ (_13444_, _13443_, _02054_);
  and _45591_ (_13445_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _45592_ (_13446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _45593_ (_13447_, _13446_, _13445_);
  and _45594_ (_13448_, _13447_, _01954_);
  and _45595_ (_13449_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and _45596_ (_13450_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _45597_ (_13451_, _13450_, _13449_);
  and _45598_ (_13452_, _13451_, _02150_);
  or _45599_ (_13453_, _13452_, _13448_);
  or _45600_ (_13454_, _13453_, _02144_);
  and _45601_ (_13455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _45602_ (_13456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _45603_ (_13457_, _13456_, _13455_);
  and _45604_ (_13458_, _13457_, _01954_);
  and _45605_ (_13459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and _45606_ (_13460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _45607_ (_13461_, _13460_, _13459_);
  and _45608_ (_13462_, _13461_, _02150_);
  or _45609_ (_13463_, _13462_, _13458_);
  or _45610_ (_13464_, _13463_, _02131_);
  and _45611_ (_13465_, _13464_, _02157_);
  and _45612_ (_13466_, _13465_, _13454_);
  or _45613_ (_13467_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _45614_ (_13468_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _45615_ (_13469_, _13468_, _02150_);
  and _45616_ (_13470_, _13469_, _13467_);
  or _45617_ (_13471_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _45618_ (_13472_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _45619_ (_13473_, _13472_, _01954_);
  and _45620_ (_13474_, _13473_, _13471_);
  or _45621_ (_13475_, _13474_, _13470_);
  or _45622_ (_13476_, _13475_, _02144_);
  or _45623_ (_13477_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _45624_ (_13478_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and _45625_ (_13479_, _13478_, _02150_);
  and _45626_ (_13480_, _13479_, _13477_);
  or _45627_ (_13481_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _45628_ (_13482_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _45629_ (_13483_, _13482_, _01954_);
  and _45630_ (_13484_, _13483_, _13481_);
  or _45631_ (_13485_, _13484_, _13480_);
  or _45632_ (_13486_, _13485_, _02131_);
  and _45633_ (_13487_, _13486_, _02077_);
  and _45634_ (_13488_, _13487_, _13476_);
  or _45635_ (_13489_, _13488_, _13466_);
  and _45636_ (_13490_, _13489_, _02194_);
  and _45637_ (_13491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _45638_ (_13492_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _45639_ (_13493_, _13492_, _13491_);
  and _45640_ (_13494_, _13493_, _01954_);
  and _45641_ (_13495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _45642_ (_13496_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _45643_ (_13497_, _13496_, _13495_);
  and _45644_ (_13498_, _13497_, _02150_);
  or _45645_ (_13499_, _13498_, _13494_);
  or _45646_ (_13500_, _13499_, _02144_);
  and _45647_ (_13501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _45648_ (_13502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _45649_ (_13503_, _13502_, _13501_);
  and _45650_ (_13504_, _13503_, _01954_);
  and _45651_ (_13505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _45652_ (_13506_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _45653_ (_13507_, _13506_, _13505_);
  and _45654_ (_13508_, _13507_, _02150_);
  or _45655_ (_13509_, _13508_, _13504_);
  or _45656_ (_13510_, _13509_, _02131_);
  and _45657_ (_13511_, _13510_, _02157_);
  and _45658_ (_13512_, _13511_, _13500_);
  or _45659_ (_13513_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _45660_ (_13514_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _45661_ (_13515_, _13514_, _13513_);
  and _45662_ (_13516_, _13515_, _01954_);
  or _45663_ (_13517_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _45664_ (_13518_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _45665_ (_13519_, _13518_, _13517_);
  and _45666_ (_13520_, _13519_, _02150_);
  or _45667_ (_13521_, _13520_, _13516_);
  or _45668_ (_13522_, _13521_, _02144_);
  or _45669_ (_13523_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _45670_ (_13524_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _45671_ (_13525_, _13524_, _13523_);
  and _45672_ (_13526_, _13525_, _01954_);
  or _45673_ (_13527_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _45674_ (_13528_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _45675_ (_13529_, _13528_, _13527_);
  and _45676_ (_13530_, _13529_, _02150_);
  or _45677_ (_13531_, _13530_, _13526_);
  or _45678_ (_13532_, _13531_, _02131_);
  and _45679_ (_13533_, _13532_, _02077_);
  and _45680_ (_13534_, _13533_, _13522_);
  or _45681_ (_13535_, _13534_, _13512_);
  and _45682_ (_13536_, _13535_, _02065_);
  or _45683_ (_13537_, _13536_, _13490_);
  and _45684_ (_13538_, _13537_, _02143_);
  or _45685_ (_13539_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _45686_ (_13540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _45687_ (_13541_, _13540_, _13539_);
  and _45688_ (_13542_, _13541_, _01954_);
  or _45689_ (_13543_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _45690_ (_13544_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _45691_ (_13545_, _13544_, _13543_);
  and _45692_ (_13546_, _13545_, _02150_);
  or _45693_ (_13547_, _13546_, _13542_);
  and _45694_ (_13548_, _13547_, _02144_);
  or _45695_ (_13549_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _45696_ (_13550_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _45697_ (_13551_, _13550_, _13549_);
  and _45698_ (_13552_, _13551_, _01954_);
  or _45699_ (_13553_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _45700_ (_13554_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _45701_ (_13555_, _13554_, _13553_);
  and _45702_ (_13556_, _13555_, _02150_);
  or _45703_ (_13557_, _13556_, _13552_);
  and _45704_ (_13558_, _13557_, _02131_);
  or _45705_ (_13559_, _13558_, _13548_);
  and _45706_ (_13560_, _13559_, _02077_);
  and _45707_ (_13561_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _45708_ (_13562_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _45709_ (_13563_, _13562_, _13561_);
  and _45710_ (_13564_, _13563_, _01954_);
  and _45711_ (_13565_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _45712_ (_13566_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _45713_ (_13567_, _13566_, _13565_);
  and _45714_ (_13568_, _13567_, _02150_);
  or _45715_ (_13569_, _13568_, _13564_);
  and _45716_ (_13570_, _13569_, _02144_);
  and _45717_ (_13571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _45718_ (_13572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _45719_ (_13573_, _13572_, _13571_);
  and _45720_ (_13574_, _13573_, _01954_);
  and _45721_ (_13575_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _45722_ (_13576_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _45723_ (_13577_, _13576_, _13575_);
  and _45724_ (_13578_, _13577_, _02150_);
  or _45725_ (_13579_, _13578_, _13574_);
  and _45726_ (_13580_, _13579_, _02131_);
  or _45727_ (_13581_, _13580_, _13570_);
  and _45728_ (_13582_, _13581_, _02157_);
  or _45729_ (_13583_, _13582_, _13560_);
  and _45730_ (_13584_, _13583_, _02065_);
  or _45731_ (_13585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _45732_ (_13586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _45733_ (_13587_, _13586_, _02150_);
  and _45734_ (_13588_, _13587_, _13585_);
  or _45735_ (_13589_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _45736_ (_13590_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _45737_ (_13591_, _13590_, _01954_);
  and _45738_ (_13592_, _13591_, _13589_);
  or _45739_ (_13593_, _13592_, _13588_);
  and _45740_ (_13594_, _13593_, _02144_);
  or _45741_ (_13595_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _45742_ (_13596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _45743_ (_13597_, _13596_, _02150_);
  and _45744_ (_13598_, _13597_, _13595_);
  or _45745_ (_13599_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _45746_ (_13600_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _45747_ (_13601_, _13600_, _01954_);
  and _45748_ (_13602_, _13601_, _13599_);
  or _45749_ (_13603_, _13602_, _13598_);
  and _45750_ (_13604_, _13603_, _02131_);
  or _45751_ (_13605_, _13604_, _13594_);
  and _45752_ (_13606_, _13605_, _02077_);
  and _45753_ (_13607_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _45754_ (_13608_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _45755_ (_13609_, _13608_, _13607_);
  and _45756_ (_13610_, _13609_, _01954_);
  and _45757_ (_13611_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _45758_ (_13612_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _45759_ (_13613_, _13612_, _13611_);
  and _45760_ (_13614_, _13613_, _02150_);
  or _45761_ (_13615_, _13614_, _13610_);
  and _45762_ (_13616_, _13615_, _02144_);
  and _45763_ (_13617_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _45764_ (_13618_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _45765_ (_13619_, _13618_, _13617_);
  and _45766_ (_13620_, _13619_, _01954_);
  and _45767_ (_13621_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _45768_ (_13622_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _45769_ (_13623_, _13622_, _13621_);
  and _45770_ (_13624_, _13623_, _02150_);
  or _45771_ (_13625_, _13624_, _13620_);
  and _45772_ (_13626_, _13625_, _02131_);
  or _45773_ (_13627_, _13626_, _13616_);
  and _45774_ (_13628_, _13627_, _02157_);
  or _45775_ (_13629_, _13628_, _13606_);
  and _45776_ (_13630_, _13629_, _02194_);
  or _45777_ (_13631_, _13630_, _13584_);
  and _45778_ (_13632_, _13631_, _02005_);
  or _45779_ (_13633_, _13632_, _13538_);
  or _45780_ (_13634_, _13633_, _02374_);
  and _45781_ (_13635_, _13634_, _13444_);
  or _45782_ (_13636_, _13635_, _01748_);
  and _45783_ (_13637_, _13636_, _13254_);
  or _45784_ (_13638_, _13637_, _02141_);
  or _45785_ (_13639_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _45786_ (_13640_, _13639_, _27355_);
  and _45787_ (_15244_, _13640_, _13638_);
  and _45788_ (_13641_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _45789_ (_13642_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _45790_ (_13643_, _13642_, _13641_);
  and _45791_ (_13644_, _13643_, _01954_);
  and _45792_ (_13645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _45793_ (_13646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _45794_ (_13647_, _13646_, _13645_);
  and _45795_ (_13648_, _13647_, _02150_);
  or _45796_ (_13649_, _13648_, _13644_);
  or _45797_ (_13650_, _13649_, _02144_);
  and _45798_ (_13651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _45799_ (_13652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _45800_ (_13653_, _13652_, _13651_);
  and _45801_ (_13654_, _13653_, _01954_);
  and _45802_ (_13655_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and _45803_ (_13656_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _45804_ (_13657_, _13656_, _13655_);
  and _45805_ (_13658_, _13657_, _02150_);
  or _45806_ (_13659_, _13658_, _13654_);
  or _45807_ (_13660_, _13659_, _02131_);
  and _45808_ (_13661_, _13660_, _02157_);
  and _45809_ (_13662_, _13661_, _13650_);
  or _45810_ (_13663_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _45811_ (_13664_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _45812_ (_13665_, _13664_, _13663_);
  and _45813_ (_13666_, _13665_, _01954_);
  or _45814_ (_13667_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _45815_ (_13668_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _45816_ (_13669_, _13668_, _13667_);
  and _45817_ (_13670_, _13669_, _02150_);
  or _45818_ (_13671_, _13670_, _13666_);
  or _45819_ (_13672_, _13671_, _02144_);
  or _45820_ (_13673_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _45821_ (_13674_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _45822_ (_13675_, _13674_, _13673_);
  and _45823_ (_13676_, _13675_, _01954_);
  or _45824_ (_13677_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _45825_ (_13678_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _45826_ (_13679_, _13678_, _13677_);
  and _45827_ (_13680_, _13679_, _02150_);
  or _45828_ (_13681_, _13680_, _13676_);
  or _45829_ (_13682_, _13681_, _02131_);
  and _45830_ (_13684_, _13682_, _02077_);
  and _45831_ (_13685_, _13684_, _13672_);
  or _45832_ (_13686_, _13685_, _13662_);
  and _45833_ (_13687_, _13686_, _02065_);
  and _45834_ (_13688_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _45835_ (_13689_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _45836_ (_13690_, _13689_, _13688_);
  and _45837_ (_13691_, _13690_, _01954_);
  and _45838_ (_13692_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _45839_ (_13693_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _45840_ (_13695_, _13693_, _13692_);
  and _45841_ (_13696_, _13695_, _02150_);
  or _45842_ (_13697_, _13696_, _13691_);
  or _45843_ (_13698_, _13697_, _02144_);
  and _45844_ (_13699_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _45845_ (_13700_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _45846_ (_13701_, _13700_, _13699_);
  and _45847_ (_13702_, _13701_, _01954_);
  and _45848_ (_13703_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _45849_ (_13704_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _45850_ (_13706_, _13704_, _13703_);
  and _45851_ (_13707_, _13706_, _02150_);
  or _45852_ (_13708_, _13707_, _13702_);
  or _45853_ (_13709_, _13708_, _02131_);
  and _45854_ (_13710_, _13709_, _02157_);
  and _45855_ (_13711_, _13710_, _13698_);
  or _45856_ (_13712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _45857_ (_13713_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and _45858_ (_13714_, _13713_, _02150_);
  and _45859_ (_13715_, _13714_, _13712_);
  or _45860_ (_13717_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _45861_ (_13718_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _45862_ (_13719_, _13718_, _01954_);
  and _45863_ (_13720_, _13719_, _13717_);
  or _45864_ (_13721_, _13720_, _13715_);
  or _45865_ (_13722_, _13721_, _02144_);
  or _45866_ (_13723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _45867_ (_13724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and _45868_ (_13725_, _13724_, _02150_);
  and _45869_ (_13726_, _13725_, _13723_);
  or _45870_ (_13728_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _45871_ (_13729_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _45872_ (_13730_, _13729_, _01954_);
  and _45873_ (_13731_, _13730_, _13728_);
  or _45874_ (_13732_, _13731_, _13726_);
  or _45875_ (_13733_, _13732_, _02131_);
  and _45876_ (_13734_, _13733_, _02077_);
  and _45877_ (_13735_, _13734_, _13722_);
  or _45878_ (_13736_, _13735_, _13711_);
  and _45879_ (_13737_, _13736_, _02194_);
  or _45880_ (_13739_, _13737_, _13687_);
  and _45881_ (_13740_, _13739_, _02143_);
  and _45882_ (_13741_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _45883_ (_13742_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _45884_ (_13743_, _13742_, _13741_);
  and _45885_ (_13744_, _13743_, _01954_);
  and _45886_ (_13745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _45887_ (_13746_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _45888_ (_13747_, _13746_, _13745_);
  and _45889_ (_13748_, _13747_, _02150_);
  or _45890_ (_13750_, _13748_, _13744_);
  and _45891_ (_13751_, _13750_, _02131_);
  and _45892_ (_13752_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _45893_ (_13753_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _45894_ (_13754_, _13753_, _13752_);
  and _45895_ (_13755_, _13754_, _01954_);
  and _45896_ (_13756_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _45897_ (_13757_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _45898_ (_13758_, _13757_, _13756_);
  and _45899_ (_13759_, _13758_, _02150_);
  or _45900_ (_13761_, _13759_, _13755_);
  and _45901_ (_13762_, _13761_, _02144_);
  or _45902_ (_13763_, _13762_, _13751_);
  and _45903_ (_13764_, _13763_, _02157_);
  or _45904_ (_13765_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _45905_ (_13766_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _45906_ (_13767_, _13766_, _02150_);
  and _45907_ (_13768_, _13767_, _13765_);
  or _45908_ (_13769_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _45909_ (_13770_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _45910_ (_13772_, _13770_, _01954_);
  and _45911_ (_13773_, _13772_, _13769_);
  or _45912_ (_13774_, _13773_, _13768_);
  and _45913_ (_13775_, _13774_, _02131_);
  or _45914_ (_13776_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _45915_ (_13777_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _45916_ (_13778_, _13777_, _02150_);
  and _45917_ (_13779_, _13778_, _13776_);
  or _45918_ (_13780_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _45919_ (_13781_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _45920_ (_13783_, _13781_, _01954_);
  and _45921_ (_13784_, _13783_, _13780_);
  or _45922_ (_13785_, _13784_, _13779_);
  and _45923_ (_13786_, _13785_, _02144_);
  or _45924_ (_13787_, _13786_, _13775_);
  and _45925_ (_13788_, _13787_, _02077_);
  or _45926_ (_13789_, _13788_, _13764_);
  and _45927_ (_13790_, _13789_, _02194_);
  and _45928_ (_13791_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _45929_ (_13792_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _45930_ (_13794_, _13792_, _13791_);
  and _45931_ (_13795_, _13794_, _01954_);
  and _45932_ (_13796_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _45933_ (_13797_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _45934_ (_13798_, _13797_, _13796_);
  and _45935_ (_13799_, _13798_, _02150_);
  or _45936_ (_13800_, _13799_, _13795_);
  and _45937_ (_13801_, _13800_, _02131_);
  and _45938_ (_13802_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _45939_ (_13803_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _45940_ (_13805_, _13803_, _13802_);
  and _45941_ (_13806_, _13805_, _01954_);
  and _45942_ (_13807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and _45943_ (_13808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _45944_ (_13809_, _13808_, _13807_);
  and _45945_ (_13810_, _13809_, _02150_);
  or _45946_ (_13811_, _13810_, _13806_);
  and _45947_ (_13812_, _13811_, _02144_);
  or _45948_ (_13813_, _13812_, _13801_);
  and _45949_ (_13814_, _13813_, _02157_);
  or _45950_ (_13816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _45951_ (_13817_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and _45952_ (_13818_, _13817_, _13816_);
  and _45953_ (_13819_, _13818_, _01954_);
  or _45954_ (_13820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _45955_ (_13821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _45956_ (_13822_, _13821_, _13820_);
  and _45957_ (_13823_, _13822_, _02150_);
  or _45958_ (_13824_, _13823_, _13819_);
  and _45959_ (_13825_, _13824_, _02131_);
  or _45960_ (_13827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _45961_ (_13828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and _45962_ (_13829_, _13828_, _13827_);
  and _45963_ (_13830_, _13829_, _01954_);
  or _45964_ (_13831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _45965_ (_13832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _45966_ (_13833_, _13832_, _13831_);
  and _45967_ (_13834_, _13833_, _02150_);
  or _45968_ (_13835_, _13834_, _13830_);
  and _45969_ (_13836_, _13835_, _02144_);
  or _45970_ (_13837_, _13836_, _13825_);
  and _45971_ (_13838_, _13837_, _02077_);
  or _45972_ (_13839_, _13838_, _13814_);
  and _45973_ (_13840_, _13839_, _02065_);
  or _45974_ (_13841_, _13840_, _13790_);
  and _45975_ (_13842_, _13841_, _02005_);
  or _45976_ (_13843_, _13842_, _13740_);
  or _45977_ (_13844_, _13843_, _02054_);
  and _45978_ (_13845_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _45979_ (_13846_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _45980_ (_13847_, _13846_, _13845_);
  and _45981_ (_13848_, _13847_, _01954_);
  and _45982_ (_13849_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _45983_ (_13850_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _45984_ (_13851_, _13850_, _13849_);
  and _45985_ (_13852_, _13851_, _02150_);
  or _45986_ (_13853_, _13852_, _13848_);
  or _45987_ (_13854_, _13853_, _02144_);
  and _45988_ (_13855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _45989_ (_13856_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _45990_ (_13857_, _13856_, _13855_);
  and _45991_ (_13858_, _13857_, _01954_);
  and _45992_ (_13859_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _45993_ (_13860_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _45994_ (_13861_, _13860_, _13859_);
  and _45995_ (_13862_, _13861_, _02150_);
  or _45996_ (_13863_, _13862_, _13858_);
  or _45997_ (_13864_, _13863_, _02131_);
  and _45998_ (_13865_, _13864_, _02157_);
  and _45999_ (_13866_, _13865_, _13854_);
  or _46000_ (_13867_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _46001_ (_13868_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _46002_ (_13869_, _13868_, _02150_);
  and _46003_ (_13870_, _13869_, _13867_);
  or _46004_ (_13871_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _46005_ (_13872_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _46006_ (_13873_, _13872_, _01954_);
  and _46007_ (_13874_, _13873_, _13871_);
  or _46008_ (_13875_, _13874_, _13870_);
  or _46009_ (_13876_, _13875_, _02144_);
  or _46010_ (_13877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _46011_ (_13878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and _46012_ (_13879_, _13878_, _02150_);
  and _46013_ (_13880_, _13879_, _13877_);
  or _46014_ (_13881_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _46015_ (_13882_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and _46016_ (_13883_, _13882_, _01954_);
  and _46017_ (_13884_, _13883_, _13881_);
  or _46018_ (_13885_, _13884_, _13880_);
  or _46019_ (_13886_, _13885_, _02131_);
  and _46020_ (_13887_, _13886_, _02077_);
  and _46021_ (_13888_, _13887_, _13876_);
  or _46022_ (_13889_, _13888_, _13866_);
  and _46023_ (_13890_, _13889_, _02194_);
  and _46024_ (_13891_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _46025_ (_13892_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _46026_ (_13893_, _13892_, _13891_);
  and _46027_ (_13894_, _13893_, _01954_);
  and _46028_ (_13895_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _46029_ (_13896_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _46030_ (_13897_, _13896_, _13895_);
  and _46031_ (_13898_, _13897_, _02150_);
  or _46032_ (_13899_, _13898_, _13894_);
  or _46033_ (_13900_, _13899_, _02144_);
  and _46034_ (_13901_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _46035_ (_13902_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _46036_ (_13903_, _13902_, _13901_);
  and _46037_ (_13904_, _13903_, _01954_);
  and _46038_ (_13905_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _46039_ (_13906_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _46040_ (_13907_, _13906_, _13905_);
  and _46041_ (_13908_, _13907_, _02150_);
  or _46042_ (_13909_, _13908_, _13904_);
  or _46043_ (_13910_, _13909_, _02131_);
  and _46044_ (_13911_, _13910_, _02157_);
  and _46045_ (_13912_, _13911_, _13900_);
  or _46046_ (_13913_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _46047_ (_13914_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _46048_ (_13915_, _13914_, _13913_);
  and _46049_ (_13916_, _13915_, _01954_);
  or _46050_ (_13917_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _46051_ (_13918_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _46052_ (_13919_, _13918_, _13917_);
  and _46053_ (_13920_, _13919_, _02150_);
  or _46054_ (_13921_, _13920_, _13916_);
  or _46055_ (_13922_, _13921_, _02144_);
  or _46056_ (_13923_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _46057_ (_13924_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _46058_ (_13925_, _13924_, _13923_);
  and _46059_ (_13926_, _13925_, _01954_);
  or _46060_ (_13927_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _46061_ (_13928_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _46062_ (_13929_, _13928_, _13927_);
  and _46063_ (_13930_, _13929_, _02150_);
  or _46064_ (_13931_, _13930_, _13926_);
  or _46065_ (_13932_, _13931_, _02131_);
  and _46066_ (_13933_, _13932_, _02077_);
  and _46067_ (_13934_, _13933_, _13922_);
  or _46068_ (_13935_, _13934_, _13912_);
  and _46069_ (_13936_, _13935_, _02065_);
  or _46070_ (_13937_, _13936_, _13890_);
  and _46071_ (_13938_, _13937_, _02143_);
  or _46072_ (_13939_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _46073_ (_13940_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and _46074_ (_13941_, _13940_, _13939_);
  and _46075_ (_13942_, _13941_, _01954_);
  or _46076_ (_13943_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _46077_ (_13944_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _46078_ (_13945_, _13944_, _13943_);
  and _46079_ (_13946_, _13945_, _02150_);
  or _46080_ (_13947_, _13946_, _13942_);
  and _46081_ (_13948_, _13947_, _02144_);
  or _46082_ (_13949_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _46083_ (_13950_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _46084_ (_13951_, _13950_, _13949_);
  and _46085_ (_13952_, _13951_, _01954_);
  or _46086_ (_13953_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _46087_ (_13954_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _46088_ (_13955_, _13954_, _13953_);
  and _46089_ (_13956_, _13955_, _02150_);
  or _46090_ (_13957_, _13956_, _13952_);
  and _46091_ (_13958_, _13957_, _02131_);
  or _46092_ (_13959_, _13958_, _13948_);
  and _46093_ (_13960_, _13959_, _02077_);
  and _46094_ (_13961_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and _46095_ (_13962_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _46096_ (_13963_, _13962_, _13961_);
  and _46097_ (_13964_, _13963_, _01954_);
  and _46098_ (_13965_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and _46099_ (_13966_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _46100_ (_13967_, _13966_, _13965_);
  and _46101_ (_13968_, _13967_, _02150_);
  or _46102_ (_13969_, _13968_, _13964_);
  and _46103_ (_13970_, _13969_, _02144_);
  and _46104_ (_13971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and _46105_ (_13972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _46106_ (_13973_, _13972_, _13971_);
  and _46107_ (_13974_, _13973_, _01954_);
  and _46108_ (_13975_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _46109_ (_13976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _46110_ (_13977_, _13976_, _13975_);
  and _46111_ (_13978_, _13977_, _02150_);
  or _46112_ (_13979_, _13978_, _13974_);
  and _46113_ (_13980_, _13979_, _02131_);
  or _46114_ (_13981_, _13980_, _13970_);
  and _46115_ (_13982_, _13981_, _02157_);
  or _46116_ (_13983_, _13982_, _13960_);
  and _46117_ (_13984_, _13983_, _02065_);
  or _46118_ (_13985_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _46119_ (_13986_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _46120_ (_13987_, _13986_, _02150_);
  and _46121_ (_13988_, _13987_, _13985_);
  or _46122_ (_13989_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _46123_ (_13990_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _46124_ (_13991_, _13990_, _01954_);
  and _46125_ (_13992_, _13991_, _13989_);
  or _46126_ (_13993_, _13992_, _13988_);
  and _46127_ (_13994_, _13993_, _02144_);
  or _46128_ (_13995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _46129_ (_13996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _46130_ (_13997_, _13996_, _02150_);
  and _46131_ (_13998_, _13997_, _13995_);
  or _46132_ (_13999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _46133_ (_14000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and _46134_ (_14001_, _14000_, _01954_);
  and _46135_ (_14002_, _14001_, _13999_);
  or _46136_ (_14003_, _14002_, _13998_);
  and _46137_ (_14004_, _14003_, _02131_);
  or _46138_ (_14005_, _14004_, _13994_);
  and _46139_ (_14006_, _14005_, _02077_);
  and _46140_ (_14007_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and _46141_ (_14008_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _46142_ (_14009_, _14008_, _14007_);
  and _46143_ (_14010_, _14009_, _01954_);
  and _46144_ (_14011_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _46145_ (_14012_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _46146_ (_14013_, _14012_, _14011_);
  and _46147_ (_14014_, _14013_, _02150_);
  or _46148_ (_14015_, _14014_, _14010_);
  and _46149_ (_14016_, _14015_, _02144_);
  and _46150_ (_14017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _46151_ (_14018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _46152_ (_14019_, _14018_, _14017_);
  and _46153_ (_14020_, _14019_, _01954_);
  and _46154_ (_14021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _46155_ (_14022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _46156_ (_14023_, _14022_, _14021_);
  and _46157_ (_14024_, _14023_, _02150_);
  or _46158_ (_14025_, _14024_, _14020_);
  and _46159_ (_14026_, _14025_, _02131_);
  or _46160_ (_14027_, _14026_, _14016_);
  and _46161_ (_14028_, _14027_, _02157_);
  or _46162_ (_14029_, _14028_, _14006_);
  and _46163_ (_14030_, _14029_, _02194_);
  or _46164_ (_14031_, _14030_, _13984_);
  and _46165_ (_14032_, _14031_, _02005_);
  or _46166_ (_14033_, _14032_, _13938_);
  or _46167_ (_14034_, _14033_, _02374_);
  and _46168_ (_14035_, _14034_, _13844_);
  or _46169_ (_14036_, _14035_, _02142_);
  and _46170_ (_14037_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and _46171_ (_14038_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _46172_ (_14039_, _14038_, _14037_);
  and _46173_ (_14040_, _14039_, _01954_);
  and _46174_ (_14041_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _46175_ (_14042_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _46176_ (_14043_, _14042_, _14041_);
  and _46177_ (_14044_, _14043_, _02150_);
  or _46178_ (_14045_, _14044_, _14040_);
  or _46179_ (_14046_, _14045_, _02144_);
  and _46180_ (_14047_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _46181_ (_14048_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _46182_ (_14049_, _14048_, _14047_);
  and _46183_ (_14050_, _14049_, _01954_);
  and _46184_ (_14051_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _46185_ (_14052_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _46186_ (_14053_, _14052_, _14051_);
  and _46187_ (_14054_, _14053_, _02150_);
  or _46188_ (_14055_, _14054_, _14050_);
  or _46189_ (_14056_, _14055_, _02131_);
  and _46190_ (_14057_, _14056_, _02157_);
  and _46191_ (_14058_, _14057_, _14046_);
  or _46192_ (_14059_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _46193_ (_14060_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _46194_ (_14061_, _14060_, _14059_);
  and _46195_ (_14062_, _14061_, _01954_);
  or _46196_ (_14063_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _46197_ (_14064_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _46198_ (_14065_, _14064_, _14063_);
  and _46199_ (_14066_, _14065_, _02150_);
  or _46200_ (_14067_, _14066_, _14062_);
  or _46201_ (_14068_, _14067_, _02144_);
  or _46202_ (_14069_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _46203_ (_14070_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and _46204_ (_14071_, _14070_, _14069_);
  and _46205_ (_14072_, _14071_, _01954_);
  or _46206_ (_14073_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _46207_ (_14074_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _46208_ (_14075_, _14074_, _14073_);
  and _46209_ (_14076_, _14075_, _02150_);
  or _46210_ (_14077_, _14076_, _14072_);
  or _46211_ (_14078_, _14077_, _02131_);
  and _46212_ (_14079_, _14078_, _02077_);
  and _46213_ (_14080_, _14079_, _14068_);
  or _46214_ (_14081_, _14080_, _14058_);
  and _46215_ (_14082_, _14081_, _02065_);
  and _46216_ (_14083_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _46217_ (_14084_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _46218_ (_14085_, _14084_, _14083_);
  and _46219_ (_14086_, _14085_, _01954_);
  and _46220_ (_14087_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _46221_ (_14088_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _46222_ (_14089_, _14088_, _14087_);
  and _46223_ (_14090_, _14089_, _02150_);
  or _46224_ (_14091_, _14090_, _14086_);
  or _46225_ (_14092_, _14091_, _02144_);
  and _46226_ (_14093_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _46227_ (_14094_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _46228_ (_14095_, _14094_, _14093_);
  and _46229_ (_14096_, _14095_, _01954_);
  and _46230_ (_14097_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _46231_ (_14098_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _46232_ (_14099_, _14098_, _14097_);
  and _46233_ (_14100_, _14099_, _02150_);
  or _46234_ (_14101_, _14100_, _14096_);
  or _46235_ (_14102_, _14101_, _02131_);
  and _46236_ (_14103_, _14102_, _02157_);
  and _46237_ (_14104_, _14103_, _14092_);
  or _46238_ (_14105_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _46239_ (_14106_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _46240_ (_14107_, _14106_, _02150_);
  and _46241_ (_14108_, _14107_, _14105_);
  or _46242_ (_14109_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _46243_ (_14110_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _46244_ (_14111_, _14110_, _01954_);
  and _46245_ (_14112_, _14111_, _14109_);
  or _46246_ (_14113_, _14112_, _14108_);
  or _46247_ (_14114_, _14113_, _02144_);
  or _46248_ (_14115_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _46249_ (_14116_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _46250_ (_14117_, _14116_, _02150_);
  and _46251_ (_14118_, _14117_, _14115_);
  or _46252_ (_14119_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _46253_ (_14120_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _46254_ (_14121_, _14120_, _01954_);
  and _46255_ (_14122_, _14121_, _14119_);
  or _46256_ (_14123_, _14122_, _14118_);
  or _46257_ (_14124_, _14123_, _02131_);
  and _46258_ (_14125_, _14124_, _02077_);
  and _46259_ (_14126_, _14125_, _14114_);
  or _46260_ (_14127_, _14126_, _14104_);
  and _46261_ (_14128_, _14127_, _02194_);
  or _46262_ (_14129_, _14128_, _14082_);
  and _46263_ (_14130_, _14129_, _02143_);
  and _46264_ (_14131_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _46265_ (_14132_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _46266_ (_14133_, _14132_, _14131_);
  and _46267_ (_14134_, _14133_, _01954_);
  and _46268_ (_14135_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _46269_ (_14136_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _46270_ (_14137_, _14136_, _14135_);
  and _46271_ (_14138_, _14137_, _02150_);
  or _46272_ (_14139_, _14138_, _14134_);
  and _46273_ (_14140_, _14139_, _02131_);
  and _46274_ (_14141_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _46275_ (_14142_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _46276_ (_14143_, _14142_, _14141_);
  and _46277_ (_14144_, _14143_, _01954_);
  and _46278_ (_14145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _46279_ (_14146_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _46280_ (_14147_, _14146_, _14145_);
  and _46281_ (_14148_, _14147_, _02150_);
  or _46282_ (_14149_, _14148_, _14144_);
  and _46283_ (_14150_, _14149_, _02144_);
  or _46284_ (_14151_, _14150_, _14140_);
  and _46285_ (_14152_, _14151_, _02157_);
  or _46286_ (_14153_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _46287_ (_14154_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _46288_ (_14155_, _14154_, _02150_);
  and _46289_ (_14156_, _14155_, _14153_);
  or _46290_ (_14157_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _46291_ (_14158_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _46292_ (_14159_, _14158_, _01954_);
  and _46293_ (_14160_, _14159_, _14157_);
  or _46294_ (_14161_, _14160_, _14156_);
  and _46295_ (_14162_, _14161_, _02131_);
  or _46296_ (_14163_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _46297_ (_14164_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _46298_ (_14165_, _14164_, _02150_);
  and _46299_ (_14166_, _14165_, _14163_);
  or _46300_ (_14167_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _46301_ (_14168_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _46302_ (_14169_, _14168_, _01954_);
  and _46303_ (_14170_, _14169_, _14167_);
  or _46304_ (_14171_, _14170_, _14166_);
  and _46305_ (_14172_, _14171_, _02144_);
  or _46306_ (_14173_, _14172_, _14162_);
  and _46307_ (_14174_, _14173_, _02077_);
  or _46308_ (_14175_, _14174_, _14152_);
  and _46309_ (_14176_, _14175_, _02194_);
  and _46310_ (_14177_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _46311_ (_14178_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _46312_ (_14179_, _14178_, _14177_);
  and _46313_ (_14180_, _14179_, _01954_);
  and _46314_ (_14181_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _46315_ (_14182_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _46316_ (_14183_, _14182_, _14181_);
  and _46317_ (_14184_, _14183_, _02150_);
  or _46318_ (_14185_, _14184_, _14180_);
  and _46319_ (_14186_, _14185_, _02131_);
  and _46320_ (_14187_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _46321_ (_14188_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _46322_ (_14189_, _14188_, _14187_);
  and _46323_ (_14190_, _14189_, _01954_);
  and _46324_ (_14191_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _46325_ (_14192_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _46326_ (_14193_, _14192_, _14191_);
  and _46327_ (_14194_, _14193_, _02150_);
  or _46328_ (_14195_, _14194_, _14190_);
  and _46329_ (_14196_, _14195_, _02144_);
  or _46330_ (_14197_, _14196_, _14186_);
  and _46331_ (_14198_, _14197_, _02157_);
  or _46332_ (_14199_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _46333_ (_14200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _46334_ (_14201_, _14200_, _14199_);
  and _46335_ (_14202_, _14201_, _01954_);
  or _46336_ (_14203_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _46337_ (_14204_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _46338_ (_14205_, _14204_, _14203_);
  and _46339_ (_14206_, _14205_, _02150_);
  or _46340_ (_14207_, _14206_, _14202_);
  and _46341_ (_14208_, _14207_, _02131_);
  or _46342_ (_14209_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _46343_ (_14210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _46344_ (_14211_, _14210_, _14209_);
  and _46345_ (_14212_, _14211_, _01954_);
  or _46346_ (_14213_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _46347_ (_14214_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _46348_ (_14215_, _14214_, _14213_);
  and _46349_ (_14216_, _14215_, _02150_);
  or _46350_ (_14217_, _14216_, _14212_);
  and _46351_ (_14218_, _14217_, _02144_);
  or _46352_ (_14219_, _14218_, _14208_);
  and _46353_ (_14220_, _14219_, _02077_);
  or _46354_ (_14221_, _14220_, _14198_);
  and _46355_ (_14222_, _14221_, _02065_);
  or _46356_ (_14223_, _14222_, _14176_);
  and _46357_ (_14224_, _14223_, _02005_);
  or _46358_ (_14225_, _14224_, _14130_);
  or _46359_ (_14226_, _14225_, _02054_);
  and _46360_ (_14227_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and _46361_ (_14228_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _46362_ (_14229_, _14228_, _14227_);
  and _46363_ (_14230_, _14229_, _01954_);
  and _46364_ (_14231_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _46365_ (_14232_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _46366_ (_14233_, _14232_, _14231_);
  and _46367_ (_14234_, _14233_, _02150_);
  or _46368_ (_14235_, _14234_, _14230_);
  or _46369_ (_14236_, _14235_, _02144_);
  and _46370_ (_14237_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _46371_ (_14238_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _46372_ (_14239_, _14238_, _14237_);
  and _46373_ (_14240_, _14239_, _01954_);
  and _46374_ (_14241_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and _46375_ (_14242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _46376_ (_14243_, _14242_, _14241_);
  and _46377_ (_14244_, _14243_, _02150_);
  or _46378_ (_14245_, _14244_, _14240_);
  or _46379_ (_14246_, _14245_, _02131_);
  and _46380_ (_14247_, _14246_, _02157_);
  and _46381_ (_14248_, _14247_, _14236_);
  or _46382_ (_14249_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _46383_ (_14250_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _46384_ (_14251_, _14250_, _02150_);
  and _46385_ (_14252_, _14251_, _14249_);
  or _46386_ (_14253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _46387_ (_14254_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _46388_ (_14255_, _14254_, _01954_);
  and _46389_ (_14256_, _14255_, _14253_);
  or _46390_ (_14257_, _14256_, _14252_);
  or _46391_ (_14258_, _14257_, _02144_);
  or _46392_ (_14259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _46393_ (_14260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and _46394_ (_14261_, _14260_, _02150_);
  and _46395_ (_14262_, _14261_, _14259_);
  or _46396_ (_14263_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _46397_ (_14264_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and _46398_ (_14265_, _14264_, _01954_);
  and _46399_ (_14266_, _14265_, _14263_);
  or _46400_ (_14267_, _14266_, _14262_);
  or _46401_ (_14268_, _14267_, _02131_);
  and _46402_ (_14269_, _14268_, _02077_);
  and _46403_ (_14270_, _14269_, _14258_);
  or _46404_ (_14271_, _14270_, _14248_);
  and _46405_ (_14272_, _14271_, _02194_);
  and _46406_ (_14273_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _46407_ (_14274_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _46408_ (_14275_, _14274_, _14273_);
  and _46409_ (_14276_, _14275_, _01954_);
  and _46410_ (_14277_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _46411_ (_14278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _46412_ (_14279_, _14278_, _14277_);
  and _46413_ (_14280_, _14279_, _02150_);
  or _46414_ (_14281_, _14280_, _14276_);
  or _46415_ (_14282_, _14281_, _02144_);
  and _46416_ (_14283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _46417_ (_14284_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _46418_ (_14285_, _14284_, _14283_);
  and _46419_ (_14286_, _14285_, _01954_);
  and _46420_ (_14287_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _46421_ (_14288_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _46422_ (_14289_, _14288_, _14287_);
  and _46423_ (_14290_, _14289_, _02150_);
  or _46424_ (_14291_, _14290_, _14286_);
  or _46425_ (_14292_, _14291_, _02131_);
  and _46426_ (_14293_, _14292_, _02157_);
  and _46427_ (_14294_, _14293_, _14282_);
  or _46428_ (_14295_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _46429_ (_14296_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _46430_ (_14297_, _14296_, _14295_);
  and _46431_ (_14298_, _14297_, _01954_);
  or _46432_ (_14299_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _46433_ (_14300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _46434_ (_14301_, _14300_, _14299_);
  and _46435_ (_14302_, _14301_, _02150_);
  or _46436_ (_14303_, _14302_, _14298_);
  or _46437_ (_14304_, _14303_, _02144_);
  or _46438_ (_14305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _46439_ (_14306_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _46440_ (_14307_, _14306_, _14305_);
  and _46441_ (_14308_, _14307_, _01954_);
  or _46442_ (_14309_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _46443_ (_14310_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _46444_ (_14311_, _14310_, _14309_);
  and _46445_ (_14312_, _14311_, _02150_);
  or _46446_ (_14313_, _14312_, _14308_);
  or _46447_ (_14314_, _14313_, _02131_);
  and _46448_ (_14315_, _14314_, _02077_);
  and _46449_ (_14316_, _14315_, _14304_);
  or _46450_ (_14317_, _14316_, _14294_);
  and _46451_ (_14318_, _14317_, _02065_);
  or _46452_ (_14319_, _14318_, _14272_);
  and _46453_ (_14320_, _14319_, _02143_);
  or _46454_ (_14321_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _46455_ (_14322_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _46456_ (_14323_, _14322_, _14321_);
  and _46457_ (_14324_, _14323_, _01954_);
  or _46458_ (_14325_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _46459_ (_14326_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _46460_ (_14327_, _14326_, _14325_);
  and _46461_ (_14328_, _14327_, _02150_);
  or _46462_ (_14329_, _14328_, _14324_);
  and _46463_ (_14330_, _14329_, _02144_);
  or _46464_ (_14331_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _46465_ (_14332_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _46466_ (_14333_, _14332_, _14331_);
  and _46467_ (_14334_, _14333_, _01954_);
  or _46468_ (_14335_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _46469_ (_14336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _46470_ (_14337_, _14336_, _14335_);
  and _46471_ (_14338_, _14337_, _02150_);
  or _46472_ (_14339_, _14338_, _14334_);
  and _46473_ (_14340_, _14339_, _02131_);
  or _46474_ (_14341_, _14340_, _14330_);
  and _46475_ (_14342_, _14341_, _02077_);
  and _46476_ (_14343_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _46477_ (_14344_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _46478_ (_14345_, _14344_, _14343_);
  and _46479_ (_14346_, _14345_, _01954_);
  and _46480_ (_14347_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _46481_ (_14348_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _46482_ (_14349_, _14348_, _14347_);
  and _46483_ (_14350_, _14349_, _02150_);
  or _46484_ (_14351_, _14350_, _14346_);
  and _46485_ (_14352_, _14351_, _02144_);
  and _46486_ (_14353_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _46487_ (_14354_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _46488_ (_14355_, _14354_, _14353_);
  and _46489_ (_14356_, _14355_, _01954_);
  and _46490_ (_14357_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _46491_ (_14358_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _46492_ (_14359_, _14358_, _14357_);
  and _46493_ (_14360_, _14359_, _02150_);
  or _46494_ (_14361_, _14360_, _14356_);
  and _46495_ (_14362_, _14361_, _02131_);
  or _46496_ (_14363_, _14362_, _14352_);
  and _46497_ (_14364_, _14363_, _02157_);
  or _46498_ (_14365_, _14364_, _14342_);
  and _46499_ (_14366_, _14365_, _02065_);
  or _46500_ (_14367_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _46501_ (_14368_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _46502_ (_14369_, _14368_, _02150_);
  and _46503_ (_14370_, _14369_, _14367_);
  or _46504_ (_14371_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _46505_ (_14372_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _46506_ (_14373_, _14372_, _01954_);
  and _46507_ (_14374_, _14373_, _14371_);
  or _46508_ (_14375_, _14374_, _14370_);
  and _46509_ (_14376_, _14375_, _02144_);
  or _46510_ (_14377_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _46511_ (_14378_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _46512_ (_14379_, _14378_, _02150_);
  and _46513_ (_14380_, _14379_, _14377_);
  or _46514_ (_14381_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _46515_ (_14382_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _46516_ (_14383_, _14382_, _01954_);
  and _46517_ (_14384_, _14383_, _14381_);
  or _46518_ (_14385_, _14384_, _14380_);
  and _46519_ (_14386_, _14385_, _02131_);
  or _46520_ (_14387_, _14386_, _14376_);
  and _46521_ (_14388_, _14387_, _02077_);
  and _46522_ (_14389_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _46523_ (_14390_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _46524_ (_14391_, _14390_, _14389_);
  and _46525_ (_14392_, _14391_, _01954_);
  and _46526_ (_14393_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _46527_ (_14394_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _46528_ (_14395_, _14394_, _14393_);
  and _46529_ (_14396_, _14395_, _02150_);
  or _46530_ (_14397_, _14396_, _14392_);
  and _46531_ (_14398_, _14397_, _02144_);
  and _46532_ (_14399_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and _46533_ (_14400_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _46534_ (_14401_, _14400_, _14399_);
  and _46535_ (_14402_, _14401_, _01954_);
  and _46536_ (_14403_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _46537_ (_14404_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _46538_ (_14405_, _14404_, _14403_);
  and _46539_ (_14406_, _14405_, _02150_);
  or _46540_ (_14407_, _14406_, _14402_);
  and _46541_ (_14408_, _14407_, _02131_);
  or _46542_ (_14409_, _14408_, _14398_);
  and _46543_ (_14410_, _14409_, _02157_);
  or _46544_ (_14411_, _14410_, _14388_);
  and _46545_ (_14412_, _14411_, _02194_);
  or _46546_ (_14413_, _14412_, _14366_);
  and _46547_ (_14414_, _14413_, _02005_);
  or _46548_ (_14415_, _14414_, _14320_);
  or _46549_ (_14416_, _14415_, _02374_);
  and _46550_ (_14417_, _14416_, _14226_);
  or _46551_ (_14418_, _14417_, _01748_);
  and _46552_ (_14419_, _14418_, _14036_);
  or _46553_ (_14420_, _14419_, _02141_);
  or _46554_ (_14421_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _46555_ (_14422_, _14421_, _27355_);
  and _46556_ (_15246_, _14422_, _14420_);
  and _46557_ (_14423_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _46558_ (_14424_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _46559_ (_14425_, _14424_, _14423_);
  and _46560_ (_14426_, _14425_, _01954_);
  and _46561_ (_14427_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _46562_ (_14428_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _46563_ (_14429_, _14428_, _14427_);
  and _46564_ (_14430_, _14429_, _02150_);
  or _46565_ (_14431_, _14430_, _14426_);
  or _46566_ (_14432_, _14431_, _02144_);
  and _46567_ (_14433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _46568_ (_14434_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _46569_ (_14435_, _14434_, _14433_);
  and _46570_ (_14436_, _14435_, _01954_);
  and _46571_ (_14437_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _46572_ (_14438_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _46573_ (_14439_, _14438_, _14437_);
  and _46574_ (_14440_, _14439_, _02150_);
  or _46575_ (_14441_, _14440_, _14436_);
  or _46576_ (_14442_, _14441_, _02131_);
  and _46577_ (_14443_, _14442_, _02157_);
  and _46578_ (_14444_, _14443_, _14432_);
  or _46579_ (_14445_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _46580_ (_14446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _46581_ (_14447_, _14446_, _14445_);
  and _46582_ (_14448_, _14447_, _01954_);
  or _46583_ (_14449_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _46584_ (_14450_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _46585_ (_14451_, _14450_, _14449_);
  and _46586_ (_14452_, _14451_, _02150_);
  or _46587_ (_14453_, _14452_, _14448_);
  or _46588_ (_14454_, _14453_, _02144_);
  or _46589_ (_14455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _46590_ (_14456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and _46591_ (_14457_, _14456_, _14455_);
  and _46592_ (_14458_, _14457_, _01954_);
  or _46593_ (_14459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _46594_ (_14460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _46595_ (_14461_, _14460_, _14459_);
  and _46596_ (_14462_, _14461_, _02150_);
  or _46597_ (_14463_, _14462_, _14458_);
  or _46598_ (_14464_, _14463_, _02131_);
  and _46599_ (_14465_, _14464_, _02077_);
  and _46600_ (_14466_, _14465_, _14454_);
  or _46601_ (_14467_, _14466_, _14444_);
  and _46602_ (_14468_, _14467_, _02065_);
  and _46603_ (_14469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _46604_ (_14470_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _46605_ (_14471_, _14470_, _14469_);
  and _46606_ (_14472_, _14471_, _01954_);
  and _46607_ (_14473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _46608_ (_14474_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _46609_ (_14475_, _14474_, _14473_);
  and _46610_ (_14476_, _14475_, _02150_);
  or _46611_ (_14477_, _14476_, _14472_);
  or _46612_ (_14478_, _14477_, _02144_);
  and _46613_ (_14479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _46614_ (_14480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _46615_ (_14481_, _14480_, _14479_);
  and _46616_ (_14482_, _14481_, _01954_);
  and _46617_ (_14483_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _46618_ (_14484_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _46619_ (_14485_, _14484_, _14483_);
  and _46620_ (_14486_, _14485_, _02150_);
  or _46621_ (_14487_, _14486_, _14482_);
  or _46622_ (_14488_, _14487_, _02131_);
  and _46623_ (_14489_, _14488_, _02157_);
  and _46624_ (_14490_, _14489_, _14478_);
  or _46625_ (_14491_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _46626_ (_14492_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _46627_ (_14493_, _14492_, _02150_);
  and _46628_ (_14494_, _14493_, _14491_);
  or _46629_ (_14495_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _46630_ (_14496_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _46631_ (_14497_, _14496_, _01954_);
  and _46632_ (_14498_, _14497_, _14495_);
  or _46633_ (_14499_, _14498_, _14494_);
  or _46634_ (_14500_, _14499_, _02144_);
  or _46635_ (_14501_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _46636_ (_14502_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _46637_ (_14503_, _14502_, _02150_);
  and _46638_ (_14504_, _14503_, _14501_);
  or _46639_ (_14505_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _46640_ (_14506_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _46641_ (_14507_, _14506_, _01954_);
  and _46642_ (_14508_, _14507_, _14505_);
  or _46643_ (_14509_, _14508_, _14504_);
  or _46644_ (_14510_, _14509_, _02131_);
  and _46645_ (_14511_, _14510_, _02077_);
  and _46646_ (_14512_, _14511_, _14500_);
  or _46647_ (_14513_, _14512_, _14490_);
  and _46648_ (_14514_, _14513_, _02194_);
  or _46649_ (_14515_, _14514_, _14468_);
  and _46650_ (_14516_, _14515_, _02143_);
  and _46651_ (_14517_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _46652_ (_14518_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _46653_ (_14519_, _14518_, _14517_);
  and _46654_ (_14520_, _14519_, _01954_);
  and _46655_ (_14521_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _46656_ (_14522_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _46657_ (_14523_, _14522_, _14521_);
  and _46658_ (_14524_, _14523_, _02150_);
  or _46659_ (_14525_, _14524_, _14520_);
  and _46660_ (_14526_, _14525_, _02131_);
  and _46661_ (_14527_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _46662_ (_14528_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _46663_ (_14529_, _14528_, _14527_);
  and _46664_ (_14530_, _14529_, _01954_);
  and _46665_ (_14531_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _46666_ (_14532_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _46667_ (_14533_, _14532_, _14531_);
  and _46668_ (_14534_, _14533_, _02150_);
  or _46669_ (_14535_, _14534_, _14530_);
  and _46670_ (_14536_, _14535_, _02144_);
  or _46671_ (_14537_, _14536_, _14526_);
  and _46672_ (_14538_, _14537_, _02157_);
  or _46673_ (_14539_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _46674_ (_14540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _46675_ (_14541_, _14540_, _02150_);
  and _46676_ (_14542_, _14541_, _14539_);
  or _46677_ (_14543_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _46678_ (_14544_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _46679_ (_14545_, _14544_, _01954_);
  and _46680_ (_14546_, _14545_, _14543_);
  or _46681_ (_14547_, _14546_, _14542_);
  and _46682_ (_14548_, _14547_, _02131_);
  or _46683_ (_14549_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _46684_ (_14550_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _46685_ (_14551_, _14550_, _02150_);
  and _46686_ (_14552_, _14551_, _14549_);
  or _46687_ (_14553_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _46688_ (_14554_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _46689_ (_14555_, _14554_, _01954_);
  and _46690_ (_14556_, _14555_, _14553_);
  or _46691_ (_14557_, _14556_, _14552_);
  and _46692_ (_14558_, _14557_, _02144_);
  or _46693_ (_14559_, _14558_, _14548_);
  and _46694_ (_14560_, _14559_, _02077_);
  or _46695_ (_14561_, _14560_, _14538_);
  and _46696_ (_14562_, _14561_, _02194_);
  and _46697_ (_14563_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and _46698_ (_14564_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _46699_ (_14565_, _14564_, _14563_);
  and _46700_ (_14566_, _14565_, _01954_);
  and _46701_ (_14567_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _46702_ (_14568_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _46703_ (_14569_, _14568_, _14567_);
  and _46704_ (_14570_, _14569_, _02150_);
  or _46705_ (_14571_, _14570_, _14566_);
  and _46706_ (_14572_, _14571_, _02131_);
  and _46707_ (_14573_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and _46708_ (_14574_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _46709_ (_14575_, _14574_, _14573_);
  and _46710_ (_14576_, _14575_, _01954_);
  and _46711_ (_14577_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and _46712_ (_14578_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _46713_ (_14579_, _14578_, _14577_);
  and _46714_ (_14580_, _14579_, _02150_);
  or _46715_ (_14581_, _14580_, _14576_);
  and _46716_ (_14582_, _14581_, _02144_);
  or _46717_ (_14583_, _14582_, _14572_);
  and _46718_ (_14584_, _14583_, _02157_);
  or _46719_ (_14585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _46720_ (_14586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and _46721_ (_14587_, _14586_, _14585_);
  and _46722_ (_14588_, _14587_, _01954_);
  or _46723_ (_14589_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _46724_ (_14590_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _46725_ (_14591_, _14590_, _14589_);
  and _46726_ (_14592_, _14591_, _02150_);
  or _46727_ (_14593_, _14592_, _14588_);
  and _46728_ (_14594_, _14593_, _02131_);
  or _46729_ (_14595_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _46730_ (_14596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and _46731_ (_14597_, _14596_, _14595_);
  and _46732_ (_14598_, _14597_, _01954_);
  or _46733_ (_14599_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _46734_ (_14600_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _46735_ (_14601_, _14600_, _14599_);
  and _46736_ (_14602_, _14601_, _02150_);
  or _46737_ (_14603_, _14602_, _14598_);
  and _46738_ (_14604_, _14603_, _02144_);
  or _46739_ (_14605_, _14604_, _14594_);
  and _46740_ (_14606_, _14605_, _02077_);
  or _46741_ (_14607_, _14606_, _14584_);
  and _46742_ (_14608_, _14607_, _02065_);
  or _46743_ (_14609_, _14608_, _14562_);
  and _46744_ (_14610_, _14609_, _02005_);
  or _46745_ (_14611_, _14610_, _14516_);
  or _46746_ (_14612_, _14611_, _02054_);
  and _46747_ (_14613_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and _46748_ (_14614_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _46749_ (_14615_, _14614_, _14613_);
  and _46750_ (_14616_, _14615_, _01954_);
  and _46751_ (_14617_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _46752_ (_14618_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _46753_ (_14619_, _14618_, _14617_);
  and _46754_ (_14620_, _14619_, _02150_);
  or _46755_ (_14621_, _14620_, _14616_);
  or _46756_ (_14622_, _14621_, _02144_);
  and _46757_ (_14623_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _46758_ (_14624_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _46759_ (_14625_, _14624_, _14623_);
  and _46760_ (_14626_, _14625_, _01954_);
  and _46761_ (_14627_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and _46762_ (_14628_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _46763_ (_14629_, _14628_, _14627_);
  and _46764_ (_14630_, _14629_, _02150_);
  or _46765_ (_14631_, _14630_, _14626_);
  or _46766_ (_14632_, _14631_, _02131_);
  and _46767_ (_14633_, _14632_, _02157_);
  and _46768_ (_14634_, _14633_, _14622_);
  or _46769_ (_14635_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _46770_ (_14636_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _46771_ (_14637_, _14636_, _02150_);
  and _46772_ (_14638_, _14637_, _14635_);
  or _46773_ (_14639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _46774_ (_14640_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _46775_ (_14641_, _14640_, _01954_);
  and _46776_ (_14642_, _14641_, _14639_);
  or _46777_ (_14643_, _14642_, _14638_);
  or _46778_ (_14644_, _14643_, _02144_);
  or _46779_ (_14645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _46780_ (_14646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _46781_ (_14647_, _14646_, _02150_);
  and _46782_ (_14648_, _14647_, _14645_);
  or _46783_ (_14649_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _46784_ (_14650_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _46785_ (_14651_, _14650_, _01954_);
  and _46786_ (_14652_, _14651_, _14649_);
  or _46787_ (_14653_, _14652_, _14648_);
  or _46788_ (_14654_, _14653_, _02131_);
  and _46789_ (_14655_, _14654_, _02077_);
  and _46790_ (_14656_, _14655_, _14644_);
  or _46791_ (_14657_, _14656_, _14634_);
  and _46792_ (_14658_, _14657_, _02194_);
  and _46793_ (_14659_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _46794_ (_14660_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _46795_ (_14661_, _14660_, _14659_);
  and _46796_ (_14662_, _14661_, _01954_);
  and _46797_ (_14663_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _46798_ (_14664_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _46799_ (_14665_, _14664_, _14663_);
  and _46800_ (_14666_, _14665_, _02150_);
  or _46801_ (_14667_, _14666_, _14662_);
  or _46802_ (_14668_, _14667_, _02144_);
  and _46803_ (_14669_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _46804_ (_14670_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _46805_ (_14671_, _14670_, _14669_);
  and _46806_ (_14672_, _14671_, _01954_);
  and _46807_ (_14673_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _46808_ (_14674_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _46809_ (_14675_, _14674_, _14673_);
  and _46810_ (_14676_, _14675_, _02150_);
  or _46811_ (_14677_, _14676_, _14672_);
  or _46812_ (_14678_, _14677_, _02131_);
  and _46813_ (_14679_, _14678_, _02157_);
  and _46814_ (_14680_, _14679_, _14668_);
  or _46815_ (_14681_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _46816_ (_14682_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _46817_ (_14683_, _14682_, _14681_);
  and _46818_ (_14684_, _14683_, _01954_);
  or _46819_ (_14685_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _46820_ (_14686_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _46821_ (_14687_, _14686_, _14685_);
  and _46822_ (_14688_, _14687_, _02150_);
  or _46823_ (_14689_, _14688_, _14684_);
  or _46824_ (_14690_, _14689_, _02144_);
  or _46825_ (_14691_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _46826_ (_14692_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _46827_ (_14693_, _14692_, _14691_);
  and _46828_ (_14694_, _14693_, _01954_);
  or _46829_ (_14695_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _46830_ (_14696_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _46831_ (_14697_, _14696_, _14695_);
  and _46832_ (_14698_, _14697_, _02150_);
  or _46833_ (_14699_, _14698_, _14694_);
  or _46834_ (_14700_, _14699_, _02131_);
  and _46835_ (_14701_, _14700_, _02077_);
  and _46836_ (_14702_, _14701_, _14690_);
  or _46837_ (_14703_, _14702_, _14680_);
  and _46838_ (_14704_, _14703_, _02065_);
  or _46839_ (_14705_, _14704_, _14658_);
  and _46840_ (_14706_, _14705_, _02143_);
  or _46841_ (_14707_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _46842_ (_14708_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _46843_ (_14709_, _14708_, _14707_);
  and _46844_ (_14710_, _14709_, _01954_);
  or _46845_ (_14711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _46846_ (_14712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and _46847_ (_14713_, _14712_, _14711_);
  and _46848_ (_14714_, _14713_, _02150_);
  or _46849_ (_14715_, _14714_, _14710_);
  and _46850_ (_14716_, _14715_, _02144_);
  or _46851_ (_14717_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _46852_ (_14718_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _46853_ (_14719_, _14718_, _14717_);
  and _46854_ (_14720_, _14719_, _01954_);
  or _46855_ (_14721_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _46856_ (_14722_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _46857_ (_14723_, _14722_, _14721_);
  and _46858_ (_14724_, _14723_, _02150_);
  or _46859_ (_14725_, _14724_, _14720_);
  and _46860_ (_14726_, _14725_, _02131_);
  or _46861_ (_14727_, _14726_, _14716_);
  and _46862_ (_14728_, _14727_, _02077_);
  and _46863_ (_14729_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _46864_ (_14730_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _46865_ (_14731_, _14730_, _14729_);
  and _46866_ (_14732_, _14731_, _01954_);
  and _46867_ (_14733_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _46868_ (_14734_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _46869_ (_14735_, _14734_, _14733_);
  and _46870_ (_14736_, _14735_, _02150_);
  or _46871_ (_14737_, _14736_, _14732_);
  and _46872_ (_14738_, _14737_, _02144_);
  and _46873_ (_14739_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _46874_ (_14740_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _46875_ (_14741_, _14740_, _14739_);
  and _46876_ (_14742_, _14741_, _01954_);
  and _46877_ (_14743_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and _46878_ (_14744_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _46879_ (_14745_, _14744_, _14743_);
  and _46880_ (_14746_, _14745_, _02150_);
  or _46881_ (_14747_, _14746_, _14742_);
  and _46882_ (_14748_, _14747_, _02131_);
  or _46883_ (_14749_, _14748_, _14738_);
  and _46884_ (_14750_, _14749_, _02157_);
  or _46885_ (_14751_, _14750_, _14728_);
  and _46886_ (_14752_, _14751_, _02065_);
  or _46887_ (_14753_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _46888_ (_14754_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _46889_ (_14755_, _14754_, _02150_);
  and _46890_ (_14756_, _14755_, _14753_);
  or _46891_ (_14757_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _46892_ (_14758_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _46893_ (_14759_, _14758_, _01954_);
  and _46894_ (_14760_, _14759_, _14757_);
  or _46895_ (_14761_, _14760_, _14756_);
  and _46896_ (_14762_, _14761_, _02144_);
  or _46897_ (_14763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _46898_ (_14764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _46899_ (_14765_, _14764_, _02150_);
  and _46900_ (_14766_, _14765_, _14763_);
  or _46901_ (_14767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _46902_ (_14768_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _46903_ (_14769_, _14768_, _01954_);
  and _46904_ (_14770_, _14769_, _14767_);
  or _46905_ (_14771_, _14770_, _14766_);
  and _46906_ (_14772_, _14771_, _02131_);
  or _46907_ (_14773_, _14772_, _14762_);
  and _46908_ (_14774_, _14773_, _02077_);
  and _46909_ (_14775_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _46910_ (_14776_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _46911_ (_14777_, _14776_, _14775_);
  and _46912_ (_14778_, _14777_, _01954_);
  and _46913_ (_14779_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _46914_ (_14780_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _46915_ (_14781_, _14780_, _14779_);
  and _46916_ (_14782_, _14781_, _02150_);
  or _46917_ (_14783_, _14782_, _14778_);
  and _46918_ (_14784_, _14783_, _02144_);
  and _46919_ (_14785_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _46920_ (_14786_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _46921_ (_14787_, _14786_, _14785_);
  and _46922_ (_14788_, _14787_, _01954_);
  and _46923_ (_14789_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _46924_ (_14790_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _46925_ (_14791_, _14790_, _14789_);
  and _46926_ (_14792_, _14791_, _02150_);
  or _46927_ (_14793_, _14792_, _14788_);
  and _46928_ (_14794_, _14793_, _02131_);
  or _46929_ (_14795_, _14794_, _14784_);
  and _46930_ (_14796_, _14795_, _02157_);
  or _46931_ (_14797_, _14796_, _14774_);
  and _46932_ (_14798_, _14797_, _02194_);
  or _46933_ (_14799_, _14798_, _14752_);
  and _46934_ (_14800_, _14799_, _02005_);
  or _46935_ (_14801_, _14800_, _14706_);
  or _46936_ (_14802_, _14801_, _02374_);
  and _46937_ (_14803_, _14802_, _14612_);
  or _46938_ (_14804_, _14803_, _02142_);
  and _46939_ (_14805_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _46940_ (_14806_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _46941_ (_14807_, _14806_, _14805_);
  and _46942_ (_14808_, _14807_, _01954_);
  and _46943_ (_14809_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _46944_ (_14810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _46945_ (_14811_, _14810_, _14809_);
  and _46946_ (_14812_, _14811_, _02150_);
  or _46947_ (_14813_, _14812_, _14808_);
  or _46948_ (_14814_, _14813_, _02144_);
  and _46949_ (_14815_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _46950_ (_14816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _46951_ (_14817_, _14816_, _14815_);
  and _46952_ (_14818_, _14817_, _01954_);
  and _46953_ (_14819_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _46954_ (_14820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _46955_ (_14821_, _14820_, _14819_);
  and _46956_ (_14822_, _14821_, _02150_);
  or _46957_ (_14823_, _14822_, _14818_);
  or _46958_ (_14824_, _14823_, _02131_);
  and _46959_ (_14825_, _14824_, _02157_);
  and _46960_ (_14826_, _14825_, _14814_);
  or _46961_ (_14827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _46962_ (_14828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _46963_ (_14829_, _14828_, _14827_);
  and _46964_ (_14830_, _14829_, _01954_);
  or _46965_ (_14831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _46966_ (_14832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _46967_ (_14833_, _14832_, _14831_);
  and _46968_ (_14834_, _14833_, _02150_);
  or _46969_ (_14835_, _14834_, _14830_);
  or _46970_ (_14836_, _14835_, _02144_);
  or _46971_ (_14837_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _46972_ (_14838_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _46973_ (_14839_, _14838_, _14837_);
  and _46974_ (_14840_, _14839_, _01954_);
  or _46975_ (_14841_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _46976_ (_14842_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _46977_ (_14843_, _14842_, _14841_);
  and _46978_ (_14844_, _14843_, _02150_);
  or _46979_ (_14845_, _14844_, _14840_);
  or _46980_ (_14846_, _14845_, _02131_);
  and _46981_ (_14847_, _14846_, _02077_);
  and _46982_ (_14848_, _14847_, _14836_);
  or _46983_ (_14849_, _14848_, _14826_);
  and _46984_ (_14850_, _14849_, _02065_);
  and _46985_ (_14851_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _46986_ (_14852_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _46987_ (_14853_, _14852_, _14851_);
  and _46988_ (_14854_, _14853_, _01954_);
  and _46989_ (_14855_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _46990_ (_14856_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _46991_ (_14857_, _14856_, _14855_);
  and _46992_ (_14858_, _14857_, _02150_);
  or _46993_ (_14859_, _14858_, _14854_);
  or _46994_ (_14860_, _14859_, _02144_);
  and _46995_ (_14861_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _46996_ (_14862_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _46997_ (_14863_, _14862_, _14861_);
  and _46998_ (_14864_, _14863_, _01954_);
  and _46999_ (_14865_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _47000_ (_14866_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _47001_ (_14867_, _14866_, _14865_);
  and _47002_ (_14868_, _14867_, _02150_);
  or _47003_ (_14869_, _14868_, _14864_);
  or _47004_ (_14870_, _14869_, _02131_);
  and _47005_ (_14871_, _14870_, _02157_);
  and _47006_ (_14872_, _14871_, _14860_);
  or _47007_ (_14873_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _47008_ (_14874_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _47009_ (_14875_, _14874_, _02150_);
  and _47010_ (_14876_, _14875_, _14873_);
  or _47011_ (_14877_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _47012_ (_14878_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _47013_ (_14879_, _14878_, _01954_);
  and _47014_ (_14880_, _14879_, _14877_);
  or _47015_ (_14881_, _14880_, _14876_);
  or _47016_ (_14882_, _14881_, _02144_);
  or _47017_ (_14883_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _47018_ (_14884_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _47019_ (_14885_, _14884_, _02150_);
  and _47020_ (_14886_, _14885_, _14883_);
  or _47021_ (_14887_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _47022_ (_14888_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _47023_ (_14889_, _14888_, _01954_);
  and _47024_ (_14890_, _14889_, _14887_);
  or _47025_ (_14891_, _14890_, _14886_);
  or _47026_ (_14892_, _14891_, _02131_);
  and _47027_ (_14893_, _14892_, _02077_);
  and _47028_ (_14894_, _14893_, _14882_);
  or _47029_ (_14895_, _14894_, _14872_);
  and _47030_ (_14896_, _14895_, _02194_);
  or _47031_ (_14897_, _14896_, _14850_);
  and _47032_ (_14898_, _14897_, _02143_);
  and _47033_ (_14899_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _47034_ (_14900_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _47035_ (_14901_, _14900_, _14899_);
  and _47036_ (_14902_, _14901_, _01954_);
  and _47037_ (_14903_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _47038_ (_14904_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _47039_ (_14905_, _14904_, _14903_);
  and _47040_ (_14906_, _14905_, _02150_);
  or _47041_ (_14907_, _14906_, _14902_);
  and _47042_ (_14908_, _14907_, _02131_);
  and _47043_ (_14909_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _47044_ (_14910_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _47045_ (_14911_, _14910_, _14909_);
  and _47046_ (_14912_, _14911_, _01954_);
  and _47047_ (_14913_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _47048_ (_14914_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _47049_ (_14915_, _14914_, _14913_);
  and _47050_ (_14916_, _14915_, _02150_);
  or _47051_ (_14917_, _14916_, _14912_);
  and _47052_ (_14918_, _14917_, _02144_);
  or _47053_ (_14919_, _14918_, _14908_);
  and _47054_ (_14920_, _14919_, _02157_);
  or _47055_ (_14921_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _47056_ (_14922_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _47057_ (_14923_, _14922_, _02150_);
  and _47058_ (_14924_, _14923_, _14921_);
  or _47059_ (_14925_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _47060_ (_14926_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _47061_ (_14927_, _14926_, _01954_);
  and _47062_ (_14928_, _14927_, _14925_);
  or _47063_ (_14929_, _14928_, _14924_);
  and _47064_ (_14930_, _14929_, _02131_);
  or _47065_ (_14931_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _47066_ (_14932_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _47067_ (_14933_, _14932_, _02150_);
  and _47068_ (_14934_, _14933_, _14931_);
  or _47069_ (_14935_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _47070_ (_14936_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _47071_ (_14937_, _14936_, _01954_);
  and _47072_ (_14938_, _14937_, _14935_);
  or _47073_ (_14939_, _14938_, _14934_);
  and _47074_ (_14940_, _14939_, _02144_);
  or _47075_ (_14941_, _14940_, _14930_);
  and _47076_ (_14942_, _14941_, _02077_);
  or _47077_ (_14943_, _14942_, _14920_);
  and _47078_ (_14944_, _14943_, _02194_);
  and _47079_ (_14945_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _47080_ (_14946_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _47081_ (_14947_, _14946_, _14945_);
  and _47082_ (_14948_, _14947_, _01954_);
  and _47083_ (_14949_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _47084_ (_14950_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _47085_ (_14951_, _14950_, _14949_);
  and _47086_ (_14952_, _14951_, _02150_);
  or _47087_ (_14953_, _14952_, _14948_);
  and _47088_ (_14954_, _14953_, _02131_);
  and _47089_ (_14955_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _47090_ (_14956_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _47091_ (_14957_, _14956_, _14955_);
  and _47092_ (_14958_, _14957_, _01954_);
  and _47093_ (_14959_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _47094_ (_14960_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _47095_ (_14961_, _14960_, _14959_);
  and _47096_ (_14962_, _14961_, _02150_);
  or _47097_ (_14963_, _14962_, _14958_);
  and _47098_ (_14964_, _14963_, _02144_);
  or _47099_ (_14965_, _14964_, _14954_);
  and _47100_ (_14966_, _14965_, _02157_);
  or _47101_ (_14967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _47102_ (_14968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _47103_ (_14969_, _14968_, _14967_);
  and _47104_ (_14970_, _14969_, _01954_);
  or _47105_ (_14971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _47106_ (_14972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _47107_ (_14973_, _14972_, _14971_);
  and _47108_ (_14974_, _14973_, _02150_);
  or _47109_ (_14975_, _14974_, _14970_);
  and _47110_ (_14976_, _14975_, _02131_);
  or _47111_ (_14977_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _47112_ (_14978_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _47113_ (_14979_, _14978_, _14977_);
  and _47114_ (_14980_, _14979_, _01954_);
  or _47115_ (_14981_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _47116_ (_14982_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _47117_ (_14983_, _14982_, _14981_);
  and _47118_ (_14984_, _14983_, _02150_);
  or _47119_ (_14985_, _14984_, _14980_);
  and _47120_ (_14986_, _14985_, _02144_);
  or _47121_ (_14987_, _14986_, _14976_);
  and _47122_ (_14988_, _14987_, _02077_);
  or _47123_ (_14989_, _14988_, _14966_);
  and _47124_ (_14990_, _14989_, _02065_);
  or _47125_ (_14991_, _14990_, _14944_);
  and _47126_ (_14992_, _14991_, _02005_);
  or _47127_ (_14993_, _14992_, _14898_);
  or _47128_ (_14994_, _14993_, _02054_);
  and _47129_ (_14995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _47130_ (_14996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _47131_ (_14997_, _14996_, _14995_);
  and _47132_ (_14998_, _14997_, _01954_);
  and _47133_ (_14999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and _47134_ (_15000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _47135_ (_15001_, _15000_, _14999_);
  and _47136_ (_15002_, _15001_, _02150_);
  or _47137_ (_15003_, _15002_, _14998_);
  or _47138_ (_15004_, _15003_, _02144_);
  and _47139_ (_15005_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _47140_ (_15006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _47141_ (_15007_, _15006_, _15005_);
  and _47142_ (_15008_, _15007_, _01954_);
  and _47143_ (_15009_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _47144_ (_15010_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _47145_ (_15011_, _15010_, _15009_);
  and _47146_ (_15012_, _15011_, _02150_);
  or _47147_ (_15013_, _15012_, _15008_);
  or _47148_ (_15014_, _15013_, _02131_);
  and _47149_ (_15015_, _15014_, _02157_);
  and _47150_ (_15016_, _15015_, _15004_);
  or _47151_ (_15017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _47152_ (_15018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _47153_ (_15019_, _15018_, _02150_);
  and _47154_ (_15020_, _15019_, _15017_);
  or _47155_ (_15021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _47156_ (_15022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _47157_ (_15023_, _15022_, _01954_);
  and _47158_ (_15024_, _15023_, _15021_);
  or _47159_ (_15025_, _15024_, _15020_);
  or _47160_ (_15026_, _15025_, _02144_);
  or _47161_ (_15027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _47162_ (_15028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _47163_ (_15029_, _15028_, _02150_);
  and _47164_ (_15030_, _15029_, _15027_);
  or _47165_ (_15031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _47166_ (_15032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _47167_ (_15033_, _15032_, _01954_);
  and _47168_ (_15034_, _15033_, _15031_);
  or _47169_ (_15035_, _15034_, _15030_);
  or _47170_ (_15036_, _15035_, _02131_);
  and _47171_ (_15037_, _15036_, _02077_);
  and _47172_ (_15038_, _15037_, _15026_);
  or _47173_ (_15039_, _15038_, _15016_);
  and _47174_ (_15040_, _15039_, _02194_);
  and _47175_ (_15041_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _47176_ (_15042_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _47177_ (_15043_, _15042_, _15041_);
  and _47178_ (_15044_, _15043_, _01954_);
  and _47179_ (_15045_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _47180_ (_15046_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _47181_ (_15047_, _15046_, _15045_);
  and _47182_ (_15048_, _15047_, _02150_);
  or _47183_ (_15049_, _15048_, _15044_);
  or _47184_ (_15050_, _15049_, _02144_);
  and _47185_ (_15051_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _47186_ (_15052_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _47187_ (_15053_, _15052_, _15051_);
  and _47188_ (_15054_, _15053_, _01954_);
  and _47189_ (_15055_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _47190_ (_15056_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _47191_ (_15057_, _15056_, _15055_);
  and _47192_ (_15058_, _15057_, _02150_);
  or _47193_ (_15059_, _15058_, _15054_);
  or _47194_ (_15060_, _15059_, _02131_);
  and _47195_ (_15061_, _15060_, _02157_);
  and _47196_ (_15062_, _15061_, _15050_);
  or _47197_ (_15063_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _47198_ (_15064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _47199_ (_15065_, _15064_, _15063_);
  and _47200_ (_15066_, _15065_, _01954_);
  or _47201_ (_15067_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _47202_ (_15068_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _47203_ (_15069_, _15068_, _15067_);
  and _47204_ (_15070_, _15069_, _02150_);
  or _47205_ (_15071_, _15070_, _15066_);
  or _47206_ (_15072_, _15071_, _02144_);
  or _47207_ (_15073_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _47208_ (_15074_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _47209_ (_15075_, _15074_, _15073_);
  and _47210_ (_15076_, _15075_, _01954_);
  or _47211_ (_15077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _47212_ (_15078_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _47213_ (_15079_, _15078_, _15077_);
  and _47214_ (_15080_, _15079_, _02150_);
  or _47215_ (_15081_, _15080_, _15076_);
  or _47216_ (_15082_, _15081_, _02131_);
  and _47217_ (_15083_, _15082_, _02077_);
  and _47218_ (_15084_, _15083_, _15072_);
  or _47219_ (_15085_, _15084_, _15062_);
  and _47220_ (_15086_, _15085_, _02065_);
  or _47221_ (_15087_, _15086_, _15040_);
  and _47222_ (_15088_, _15087_, _02143_);
  or _47223_ (_15089_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _47224_ (_15090_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _47225_ (_15091_, _15090_, _15089_);
  and _47226_ (_15092_, _15091_, _01954_);
  or _47227_ (_15093_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _47228_ (_15094_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _47229_ (_15095_, _15094_, _15093_);
  and _47230_ (_15096_, _15095_, _02150_);
  or _47231_ (_15097_, _15096_, _15092_);
  and _47232_ (_15098_, _15097_, _02144_);
  or _47233_ (_15099_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _47234_ (_15100_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _47235_ (_15101_, _15100_, _15099_);
  and _47236_ (_15102_, _15101_, _01954_);
  or _47237_ (_15103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _47238_ (_15104_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _47239_ (_15105_, _15104_, _15103_);
  and _47240_ (_15106_, _15105_, _02150_);
  or _47241_ (_15107_, _15106_, _15102_);
  and _47242_ (_15108_, _15107_, _02131_);
  or _47243_ (_15109_, _15108_, _15098_);
  and _47244_ (_15110_, _15109_, _02077_);
  and _47245_ (_15111_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _47246_ (_15112_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _47247_ (_15113_, _15112_, _15111_);
  and _47248_ (_15114_, _15113_, _01954_);
  and _47249_ (_15115_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _47250_ (_15116_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _47251_ (_15117_, _15116_, _15115_);
  and _47252_ (_15118_, _15117_, _02150_);
  or _47253_ (_15119_, _15118_, _15114_);
  and _47254_ (_15120_, _15119_, _02144_);
  and _47255_ (_15121_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _47256_ (_15122_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _47257_ (_15123_, _15122_, _15121_);
  and _47258_ (_15124_, _15123_, _01954_);
  and _47259_ (_15125_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _47260_ (_15126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _47261_ (_15127_, _15126_, _15125_);
  and _47262_ (_15128_, _15127_, _02150_);
  or _47263_ (_15129_, _15128_, _15124_);
  and _47264_ (_15130_, _15129_, _02131_);
  or _47265_ (_15131_, _15130_, _15120_);
  and _47266_ (_15132_, _15131_, _02157_);
  or _47267_ (_15133_, _15132_, _15110_);
  and _47268_ (_15134_, _15133_, _02065_);
  or _47269_ (_15135_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _47270_ (_15136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _47271_ (_15137_, _15136_, _02150_);
  and _47272_ (_15138_, _15137_, _15135_);
  or _47273_ (_15139_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _47274_ (_15140_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _47275_ (_15141_, _15140_, _01954_);
  and _47276_ (_15142_, _15141_, _15139_);
  or _47277_ (_15143_, _15142_, _15138_);
  and _47278_ (_15144_, _15143_, _02144_);
  or _47279_ (_15145_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _47280_ (_15146_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _47281_ (_15147_, _15146_, _02150_);
  and _47282_ (_15148_, _15147_, _15145_);
  or _47283_ (_15149_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _47284_ (_15150_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _47285_ (_15151_, _15150_, _01954_);
  and _47286_ (_15152_, _15151_, _15149_);
  or _47287_ (_15153_, _15152_, _15148_);
  and _47288_ (_15154_, _15153_, _02131_);
  or _47289_ (_15155_, _15154_, _15144_);
  and _47290_ (_15156_, _15155_, _02077_);
  and _47291_ (_15157_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _47292_ (_15158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _47293_ (_15159_, _15158_, _15157_);
  and _47294_ (_15160_, _15159_, _01954_);
  and _47295_ (_15161_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _47296_ (_15162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _47297_ (_15163_, _15162_, _15161_);
  and _47298_ (_15164_, _15163_, _02150_);
  or _47299_ (_15165_, _15164_, _15160_);
  and _47300_ (_15166_, _15165_, _02144_);
  and _47301_ (_15167_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _47302_ (_15168_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _47303_ (_15169_, _15168_, _15167_);
  and _47304_ (_15170_, _15169_, _01954_);
  and _47305_ (_15171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _47306_ (_15172_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _47307_ (_15173_, _15172_, _15171_);
  and _47308_ (_15174_, _15173_, _02150_);
  or _47309_ (_15175_, _15174_, _15170_);
  and _47310_ (_15176_, _15175_, _02131_);
  or _47311_ (_15177_, _15176_, _15166_);
  and _47312_ (_15178_, _15177_, _02157_);
  or _47313_ (_15179_, _15178_, _15156_);
  and _47314_ (_15180_, _15179_, _02194_);
  or _47315_ (_15181_, _15180_, _15134_);
  and _47316_ (_15182_, _15181_, _02005_);
  or _47317_ (_15183_, _15182_, _15088_);
  or _47318_ (_15184_, _15183_, _02374_);
  and _47319_ (_15185_, _15184_, _14994_);
  or _47320_ (_15186_, _15185_, _01748_);
  and _47321_ (_15187_, _15186_, _14804_);
  or _47322_ (_15188_, _15187_, _02141_);
  or _47323_ (_15189_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _47324_ (_15190_, _15189_, _27355_);
  and _47325_ (_15248_, _15190_, _15188_);
  and _47326_ (pc_log_change, _25988_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  nor _47327_ (_18890_, _26452_, rst);
  and _47328_ (_15191_, _26350_, _26286_);
  and _47329_ (_15192_, _15191_, _26269_);
  not _47330_ (_15193_, _15192_);
  and _47331_ (_15194_, _26335_, _26413_);
  and _47332_ (_15195_, _26351_, _26155_);
  nor _47333_ (_15196_, _15195_, _15194_);
  and _47334_ (_15197_, _15196_, _15193_);
  and _47335_ (_15198_, _26350_, _26181_);
  or _47336_ (_15199_, _26286_, _26155_);
  nand _47337_ (_15200_, _15199_, _15198_);
  and _47338_ (_15201_, _15200_, _15197_);
  and _47339_ (_15202_, _25987_, _27355_);
  not _47340_ (_15203_, _15202_);
  or _47341_ (_15204_, _15203_, _15194_);
  or _47342_ (_18893_, _15204_, _15201_);
  not _47343_ (_15205_, _26121_);
  nor _47344_ (_15206_, _15205_, _26079_);
  and _47345_ (_15207_, _15206_, _26149_);
  and _47346_ (_15208_, _15207_, _26028_);
  nor _47347_ (_15209_, _26259_, _26204_);
  not _47348_ (_15210_, _26177_);
  nor _47349_ (_15211_, _26232_, _15210_);
  and _47350_ (_15212_, _15211_, _15209_);
  and _47351_ (_15213_, _15212_, _15208_);
  and _47352_ (_15214_, _26232_, _26177_);
  and _47353_ (_15215_, _26259_, _26204_);
  and _47354_ (_15216_, _15215_, _15214_);
  and _47355_ (_15217_, _15216_, _15207_);
  nor _47356_ (_15218_, _26149_, _26079_);
  and _47357_ (_15219_, _15218_, _15205_);
  not _47358_ (_15220_, _26204_);
  nor _47359_ (_15221_, _26259_, _15220_);
  and _47360_ (_15223_, _15221_, _15214_);
  and _47361_ (_15224_, _15223_, _15219_);
  and _47362_ (_15225_, _26149_, _15205_);
  or _47363_ (_15226_, _15225_, _26079_);
  and _47364_ (_15227_, _15226_, _15223_);
  or _47365_ (_15228_, _15227_, _15224_);
  or _47366_ (_15229_, _15228_, _15217_);
  or _47367_ (_15230_, _15229_, _15213_);
  not _47368_ (_15231_, _26232_);
  and _47369_ (_15232_, _15209_, _15231_);
  and _47370_ (_15233_, _15232_, _15208_);
  and _47371_ (_15234_, _15233_, _15210_);
  and _47372_ (_15235_, _15209_, _26232_);
  and _47373_ (_15237_, _15235_, _15208_);
  and _47374_ (_15239_, _15221_, _15231_);
  not _47375_ (_15241_, _26028_);
  and _47376_ (_15243_, _15207_, _15241_);
  and _47377_ (_15245_, _15243_, _15239_);
  or _47378_ (_15247_, _15245_, _15237_);
  or _47379_ (_15249_, _15247_, _15234_);
  or _47380_ (_15250_, _15249_, _15230_);
  and _47381_ (_15251_, _26232_, _15210_);
  and _47382_ (_15252_, _26259_, _15220_);
  and _47383_ (_15253_, _15252_, _15251_);
  nor _47384_ (_15254_, _15253_, _15241_);
  not _47385_ (_15255_, _26149_);
  and _47386_ (_15256_, _15206_, _15255_);
  not _47387_ (_15257_, _15256_);
  nor _47388_ (_15258_, _15257_, _15254_);
  not _47389_ (_15259_, _15258_);
  and _47390_ (_15260_, _15214_, _15209_);
  and _47391_ (_15261_, _15255_, _26028_);
  and _47392_ (_15262_, _15261_, _15206_);
  and _47393_ (_15263_, _15262_, _15260_);
  nor _47394_ (_15264_, _26232_, _26177_);
  and _47395_ (_15265_, _15252_, _15264_);
  and _47396_ (_15266_, _15265_, _15262_);
  nor _47397_ (_15267_, _15266_, _15263_);
  and _47398_ (_15268_, _15267_, _15259_);
  and _47399_ (_15269_, _15252_, _15214_);
  and _47400_ (_15270_, _15269_, _15243_);
  and _47401_ (_15271_, _15215_, _15211_);
  and _47402_ (_15272_, _15219_, _15241_);
  and _47403_ (_15273_, _15272_, _15271_);
  or _47404_ (_15274_, _15273_, _15270_);
  and _47405_ (_15275_, _15252_, _26177_);
  and _47406_ (_15276_, _15275_, _15262_);
  and _47407_ (_15277_, _15215_, _26232_);
  and _47408_ (_15278_, _15262_, _15277_);
  or _47409_ (_15279_, _15278_, _15276_);
  or _47410_ (_15280_, _15279_, _15274_);
  and _47411_ (_15281_, _15251_, _15209_);
  or _47412_ (_15282_, _15281_, _15212_);
  and _47413_ (_15283_, _15282_, _15262_);
  and _47414_ (_15284_, _15271_, _26079_);
  and _47415_ (_15285_, _15251_, _15215_);
  and _47416_ (_15286_, _15285_, _15207_);
  or _47417_ (_15287_, _15286_, _15284_);
  or _47418_ (_15288_, _15287_, _15283_);
  and _47419_ (_15289_, _15219_, _26028_);
  and _47420_ (_15290_, _15221_, _15210_);
  and _47421_ (_15291_, _15290_, _15289_);
  and _47422_ (_15292_, _15264_, _15221_);
  and _47423_ (_15293_, _15262_, _15292_);
  or _47424_ (_15294_, _15293_, _15291_);
  or _47425_ (_15295_, _15294_, _15288_);
  nor _47426_ (_15296_, _15295_, _15280_);
  nand _47427_ (_15297_, _15296_, _15268_);
  or _47428_ (_15298_, _15297_, _15250_);
  and _47429_ (_15299_, _15298_, _25988_);
  not _47430_ (_15300_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _47431_ (_15301_, _25986_, _23914_);
  and _47432_ (_15302_, _15301_, _26370_);
  nor _47433_ (_15303_, _15302_, _15300_);
  or _47434_ (_15304_, _15303_, rst);
  or _47435_ (_18896_, _15304_, _15299_);
  not _47436_ (_15305_, _25982_);
  or _47437_ (_15306_, _26204_, _15305_);
  or _47438_ (_15307_, _25982_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _47439_ (_15308_, _15307_, _27355_);
  and _47440_ (_18899_, _15308_, _15306_);
  and _47441_ (_15309_, \oc8051_top_1.oc8051_sfr1.wait_data , _27355_);
  and _47442_ (_15310_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _47443_ (_15311_, _26272_, _26413_);
  or _47444_ (_15312_, _26306_, _26274_);
  or _47445_ (_15313_, _15312_, _15311_);
  and _47446_ (_15314_, _26438_, _26351_);
  and _47447_ (_15315_, _15194_, _26269_);
  or _47448_ (_15316_, _15315_, _15314_);
  and _47449_ (_15317_, _26336_, _26286_);
  nor _47450_ (_15318_, _15317_, _26375_);
  not _47451_ (_15319_, _15318_);
  or _47452_ (_15320_, _15319_, _15316_);
  or _47453_ (_15321_, _15320_, _15313_);
  or _47454_ (_15322_, _15321_, _26318_);
  and _47455_ (_15323_, _15322_, _15202_);
  or _47456_ (_18902_, _15323_, _15310_);
  and _47457_ (_15324_, _26359_, _26286_);
  or _47458_ (_15325_, _15324_, _26414_);
  nor _47459_ (_15326_, _26181_, _26087_);
  and _47460_ (_15327_, _15326_, _26271_);
  or _47461_ (_15328_, _15327_, _26405_);
  and _47462_ (_15329_, _26277_, _26278_);
  and _47463_ (_15330_, _15329_, _26272_);
  or _47464_ (_15331_, _15330_, _15328_);
  or _47465_ (_15332_, _15331_, _15325_);
  and _47466_ (_15333_, _15332_, _25987_);
  and _47467_ (_15334_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47468_ (_15335_, _26382_, _15300_);
  not _47469_ (_15336_, _26441_);
  and _47470_ (_15337_, _15336_, _15335_);
  or _47471_ (_15338_, _15337_, _15334_);
  or _47472_ (_15339_, _15338_, _15333_);
  and _47473_ (_18905_, _15339_, _27355_);
  and _47474_ (_15340_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _47475_ (_15341_, _26438_, _26320_);
  not _47476_ (_15342_, _26280_);
  nor _47477_ (_15343_, _26320_, _26289_);
  nor _47478_ (_15344_, _15343_, _15342_);
  or _47479_ (_15345_, _15344_, _15341_);
  and _47480_ (_15346_, _15329_, _26294_);
  or _47481_ (_15347_, _15346_, _15345_);
  not _47482_ (_15348_, _26400_);
  nor _47483_ (_15349_, _15343_, _26087_);
  nor _47484_ (_15350_, _26269_, _26087_);
  and _47485_ (_15351_, _15350_, _26293_);
  or _47486_ (_15352_, _15351_, _15349_);
  or _47487_ (_15353_, _15352_, _15348_);
  and _47488_ (_15354_, _26438_, _26362_);
  and _47489_ (_15355_, _15350_, _26265_);
  or _47490_ (_15356_, _15355_, _15325_);
  or _47491_ (_15357_, _15356_, _15354_);
  or _47492_ (_15358_, _15357_, _15353_);
  or _47493_ (_15359_, _15358_, _15347_);
  and _47494_ (_15360_, _15359_, _15202_);
  or _47495_ (_18908_, _15360_, _15340_);
  and _47496_ (_15361_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47497_ (_15362_, _26357_, _25987_);
  or _47498_ (_15363_, _15362_, _15361_);
  or _47499_ (_15364_, _15363_, _15337_);
  and _47500_ (_18911_, _15364_, _27355_);
  not _47501_ (_15365_, _15197_);
  and _47502_ (_15366_, _15365_, _15335_);
  or _47503_ (_15367_, _15366_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47504_ (_15368_, _26279_, _26284_);
  and _47505_ (_15369_, _15368_, _26181_);
  and _47506_ (_15370_, _26087_, _26034_);
  and _47507_ (_15371_, _15370_, _26154_);
  and _47508_ (_15372_, _26294_, _15371_);
  or _47509_ (_15373_, _15372_, _15369_);
  and _47510_ (_15374_, _15373_, _26372_);
  or _47511_ (_15375_, _15374_, _25983_);
  and _47512_ (_15376_, _26293_, _26273_);
  nor _47513_ (_15377_, _15376_, _15368_);
  nor _47514_ (_15378_, _15377_, _26269_);
  or _47515_ (_15379_, _15378_, _15315_);
  and _47516_ (_15380_, _15379_, _15375_);
  or _47517_ (_15381_, _15380_, _15367_);
  or _47518_ (_15382_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _23914_);
  and _47519_ (_15383_, _15382_, _27355_);
  and _47520_ (_18914_, _15383_, _15381_);
  and _47521_ (_15384_, _15309_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _47522_ (_15385_, _15327_, _26348_);
  or _47523_ (_15386_, _26309_, _26306_);
  or _47524_ (_15387_, _15386_, _26268_);
  or _47525_ (_15388_, _15387_, _15385_);
  and _47526_ (_15389_, _15350_, _26271_);
  or _47527_ (_15390_, _15389_, _15351_);
  or _47528_ (_15391_, _26414_, _26290_);
  or _47529_ (_15392_, _15391_, _15390_);
  and _47530_ (_15393_, _26326_, _26294_);
  and _47531_ (_15394_, _26326_, _26272_);
  or _47532_ (_15395_, _15394_, _15346_);
  or _47533_ (_15396_, _15395_, _15393_);
  or _47534_ (_15397_, _15396_, _15392_);
  or _47535_ (_15398_, _15397_, _15388_);
  and _47536_ (_15399_, _15398_, _15202_);
  or _47537_ (_18917_, _15399_, _15384_);
  and _47538_ (_15400_, _15309_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _47539_ (_15401_, _15329_, _26341_);
  and _47540_ (_15402_, _26263_, _26208_);
  and _47541_ (_15403_, _15402_, _26413_);
  or _47542_ (_15404_, _15403_, _15330_);
  or _47543_ (_15405_, _15404_, _15401_);
  or _47544_ (_15406_, _15405_, _15352_);
  not _47545_ (_15407_, _26302_);
  and _47546_ (_15408_, _26438_, _26282_);
  or _47547_ (_15409_, _15408_, _15407_);
  and _47548_ (_15410_, _26326_, _26289_);
  not _47549_ (_15411_, _26425_);
  and _47550_ (_15412_, _26327_, _26270_);
  or _47551_ (_15413_, _15412_, _15411_);
  or _47552_ (_15414_, _15413_, _15410_);
  or _47553_ (_15415_, _15414_, _15409_);
  or _47554_ (_15416_, _15415_, _15406_);
  and _47555_ (_15417_, _15326_, _26270_);
  and _47556_ (_15418_, _15326_, _26298_);
  or _47557_ (_15419_, _15418_, _15417_);
  nor _47558_ (_15420_, _26399_, _26342_);
  not _47559_ (_15421_, _15420_);
  or _47560_ (_15422_, _15421_, _26288_);
  or _47561_ (_15423_, _15422_, _15419_);
  or _47562_ (_15424_, _15423_, _15347_);
  or _47563_ (_15425_, _15424_, _15416_);
  and _47564_ (_15426_, _15425_, _15202_);
  or _47565_ (_18920_, _15426_, _15400_);
  and _47566_ (_15427_, _15350_, _26335_);
  and _47567_ (_15428_, _15329_, _26311_);
  or _47568_ (_15429_, _15428_, _26403_);
  or _47569_ (_15430_, _15429_, _15427_);
  not _47570_ (_15431_, _26407_);
  and _47571_ (_15432_, _26311_, _26322_);
  or _47572_ (_15433_, _15432_, _15431_);
  or _47573_ (_15434_, _15433_, _15430_);
  and _47574_ (_15435_, _15329_, _26359_);
  or _47575_ (_15436_, _15435_, _15434_);
  and _47576_ (_15437_, _15436_, _25987_);
  nand _47577_ (_15438_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand _47578_ (_15439_, _15438_, _26449_);
  or _47579_ (_15440_, _15439_, _15437_);
  and _47580_ (_18923_, _15440_, _27355_);
  not _47581_ (_15441_, _26361_);
  or _47582_ (_15442_, _15441_, _26344_);
  or _47583_ (_15443_, _15442_, _15344_);
  or _47584_ (_15444_, _26348_, _26307_);
  and _47585_ (_15445_, _26297_, _26181_);
  and _47586_ (_15446_, _15445_, _26280_);
  or _47587_ (_15447_, _15446_, _26301_);
  and _47588_ (_15448_, _26294_, _26273_);
  or _47589_ (_15449_, _15448_, _26295_);
  or _47590_ (_15450_, _15449_, _15447_);
  or _47591_ (_15451_, _15450_, _26275_);
  or _47592_ (_15452_, _15451_, _15444_);
  or _47593_ (_15453_, _15452_, _15443_);
  and _47594_ (_15454_, _15350_, _26297_);
  or _47595_ (_15455_, _15454_, _26323_);
  and _47596_ (_15456_, _15326_, _26335_);
  or _47597_ (_15457_, _15456_, _15369_);
  or _47598_ (_15458_, _15457_, _15328_);
  or _47599_ (_15459_, _15458_, _15455_);
  and _47600_ (_15460_, _15445_, _26326_);
  nor _47601_ (_15461_, _15460_, _26399_);
  nand _47602_ (_15462_, _15461_, _26328_);
  or _47603_ (_15463_, _26420_, _26334_);
  or _47604_ (_15464_, _15463_, _15462_);
  or _47605_ (_15465_, _15464_, _15459_);
  or _47606_ (_15466_, _15465_, _15352_);
  or _47607_ (_15467_, _15466_, _15453_);
  and _47608_ (_15468_, _15467_, _25987_);
  and _47609_ (_15469_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47610_ (_15470_, _26372_, _26316_);
  or _47611_ (_15471_, _15374_, _15337_);
  or _47612_ (_15472_, _15471_, _15470_);
  or _47613_ (_15473_, _15472_, _15469_);
  or _47614_ (_15474_, _15473_, _15468_);
  and _47615_ (_18926_, _15474_, _27355_);
  nor _47616_ (_18984_, _26434_, rst);
  and _47617_ (_18986_, _26387_, _27355_);
  or _47618_ (_18989_, _15203_, _15197_);
  nor _47619_ (_15475_, _15194_, _15191_);
  or _47620_ (_18992_, _15475_, _15203_);
  or _47621_ (_15476_, _15291_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _47622_ (_15477_, _15476_, _15247_);
  and _47623_ (_15478_, _15477_, _15302_);
  nor _47624_ (_15479_, _15301_, _26370_);
  or _47625_ (_15480_, _15479_, rst);
  or _47626_ (_18995_, _15480_, _15478_);
  nand _47627_ (_15481_, _26028_, _25982_);
  or _47628_ (_15482_, _25982_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _47629_ (_15483_, _15482_, _27355_);
  and _47630_ (_18998_, _15483_, _15481_);
  or _47631_ (_15484_, _26149_, _15305_);
  or _47632_ (_15485_, _25982_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _47633_ (_15486_, _15485_, _27355_);
  and _47634_ (_19001_, _15486_, _15484_);
  nand _47635_ (_15487_, _26121_, _25982_);
  or _47636_ (_15488_, _25982_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _47637_ (_15489_, _15488_, _27355_);
  and _47638_ (_19004_, _15489_, _15487_);
  or _47639_ (_15490_, _26079_, _15305_);
  or _47640_ (_15491_, _25982_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _47641_ (_15492_, _15491_, _27355_);
  and _47642_ (_19007_, _15492_, _15490_);
  or _47643_ (_15493_, _26177_, _15305_);
  or _47644_ (_15494_, _25982_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _47645_ (_15495_, _15494_, _27355_);
  and _47646_ (_19010_, _15495_, _15493_);
  or _47647_ (_15496_, _26232_, _15305_);
  or _47648_ (_15497_, _25982_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _47649_ (_15498_, _15497_, _27355_);
  and _47650_ (_19013_, _15498_, _15496_);
  or _47651_ (_15499_, _26259_, _15305_);
  or _47652_ (_15500_, _25982_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _47653_ (_15501_, _15500_, _27355_);
  and _47654_ (_19016_, _15501_, _15499_);
  or _47655_ (_15502_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _23914_);
  and _47656_ (_15503_, _15502_, _27355_);
  and _47657_ (_15504_, _15503_, _15367_);
  and _47658_ (_15505_, _26438_, _26294_);
  and _47659_ (_15506_, _26438_, _26289_);
  or _47660_ (_15507_, _15506_, _15505_);
  or _47661_ (_15508_, _15507_, _15341_);
  and _47662_ (_15509_, _15350_, _26281_);
  or _47663_ (_15510_, _15509_, _15432_);
  and _47664_ (_15511_, _15329_, _26282_);
  or _47665_ (_15512_, _15511_, _15324_);
  or _47666_ (_15513_, _15512_, _15510_);
  or _47667_ (_15514_, _15513_, _15508_);
  nor _47668_ (_15515_, _15418_, _15431_);
  nand _47669_ (_15516_, _15515_, _26426_);
  or _47670_ (_15517_, _15403_, _26414_);
  or _47671_ (_15518_, _15517_, _15430_);
  or _47672_ (_15519_, _15518_, _15516_);
  not _47673_ (_15520_, _15326_);
  nor _47674_ (_15521_, _26423_, _15520_);
  and _47675_ (_15522_, _15329_, _26351_);
  or _47676_ (_15523_, _15522_, _15521_);
  and _47677_ (_15524_, _15198_, _26438_);
  and _47678_ (_15525_, _26333_, _26326_);
  or _47679_ (_15526_, _15525_, _15524_);
  or _47680_ (_15527_, _15526_, _15523_);
  or _47681_ (_15528_, _15435_, _15401_);
  and _47682_ (_15529_, _26438_, _26299_);
  and _47683_ (_15530_, _15329_, _26333_);
  or _47684_ (_15531_, _15530_, _15529_);
  or _47685_ (_15532_, _15531_, _15528_);
  or _47686_ (_15533_, _15532_, _15527_);
  or _47687_ (_15534_, _15533_, _15519_);
  or _47688_ (_15535_, _15534_, _15514_);
  and _47689_ (_15536_, _15535_, _15202_);
  or _47690_ (_19019_, _15536_, _15504_);
  and _47691_ (_15537_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _47692_ (_15538_, _26438_, _26339_);
  nor _47693_ (_15539_, _15355_, _26398_);
  or _47694_ (_15540_, _26341_, _26282_);
  nand _47695_ (_15541_, _15540_, _26273_);
  nand _47696_ (_15542_, _15541_, _15539_);
  or _47697_ (_15543_, _15542_, _15538_);
  or _47698_ (_15544_, _15354_, _15316_);
  or _47699_ (_15545_, _15512_, _15419_);
  or _47700_ (_15546_, _15545_, _15544_);
  not _47701_ (_15547_, _26349_);
  and _47702_ (_15548_, _26438_, _26341_);
  or _47703_ (_15549_, _15548_, _15547_);
  or _47704_ (_15550_, _15549_, _15414_);
  or _47705_ (_15551_, _15550_, _15546_);
  or _47706_ (_15552_, _15551_, _15543_);
  and _47707_ (_15553_, _15552_, _15202_);
  or _47708_ (_23904_, _15553_, _15537_);
  or _47709_ (_15554_, _15463_, _15457_);
  or _47710_ (_15555_, _15554_, _15453_);
  and _47711_ (_15556_, _15555_, _25987_);
  and _47712_ (_15557_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47713_ (_15558_, _15557_, _15472_);
  or _47714_ (_15559_, _15558_, _15556_);
  and _47715_ (_23905_, _15559_, _27355_);
  and _47716_ (_15560_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47717_ (_15561_, _15560_, _15471_);
  and _47718_ (_15562_, _15561_, _27355_);
  and _47719_ (_15563_, _26343_, _26269_);
  or _47720_ (_15564_, _15563_, _26405_);
  or _47721_ (_15565_, _15564_, _15378_);
  or _47722_ (_15566_, _15565_, _15462_);
  and _47723_ (_15567_, _15566_, _15202_);
  or _47724_ (_23906_, _15567_, _15562_);
  and _47725_ (_15568_, _26438_, _26272_);
  or _47726_ (_15569_, _15435_, _15568_);
  or _47727_ (_15570_, _15524_, _26439_);
  and _47728_ (_15571_, _15329_, _26266_);
  or _47729_ (_15572_, _15571_, _15314_);
  or _47730_ (_15573_, _15572_, _15570_);
  or _47731_ (_15574_, _15573_, _15508_);
  or _47732_ (_15575_, _15574_, _15569_);
  or _47733_ (_15576_, _15408_, _15431_);
  or _47734_ (_15577_, _15529_, _15548_);
  or _47735_ (_15578_, _15577_, _15576_);
  nor _47736_ (_15579_, _15460_, _15454_);
  nand _47737_ (_15580_, _15579_, _26417_);
  or _47738_ (_15581_, _15580_, _15378_);
  or _47739_ (_15582_, _15581_, _15578_);
  or _47740_ (_15583_, _15194_, _26440_);
  and _47741_ (_15584_, _15428_, _26181_);
  or _47742_ (_15585_, _15584_, _15530_);
  or _47743_ (_15586_, _15585_, _15583_);
  and _47744_ (_15587_, _26333_, _26273_);
  and _47745_ (_15588_, _15198_, _26280_);
  and _47746_ (_15589_, _15428_, _26269_);
  or _47747_ (_15590_, _15589_, _15588_);
  or _47748_ (_15591_, _15590_, _15587_);
  or _47749_ (_15592_, _15591_, _15586_);
  or _47750_ (_15593_, _15427_, _26404_);
  or _47751_ (_15594_, _15510_, _15403_);
  or _47752_ (_15595_, _15594_, _15593_);
  or _47753_ (_15596_, _15595_, _15592_);
  or _47754_ (_15597_, _15596_, _15582_);
  or _47755_ (_15598_, _15597_, _15575_);
  and _47756_ (_15599_, _15598_, _25987_);
  and _47757_ (_15600_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47758_ (_15601_, _15366_, _26450_);
  or _47759_ (_15602_, _15601_, _15600_);
  or _47760_ (_15603_, _15602_, _15599_);
  and _47761_ (_23907_, _15603_, _27355_);
  and _47762_ (_15604_, _15350_, _26350_);
  nor _47763_ (_15605_, _15604_, _15446_);
  and _47764_ (_15606_, _15605_, _26407_);
  nand _47765_ (_15607_, _15606_, _26418_);
  and _47766_ (_15608_, _15540_, _26413_);
  or _47767_ (_15609_, _15608_, _26340_);
  or _47768_ (_15610_, _15609_, _15607_);
  or _47769_ (_15611_, _26440_, _26334_);
  and _47770_ (_15612_, _15198_, _26326_);
  or _47771_ (_15613_, _15612_, _15324_);
  or _47772_ (_15614_, _15613_, _15611_);
  or _47773_ (_15615_, _15614_, _15594_);
  or _47774_ (_15616_, _15615_, _15593_);
  or _47775_ (_15617_, _15616_, _15610_);
  or _47776_ (_15618_, _15617_, _15575_);
  and _47777_ (_15619_, _15618_, _25987_);
  and _47778_ (_15620_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47779_ (_15621_, _15620_, _15601_);
  or _47780_ (_15622_, _15621_, _15619_);
  and _47781_ (_23908_, _15622_, _27355_);
  and _47782_ (_15623_, _15309_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _47783_ (_15624_, _26312_, _26413_);
  or _47784_ (_15625_, _15584_, _15624_);
  and _47785_ (_15626_, _26397_, _26311_);
  and _47786_ (_15627_, _15350_, _26264_);
  and _47787_ (_15628_, _15627_, _26208_);
  or _47788_ (_15629_, _15628_, _15626_);
  or _47789_ (_15630_, _15629_, _15625_);
  or _47790_ (_15631_, _15630_, _15392_);
  or _47791_ (_15632_, _15435_, _01750_);
  or _47792_ (_15633_, _15632_, _15444_);
  or _47793_ (_15634_, _15633_, _15631_);
  or _47794_ (_15635_, _15506_, _15346_);
  and _47795_ (_15636_, _26289_, _26413_);
  and _47796_ (_15637_, _26294_, _26413_);
  or _47797_ (_15638_, _15637_, _15636_);
  or _47798_ (_15639_, _15427_, _15327_);
  or _47799_ (_15640_, _15639_, _15638_);
  or _47800_ (_15641_, _15640_, _15635_);
  nand _47801_ (_15642_, _26407_, _26360_);
  or _47802_ (_15643_, _15394_, _15393_);
  or _47803_ (_15644_, _15643_, _15642_);
  and _47804_ (_15645_, _26266_, _26413_);
  or _47805_ (_15646_, _15645_, _01753_);
  or _47806_ (_15647_, _15646_, _15644_);
  or _47807_ (_15648_, _15647_, _15641_);
  or _47808_ (_15649_, _15648_, _15634_);
  and _47809_ (_15650_, _15649_, _15202_);
  or _47810_ (_23909_, _15650_, _15623_);
  or _47811_ (_15651_, _15589_, _15410_);
  or _47812_ (_15652_, _15651_, _15637_);
  or _47813_ (_15653_, _15652_, _15409_);
  or _47814_ (_15654_, _15653_, _15586_);
  or _47815_ (_15655_, _15506_, _15624_);
  not _47816_ (_15656_, _26338_);
  or _47817_ (_15657_, _15510_, _15656_);
  or _47818_ (_15658_, _15657_, _15655_);
  not _47819_ (_15659_, _26417_);
  or _47820_ (_15660_, _15659_, _26283_);
  or _47821_ (_15661_, _15412_, _15330_);
  or _47822_ (_15662_, _15661_, _15660_);
  or _47823_ (_15663_, _15417_, _26414_);
  or _47824_ (_15664_, _15663_, _26404_);
  or _47825_ (_15665_, _15664_, _15662_);
  or _47826_ (_15666_, _15665_, _15658_);
  or _47827_ (_15667_, _15666_, _15654_);
  and _47828_ (_15668_, _15667_, _15202_);
  and _47829_ (_15669_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47830_ (_15670_, _26440_, _26393_);
  or _47831_ (_15671_, _15670_, _15669_);
  and _47832_ (_15672_, _15671_, _27355_);
  or _47833_ (_23910_, _15672_, _15668_);
  nor _47834_ (_15673_, _15530_, _15656_);
  or _47835_ (_15674_, _15435_, _15314_);
  or _47836_ (_15675_, _15674_, _15571_);
  and _47837_ (_15676_, _26311_, _26413_);
  or _47838_ (_15677_, _15676_, _01752_);
  or _47839_ (_15678_, _15355_, _15330_);
  or _47840_ (_15679_, _15678_, _15677_);
  nor _47841_ (_15680_, _15679_, _15675_);
  nand _47842_ (_15681_, _15680_, _15673_);
  or _47843_ (_15682_, _15639_, _26409_);
  or _47844_ (_15683_, _15524_, _26267_);
  or _47845_ (_15684_, _15509_, _26402_);
  or _47846_ (_15685_, _15684_, _15683_);
  or _47847_ (_15686_, _15685_, _15682_);
  or _47848_ (_15687_, _15686_, _15353_);
  or _47849_ (_15688_, _15687_, _15347_);
  or _47850_ (_15689_, _15688_, _15681_);
  and _47851_ (_15690_, _15689_, _25987_);
  and _47852_ (_15691_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47853_ (_15692_, _15691_, _26447_);
  or _47854_ (_15693_, _15692_, _15690_);
  and _47855_ (_23911_, _15693_, _27355_);
  or _47856_ (_15694_, _15683_, _15635_);
  or _47857_ (_15695_, _15694_, _15684_);
  and _47858_ (_15696_, _26293_, _26413_);
  or _47859_ (_15697_, _26405_, _26399_);
  or _47860_ (_15698_, _15697_, _15696_);
  or _47861_ (_15699_, _15530_, _26334_);
  or _47862_ (_15700_, _15699_, _15698_);
  or _47863_ (_15701_, _15385_, _01750_);
  or _47864_ (_15702_, _15701_, _15700_);
  or _47865_ (_15703_, _15352_, _15345_);
  or _47866_ (_15704_, _15703_, _15702_);
  or _47867_ (_15705_, _15704_, _15695_);
  and _47868_ (_15706_, _15705_, _25987_);
  and _47869_ (_15707_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _47870_ (_15708_, _15707_, _26448_);
  or _47871_ (_15709_, _15708_, _15706_);
  and _47872_ (_23912_, _15709_, _27355_);
  and _47873_ (_15710_, _15309_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _47874_ (_15711_, _15655_, _15638_);
  or _47875_ (_15712_, _15711_, _15646_);
  not _47876_ (_15713_, _26284_);
  and _47877_ (_15714_, _26266_, _15713_);
  or _47878_ (_15715_, _15311_, _26309_);
  or _47879_ (_15716_, _15715_, _15714_);
  or _47880_ (_15717_, _15716_, _15434_);
  or _47881_ (_15718_, _15717_, _15632_);
  or _47882_ (_15719_, _15718_, _15712_);
  and _47883_ (_15720_, _15719_, _15202_);
  or _47884_ (_23913_, _15720_, _15710_);
  and _47885_ (_24306_, _26204_, _27355_);
  nor _47886_ (_24307_, _01743_, rst);
  and _47887_ (_15721_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _47888_ (_15722_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _47889_ (_15723_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _47890_ (_15724_, _26002_, _26193_);
  nor _47891_ (_15725_, _15724_, _15723_);
  nor _47892_ (_15726_, _25996_, _01735_);
  and _47893_ (_15727_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _47894_ (_15728_, _15727_, _15726_);
  not _47895_ (_15729_, _26009_);
  and _47896_ (_15730_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _47897_ (_15731_, _26018_, _26190_);
  nor _47898_ (_15732_, _15731_, _15730_);
  and _47899_ (_15733_, _15732_, _15728_);
  and _47900_ (_15734_, _15733_, _15725_);
  nor _47901_ (_15735_, _15734_, _25992_);
  nor _47902_ (_15736_, _15735_, _15722_);
  nor _47903_ (_15737_, _15736_, _01726_);
  nor _47904_ (_15738_, _15737_, _15721_);
  nor _47905_ (_24308_, _15738_, rst);
  nor _47906_ (_24320_, _26028_, rst);
  and _47907_ (_24321_, _26149_, _27355_);
  nor _47908_ (_24322_, _26121_, rst);
  and _47909_ (_24323_, _26079_, _27355_);
  and _47910_ (_24324_, _26177_, _27355_);
  and _47911_ (_24325_, _26232_, _27355_);
  and _47912_ (_24327_, _26259_, _27355_);
  nor _47913_ (_24328_, _01847_, rst);
  nor _47914_ (_24329_, _01947_, rst);
  nor _47915_ (_24330_, _02124_, rst);
  nor _47916_ (_24331_, _01806_, rst);
  nor _47917_ (_24333_, _01902_, rst);
  nor _47918_ (_24334_, _01980_, rst);
  nor _47919_ (_24335_, _02047_, rst);
  and _47920_ (_15739_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _47921_ (_15740_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _47922_ (_15741_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _47923_ (_15742_, _26002_, _25994_);
  nor _47924_ (_15743_, _15742_, _15741_);
  nor _47925_ (_15744_, _25996_, _01841_);
  and _47926_ (_15745_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _47927_ (_15746_, _15745_, _15744_);
  and _47928_ (_15747_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _47929_ (_15748_, _26018_, _26008_);
  nor _47930_ (_15749_, _15748_, _15747_);
  and _47931_ (_15750_, _15749_, _15746_);
  and _47932_ (_15751_, _15750_, _15743_);
  nor _47933_ (_15752_, _15751_, _25992_);
  nor _47934_ (_15753_, _15752_, _15740_);
  nor _47935_ (_15754_, _15753_, _01726_);
  nor _47936_ (_15755_, _15754_, _15739_);
  nor _47937_ (_24336_, _15755_, rst);
  and _47938_ (_15756_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _47939_ (_15757_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  nor _47940_ (_15758_, _25996_, _01935_);
  nor _47941_ (_15759_, _26002_, _26129_);
  nor _47942_ (_15760_, _15759_, _15758_);
  and _47943_ (_15761_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _47944_ (_15762_, _26018_, _26127_);
  nor _47945_ (_15763_, _15762_, _15761_);
  and _47946_ (_15764_, _15763_, _15760_);
  and _47947_ (_15765_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _47948_ (_15766_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _47949_ (_15767_, _15766_, _15765_);
  and _47950_ (_15768_, _15767_, _15764_);
  nor _47951_ (_15769_, _15768_, _25992_);
  nor _47952_ (_15770_, _15769_, _15757_);
  nor _47953_ (_15771_, _15770_, _01726_);
  nor _47954_ (_15772_, _15771_, _15756_);
  nor _47955_ (_24337_, _15772_, rst);
  and _47956_ (_15773_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _47957_ (_15774_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor _47958_ (_15775_, _25996_, _02112_);
  nor _47959_ (_15776_, _26002_, _26111_);
  nor _47960_ (_15777_, _15776_, _15775_);
  and _47961_ (_15778_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _47962_ (_15779_, _26018_, _26105_);
  nor _47963_ (_15780_, _15779_, _15778_);
  and _47964_ (_15781_, _15780_, _15777_);
  and _47965_ (_15782_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _47966_ (_15783_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _47967_ (_15784_, _15783_, _15782_);
  and _47968_ (_15785_, _15784_, _15781_);
  nor _47969_ (_15786_, _15785_, _25992_);
  nor _47970_ (_15787_, _15786_, _15774_);
  nor _47971_ (_15788_, _15787_, _01726_);
  nor _47972_ (_15789_, _15788_, _15773_);
  nor _47973_ (_24339_, _15789_, rst);
  and _47974_ (_15790_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _47975_ (_15791_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _47976_ (_15792_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _47977_ (_15793_, _26002_, _26057_);
  nor _47978_ (_15794_, _15793_, _15792_);
  nor _47979_ (_15795_, _25996_, _01794_);
  and _47980_ (_15796_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _47981_ (_15797_, _15796_, _15795_);
  and _47982_ (_15798_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _47983_ (_15799_, _26018_, _26051_);
  nor _47984_ (_15800_, _15799_, _15798_);
  and _47985_ (_15801_, _15800_, _15797_);
  and _47986_ (_15802_, _15801_, _15794_);
  nor _47987_ (_15803_, _15802_, _25992_);
  nor _47988_ (_15804_, _15803_, _15791_);
  nor _47989_ (_15805_, _15804_, _01726_);
  nor _47990_ (_15806_, _15805_, _15790_);
  nor _47991_ (_24340_, _15806_, rst);
  and _47992_ (_15807_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _47993_ (_15808_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  nor _47994_ (_15809_, _25996_, _01892_);
  nor _47995_ (_15810_, _26002_, _26159_);
  nor _47996_ (_15811_, _15810_, _15809_);
  and _47997_ (_15812_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _47998_ (_15813_, _26018_, _26157_);
  nor _47999_ (_15814_, _15813_, _15812_);
  and _48000_ (_15815_, _15814_, _15811_);
  and _48001_ (_15816_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _48002_ (_15817_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _48003_ (_15818_, _15817_, _15816_);
  and _48004_ (_15819_, _15818_, _15815_);
  nor _48005_ (_15820_, _15819_, _25992_);
  nor _48006_ (_15821_, _15820_, _15808_);
  nor _48007_ (_15822_, _15821_, _01726_);
  nor _48008_ (_15823_, _15822_, _15807_);
  nor _48009_ (_24341_, _15823_, rst);
  and _48010_ (_15824_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _48011_ (_15825_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _48012_ (_15826_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _48013_ (_15827_, _26002_, _26212_);
  nor _48014_ (_15828_, _15827_, _15826_);
  nor _48015_ (_15829_, _25996_, _01971_);
  and _48016_ (_15830_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _48017_ (_15831_, _15830_, _15829_);
  and _48018_ (_15832_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _48019_ (_15833_, _26018_, _26218_);
  nor _48020_ (_15834_, _15833_, _15832_);
  and _48021_ (_15835_, _15834_, _15831_);
  and _48022_ (_15836_, _15835_, _15828_);
  nor _48023_ (_15837_, _15836_, _25992_);
  nor _48024_ (_15838_, _15837_, _15825_);
  nor _48025_ (_15839_, _15838_, _01726_);
  nor _48026_ (_15840_, _15839_, _15824_);
  nor _48027_ (_24342_, _15840_, rst);
  and _48028_ (_15841_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _48029_ (_15842_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _48030_ (_15843_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _48031_ (_15844_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _48032_ (_15845_, _15844_, _15843_);
  and _48033_ (_15846_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _48034_ (_15847_, _26018_, _26251_);
  nor _48035_ (_15848_, _15847_, _15846_);
  nor _48036_ (_15849_, _26002_, _26245_);
  nor _48037_ (_15850_, _25996_, _02035_);
  nor _48038_ (_15851_, _15850_, _15849_);
  and _48039_ (_15852_, _15851_, _15848_);
  and _48040_ (_15853_, _15852_, _15845_);
  nor _48041_ (_15854_, _15853_, _25992_);
  nor _48042_ (_15855_, _15854_, _15842_);
  nor _48043_ (_15856_, _15855_, _01726_);
  nor _48044_ (_15857_, _15856_, _15841_);
  nor _48045_ (_24343_, _15857_, rst);
  and _48046_ (_15858_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _48047_ (_15859_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _48048_ (_15860_, pc_log_change, _15859_);
  or _48049_ (_15861_, _15860_, _15858_);
  and _48050_ (_24370_, _15861_, _27355_);
  or _48051_ (_15862_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand _48052_ (_15863_, pc_log_change, _15859_);
  and _48053_ (_15864_, _15863_, _27355_);
  and _48054_ (_24372_, _15864_, _15862_);
  nor _48055_ (_24404_, _01748_, rst);
  nor _48056_ (_24405_, _01639_, rst);
  and _48057_ (_24406_, _01721_, _27355_);
  and _48058_ (_15865_, _26383_, _26353_);
  not _48059_ (_15866_, _15865_);
  nor _48060_ (_15867_, _02004_, _26922_);
  and _48061_ (_15868_, _02004_, _26922_);
  nor _48062_ (_15869_, _15868_, _15867_);
  nor _48063_ (_15870_, _01907_, _01637_);
  and _48064_ (_15871_, _01907_, _01637_);
  nor _48065_ (_15872_, _15871_, _15870_);
  and _48066_ (_15873_, _15872_, _15869_);
  nor _48067_ (_15874_, _01811_, _25116_);
  and _48068_ (_15875_, _01811_, _25116_);
  nor _48069_ (_15876_, _15875_, _15874_);
  nor _48070_ (_15877_, _02053_, _26458_);
  and _48071_ (_15878_, _02053_, _26458_);
  nor _48072_ (_15879_, _15878_, _15877_);
  and _48073_ (_15880_, _15879_, _02062_);
  and _48074_ (_15881_, _15880_, _15876_);
  and _48075_ (_15882_, _15881_, _15873_);
  nor _48076_ (_15883_, _01854_, _25053_);
  and _48077_ (_15884_, _01854_, _25053_);
  nor _48078_ (_15885_, _15884_, _15883_);
  nor _48079_ (_15886_, _15885_, _27160_);
  and _48080_ (_15887_, _01952_, _25714_);
  nor _48081_ (_15888_, _01952_, _25714_);
  or _48082_ (_15889_, _15888_, _15887_);
  nor _48083_ (_15890_, _02129_, _25020_);
  and _48084_ (_15891_, _02129_, _25020_);
  nor _48085_ (_15892_, _15891_, _15890_);
  nor _48086_ (_15893_, _15892_, _15889_);
  and _48087_ (_15894_, _15893_, _15886_);
  and _48088_ (_15895_, _15894_, _15882_);
  nor _48089_ (_15896_, _25101_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _48090_ (_15897_, _15896_, _15895_);
  not _48091_ (_15898_, _15897_);
  nor _48092_ (_15899_, _26319_, _26382_);
  nor _48093_ (_15900_, _25517_, _27575_);
  and _48094_ (_15901_, _15900_, _15882_);
  and _48095_ (_15902_, _15901_, _15899_);
  nor _48096_ (_15903_, _15377_, _26393_);
  nor _48097_ (_15904_, _15865_, _26372_);
  and _48098_ (_15905_, _26311_, _15371_);
  or _48099_ (_15906_, _15317_, _15659_);
  and _48100_ (_15907_, _15899_, _25193_);
  not _48101_ (_15908_, _15907_);
  nor _48102_ (_15909_, _15899_, _26446_);
  and _48103_ (_15910_, _25675_, _25530_);
  nand _48104_ (_15911_, _15910_, _25760_);
  nor _48105_ (_15912_, _15911_, _25792_);
  and _48106_ (_15913_, _15912_, _25857_);
  and _48107_ (_15914_, _15913_, _25335_);
  and _48108_ (_15915_, _15914_, _25918_);
  and _48109_ (_15916_, _15915_, _15909_);
  and _48110_ (_15917_, _15916_, _25351_);
  and _48111_ (_15918_, _26376_, _26291_);
  and _48112_ (_15919_, _15918_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _48113_ (_15920_, _15919_, _15917_);
  nor _48114_ (_15921_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _48115_ (_15922_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _48116_ (_15923_, _15922_, _15921_);
  nor _48117_ (_15924_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _48118_ (_15925_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _48119_ (_15926_, _15925_, _15924_);
  and _48120_ (_15927_, _15926_, _15923_);
  nand _48121_ (_15928_, _15927_, _26432_);
  and _48122_ (_15929_, _15928_, _15920_);
  and _48123_ (_15930_, _15929_, _15908_);
  not _48124_ (_15931_, _26286_);
  or _48125_ (_15932_, _26312_, _26299_);
  nor _48126_ (_15933_, _15932_, _26333_);
  nor _48127_ (_15934_, _15933_, _15931_);
  not _48128_ (_15935_, _15934_);
  or _48129_ (_15936_, _15571_, _26290_);
  nor _48130_ (_15937_, _15936_, _15389_);
  and _48131_ (_15938_, _15937_, _15539_);
  and _48132_ (_15939_, _15938_, _15935_);
  not _48133_ (_15940_, _15939_);
  and _48134_ (_15941_, _15940_, _15930_);
  and _48135_ (_15942_, _26375_, _26269_);
  nor _48136_ (_15943_, _15942_, _26317_);
  nor _48137_ (_15944_, _15943_, _15930_);
  or _48138_ (_15945_, _15944_, _15941_);
  or _48139_ (_15946_, _15945_, _15906_);
  nor _48140_ (_15947_, _15946_, _15905_);
  nor _48141_ (_15948_, _15947_, _15904_);
  nor _48142_ (_15949_, _15948_, _15903_);
  not _48143_ (_15950_, _26446_);
  nor _48144_ (_15951_, _15899_, _26281_);
  nor _48145_ (_15952_, _15951_, _15950_);
  nor _48146_ (_15953_, _26942_, _26933_);
  and _48147_ (_15954_, _15953_, _26998_);
  not _48148_ (_15955_, _15954_);
  and _48149_ (_15956_, _15955_, _15952_);
  and _48150_ (_15957_, _26446_, _26236_);
  not _48151_ (_15958_, _27102_);
  and _48152_ (_15959_, _15958_, _15957_);
  nor _48153_ (_15960_, _15959_, _15956_);
  not _48154_ (_15961_, _15960_);
  nor _48155_ (_15962_, _15961_, _15949_);
  not _48156_ (_15963_, _15962_);
  nor _48157_ (_15964_, _15963_, _15902_);
  and _48158_ (_15965_, _15964_, _15898_);
  and _48159_ (_15966_, _15965_, _15866_);
  and _48160_ (_24410_, _15966_, _27355_);
  and _48161_ (_24411_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _27355_);
  and _48162_ (_24412_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _27355_);
  and _48163_ (_15967_, _25995_, _25999_);
  nor _48164_ (_15968_, _15967_, _01726_);
  nor _48165_ (_15969_, _15968_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _48166_ (_15970_, _15969_);
  and _48167_ (_15971_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _48168_ (_15972_, _15971_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _48169_ (_15973_, _15972_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _48170_ (_15974_, _15973_, _15970_);
  and _48171_ (_15975_, _15974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _48172_ (_15976_, _15975_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _48173_ (_15977_, _15976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _48174_ (_15978_, _15977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _48175_ (_15979_, _15978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _48176_ (_15980_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _48177_ (_15981_, _15980_, _15979_);
  and _48178_ (_15982_, _15981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _48179_ (_15983_, _15982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _48180_ (_15984_, _15983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _48181_ (_15985_, _15983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _48182_ (_15986_, _15985_, _15984_);
  or _48183_ (_15987_, _15986_, _15965_);
  and _48184_ (_15988_, _15987_, _27355_);
  and _48185_ (_15989_, _26286_, _25983_);
  and _48186_ (_15990_, _15989_, _26311_);
  not _48187_ (_15991_, _15990_);
  nand _48188_ (_15992_, _15539_, _26319_);
  or _48189_ (_15993_, _15992_, _15936_);
  nand _48190_ (_15994_, _15993_, _26372_);
  and _48191_ (_15995_, _26383_, _15905_);
  and _48192_ (_15996_, _26293_, _15371_);
  and _48193_ (_15997_, _15996_, _25983_);
  nor _48194_ (_15998_, _15997_, _15995_);
  and _48195_ (_15999_, _15998_, _15994_);
  and _48196_ (_16000_, _15999_, _15991_);
  and _48197_ (_16001_, _16000_, _01743_);
  nand _48198_ (_16002_, _15999_, _15991_);
  and _48199_ (_16003_, _16002_, _15738_);
  nor _48200_ (_16004_, _16003_, _16001_);
  and _48201_ (_16005_, _16004_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _48202_ (_16006_, _16005_);
  nor _48203_ (_16007_, _16004_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _48204_ (_16008_, _16007_, _16005_);
  not _48205_ (_16009_, _16008_);
  and _48206_ (_16010_, _16000_, _02047_);
  and _48207_ (_16011_, _16002_, _15857_);
  nor _48208_ (_16012_, _16011_, _16010_);
  and _48209_ (_16013_, _16012_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _48210_ (_16014_, _16013_);
  nor _48211_ (_16015_, _16012_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _48212_ (_16016_, _16015_, _16013_);
  and _48213_ (_16017_, _16000_, _01980_);
  and _48214_ (_16018_, _16002_, _15840_);
  nor _48215_ (_16019_, _16018_, _16017_);
  nor _48216_ (_16020_, _16019_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _48217_ (_16021_, _16019_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _48218_ (_16022_, _16000_, _01902_);
  and _48219_ (_16023_, _16002_, _15823_);
  nor _48220_ (_16024_, _16023_, _16022_);
  nand _48221_ (_16025_, _16024_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _48222_ (_16026_, _16000_, _01806_);
  and _48223_ (_16027_, _16002_, _15806_);
  nor _48224_ (_16028_, _16027_, _16026_);
  nor _48225_ (_16029_, _16028_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _48226_ (_16030_, _16028_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _48227_ (_16031_, _16002_, _02125_);
  not _48228_ (_16032_, _15789_);
  or _48229_ (_16033_, _16000_, _16032_);
  and _48230_ (_16034_, _16033_, _16031_);
  and _48231_ (_16035_, _16034_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _48232_ (_16036_, _16002_, _01948_);
  not _48233_ (_16037_, _15772_);
  or _48234_ (_16038_, _16000_, _16037_);
  and _48235_ (_16039_, _16038_, _16036_);
  nand _48236_ (_16040_, _16039_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _48237_ (_16041_, _16040_);
  or _48238_ (_16042_, _16002_, _01848_);
  not _48239_ (_16043_, _15755_);
  or _48240_ (_16044_, _16000_, _16043_);
  and _48241_ (_16045_, _16044_, _16042_);
  and _48242_ (_16046_, _16045_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _48243_ (_16047_, _16039_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _48244_ (_16048_, _16047_, _16040_);
  and _48245_ (_16049_, _16048_, _16046_);
  or _48246_ (_16050_, _16049_, _16041_);
  not _48247_ (_16051_, _16035_);
  or _48248_ (_16052_, _16034_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _48249_ (_16053_, _16052_, _16051_);
  and _48250_ (_16054_, _16053_, _16050_);
  or _48251_ (_16055_, _16054_, _16035_);
  nor _48252_ (_16056_, _16055_, _16030_);
  nor _48253_ (_16057_, _16056_, _16029_);
  or _48254_ (_16058_, _16024_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _48255_ (_16059_, _16058_, _16025_);
  nand _48256_ (_16060_, _16059_, _16057_);
  nand _48257_ (_16061_, _16060_, _16025_);
  nor _48258_ (_16062_, _16061_, _16021_);
  nor _48259_ (_16063_, _16062_, _16020_);
  nand _48260_ (_16064_, _16063_, _16016_);
  and _48261_ (_16065_, _16064_, _16014_);
  or _48262_ (_16066_, _16065_, _16009_);
  and _48263_ (_16067_, _16066_, _16006_);
  nand _48264_ (_16068_, _16067_, _24240_);
  or _48265_ (_16069_, _16068_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _48266_ (_16070_, _16069_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _48267_ (_16071_, _16070_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _48268_ (_16072_, _16071_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _48269_ (_16073_, _16072_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _48270_ (_16074_, _16073_, _24129_);
  nand _48271_ (_16075_, _16074_, _16004_);
  not _48272_ (_16076_, _16004_);
  nor _48273_ (_16077_, _16067_, _24240_);
  and _48274_ (_16078_, _16077_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _48275_ (_16079_, _16078_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _48276_ (_16080_, _16079_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _48277_ (_16081_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _48278_ (_16082_, _16081_, _16080_);
  nand _48279_ (_16083_, _16082_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _48280_ (_16084_, _16083_, _16076_);
  nand _48281_ (_16085_, _16084_, _16075_);
  nand _48282_ (_16086_, _16085_, _24158_);
  or _48283_ (_16087_, _16085_, _24158_);
  and _48284_ (_16088_, _16087_, _16086_);
  not _48285_ (_16089_, _26372_);
  not _48286_ (_16090_, _15992_);
  and _48287_ (_16091_, _15318_, _26417_);
  and _48288_ (_16092_, _16091_, _15937_);
  and _48289_ (_16093_, _16092_, _16090_);
  nor _48290_ (_16094_, _16093_, _16089_);
  nor _48291_ (_16095_, _16094_, _15990_);
  nor _48292_ (_16096_, _26417_, _16089_);
  nor _48293_ (_16097_, _16096_, _15903_);
  not _48294_ (_16098_, _16097_);
  and _48295_ (_16099_, _16098_, _16000_);
  nor _48296_ (_16100_, _16099_, _16095_);
  and _48297_ (_16101_, _16100_, _16088_);
  and _48298_ (_16102_, _15895_, _25102_);
  and _48299_ (_16103_, _16102_, _25444_);
  nor _48300_ (_16104_, _16103_, _15902_);
  and _48301_ (_16105_, _15958_, _26432_);
  not _48302_ (_16106_, _16105_);
  and _48303_ (_16107_, _15955_, _15918_);
  nor _48304_ (_16108_, _16107_, _15949_);
  and _48305_ (_16109_, _16108_, _16106_);
  and _48306_ (_16110_, _16109_, _16104_);
  and _48307_ (_16111_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _48308_ (_16112_, _16111_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _48309_ (_16113_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _48310_ (_16114_, _16113_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _48311_ (_16115_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _48312_ (_16116_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _48313_ (_16117_, _16116_, _16115_);
  and _48314_ (_16118_, _16117_, _16114_);
  and _48315_ (_16119_, _16118_, _16112_);
  and _48316_ (_16120_, _16119_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _48317_ (_16121_, _16120_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _48318_ (_16122_, _16121_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _48319_ (_16123_, _16122_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _48320_ (_16124_, _16123_, _24158_);
  or _48321_ (_16125_, _16123_, _24158_);
  and _48322_ (_16126_, _16125_, _16124_);
  and _48323_ (_16127_, _15999_, _15903_);
  and _48324_ (_16128_, _16127_, _16126_);
  and _48325_ (_16129_, _15995_, _25441_);
  and _48326_ (_16130_, _16096_, _26678_);
  and _48327_ (_16131_, _16097_, _15999_);
  and _48328_ (_16132_, _16131_, _16095_);
  and _48329_ (_16133_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _48330_ (_16134_, _15376_, _25983_);
  and _48331_ (_16135_, _16134_, _01744_);
  or _48332_ (_16136_, _16135_, _16133_);
  or _48333_ (_16137_, _16136_, _16130_);
  or _48334_ (_16138_, _16137_, _16129_);
  nor _48335_ (_16139_, _16138_, _16128_);
  nand _48336_ (_16140_, _16139_, _16110_);
  or _48337_ (_16141_, _16140_, _16101_);
  and _48338_ (_24414_, _16141_, _15988_);
  and _48339_ (_16142_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _27355_);
  and _48340_ (_16143_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _48341_ (_16144_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _48342_ (_16145_, _25987_, _16144_);
  not _48343_ (_16146_, _16145_);
  not _48344_ (_16147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _48345_ (_16148_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _48346_ (_16149_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _48347_ (_16150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _48348_ (_16151_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _48349_ (_16152_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _48350_ (_16153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _48351_ (_16154_, _16153_, _16151_);
  and _48352_ (_16155_, _16154_, _16152_);
  nor _48353_ (_16156_, _16155_, _16151_);
  nor _48354_ (_16157_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _48355_ (_16158_, _16157_, _16150_);
  not _48356_ (_16159_, _16158_);
  nor _48357_ (_16160_, _16159_, _16156_);
  nor _48358_ (_16161_, _16160_, _16150_);
  not _48359_ (_16162_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _48360_ (_16163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _48361_ (_16164_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _48362_ (_16165_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _48363_ (_16166_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _48364_ (_16167_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _48365_ (_16168_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _48366_ (_16169_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _48367_ (_16170_, _16169_, _16168_);
  and _48368_ (_16171_, _16170_, _16167_);
  and _48369_ (_16172_, _16171_, _16166_);
  and _48370_ (_16173_, _16172_, _16165_);
  and _48371_ (_16174_, _16173_, _16164_);
  and _48372_ (_16175_, _16174_, _16163_);
  and _48373_ (_16176_, _16175_, _16162_);
  and _48374_ (_16177_, _16176_, _16161_);
  and _48375_ (_16178_, _16177_, _16149_);
  and _48376_ (_16179_, _16178_, _16148_);
  and _48377_ (_16180_, _16179_, _16147_);
  nor _48378_ (_16181_, _16180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _48379_ (_16182_, _16180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _48380_ (_16183_, _16182_, _16181_);
  nor _48381_ (_16184_, _16179_, _16147_);
  nor _48382_ (_16185_, _16184_, _16180_);
  not _48383_ (_16186_, _16185_);
  nor _48384_ (_16187_, _16178_, _16148_);
  nor _48385_ (_16188_, _16187_, _16179_);
  not _48386_ (_16189_, _16188_);
  nor _48387_ (_16190_, _16177_, _16149_);
  nor _48388_ (_16191_, _16190_, _16178_);
  not _48389_ (_16192_, _16191_);
  and _48390_ (_16193_, _16161_, _16175_);
  nor _48391_ (_16194_, _16193_, _16162_);
  nor _48392_ (_16195_, _16194_, _16177_);
  not _48393_ (_16196_, _16195_);
  and _48394_ (_16197_, _16161_, _16173_);
  and _48395_ (_16198_, _16197_, _16164_);
  nor _48396_ (_16199_, _16198_, _16163_);
  or _48397_ (_16200_, _16199_, _16193_);
  nor _48398_ (_16201_, _16197_, _16164_);
  nor _48399_ (_16202_, _16201_, _16198_);
  not _48400_ (_16203_, _16202_);
  and _48401_ (_16204_, _16161_, _16171_);
  nor _48402_ (_16205_, _16204_, _16166_);
  and _48403_ (_16206_, _16161_, _16172_);
  or _48404_ (_16207_, _16206_, _16205_);
  and _48405_ (_16208_, _16161_, _16170_);
  nor _48406_ (_16209_, _16208_, _16167_);
  nor _48407_ (_16210_, _16209_, _16204_);
  not _48408_ (_16211_, _16210_);
  and _48409_ (_16212_, _16161_, _16169_);
  nor _48410_ (_16213_, _16212_, _16168_);
  nor _48411_ (_16214_, _16213_, _16208_);
  not _48412_ (_16215_, _16214_);
  not _48413_ (_16216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _48414_ (_16217_, _16161_, _16216_);
  nor _48415_ (_16218_, _16161_, _16216_);
  nor _48416_ (_16219_, _16218_, _16217_);
  not _48417_ (_16220_, _16219_);
  and _48418_ (_16221_, _15265_, _15243_);
  and _48419_ (_16222_, _15221_, _15211_);
  and _48420_ (_16223_, _15262_, _16222_);
  and _48421_ (_16224_, _15262_, _15223_);
  or _48422_ (_16225_, _16224_, _16223_);
  nor _48423_ (_16226_, _16225_, _16221_);
  and _48424_ (_16227_, _15289_, _15281_);
  and _48425_ (_16228_, _15272_, _15235_);
  nor _48426_ (_16229_, _16228_, _16227_);
  and _48427_ (_16230_, _16229_, _16226_);
  nor _48428_ (_16231_, _15293_, _15276_);
  not _48429_ (_16232_, _26079_);
  and _48430_ (_16233_, _15251_, _15221_);
  nor _48431_ (_16234_, _16233_, _15269_);
  nor _48432_ (_16235_, _16234_, _16232_);
  not _48433_ (_16236_, _15272_);
  nor _48434_ (_16237_, _15269_, _15292_);
  nor _48435_ (_16238_, _16237_, _16236_);
  nor _48436_ (_16239_, _16238_, _16235_);
  and _48437_ (_16240_, _16239_, _16231_);
  and _48438_ (_16241_, _16240_, _16230_);
  not _48439_ (_16242_, _15262_);
  and _48440_ (_16243_, _15215_, _15231_);
  nor _48441_ (_16244_, _16233_, _16243_);
  nor _48442_ (_16245_, _16244_, _16242_);
  not _48443_ (_16246_, _16245_);
  and _48444_ (_16247_, _15285_, _15272_);
  not _48445_ (_16248_, _15208_);
  nor _48446_ (_16249_, _15271_, _15269_);
  nor _48447_ (_16250_, _16249_, _16248_);
  nor _48448_ (_16251_, _16250_, _16247_);
  and _48449_ (_16252_, _16251_, _16246_);
  and _48450_ (_16253_, _16252_, _15268_);
  and _48451_ (_16254_, _16253_, _16241_);
  not _48452_ (_16255_, _15292_);
  nor _48453_ (_16256_, _15208_, _26079_);
  nor _48454_ (_16257_, _16256_, _16255_);
  not _48455_ (_16258_, _16257_);
  and _48456_ (_16259_, _15264_, _15215_);
  nor _48457_ (_16260_, _16259_, _16222_);
  nor _48458_ (_16261_, _15265_, _15216_);
  and _48459_ (_16262_, _16261_, _16260_);
  nor _48460_ (_16263_, _16262_, _16236_);
  not _48461_ (_16264_, _15232_);
  nor _48462_ (_16265_, _15272_, _15208_);
  nor _48463_ (_16266_, _16265_, _16264_);
  nor _48464_ (_16267_, _16266_, _16263_);
  and _48465_ (_16268_, _16267_, _16258_);
  or _48466_ (_16269_, _16233_, _16222_);
  not _48467_ (_16270_, _16269_);
  nor _48468_ (_16271_, _16259_, _15223_);
  and _48469_ (_16272_, _16271_, _16270_);
  nor _48470_ (_16273_, _16272_, _16248_);
  and _48471_ (_16274_, _15225_, _16232_);
  and _48472_ (_16275_, _15290_, _16274_);
  not _48473_ (_16276_, _16275_);
  nor _48474_ (_16277_, _15284_, _15227_);
  and _48475_ (_16278_, _16277_, _16276_);
  not _48476_ (_16279_, _16278_);
  nor _48477_ (_16280_, _16279_, _16273_);
  and _48478_ (_16281_, _15252_, _15211_);
  not _48479_ (_16282_, _16281_);
  nor _48480_ (_16283_, _15219_, _15208_);
  nor _48481_ (_16284_, _16283_, _16282_);
  nor _48482_ (_16285_, _15219_, _15207_);
  and _48483_ (_16286_, _15265_, _26028_);
  nor _48484_ (_16287_, _16286_, _15253_);
  nor _48485_ (_16288_, _16287_, _16285_);
  nor _48486_ (_16289_, _16288_, _16284_);
  and _48487_ (_16290_, _16289_, _16280_);
  and _48488_ (_16291_, _16290_, _16268_);
  nor _48489_ (_16292_, _15283_, _15273_);
  nand _48490_ (_16293_, _15224_, _15241_);
  and _48491_ (_16294_, _15289_, _15223_);
  and _48492_ (_16295_, _16281_, _15243_);
  nor _48493_ (_16296_, _16295_, _16294_);
  and _48494_ (_16297_, _16296_, _16293_);
  and _48495_ (_16298_, _16297_, _16292_);
  not _48496_ (_16299_, _16298_);
  nor _48497_ (_16300_, _15289_, _16274_);
  not _48498_ (_16301_, _15289_);
  nor _48499_ (_16302_, _16222_, _15260_);
  nor _48500_ (_16303_, _16302_, _16301_);
  nor _48501_ (_16304_, _16303_, _15269_);
  nor _48502_ (_16305_, _16304_, _16300_);
  nor _48503_ (_16306_, _16305_, _16299_);
  and _48504_ (_16307_, _16306_, _16291_);
  and _48505_ (_16308_, _16307_, _16254_);
  nor _48506_ (_16309_, _16154_, _16152_);
  nor _48507_ (_16310_, _16309_, _16155_);
  not _48508_ (_16311_, _16310_);
  nor _48509_ (_16312_, _16311_, _16308_);
  not _48510_ (_16313_, _16312_);
  and _48511_ (_16314_, _15253_, _15243_);
  or _48512_ (_16315_, _16223_, _16221_);
  or _48513_ (_16316_, _16315_, _16314_);
  or _48514_ (_16317_, _15263_, _15227_);
  or _48515_ (_16318_, _16238_, _15233_);
  or _48516_ (_16319_, _16318_, _16317_);
  or _48517_ (_16320_, _16319_, _16316_);
  or _48518_ (_16321_, _16320_, _16299_);
  nor _48519_ (_16322_, _16321_, _16308_);
  not _48520_ (_16323_, _16322_);
  nor _48521_ (_16324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _48522_ (_16325_, _16324_, _16152_);
  and _48523_ (_16326_, _16325_, _16323_);
  and _48524_ (_16327_, _16311_, _16308_);
  nor _48525_ (_16328_, _16327_, _16312_);
  nand _48526_ (_16329_, _16328_, _16326_);
  and _48527_ (_16330_, _16329_, _16313_);
  not _48528_ (_16331_, _16330_);
  and _48529_ (_16332_, _16159_, _16156_);
  nor _48530_ (_16333_, _16332_, _16160_);
  and _48531_ (_16334_, _16333_, _16331_);
  and _48532_ (_16335_, _16334_, _16220_);
  not _48533_ (_16336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _48534_ (_16337_, _16217_, _16336_);
  or _48535_ (_16338_, _16337_, _16212_);
  and _48536_ (_16339_, _16338_, _16335_);
  and _48537_ (_16340_, _16339_, _16215_);
  and _48538_ (_16341_, _16340_, _16211_);
  and _48539_ (_16342_, _16341_, _16207_);
  nor _48540_ (_16343_, _16206_, _16165_);
  or _48541_ (_16344_, _16343_, _16197_);
  and _48542_ (_16345_, _16344_, _16342_);
  and _48543_ (_16346_, _16345_, _16203_);
  and _48544_ (_16347_, _16346_, _16200_);
  and _48545_ (_16348_, _16347_, _16196_);
  and _48546_ (_16349_, _16348_, _16192_);
  and _48547_ (_16350_, _16349_, _16189_);
  and _48548_ (_16351_, _16350_, _16186_);
  or _48549_ (_16352_, _16351_, _16183_);
  nand _48550_ (_16353_, _16351_, _16183_);
  and _48551_ (_16354_, _16353_, _16352_);
  or _48552_ (_16355_, _16354_, _16146_);
  or _48553_ (_16356_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _48554_ (_16357_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _48555_ (_16358_, _16357_, _16356_);
  and _48556_ (_16359_, _16358_, _16355_);
  or _48557_ (_24415_, _16359_, _16143_);
  nor _48558_ (_16360_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _48559_ (_24416_, _16360_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _48560_ (_24417_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _27355_);
  nor _48561_ (_16361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _48562_ (_16362_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48563_ (_16363_, _16362_, _16361_);
  nor _48564_ (_16364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _48565_ (_16365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _48566_ (_16366_, _16365_, _16364_);
  and _48567_ (_16367_, _16366_, _16363_);
  nor _48568_ (_16368_, _16367_, rst);
  and _48569_ (_16369_, \oc8051_top_1.oc8051_rom1.ea_int , _25984_);
  nand _48570_ (_16370_, _16369_, _25987_);
  and _48571_ (_16371_, _16370_, _24417_);
  or _48572_ (_24418_, _16371_, _16368_);
  and _48573_ (_16372_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _48574_ (_16373_, _16372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _48575_ (_24419_, _16373_, _27355_);
  nor _48576_ (_16374_, _15969_, _01726_);
  nor _48577_ (_16375_, _16308_, _26000_);
  not _48578_ (_16376_, _16375_);
  nor _48579_ (_16377_, _16322_, _26016_);
  and _48580_ (_16378_, _16308_, _26000_);
  nor _48581_ (_16379_, _16378_, _16375_);
  nand _48582_ (_16380_, _16379_, _16377_);
  and _48583_ (_16381_, _16380_, _16376_);
  nor _48584_ (_16382_, _16381_, _01726_);
  and _48585_ (_16383_, _16382_, _25999_);
  nor _48586_ (_16384_, _16382_, _25999_);
  nor _48587_ (_16385_, _16384_, _16383_);
  nor _48588_ (_16386_, _16385_, _16374_);
  and _48589_ (_16387_, _26001_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _48590_ (_16388_, _16387_, _16374_);
  and _48591_ (_16389_, _16388_, _16321_);
  or _48592_ (_16390_, _16389_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _48593_ (_16391_, _16390_, _16386_);
  and _48594_ (_24420_, _16391_, _27355_);
  and _48595_ (_16392_, _26200_, _26023_);
  and _48596_ (_16393_, _16392_, _26071_);
  and _48597_ (_16394_, _26255_, _26142_);
  and _48598_ (_16395_, _16394_, _26115_);
  and _48599_ (_16396_, _25988_, _27355_);
  and _48600_ (_16397_, _16396_, _26171_);
  and _48601_ (_16398_, _16397_, _26227_);
  and _48602_ (_16399_, _16398_, _16395_);
  and _48603_ (_24423_, _16399_, _16393_);
  nor _48604_ (_16400_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _48605_ (_16401_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _48606_ (_16402_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _48607_ (_24426_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _27355_);
  and _48608_ (_16403_, _24426_, _16402_);
  or _48609_ (_24424_, _16403_, _16401_);
  not _48610_ (_16404_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _48611_ (_16405_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _48612_ (_16406_, _16405_, _16404_);
  and _48613_ (_16407_, _16405_, _16404_);
  nor _48614_ (_16408_, _16407_, _16406_);
  not _48615_ (_16409_, _16408_);
  and _48616_ (_16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _48617_ (_16411_, _16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _48618_ (_16412_, _16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _48619_ (_16413_, _16412_, _16411_);
  or _48620_ (_16414_, _16413_, _16405_);
  and _48621_ (_16415_, _16414_, _16409_);
  nor _48622_ (_16416_, _16406_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _48623_ (_16417_, _16406_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _48624_ (_16418_, _16417_, _16416_);
  or _48625_ (_16419_, _16411_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _48626_ (_24428_, _16419_, _27355_);
  and _48627_ (_16420_, _24428_, _16418_);
  and _48628_ (_24427_, _16420_, _16415_);
  not _48629_ (_16421_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _48630_ (_16422_, _15969_, _16421_);
  and _48631_ (_16423_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _48632_ (_16424_, _16422_);
  and _48633_ (_16425_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _48634_ (_16426_, _16425_, _16423_);
  and _48635_ (_24429_, _16426_, _27355_);
  and _48636_ (_16427_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _48637_ (_16428_, _16422_, _26193_);
  or _48638_ (_16429_, _16428_, _16427_);
  and _48639_ (_24430_, _16429_, _27355_);
  and _48640_ (_16430_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _48641_ (_16431_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _48642_ (_16432_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _16431_);
  and _48643_ (_16433_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _48644_ (_16434_, _16433_, _16430_);
  and _48645_ (_24431_, _16434_, _27355_);
  and _48646_ (_16435_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  or _48647_ (_16436_, _16435_, _16432_);
  and _48648_ (_24433_, _16436_, _27355_);
  or _48649_ (_16437_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _48650_ (_24434_, _16437_, _27355_);
  not _48651_ (_16438_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _48652_ (_16439_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _48653_ (_16440_, _16439_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _48654_ (_16441_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _48655_ (_16442_, _16441_, _27355_);
  and _48656_ (_24435_, _16442_, _16440_);
  or _48657_ (_16443_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _48658_ (_24436_, _16443_, _27355_);
  nor _48659_ (_16444_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _48660_ (_16445_, _16444_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _48661_ (_16446_, _16445_, _27355_);
  and _48662_ (_16447_, _24426_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _48663_ (_24437_, _16447_, _16446_);
  and _48664_ (_16448_, _16421_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _48665_ (_16449_, _16448_, _16445_);
  and _48666_ (_24438_, _16449_, _27355_);
  not _48667_ (_16450_, _16445_);
  or _48668_ (_16451_, _16450_, _26678_);
  or _48669_ (_16452_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _48670_ (_16453_, _16452_, _27355_);
  and _48671_ (_24439_, _16453_, _16451_);
  and _48672_ (_16454_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _48673_ (_16455_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _48674_ (_16456_, pc_log_change, _16455_);
  or _48675_ (_16457_, _16456_, _16454_);
  and _48676_ (_24470_, _16457_, _27355_);
  and _48677_ (_16458_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _48678_ (_16459_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _48679_ (_16460_, pc_log_change, _16459_);
  or _48680_ (_16461_, _16460_, _16458_);
  and _48681_ (_24472_, _16461_, _27355_);
  and _48682_ (_16462_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _48683_ (_16463_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _48684_ (_16464_, pc_log_change, _16463_);
  or _48685_ (_16465_, _16464_, _16462_);
  and _48686_ (_24473_, _16465_, _27355_);
  and _48687_ (_16466_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _48688_ (_16467_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _48689_ (_16468_, pc_log_change, _16467_);
  or _48690_ (_16469_, _16468_, _16466_);
  and _48691_ (_24474_, _16469_, _27355_);
  and _48692_ (_16470_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _48693_ (_16471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _48694_ (_16472_, pc_log_change, _16471_);
  or _48695_ (_16473_, _16472_, _16470_);
  and _48696_ (_24475_, _16473_, _27355_);
  and _48697_ (_16474_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _48698_ (_16475_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _48699_ (_16476_, pc_log_change, _16475_);
  or _48700_ (_16477_, _16476_, _16474_);
  and _48701_ (_24476_, _16477_, _27355_);
  and _48702_ (_16478_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _48703_ (_16479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _48704_ (_16480_, pc_log_change, _16479_);
  or _48705_ (_16481_, _16480_, _16478_);
  and _48706_ (_24477_, _16481_, _27355_);
  and _48707_ (_16482_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _48708_ (_16483_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _48709_ (_16484_, pc_log_change, _16483_);
  or _48710_ (_16485_, _16484_, _16482_);
  and _48711_ (_24478_, _16485_, _27355_);
  and _48712_ (_16486_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not _48713_ (_16487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _48714_ (_16488_, pc_log_change, _16487_);
  or _48715_ (_16489_, _16488_, _16486_);
  and _48716_ (_24479_, _16489_, _27355_);
  and _48717_ (_16490_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not _48718_ (_16491_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _48719_ (_16492_, pc_log_change, _16491_);
  or _48720_ (_16493_, _16492_, _16490_);
  and _48721_ (_24480_, _16493_, _27355_);
  and _48722_ (_16494_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not _48723_ (_16495_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _48724_ (_16496_, pc_log_change, _16495_);
  or _48725_ (_16497_, _16496_, _16494_);
  and _48726_ (_24481_, _16497_, _27355_);
  and _48727_ (_16498_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _48728_ (_16499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _48729_ (_16500_, pc_log_change, _16499_);
  or _48730_ (_16501_, _16500_, _16498_);
  and _48731_ (_24483_, _16501_, _27355_);
  and _48732_ (_16502_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not _48733_ (_16503_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _48734_ (_16504_, pc_log_change, _16503_);
  or _48735_ (_16505_, _16504_, _16502_);
  and _48736_ (_24484_, _16505_, _27355_);
  and _48737_ (_16506_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _48738_ (_16507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _48739_ (_16508_, pc_log_change, _16507_);
  or _48740_ (_16509_, _16508_, _16506_);
  and _48741_ (_24485_, _16509_, _27355_);
  and _48742_ (_16510_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _48743_ (_16511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _48744_ (_16512_, pc_log_change, _16511_);
  or _48745_ (_16513_, _16512_, _16510_);
  and _48746_ (_24486_, _16513_, _27355_);
  and _48747_ (_16514_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _48748_ (_16515_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _48749_ (_16516_, pc_log_change, _16515_);
  or _48750_ (_16517_, _16516_, _16514_);
  and _48751_ (_24490_, _16517_, _27355_);
  and _48752_ (_16518_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _48753_ (_16519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _48754_ (_16520_, pc_log_change, _16519_);
  or _48755_ (_16521_, _16520_, _16518_);
  and _48756_ (_24491_, _16521_, _27355_);
  and _48757_ (_16522_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _48758_ (_16523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _48759_ (_16524_, pc_log_change, _16523_);
  or _48760_ (_16525_, _16524_, _16522_);
  and _48761_ (_24492_, _16525_, _27355_);
  and _48762_ (_16526_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _48763_ (_16527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _48764_ (_16528_, pc_log_change, _16527_);
  or _48765_ (_16529_, _16528_, _16526_);
  and _48766_ (_24493_, _16529_, _27355_);
  or _48767_ (_16530_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand _48768_ (_16531_, pc_log_change, _16471_);
  and _48769_ (_16532_, _16531_, _27355_);
  and _48770_ (_24494_, _16532_, _16530_);
  or _48771_ (_16533_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand _48772_ (_16534_, pc_log_change, _16475_);
  and _48773_ (_16535_, _16534_, _27355_);
  and _48774_ (_24495_, _16535_, _16533_);
  or _48775_ (_16536_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand _48776_ (_16537_, pc_log_change, _16479_);
  and _48777_ (_16538_, _16537_, _27355_);
  and _48778_ (_24497_, _16538_, _16536_);
  and _48779_ (_16539_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _48780_ (_16540_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _48781_ (_16541_, pc_log_change, _16540_);
  or _48782_ (_16542_, _16541_, _16539_);
  and _48783_ (_24498_, _16542_, _27355_);
  or _48784_ (_16543_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand _48785_ (_16544_, pc_log_change, _16487_);
  and _48786_ (_16545_, _16544_, _27355_);
  and _48787_ (_24499_, _16545_, _16543_);
  and _48788_ (_16546_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not _48789_ (_16547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _48790_ (_16548_, pc_log_change, _16547_);
  or _48791_ (_16549_, _16548_, _16546_);
  and _48792_ (_24500_, _16549_, _27355_);
  and _48793_ (_16550_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not _48794_ (_16551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _48795_ (_16552_, pc_log_change, _16551_);
  or _48796_ (_16553_, _16552_, _16550_);
  and _48797_ (_24501_, _16553_, _27355_);
  or _48798_ (_16554_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand _48799_ (_16555_, pc_log_change, _16499_);
  and _48800_ (_16556_, _16555_, _27355_);
  and _48801_ (_24502_, _16556_, _16554_);
  and _48802_ (_16557_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  not _48803_ (_16558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _48804_ (_16559_, pc_log_change, _16558_);
  or _48805_ (_16560_, _16559_, _16557_);
  and _48806_ (_24503_, _16560_, _27355_);
  or _48807_ (_16561_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand _48808_ (_16562_, pc_log_change, _16507_);
  and _48809_ (_16563_, _16562_, _27355_);
  and _48810_ (_24504_, _16563_, _16561_);
  or _48811_ (_16564_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand _48812_ (_16565_, pc_log_change, _16511_);
  and _48813_ (_16566_, _16565_, _27355_);
  and _48814_ (_24505_, _16566_, _16564_);
  and _48815_ (_24692_, _26033_, _27355_);
  and _48816_ (_24693_, _26153_, _27355_);
  and _48817_ (_24695_, _26125_, _27355_);
  nor _48818_ (_24696_, _01632_, rst);
  nor _48819_ (_16567_, _16422_, _26008_);
  and _48820_ (_16568_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _48821_ (_16569_, _16568_, _16422_);
  or _48822_ (_16570_, _16569_, _16567_);
  and _48823_ (_24697_, _16570_, _27355_);
  nor _48824_ (_16571_, _16422_, _26127_);
  and _48825_ (_16572_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _48826_ (_16573_, _16572_, _16422_);
  or _48827_ (_16574_, _16573_, _16571_);
  and _48828_ (_24698_, _16574_, _27355_);
  nor _48829_ (_16575_, _16422_, _26105_);
  and _48830_ (_16576_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _48831_ (_16577_, _16576_, _16575_);
  and _48832_ (_24699_, _16577_, _27355_);
  nor _48833_ (_16578_, _16422_, _26051_);
  and _48834_ (_16579_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _48835_ (_16580_, _16579_, _16578_);
  and _48836_ (_24700_, _16580_, _27355_);
  nor _48837_ (_16581_, _16422_, _26157_);
  and _48838_ (_16582_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _48839_ (_16583_, _16582_, _16581_);
  and _48840_ (_24701_, _16583_, _27355_);
  nor _48841_ (_16584_, _16422_, _26218_);
  and _48842_ (_16585_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _48843_ (_16586_, _16585_, _16422_);
  or _48844_ (_16587_, _16586_, _16584_);
  and _48845_ (_24702_, _16587_, _27355_);
  nor _48846_ (_16588_, _16422_, _26251_);
  and _48847_ (_16589_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _48848_ (_16590_, _16589_, _16588_);
  and _48849_ (_24703_, _16590_, _27355_);
  nor _48850_ (_16591_, _16422_, _26190_);
  and _48851_ (_16592_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _48852_ (_16593_, _16592_, _16591_);
  and _48853_ (_24704_, _16593_, _27355_);
  and _48854_ (_16594_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nor _48855_ (_16595_, _16422_, _01841_);
  or _48856_ (_16596_, _16595_, _16594_);
  and _48857_ (_24706_, _16596_, _27355_);
  and _48858_ (_16597_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nor _48859_ (_16598_, _16422_, _01935_);
  or _48860_ (_16599_, _16598_, _16597_);
  and _48861_ (_24707_, _16599_, _27355_);
  and _48862_ (_16600_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nor _48863_ (_16601_, _16422_, _02112_);
  or _48864_ (_16602_, _16601_, _16600_);
  and _48865_ (_24708_, _16602_, _27355_);
  and _48866_ (_16603_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nor _48867_ (_16604_, _16422_, _01794_);
  or _48868_ (_16605_, _16604_, _16603_);
  and _48869_ (_24709_, _16605_, _27355_);
  and _48870_ (_16606_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nor _48871_ (_16607_, _16422_, _01892_);
  or _48872_ (_16608_, _16607_, _16606_);
  and _48873_ (_24710_, _16608_, _27355_);
  and _48874_ (_16609_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nor _48875_ (_16610_, _16422_, _01971_);
  or _48876_ (_16611_, _16610_, _16609_);
  and _48877_ (_24711_, _16611_, _27355_);
  and _48878_ (_16612_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nor _48879_ (_16613_, _16422_, _02035_);
  or _48880_ (_16614_, _16613_, _16612_);
  and _48881_ (_24712_, _16614_, _27355_);
  and _48882_ (_16615_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nor _48883_ (_16616_, _16422_, _01735_);
  or _48884_ (_16617_, _16616_, _16615_);
  and _48885_ (_24713_, _16617_, _27355_);
  and _48886_ (_16618_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _48887_ (_16619_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _48888_ (_16620_, _16619_, _16618_);
  and _48889_ (_24714_, _16620_, _27355_);
  and _48890_ (_16621_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _48891_ (_16622_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _48892_ (_16623_, _16622_, _16621_);
  and _48893_ (_24715_, _16623_, _27355_);
  and _48894_ (_16624_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _48895_ (_16625_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _48896_ (_16626_, _16625_, _16624_);
  and _48897_ (_24717_, _16626_, _27355_);
  and _48898_ (_16627_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _48899_ (_16628_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _48900_ (_16629_, _16628_, _16627_);
  and _48901_ (_24718_, _16629_, _27355_);
  and _48902_ (_16630_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _48903_ (_16631_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _48904_ (_16632_, _16631_, _16630_);
  and _48905_ (_24719_, _16632_, _27355_);
  and _48906_ (_16633_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _48907_ (_16634_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _48908_ (_16635_, _16634_, _16633_);
  and _48909_ (_24720_, _16635_, _27355_);
  and _48910_ (_16636_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _48911_ (_16637_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _48912_ (_16638_, _16637_, _16636_);
  and _48913_ (_24721_, _16638_, _27355_);
  and _48914_ (_16639_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _48915_ (_16640_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _48916_ (_16641_, _16640_, _16639_);
  and _48917_ (_24722_, _16641_, _27355_);
  and _48918_ (_16642_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _48919_ (_16643_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _48920_ (_16644_, _16643_, _16642_);
  and _48921_ (_24723_, _16644_, _27355_);
  and _48922_ (_16645_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _48923_ (_16646_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _48924_ (_16647_, _16646_, _16645_);
  and _48925_ (_24724_, _16647_, _27355_);
  and _48926_ (_16648_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _48927_ (_16649_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _48928_ (_16650_, _16649_, _16648_);
  and _48929_ (_24725_, _16650_, _27355_);
  and _48930_ (_16651_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _48931_ (_16652_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _48932_ (_16653_, _16652_, _16651_);
  and _48933_ (_24726_, _16653_, _27355_);
  and _48934_ (_16654_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _48935_ (_16655_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _48936_ (_16656_, _16655_, _16654_);
  and _48937_ (_24728_, _16656_, _27355_);
  and _48938_ (_16657_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _48939_ (_16658_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _48940_ (_16659_, _16658_, _16657_);
  and _48941_ (_24729_, _16659_, _27355_);
  and _48942_ (_16660_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _48943_ (_16661_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _48944_ (_16662_, _16661_, _16660_);
  and _48945_ (_24730_, _16662_, _27355_);
  and _48946_ (_24731_, _01830_, _27355_);
  and _48947_ (_24732_, _01926_, _27355_);
  and _48948_ (_24733_, _02104_, _27355_);
  and _48949_ (_24735_, _01784_, _27355_);
  and _48950_ (_24736_, _01880_, _27355_);
  and _48951_ (_24737_, _02000_, _27355_);
  and _48952_ (_24738_, _02029_, _27355_);
  and _48953_ (_24755_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _27355_);
  and _48954_ (_24756_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _27355_);
  and _48955_ (_24757_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _27355_);
  and _48956_ (_24758_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _27355_);
  and _48957_ (_24759_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _27355_);
  and _48958_ (_24760_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _27355_);
  and _48959_ (_24761_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _27355_);
  not _48960_ (_16663_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _48961_ (_16664_, _15966_, _16663_);
  or _48962_ (_16665_, _16132_, _16096_);
  and _48963_ (_16666_, _16665_, _25563_);
  or _48964_ (_16667_, _16045_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _48965_ (_16668_, _16046_);
  and _48966_ (_16669_, _26311_, _25983_);
  and _48967_ (_16670_, _16669_, _26286_);
  nor _48968_ (_16671_, _16094_, _16670_);
  not _48969_ (_16672_, _16670_);
  nor _48970_ (_16673_, _16134_, _15865_);
  and _48971_ (_16674_, _16673_, _15994_);
  and _48972_ (_16675_, _16674_, _16672_);
  and _48973_ (_16676_, _16098_, _16675_);
  nor _48974_ (_16677_, _16676_, _16671_);
  and _48975_ (_16678_, _16677_, _16668_);
  and _48976_ (_16679_, _16678_, _16667_);
  and _48977_ (_16680_, _16134_, _16043_);
  not _48978_ (_16681_, _16094_);
  and _48979_ (_16682_, _16676_, _16681_);
  and _48980_ (_16683_, _16682_, _01848_);
  or _48981_ (_16684_, _16683_, _16680_);
  or _48982_ (_16685_, _16684_, _16679_);
  or _48983_ (_16686_, _16685_, _16666_);
  and _48984_ (_16687_, _16686_, _16110_);
  or _48985_ (_16688_, _16687_, _16664_);
  and _48986_ (_24762_, _16688_, _27355_);
  not _48987_ (_16689_, _15965_);
  and _48988_ (_16690_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _48989_ (_16691_, _16665_, _25639_);
  or _48990_ (_16692_, _16048_, _16046_);
  not _48991_ (_16693_, _16049_);
  and _48992_ (_16694_, _16677_, _16693_);
  and _48993_ (_16695_, _16694_, _16692_);
  and _48994_ (_16696_, _16682_, _01948_);
  and _48995_ (_16697_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _48996_ (_16698_, _16134_, _16037_);
  or _48997_ (_16699_, _16698_, _16697_);
  or _48998_ (_16700_, _16699_, _16696_);
  or _48999_ (_16701_, _16700_, _16695_);
  or _49000_ (_16702_, _16701_, _16691_);
  and _49001_ (_16703_, _16702_, _15965_);
  or _49002_ (_16704_, _16703_, _16690_);
  and _49003_ (_24763_, _16704_, _27355_);
  not _49004_ (_16705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _49005_ (_16706_, _15969_, _16705_);
  and _49006_ (_16707_, _15969_, _16705_);
  nor _49007_ (_16708_, _16707_, _16706_);
  and _49008_ (_16709_, _16708_, _16689_);
  and _49009_ (_16710_, _16665_, _25705_);
  or _49010_ (_16711_, _16053_, _16050_);
  not _49011_ (_16712_, _16054_);
  and _49012_ (_16713_, _16677_, _16712_);
  and _49013_ (_16714_, _16713_, _16711_);
  and _49014_ (_16715_, _16682_, _02125_);
  and _49015_ (_16716_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _49016_ (_16717_, _16134_, _16032_);
  or _49017_ (_16718_, _16717_, _16716_);
  or _49018_ (_16719_, _16718_, _16715_);
  or _49019_ (_16720_, _16719_, _16714_);
  or _49020_ (_16721_, _16720_, _16710_);
  and _49021_ (_16722_, _16721_, _15965_);
  or _49022_ (_16723_, _16722_, _16709_);
  and _49023_ (_24765_, _16723_, _27355_);
  and _49024_ (_16724_, _16706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _49025_ (_16725_, _16706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _49026_ (_16726_, _16725_, _16724_);
  or _49027_ (_16727_, _16726_, _15965_);
  and _49028_ (_16728_, _16727_, _27355_);
  and _49029_ (_16729_, _16665_, _25770_);
  and _49030_ (_16730_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not _49031_ (_16731_, _15806_);
  and _49032_ (_16732_, _15997_, _16731_);
  and _49033_ (_16733_, _16127_, _01807_);
  or _49034_ (_16734_, _16733_, _16732_);
  or _49035_ (_16735_, _16734_, _16730_);
  or _49036_ (_16736_, _16029_, _16030_);
  and _49037_ (_16737_, _16736_, _16055_);
  nor _49038_ (_16738_, _16736_, _16055_);
  or _49039_ (_16739_, _16738_, _16737_);
  and _49040_ (_16740_, _16739_, _16100_);
  or _49041_ (_16741_, _16740_, _16735_);
  nor _49042_ (_16742_, _16741_, _16729_);
  nand _49043_ (_16743_, _16742_, _16110_);
  and _49044_ (_24766_, _16743_, _16728_);
  and _49045_ (_16744_, _15972_, _15970_);
  nor _49046_ (_16745_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _49047_ (_16746_, _16745_, _16744_);
  or _49048_ (_16747_, _16746_, _15965_);
  and _49049_ (_16748_, _16747_, _27355_);
  and _49050_ (_16749_, _16665_, _25830_);
  or _49051_ (_16750_, _16059_, _16057_);
  and _49052_ (_16751_, _16677_, _16060_);
  and _49053_ (_16752_, _16751_, _16750_);
  and _49054_ (_16753_, _16682_, _01903_);
  and _49055_ (_16754_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not _49056_ (_16755_, _15823_);
  and _49057_ (_16756_, _16134_, _16755_);
  or _49058_ (_16757_, _16756_, _16754_);
  or _49059_ (_16758_, _16757_, _16753_);
  nor _49060_ (_16759_, _16758_, _16752_);
  nand _49061_ (_16760_, _16759_, _15965_);
  or _49062_ (_16761_, _16760_, _16749_);
  and _49063_ (_24767_, _16761_, _16748_);
  nor _49064_ (_16762_, _16744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _49065_ (_16763_, _16762_, _15974_);
  nor _49066_ (_16764_, _16763_, _15965_);
  and _49067_ (_16765_, _16665_, _25898_);
  not _49068_ (_16766_, _16061_);
  or _49069_ (_16767_, _16021_, _16020_);
  nand _49070_ (_16768_, _16767_, _16766_);
  or _49071_ (_16769_, _16767_, _16766_);
  and _49072_ (_16770_, _16769_, _16677_);
  and _49073_ (_16771_, _16770_, _16768_);
  and _49074_ (_16772_, _16682_, _01981_);
  and _49075_ (_16773_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not _49076_ (_16774_, _15840_);
  and _49077_ (_16775_, _16134_, _16774_);
  or _49078_ (_16776_, _16775_, _16773_);
  or _49079_ (_16777_, _16776_, _16772_);
  or _49080_ (_16778_, _16777_, _16771_);
  or _49081_ (_16779_, _16778_, _16765_);
  and _49082_ (_16780_, _16779_, _15965_);
  or _49083_ (_16781_, _16780_, _16764_);
  and _49084_ (_24768_, _16781_, _27355_);
  nor _49085_ (_16782_, _15974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _49086_ (_16783_, _16782_, _15975_);
  or _49087_ (_16784_, _16783_, _15965_);
  and _49088_ (_16785_, _16784_, _27355_);
  or _49089_ (_16786_, _16063_, _16016_);
  and _49090_ (_16787_, _16786_, _16064_);
  and _49091_ (_16788_, _16787_, _16100_);
  and _49092_ (_16789_, _16665_, _25964_);
  and _49093_ (_16790_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _49094_ (_16791_, _15857_);
  and _49095_ (_16792_, _15997_, _16791_);
  and _49096_ (_16793_, _16127_, _02048_);
  or _49097_ (_16794_, _16793_, _16792_);
  or _49098_ (_16795_, _16794_, _16790_);
  or _49099_ (_16796_, _16795_, _16789_);
  nor _49100_ (_16797_, _16796_, _16788_);
  nand _49101_ (_16798_, _16797_, _16110_);
  and _49102_ (_24769_, _16798_, _16785_);
  nor _49103_ (_16799_, _15975_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _49104_ (_16800_, _16799_, _15976_);
  or _49105_ (_16801_, _16800_, _15965_);
  and _49106_ (_16802_, _16801_, _27355_);
  and _49107_ (_16803_, _16665_, _25441_);
  and _49108_ (_16804_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _49109_ (_16805_, _15738_);
  and _49110_ (_16806_, _15997_, _16805_);
  and _49111_ (_16807_, _16127_, _01744_);
  or _49112_ (_16808_, _16807_, _16806_);
  or _49113_ (_16809_, _16808_, _16804_);
  nand _49114_ (_16810_, _16065_, _16009_);
  and _49115_ (_16811_, _16100_, _16066_);
  and _49116_ (_16812_, _16811_, _16810_);
  or _49117_ (_16813_, _16812_, _16809_);
  nor _49118_ (_16814_, _16813_, _16803_);
  nand _49119_ (_16815_, _16814_, _16110_);
  and _49120_ (_24770_, _16815_, _16802_);
  nor _49121_ (_16816_, _15976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _49122_ (_16817_, _16816_, _15977_);
  or _49123_ (_16818_, _16817_, _15965_);
  and _49124_ (_16819_, _16818_, _27355_);
  nor _49125_ (_16820_, _16067_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _49126_ (_16821_, _16067_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _49127_ (_16822_, _16821_, _16820_);
  nor _49128_ (_16823_, _16822_, _16004_);
  and _49129_ (_16824_, _16822_, _16004_);
  or _49130_ (_16825_, _16824_, _16823_);
  and _49131_ (_16826_, _16825_, _16677_);
  nor _49132_ (_16827_, _15866_, _25562_);
  and _49133_ (_16828_, _16096_, _26713_);
  and _49134_ (_16829_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _49135_ (_16830_, _16134_, _01848_);
  or _49136_ (_16831_, _16830_, _16829_);
  and _49137_ (_16832_, _16682_, _26232_);
  nor _49138_ (_16833_, _16832_, _16831_);
  nand _49139_ (_16834_, _16833_, _15965_);
  or _49140_ (_16835_, _16834_, _16828_);
  or _49141_ (_16836_, _16835_, _16827_);
  or _49142_ (_16837_, _16836_, _16826_);
  and _49143_ (_24771_, _16837_, _16819_);
  nor _49144_ (_16838_, _15977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _49145_ (_16839_, _16838_, _15978_);
  or _49146_ (_16840_, _16839_, _15965_);
  and _49147_ (_16841_, _16840_, _27355_);
  nor _49148_ (_16842_, _16068_, _16076_);
  and _49149_ (_16843_, _16077_, _16076_);
  nor _49150_ (_16844_, _16843_, _16842_);
  nand _49151_ (_16845_, _16844_, _24188_);
  or _49152_ (_16846_, _16844_, _24188_);
  and _49153_ (_16847_, _16846_, _16845_);
  and _49154_ (_16848_, _16847_, _16100_);
  and _49155_ (_16849_, _16127_, _26259_);
  and _49156_ (_16850_, _15995_, _25639_);
  not _49157_ (_16851_, _16096_);
  nor _49158_ (_16852_, _16851_, _26745_);
  and _49159_ (_16853_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _49160_ (_16854_, _16134_, _01948_);
  or _49161_ (_16855_, _16854_, _16853_);
  or _49162_ (_16856_, _16855_, _16852_);
  or _49163_ (_16857_, _16856_, _16850_);
  nor _49164_ (_16858_, _16857_, _16849_);
  nand _49165_ (_16859_, _16858_, _16110_);
  or _49166_ (_16860_, _16859_, _16848_);
  and _49167_ (_24772_, _16860_, _16841_);
  nor _49168_ (_16861_, _15978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _49169_ (_16862_, _16861_, _15979_);
  or _49170_ (_16863_, _16862_, _15965_);
  and _49171_ (_16864_, _16863_, _27355_);
  and _49172_ (_16865_, _16842_, _24188_);
  and _49173_ (_16866_, _16078_, _16076_);
  nor _49174_ (_16867_, _16866_, _16865_);
  nand _49175_ (_16868_, _16867_, _24204_);
  or _49176_ (_16869_, _16867_, _24204_);
  and _49177_ (_16870_, _16869_, _16677_);
  and _49178_ (_16871_, _16870_, _16868_);
  nor _49179_ (_16872_, _15866_, _25704_);
  nor _49180_ (_16873_, _16851_, _26775_);
  and _49181_ (_16874_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _49182_ (_16875_, _16134_, _02125_);
  or _49183_ (_16876_, _16875_, _16874_);
  and _49184_ (_16877_, _16127_, _26204_);
  or _49185_ (_16878_, _16877_, _16876_);
  nor _49186_ (_16879_, _16878_, _16873_);
  nand _49187_ (_16880_, _16879_, _15965_);
  or _49188_ (_16881_, _16880_, _16872_);
  or _49189_ (_16882_, _16881_, _16871_);
  and _49190_ (_24773_, _16882_, _16864_);
  nor _49191_ (_16883_, _15979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _49192_ (_16884_, _15979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _49193_ (_16885_, _16884_, _16883_);
  or _49194_ (_16886_, _16885_, _15965_);
  and _49195_ (_16887_, _16886_, _27355_);
  nand _49196_ (_16888_, _16079_, _16076_);
  or _49197_ (_16889_, _16070_, _16076_);
  nand _49198_ (_16890_, _16889_, _16888_);
  nand _49199_ (_16891_, _16890_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _49200_ (_16892_, _16890_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _49201_ (_16893_, _16892_, _16677_);
  and _49202_ (_16894_, _16893_, _16891_);
  nor _49203_ (_16895_, _15866_, _25769_);
  nor _49204_ (_16896_, _16851_, _26808_);
  and _49205_ (_16897_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _49206_ (_16898_, _16134_, _01807_);
  or _49207_ (_16899_, _16898_, _16897_);
  nor _49208_ (_16900_, _16119_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _49209_ (_16901_, _16900_, _16120_);
  and _49210_ (_16902_, _16901_, _16682_);
  or _49211_ (_16903_, _16902_, _16899_);
  nor _49212_ (_16904_, _16903_, _16896_);
  nand _49213_ (_16905_, _16904_, _15965_);
  or _49214_ (_16906_, _16905_, _16895_);
  or _49215_ (_16907_, _16906_, _16894_);
  and _49216_ (_24774_, _16907_, _16887_);
  nor _49217_ (_16908_, _16884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _49218_ (_16909_, _16908_, _15981_);
  or _49219_ (_16910_, _16909_, _15965_);
  and _49220_ (_16911_, _16910_, _27355_);
  nor _49221_ (_16912_, _16071_, _16076_);
  and _49222_ (_16913_, _16080_, _16076_);
  nor _49223_ (_16914_, _16913_, _16912_);
  nand _49224_ (_16915_, _16914_, _23940_);
  or _49225_ (_16916_, _16914_, _23940_);
  and _49226_ (_16917_, _16916_, _16915_);
  and _49227_ (_16918_, _16917_, _16100_);
  nor _49228_ (_16919_, _16120_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _49229_ (_16920_, _16919_, _16121_);
  and _49230_ (_16921_, _16920_, _16127_);
  and _49231_ (_16922_, _15995_, _25830_);
  and _49232_ (_16923_, _16096_, _26837_);
  and _49233_ (_16924_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _49234_ (_16925_, _16134_, _01903_);
  or _49235_ (_16926_, _16925_, _16924_);
  or _49236_ (_16927_, _16926_, _16923_);
  or _49237_ (_16928_, _16927_, _16922_);
  nor _49238_ (_16929_, _16928_, _16921_);
  nand _49239_ (_16930_, _16929_, _16110_);
  or _49240_ (_16931_, _16930_, _16918_);
  and _49241_ (_24776_, _16931_, _16911_);
  not _49242_ (_16932_, _16110_);
  or _49243_ (_16933_, _16072_, _16076_);
  nand _49244_ (_16934_, _16913_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _49245_ (_16935_, _16934_, _16933_);
  nor _49246_ (_16936_, _16935_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _49247_ (_16937_, _16935_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _49248_ (_16938_, _16937_, _16936_);
  and _49249_ (_16939_, _16938_, _16677_);
  and _49250_ (_16940_, _15865_, _25898_);
  and _49251_ (_16941_, _16096_, _26867_);
  and _49252_ (_16942_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _49253_ (_16943_, _16134_, _01981_);
  or _49254_ (_16944_, _16943_, _16942_);
  nor _49255_ (_16945_, _16121_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _49256_ (_16946_, _16945_, _16122_);
  and _49257_ (_16947_, _16946_, _16682_);
  or _49258_ (_16948_, _16947_, _16944_);
  or _49259_ (_16949_, _16948_, _16941_);
  or _49260_ (_16950_, _16949_, _16940_);
  or _49261_ (_16951_, _16950_, _16939_);
  or _49262_ (_16952_, _16951_, _16932_);
  nor _49263_ (_16953_, _15981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _49264_ (_16954_, _16953_, _15982_);
  or _49265_ (_16955_, _16954_, _16110_);
  and _49266_ (_16956_, _16955_, _27355_);
  and _49267_ (_24777_, _16956_, _16952_);
  or _49268_ (_16957_, _16082_, _16004_);
  or _49269_ (_16958_, _16073_, _16076_);
  and _49270_ (_16959_, _16958_, _16957_);
  nor _49271_ (_16960_, _16959_, _24129_);
  and _49272_ (_16961_, _16959_, _24129_);
  or _49273_ (_16962_, _16961_, _16960_);
  and _49274_ (_16963_, _16962_, _16677_);
  nor _49275_ (_16964_, _15866_, _25963_);
  nor _49276_ (_16965_, _16851_, _26898_);
  and _49277_ (_16966_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _49278_ (_16967_, _16134_, _02048_);
  or _49279_ (_16968_, _16967_, _16966_);
  or _49280_ (_16969_, _16122_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _49281_ (_16970_, _16969_, _16123_);
  and _49282_ (_16971_, _16970_, _16682_);
  or _49283_ (_16972_, _16971_, _16968_);
  or _49284_ (_16973_, _16972_, _16965_);
  or _49285_ (_16974_, _16973_, _16964_);
  or _49286_ (_16975_, _16974_, _16963_);
  or _49287_ (_16976_, _16975_, _16932_);
  nor _49288_ (_16977_, _15982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _49289_ (_16978_, _16977_, _15983_);
  or _49290_ (_16979_, _16978_, _16110_);
  and _49291_ (_16980_, _16979_, _27355_);
  and _49292_ (_24778_, _16980_, _16976_);
  and _49293_ (_16981_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _49294_ (_16982_, _16325_, _16323_);
  nor _49295_ (_16983_, _16982_, _16326_);
  or _49296_ (_16984_, _16983_, _16146_);
  or _49297_ (_16985_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _49298_ (_16986_, _16985_, _16357_);
  and _49299_ (_16987_, _16986_, _16984_);
  or _49300_ (_24779_, _16987_, _16981_);
  or _49301_ (_16988_, _16328_, _16326_);
  and _49302_ (_16989_, _16988_, _16329_);
  or _49303_ (_16990_, _16989_, _16146_);
  or _49304_ (_16991_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _49305_ (_16992_, _16991_, _16357_);
  and _49306_ (_16993_, _16992_, _16990_);
  and _49307_ (_16994_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _49308_ (_24780_, _16994_, _16993_);
  nor _49309_ (_16995_, _16333_, _16331_);
  nor _49310_ (_16996_, _16995_, _16334_);
  or _49311_ (_16997_, _16996_, _16146_);
  or _49312_ (_16998_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _49313_ (_16999_, _16998_, _16357_);
  and _49314_ (_17000_, _16999_, _16997_);
  and _49315_ (_17001_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _49316_ (_24781_, _17001_, _17000_);
  nor _49317_ (_17002_, _16334_, _16220_);
  nor _49318_ (_17003_, _17002_, _16335_);
  or _49319_ (_17004_, _17003_, _16146_);
  or _49320_ (_17005_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _49321_ (_17006_, _17005_, _16357_);
  and _49322_ (_17007_, _17006_, _17004_);
  and _49323_ (_17008_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _49324_ (_24782_, _17008_, _17007_);
  and _49325_ (_17009_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _49326_ (_17010_, _16338_, _16335_);
  nor _49327_ (_17011_, _17010_, _16339_);
  or _49328_ (_17012_, _17011_, _16146_);
  or _49329_ (_17013_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _49330_ (_17014_, _17013_, _16357_);
  and _49331_ (_17015_, _17014_, _17012_);
  or _49332_ (_24783_, _17015_, _17009_);
  and _49333_ (_17016_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _49334_ (_17017_, _16339_, _16215_);
  nor _49335_ (_17018_, _17017_, _16340_);
  or _49336_ (_17019_, _17018_, _16146_);
  or _49337_ (_17020_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _49338_ (_17021_, _17020_, _16357_);
  and _49339_ (_17022_, _17021_, _17019_);
  or _49340_ (_24784_, _17022_, _17016_);
  and _49341_ (_17023_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _49342_ (_17024_, _16340_, _16211_);
  nor _49343_ (_17025_, _17024_, _16341_);
  or _49344_ (_17026_, _17025_, _16146_);
  or _49345_ (_17027_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _49346_ (_17028_, _17027_, _16357_);
  and _49347_ (_17029_, _17028_, _17026_);
  or _49348_ (_24785_, _17029_, _17023_);
  or _49349_ (_17030_, _16341_, _16207_);
  nor _49350_ (_17031_, _16342_, _16146_);
  and _49351_ (_17032_, _17031_, _17030_);
  nor _49352_ (_17033_, _16145_, _24160_);
  or _49353_ (_17034_, _17033_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _49354_ (_17035_, _17034_, _17032_);
  or _49355_ (_17036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _25984_);
  and _49356_ (_17037_, _17036_, _27355_);
  and _49357_ (_24787_, _17037_, _17035_);
  nor _49358_ (_17038_, _16344_, _16342_);
  nor _49359_ (_17039_, _17038_, _16345_);
  or _49360_ (_17040_, _17039_, _16146_);
  or _49361_ (_17041_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _49362_ (_17042_, _17041_, _16357_);
  and _49363_ (_17043_, _17042_, _17040_);
  and _49364_ (_17044_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _49365_ (_24788_, _17044_, _17043_);
  nor _49366_ (_17045_, _16345_, _16203_);
  nor _49367_ (_17046_, _17045_, _16346_);
  or _49368_ (_17047_, _17046_, _16146_);
  or _49369_ (_17048_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _49370_ (_17049_, _17048_, _16357_);
  and _49371_ (_17050_, _17049_, _17047_);
  and _49372_ (_17051_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _49373_ (_24789_, _17051_, _17050_);
  nor _49374_ (_17052_, _16346_, _16200_);
  nor _49375_ (_17053_, _17052_, _16347_);
  or _49376_ (_17054_, _17053_, _16146_);
  or _49377_ (_17055_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _49378_ (_17056_, _17055_, _16357_);
  and _49379_ (_17057_, _17056_, _17054_);
  and _49380_ (_17058_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _49381_ (_24790_, _17058_, _17057_);
  nor _49382_ (_17059_, _16347_, _16196_);
  nor _49383_ (_17060_, _17059_, _16348_);
  or _49384_ (_17061_, _17060_, _16146_);
  or _49385_ (_17062_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _49386_ (_17063_, _17062_, _16357_);
  and _49387_ (_17064_, _17063_, _17061_);
  and _49388_ (_17065_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _49389_ (_24791_, _17065_, _17064_);
  nor _49390_ (_17066_, _16348_, _16192_);
  nor _49391_ (_17067_, _17066_, _16349_);
  or _49392_ (_17068_, _17067_, _16146_);
  or _49393_ (_17069_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _49394_ (_17070_, _17069_, _16357_);
  and _49395_ (_17071_, _17070_, _17068_);
  and _49396_ (_17072_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _49397_ (_24792_, _17072_, _17071_);
  nor _49398_ (_17073_, _16349_, _16189_);
  nor _49399_ (_17074_, _17073_, _16350_);
  or _49400_ (_17075_, _17074_, _16146_);
  or _49401_ (_17076_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _49402_ (_17077_, _17076_, _16357_);
  and _49403_ (_17078_, _17077_, _17075_);
  and _49404_ (_17079_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _49405_ (_24793_, _17079_, _17078_);
  and _49406_ (_17080_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _49407_ (_17081_, _16350_, _16186_);
  nor _49408_ (_17082_, _17081_, _16351_);
  or _49409_ (_17083_, _17082_, _16146_);
  or _49410_ (_17084_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _49411_ (_17085_, _17084_, _16357_);
  and _49412_ (_17086_, _17085_, _17083_);
  or _49413_ (_24794_, _17086_, _17080_);
  and _49414_ (_17087_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _49415_ (_17088_, _17087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _49416_ (_24795_, _17088_, _27355_);
  and _49417_ (_17089_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _49418_ (_17090_, _17089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _49419_ (_24796_, _17090_, _27355_);
  and _49420_ (_17091_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _49421_ (_17092_, _17091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _49422_ (_24798_, _17092_, _27355_);
  and _49423_ (_17093_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _49424_ (_17094_, _17093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _49425_ (_24799_, _17094_, _27355_);
  and _49426_ (_17095_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _49427_ (_17096_, _17095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _49428_ (_24800_, _17096_, _27355_);
  and _49429_ (_17097_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _49430_ (_17098_, _17097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _49431_ (_24801_, _17098_, _27355_);
  and _49432_ (_17099_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _49433_ (_17100_, _17099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _49434_ (_24802_, _17100_, _27355_);
  nor _49435_ (_17101_, _16322_, _01726_);
  nand _49436_ (_17102_, _17101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _49437_ (_17103_, _17101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _49438_ (_17104_, _17103_, _16357_);
  and _49439_ (_24803_, _17104_, _17102_);
  or _49440_ (_17105_, _16379_, _16377_);
  and _49441_ (_17106_, _17105_, _16380_);
  or _49442_ (_17107_, _17106_, _01726_);
  or _49443_ (_17108_, _25987_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _49444_ (_17109_, _17108_, _16357_);
  and _49445_ (_24804_, _17109_, _17107_);
  and _49446_ (_17110_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _49447_ (_17111_, _16568_, _24426_);
  or _49448_ (_24821_, _17111_, _17110_);
  and _49449_ (_17112_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _49450_ (_17113_, _16572_, _24426_);
  or _49451_ (_24822_, _17113_, _17112_);
  and _49452_ (_17114_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _49453_ (_17115_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _49454_ (_17116_, _17115_, _24426_);
  or _49455_ (_24823_, _17116_, _17114_);
  and _49456_ (_17117_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _49457_ (_17118_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _49458_ (_17119_, _17118_, _24426_);
  or _49459_ (_24824_, _17119_, _17117_);
  and _49460_ (_17120_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _49461_ (_17121_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _49462_ (_17122_, _17121_, _24426_);
  or _49463_ (_24825_, _17122_, _17120_);
  and _49464_ (_17123_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _49465_ (_17124_, _16585_, _24426_);
  or _49466_ (_24826_, _17124_, _17123_);
  and _49467_ (_17125_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _49468_ (_17126_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _49469_ (_17127_, _17126_, _24426_);
  or _49470_ (_24827_, _17127_, _17125_);
  and _49471_ (_24828_, _16408_, _27355_);
  nor _49472_ (_24829_, _16418_, rst);
  and _49473_ (_24831_, _16414_, _27355_);
  or _49474_ (_17128_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand _49475_ (_17129_, _16422_, _26008_);
  and _49476_ (_17130_, _17129_, _27355_);
  and _49477_ (_24832_, _17130_, _17128_);
  or _49478_ (_17131_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand _49479_ (_17132_, _16422_, _26127_);
  and _49480_ (_17133_, _17132_, _27355_);
  and _49481_ (_24833_, _17133_, _17131_);
  or _49482_ (_17134_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _49483_ (_17135_, _16422_, _26105_);
  and _49484_ (_17136_, _17135_, _27355_);
  and _49485_ (_24834_, _17136_, _17134_);
  or _49486_ (_17137_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _49487_ (_17138_, _16422_, _26051_);
  and _49488_ (_17139_, _17138_, _27355_);
  and _49489_ (_24835_, _17139_, _17137_);
  or _49490_ (_17140_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand _49491_ (_17141_, _16422_, _26157_);
  and _49492_ (_17142_, _17141_, _27355_);
  and _49493_ (_24836_, _17142_, _17140_);
  or _49494_ (_17143_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _49495_ (_17144_, _16422_, _26218_);
  and _49496_ (_17145_, _17144_, _27355_);
  and _49497_ (_24837_, _17145_, _17143_);
  or _49498_ (_17146_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _49499_ (_17147_, _16422_, _26251_);
  and _49500_ (_17148_, _17147_, _27355_);
  and _49501_ (_24838_, _17148_, _17146_);
  or _49502_ (_17149_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _49503_ (_17150_, _16422_, _26190_);
  and _49504_ (_17151_, _17150_, _27355_);
  and _49505_ (_24839_, _17151_, _17149_);
  and _49506_ (_17152_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _49507_ (_17153_, _16422_, _25998_);
  or _49508_ (_17154_, _17153_, _17152_);
  and _49509_ (_24840_, _17154_, _27355_);
  and _49510_ (_17155_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _49511_ (_17156_, _16422_, _26135_);
  or _49512_ (_17157_, _17156_, _17155_);
  and _49513_ (_24842_, _17157_, _27355_);
  and _49514_ (_17158_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _49515_ (_17159_, _16422_, _26093_);
  or _49516_ (_17160_, _17159_, _17158_);
  and _49517_ (_24843_, _17160_, _27355_);
  and _49518_ (_17161_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _49519_ (_17162_, _16422_, _26061_);
  or _49520_ (_17163_, _17162_, _17161_);
  and _49521_ (_24844_, _17163_, _27355_);
  and _49522_ (_17164_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _49523_ (_17165_, _16422_, _26163_);
  or _49524_ (_17166_, _17165_, _17164_);
  and _49525_ (_24845_, _17166_, _27355_);
  and _49526_ (_17167_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _49527_ (_17168_, _16422_, _26214_);
  or _49528_ (_17169_, _17168_, _17167_);
  and _49529_ (_24846_, _17169_, _27355_);
  and _49530_ (_17170_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _49531_ (_17171_, _16422_, _26242_);
  or _49532_ (_17172_, _17171_, _17170_);
  and _49533_ (_24847_, _17172_, _27355_);
  and _49534_ (_17173_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _49535_ (_17174_, _16422_, _26195_);
  or _49536_ (_17175_, _17174_, _17173_);
  and _49537_ (_24848_, _17175_, _27355_);
  and _49538_ (_17176_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _49539_ (_17177_, _16422_, _26015_);
  or _49540_ (_17178_, _17177_, _17176_);
  and _49541_ (_24849_, _17178_, _27355_);
  and _49542_ (_17179_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _49543_ (_17180_, _16422_, _26132_);
  or _49544_ (_17181_, _17180_, _17179_);
  and _49545_ (_24850_, _17181_, _27355_);
  and _49546_ (_17182_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _49547_ (_17183_, _16422_, _26097_);
  or _49548_ (_17184_, _17183_, _17182_);
  and _49549_ (_24851_, _17184_, _27355_);
  and _49550_ (_17185_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _49551_ (_17186_, _16422_, _26043_);
  or _49552_ (_17187_, _17186_, _17185_);
  and _49553_ (_24853_, _17187_, _27355_);
  and _49554_ (_17188_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _49555_ (_17189_, _16422_, _26167_);
  or _49556_ (_17190_, _17189_, _17188_);
  and _49557_ (_24854_, _17190_, _27355_);
  and _49558_ (_17191_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _49559_ (_17192_, _16422_, _26222_);
  or _49560_ (_17193_, _17192_, _17191_);
  and _49561_ (_24855_, _17193_, _27355_);
  and _49562_ (_17194_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _49563_ (_17195_, _16422_, _26247_);
  or _49564_ (_17196_, _17195_, _17194_);
  and _49565_ (_24856_, _17196_, _27355_);
  and _49566_ (_17197_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _49567_ (_17198_, _16422_, _26186_);
  or _49568_ (_17199_, _17198_, _17197_);
  and _49569_ (_24857_, _17199_, _27355_);
  and _49570_ (_17200_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _49571_ (_17201_, _16422_, _25994_);
  or _49572_ (_17202_, _17201_, _17200_);
  and _49573_ (_24858_, _17202_, _27355_);
  and _49574_ (_17203_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _49575_ (_17204_, _16422_, _26129_);
  or _49576_ (_17205_, _17204_, _17203_);
  and _49577_ (_24859_, _17205_, _27355_);
  and _49578_ (_17206_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor _49579_ (_17207_, _16422_, _26111_);
  or _49580_ (_17208_, _17207_, _17206_);
  and _49581_ (_24860_, _17208_, _27355_);
  and _49582_ (_17209_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _49583_ (_17210_, _16422_, _26057_);
  or _49584_ (_17211_, _17210_, _17209_);
  and _49585_ (_24861_, _17211_, _27355_);
  and _49586_ (_17212_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _49587_ (_17213_, _16422_, _26159_);
  or _49588_ (_17214_, _17213_, _17212_);
  and _49589_ (_24862_, _17214_, _27355_);
  and _49590_ (_17215_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _49591_ (_17216_, _16422_, _26212_);
  or _49592_ (_17217_, _17216_, _17215_);
  and _49593_ (_24864_, _17217_, _27355_);
  and _49594_ (_17218_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _49595_ (_17219_, _16422_, _26245_);
  or _49596_ (_17220_, _17219_, _17218_);
  and _49597_ (_24865_, _17220_, _27355_);
  and _49598_ (_17221_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49599_ (_17222_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _49600_ (_17223_, _17222_, _17221_);
  and _49601_ (_24866_, _17223_, _27355_);
  and _49602_ (_17224_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49603_ (_17225_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _49604_ (_17226_, _17225_, _17224_);
  and _49605_ (_24867_, _17226_, _27355_);
  and _49606_ (_17227_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49607_ (_17228_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _49608_ (_17229_, _17228_, _17227_);
  and _49609_ (_24868_, _17229_, _27355_);
  and _49610_ (_17230_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49611_ (_17231_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _49612_ (_17232_, _17231_, _17230_);
  and _49613_ (_24869_, _17232_, _27355_);
  and _49614_ (_17233_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49615_ (_17234_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _49616_ (_17235_, _17234_, _17233_);
  and _49617_ (_24870_, _17235_, _27355_);
  and _49618_ (_17236_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49619_ (_17237_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _49620_ (_17238_, _17237_, _17236_);
  and _49621_ (_24871_, _17238_, _27355_);
  and _49622_ (_17239_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _49623_ (_17240_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _49624_ (_17241_, _17240_, _17239_);
  and _49625_ (_24872_, _17241_, _27355_);
  and _49626_ (_17242_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49627_ (_17243_, _01830_, _16438_);
  or _49628_ (_17244_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _49629_ (_17245_, _17244_, _16431_);
  and _49630_ (_17246_, _17245_, _17243_);
  or _49631_ (_17247_, _17246_, _17242_);
  and _49632_ (_24873_, _17247_, _27355_);
  and _49633_ (_17248_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49634_ (_17249_, _01926_, _16438_);
  or _49635_ (_17250_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _49636_ (_17251_, _17250_, _16431_);
  and _49637_ (_17252_, _17251_, _17249_);
  or _49638_ (_17253_, _17252_, _17248_);
  and _49639_ (_24875_, _17253_, _27355_);
  and _49640_ (_17254_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49641_ (_17255_, _02104_, _16438_);
  or _49642_ (_17256_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _49643_ (_17257_, _17256_, _16431_);
  and _49644_ (_17258_, _17257_, _17255_);
  or _49645_ (_17259_, _17258_, _17254_);
  and _49646_ (_24876_, _17259_, _27355_);
  and _49647_ (_17260_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49648_ (_17261_, _01784_, _16438_);
  or _49649_ (_17262_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _49650_ (_17263_, _17262_, _16431_);
  and _49651_ (_17264_, _17263_, _17261_);
  or _49652_ (_17265_, _17264_, _17260_);
  and _49653_ (_24877_, _17265_, _27355_);
  and _49654_ (_17266_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49655_ (_17267_, _01880_, _16438_);
  or _49656_ (_17268_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _49657_ (_17269_, _17268_, _16431_);
  and _49658_ (_17270_, _17269_, _17267_);
  or _49659_ (_17271_, _17270_, _17266_);
  and _49660_ (_24878_, _17271_, _27355_);
  and _49661_ (_17272_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49662_ (_17273_, _02000_, _16438_);
  or _49663_ (_17274_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _49664_ (_17275_, _17274_, _16431_);
  and _49665_ (_17276_, _17275_, _17273_);
  or _49666_ (_17277_, _17276_, _17272_);
  and _49667_ (_24879_, _17277_, _27355_);
  and _49668_ (_17278_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49669_ (_17279_, _02029_, _16438_);
  or _49670_ (_17280_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _49671_ (_17281_, _17280_, _16431_);
  and _49672_ (_17282_, _17281_, _17279_);
  or _49673_ (_17283_, _17282_, _17278_);
  and _49674_ (_24880_, _17283_, _27355_);
  and _49675_ (_17284_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49676_ (_17285_, _01721_, _16438_);
  or _49677_ (_17286_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _49678_ (_17287_, _17286_, _16431_);
  and _49679_ (_17289_, _17287_, _17285_);
  or _49680_ (_17290_, _17289_, _17284_);
  and _49681_ (_24881_, _17290_, _27355_);
  and _49682_ (_17291_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _49683_ (_17292_, _17291_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49684_ (_17293_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _16431_);
  and _49685_ (_17294_, _17293_, _27355_);
  and _49686_ (_24882_, _17294_, _17292_);
  and _49687_ (_17295_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _49688_ (_17296_, _17295_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49689_ (_17298_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _16431_);
  and _49690_ (_17299_, _17298_, _27355_);
  and _49691_ (_24883_, _17299_, _17296_);
  and _49692_ (_17300_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _49693_ (_17301_, _17300_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49694_ (_17302_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _16431_);
  and _49695_ (_17303_, _17302_, _27355_);
  and _49696_ (_24884_, _17303_, _17301_);
  and _49697_ (_17304_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _49698_ (_17305_, _17304_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49699_ (_17307_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _16431_);
  and _49700_ (_17308_, _17307_, _27355_);
  and _49701_ (_24886_, _17308_, _17305_);
  and _49702_ (_17309_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _49703_ (_17310_, _17309_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49704_ (_17311_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _16431_);
  and _49705_ (_17312_, _17311_, _27355_);
  and _49706_ (_24887_, _17312_, _17310_);
  and _49707_ (_17313_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _49708_ (_17314_, _17313_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49709_ (_17316_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _16431_);
  and _49710_ (_17317_, _17316_, _27355_);
  and _49711_ (_24888_, _17317_, _17314_);
  and _49712_ (_17318_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _49713_ (_17319_, _17318_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _49714_ (_17320_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _16431_);
  and _49715_ (_17321_, _17320_, _27355_);
  and _49716_ (_24889_, _17321_, _17319_);
  nand _49717_ (_17322_, _16445_, _25562_);
  or _49718_ (_17323_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _49719_ (_17325_, _17323_, _27355_);
  and _49720_ (_24890_, _17325_, _17322_);
  or _49721_ (_17326_, _16450_, _25639_);
  or _49722_ (_17327_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _49723_ (_17328_, _17327_, _27355_);
  and _49724_ (_24891_, _17328_, _17326_);
  nand _49725_ (_17329_, _16445_, _25704_);
  or _49726_ (_17330_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _49727_ (_17331_, _17330_, _27355_);
  and _49728_ (_24892_, _17331_, _17329_);
  nand _49729_ (_17333_, _16445_, _25769_);
  or _49730_ (_17334_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _49731_ (_17335_, _17334_, _27355_);
  and _49732_ (_24893_, _17335_, _17333_);
  or _49733_ (_17336_, _16450_, _25830_);
  or _49734_ (_17337_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _49735_ (_17338_, _17337_, _27355_);
  and _49736_ (_24894_, _17338_, _17336_);
  or _49737_ (_17339_, _16450_, _25898_);
  or _49738_ (_17340_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _49739_ (_17341_, _17340_, _27355_);
  and _49740_ (_24895_, _17341_, _17339_);
  nand _49741_ (_17342_, _16445_, _25963_);
  or _49742_ (_17343_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _49743_ (_17344_, _17343_, _27355_);
  and _49744_ (_24897_, _17344_, _17342_);
  or _49745_ (_17345_, _16450_, _25441_);
  or _49746_ (_17346_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _49747_ (_17347_, _17346_, _27355_);
  and _49748_ (_24898_, _17347_, _17345_);
  or _49749_ (_17348_, _16450_, _26713_);
  or _49750_ (_17349_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _49751_ (_17350_, _17349_, _27355_);
  and _49752_ (_24899_, _17350_, _17348_);
  nand _49753_ (_17351_, _16445_, _26745_);
  or _49754_ (_17352_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _49755_ (_17353_, _17352_, _27355_);
  and _49756_ (_24900_, _17353_, _17351_);
  nand _49757_ (_17354_, _16445_, _26775_);
  or _49758_ (_17355_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _49759_ (_17356_, _17355_, _27355_);
  and _49760_ (_24901_, _17356_, _17354_);
  nand _49761_ (_17357_, _16445_, _26808_);
  or _49762_ (_17358_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _49763_ (_17359_, _17358_, _27355_);
  and _49764_ (_24902_, _17359_, _17357_);
  or _49765_ (_17360_, _16450_, _26837_);
  or _49766_ (_17361_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _49767_ (_17362_, _17361_, _27355_);
  and _49768_ (_24903_, _17362_, _17360_);
  or _49769_ (_17363_, _16450_, _26867_);
  or _49770_ (_17364_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _49771_ (_17365_, _17364_, _27355_);
  and _49772_ (_24904_, _17365_, _17363_);
  nand _49773_ (_17366_, _16445_, _26898_);
  or _49774_ (_17367_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _49775_ (_17368_, _17367_, _27355_);
  and _49776_ (_24905_, _17368_, _17366_);
  nor _49777_ (_25154_, _01762_, rst);
  and _49778_ (_17369_, _01671_, _01654_);
  nand _49779_ (_17370_, _17369_, _26543_);
  or _49780_ (_17371_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _49781_ (_17372_, _17371_, _27355_);
  and _49782_ (_25156_, _17372_, _17370_);
  not _49783_ (_17373_, _01672_);
  nor _49784_ (_17374_, _17373_, _26543_);
  and _49785_ (_17375_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _49786_ (_17376_, _17375_, _01656_);
  or _49787_ (_17377_, _17376_, _17374_);
  or _49788_ (_17378_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _49789_ (_17379_, _17378_, _27355_);
  and _49790_ (_25157_, _17379_, _17377_);
  and _49791_ (_17380_, _01668_, _01654_);
  not _49792_ (_17381_, _17380_);
  nor _49793_ (_17382_, _17381_, _26543_);
  and _49794_ (_17383_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _49795_ (_17384_, _17383_, _17382_);
  and _49796_ (_25158_, _17384_, _27355_);
  and _49797_ (_17385_, _01676_, _01654_);
  not _49798_ (_17386_, _17385_);
  and _49799_ (_17387_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _49800_ (_17388_, _17386_, _26543_);
  or _49801_ (_17389_, _17388_, _17387_);
  and _49802_ (_25159_, _17389_, _27355_);
  and _49803_ (_17390_, _01678_, _01654_);
  not _49804_ (_17391_, _17390_);
  nor _49805_ (_17392_, _17391_, _26543_);
  and _49806_ (_17393_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _49807_ (_17394_, _17393_, _17392_);
  and _49808_ (_25160_, _17394_, _27355_);
  nand _49809_ (_17395_, _01673_, _01654_);
  or _49810_ (_17396_, _17395_, _01682_);
  or _49811_ (_17397_, _01676_, _01668_);
  or _49812_ (_17398_, _17397_, _01678_);
  and _49813_ (_17399_, _17398_, _01654_);
  or _49814_ (_17400_, _17399_, _17396_);
  and _49815_ (_17401_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  not _49816_ (_17402_, _26543_);
  and _49817_ (_17403_, _01679_, _01654_);
  and _49818_ (_17404_, _17403_, _17402_);
  or _49819_ (_17405_, _17404_, _17401_);
  and _49820_ (_25161_, _17405_, _27355_);
  and _49821_ (_17406_, _01663_, _01654_);
  not _49822_ (_17407_, _17406_);
  and _49823_ (_17408_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _49824_ (_17409_, _17407_, _26543_);
  or _49825_ (_17410_, _17409_, _17408_);
  and _49826_ (_25162_, _17410_, _27355_);
  and _49827_ (_17411_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  not _49828_ (_17412_, _01651_);
  nor _49829_ (_17413_, _17412_, _00755_);
  and _49830_ (_17414_, _17413_, _01654_);
  not _49831_ (_17415_, _17414_);
  nor _49832_ (_17416_, _17415_, _26543_);
  or _49833_ (_17417_, _17416_, _17411_);
  and _49834_ (_25163_, _17417_, _27355_);
  nand _49835_ (_17418_, _17369_, _26521_);
  or _49836_ (_17419_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _49837_ (_17420_, _17419_, _17418_);
  and _49838_ (_25261_, _17420_, _27355_);
  nand _49839_ (_17421_, _17369_, _26512_);
  or _49840_ (_17422_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _49841_ (_17423_, _17422_, _27355_);
  and _49842_ (_25262_, _17423_, _17421_);
  nand _49843_ (_17424_, _17369_, _26505_);
  or _49844_ (_17425_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _49845_ (_17426_, _17425_, _27355_);
  and _49846_ (_25263_, _17426_, _17424_);
  nand _49847_ (_17427_, _17369_, _26497_);
  or _49848_ (_17428_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _49849_ (_17429_, _17428_, _27355_);
  and _49850_ (_25264_, _17429_, _17427_);
  nand _49851_ (_17430_, _17369_, _26489_);
  or _49852_ (_17431_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _49853_ (_17432_, _17431_, _27355_);
  and _49854_ (_25265_, _17432_, _17430_);
  nand _49855_ (_17433_, _17369_, _26482_);
  or _49856_ (_17434_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _49857_ (_17435_, _17434_, _27355_);
  and _49858_ (_25267_, _17435_, _17433_);
  nand _49859_ (_17436_, _17369_, _26475_);
  or _49860_ (_17437_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _49861_ (_17438_, _17437_, _27355_);
  and _49862_ (_25268_, _17438_, _17436_);
  nor _49863_ (_17439_, _01656_, _26521_);
  and _49864_ (_17440_, _17439_, _01672_);
  nand _49865_ (_17441_, _01672_, _01654_);
  and _49866_ (_17442_, _17441_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _49867_ (_17443_, _17442_, _17440_);
  and _49868_ (_25269_, _17443_, _27355_);
  nor _49869_ (_17444_, _17373_, _26512_);
  and _49870_ (_17445_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _49871_ (_17446_, _17445_, _01656_);
  or _49872_ (_17447_, _17446_, _17444_);
  or _49873_ (_17448_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _49874_ (_17449_, _17448_, _27355_);
  and _49875_ (_25270_, _17449_, _17447_);
  nor _49876_ (_17450_, _17373_, _26505_);
  and _49877_ (_17451_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _49878_ (_17452_, _17451_, _01656_);
  or _49879_ (_17453_, _17452_, _17450_);
  or _49880_ (_17454_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _49881_ (_17455_, _17454_, _27355_);
  and _49882_ (_25271_, _17455_, _17453_);
  nor _49883_ (_17456_, _17373_, _26497_);
  and _49884_ (_17457_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _49885_ (_17458_, _17457_, _01656_);
  or _49886_ (_17459_, _17458_, _17456_);
  or _49887_ (_17460_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _49888_ (_17461_, _17460_, _27355_);
  and _49889_ (_25272_, _17461_, _17459_);
  nor _49890_ (_17462_, _17373_, _26489_);
  and _49891_ (_17463_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _49892_ (_17464_, _17463_, _01656_);
  or _49893_ (_17465_, _17464_, _17462_);
  or _49894_ (_17466_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _49895_ (_17467_, _17466_, _27355_);
  and _49896_ (_25273_, _17467_, _17465_);
  nor _49897_ (_17468_, _17373_, _26482_);
  and _49898_ (_17469_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _49899_ (_17470_, _17469_, _01656_);
  or _49900_ (_17471_, _17470_, _17468_);
  or _49901_ (_17472_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _49902_ (_17473_, _17472_, _27355_);
  and _49903_ (_25274_, _17473_, _17471_);
  nor _49904_ (_17474_, _17373_, _26475_);
  and _49905_ (_17475_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _49906_ (_17476_, _17475_, _01656_);
  or _49907_ (_17477_, _17476_, _17474_);
  or _49908_ (_17478_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _49909_ (_17479_, _17478_, _27355_);
  and _49910_ (_25275_, _17479_, _17477_);
  or _49911_ (_17480_, _01674_, _01656_);
  and _49912_ (_17481_, _17480_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand _49913_ (_17482_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _49914_ (_17483_, _17482_, _01673_);
  and _49915_ (_17484_, _17380_, _26522_);
  or _49916_ (_17485_, _17484_, _17483_);
  or _49917_ (_17486_, _17485_, _17481_);
  and _49918_ (_25276_, _17486_, _27355_);
  nor _49919_ (_17487_, _17381_, _26512_);
  and _49920_ (_17488_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _49921_ (_17489_, _17488_, _17487_);
  and _49922_ (_25278_, _17489_, _27355_);
  and _49923_ (_17490_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _49924_ (_17491_, _17381_, _26505_);
  or _49925_ (_17492_, _17491_, _17490_);
  and _49926_ (_25279_, _17492_, _27355_);
  nor _49927_ (_17493_, _17381_, _26497_);
  and _49928_ (_17494_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _49929_ (_17495_, _17494_, _17493_);
  and _49930_ (_25280_, _17495_, _27355_);
  and _49931_ (_17496_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _49932_ (_17497_, _17381_, _26489_);
  or _49933_ (_17498_, _17497_, _17496_);
  and _49934_ (_25281_, _17498_, _27355_);
  nor _49935_ (_17499_, _17381_, _26482_);
  and _49936_ (_17500_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _49937_ (_17501_, _17500_, _17499_);
  and _49938_ (_25282_, _17501_, _27355_);
  nor _49939_ (_17502_, _17381_, _26475_);
  and _49940_ (_17503_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _49941_ (_17504_, _17503_, _17502_);
  and _49942_ (_25283_, _17504_, _27355_);
  and _49943_ (_17505_, _17439_, _01676_);
  and _49944_ (_17506_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _49945_ (_17507_, _17506_, _17505_);
  and _49946_ (_25284_, _17507_, _27355_);
  nor _49947_ (_17508_, _17386_, _26512_);
  and _49948_ (_17509_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _49949_ (_17510_, _17509_, _17508_);
  and _49950_ (_25285_, _17510_, _27355_);
  nor _49951_ (_17511_, _17386_, _26505_);
  and _49952_ (_17512_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _49953_ (_17513_, _17512_, _17511_);
  and _49954_ (_25286_, _17513_, _27355_);
  nor _49955_ (_17514_, _17386_, _26497_);
  and _49956_ (_17515_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _49957_ (_17516_, _17515_, _17514_);
  and _49958_ (_25287_, _17516_, _27355_);
  nor _49959_ (_17517_, _17386_, _26489_);
  and _49960_ (_17518_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _49961_ (_17519_, _17518_, _17517_);
  and _49962_ (_25289_, _17519_, _27355_);
  nor _49963_ (_17520_, _17386_, _26482_);
  and _49964_ (_17521_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _49965_ (_17522_, _17521_, _17520_);
  and _49966_ (_25290_, _17522_, _27355_);
  nor _49967_ (_17523_, _17386_, _26475_);
  and _49968_ (_17524_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _49969_ (_17525_, _17524_, _17523_);
  and _49970_ (_25291_, _17525_, _27355_);
  and _49971_ (_17526_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _49972_ (_17527_, _17439_, _01678_);
  or _49973_ (_17528_, _17527_, _17526_);
  and _49974_ (_25292_, _17528_, _27355_);
  and _49975_ (_17529_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _49976_ (_17530_, _17391_, _26512_);
  or _49977_ (_17531_, _17530_, _17529_);
  and _49978_ (_25293_, _17531_, _27355_);
  and _49979_ (_17532_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _49980_ (_17533_, _17391_, _26505_);
  or _49981_ (_17534_, _17533_, _17532_);
  and _49982_ (_25294_, _17534_, _27355_);
  nor _49983_ (_17535_, _17391_, _26497_);
  and _49984_ (_17536_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _49985_ (_17537_, _17536_, _17535_);
  and _49986_ (_25295_, _17537_, _27355_);
  nor _49987_ (_17538_, _17391_, _26489_);
  and _49988_ (_17539_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _49989_ (_17540_, _17539_, _17538_);
  and _49990_ (_25296_, _17540_, _27355_);
  nor _49991_ (_17541_, _17391_, _26482_);
  and _49992_ (_17542_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _49993_ (_17543_, _17542_, _17541_);
  and _49994_ (_25297_, _17543_, _27355_);
  nor _49995_ (_17544_, _17391_, _26475_);
  and _49996_ (_17545_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or _49997_ (_17546_, _17545_, _17544_);
  and _49998_ (_25298_, _17546_, _27355_);
  and _49999_ (_17547_, _17396_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _50000_ (_17548_, _17439_, _01679_);
  and _50001_ (_17549_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _50002_ (_17550_, _17549_, _17398_);
  or _50003_ (_17551_, _17550_, _17548_);
  or _50004_ (_17552_, _17551_, _17547_);
  and _50005_ (_25300_, _17552_, _27355_);
  and _50006_ (_17553_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  not _50007_ (_17554_, _26512_);
  and _50008_ (_17555_, _17403_, _17554_);
  or _50009_ (_17556_, _17555_, _17553_);
  and _50010_ (_25301_, _17556_, _27355_);
  and _50011_ (_17557_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _50012_ (_17558_, _17403_, _27805_);
  or _50013_ (_17559_, _17558_, _17557_);
  and _50014_ (_25302_, _17559_, _27355_);
  and _50015_ (_17560_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _50016_ (_17561_, _17403_, _27827_);
  or _50017_ (_17562_, _17561_, _17560_);
  and _50018_ (_25303_, _17562_, _27355_);
  and _50019_ (_17563_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _50020_ (_17564_, _17403_, _27829_);
  or _50021_ (_17565_, _17564_, _17563_);
  and _50022_ (_25304_, _17565_, _27355_);
  and _50023_ (_17566_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _50024_ (_17567_, _17403_, _27840_);
  or _50025_ (_17568_, _17567_, _17566_);
  and _50026_ (_25305_, _17568_, _27355_);
  and _50027_ (_17569_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _50028_ (_17570_, _17403_, _27852_);
  or _50029_ (_17571_, _17570_, _17569_);
  and _50030_ (_25306_, _17571_, _27355_);
  and _50031_ (_17572_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _50032_ (_17573_, _17439_, _01663_);
  or _50033_ (_17574_, _17573_, _17572_);
  and _50034_ (_25307_, _17574_, _27355_);
  not _50035_ (_17575_, _01674_);
  or _50036_ (_17576_, _01684_, _17575_);
  and _50037_ (_17577_, _17576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _50038_ (_17578_, _17407_, _26512_);
  nand _50039_ (_17579_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _50040_ (_17580_, _17579_, _01681_);
  or _50041_ (_17581_, _17580_, _17578_);
  or _50042_ (_17582_, _17581_, _17577_);
  and _50043_ (_25308_, _17582_, _27355_);
  and _50044_ (_17583_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _50045_ (_17584_, _17407_, _26505_);
  or _50046_ (_17585_, _17584_, _17583_);
  and _50047_ (_25309_, _17585_, _27355_);
  nor _50048_ (_17586_, _17407_, _26497_);
  nor _50049_ (_17587_, _01681_, _01656_);
  or _50050_ (_17588_, _17587_, _17576_);
  and _50051_ (_17589_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _50052_ (_17590_, _17589_, _17586_);
  and _50053_ (_25311_, _17590_, _27355_);
  and _50054_ (_17591_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor _50055_ (_17592_, _17407_, _26489_);
  or _50056_ (_17593_, _17592_, _17591_);
  and _50057_ (_25312_, _17593_, _27355_);
  nor _50058_ (_17594_, _17407_, _26482_);
  and _50059_ (_17595_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _50060_ (_17596_, _17595_, _17594_);
  and _50061_ (_25313_, _17596_, _27355_);
  nor _50062_ (_17597_, _17407_, _26475_);
  and _50063_ (_17598_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _50064_ (_17599_, _17598_, _17597_);
  and _50065_ (_25314_, _17599_, _27355_);
  nand _50066_ (_17600_, _01677_, _01674_);
  or _50067_ (_17601_, _01685_, _17600_);
  and _50068_ (_17602_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _50069_ (_17603_, _01660_, _26521_);
  nand _50070_ (_17604_, _01680_, _01665_);
  and _50071_ (_17605_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _50072_ (_17606_, _17605_, _17604_);
  or _50073_ (_17607_, _17606_, _17603_);
  or _50074_ (_17608_, _17607_, _17602_);
  and _50075_ (_25315_, _17608_, _27355_);
  and _50076_ (_17609_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _50077_ (_17610_, _17415_, _26512_);
  or _50078_ (_17611_, _17610_, _17609_);
  and _50079_ (_25316_, _17611_, _27355_);
  nor _50080_ (_17612_, _01660_, _26505_);
  and _50081_ (_17613_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _50082_ (_17614_, _17613_, _17612_);
  and _50083_ (_25317_, _17614_, _27355_);
  and _50084_ (_17615_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _50085_ (_17616_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _50086_ (_17617_, _17616_, _17604_);
  nor _50087_ (_17618_, _01660_, _26497_);
  or _50088_ (_17619_, _17618_, _17617_);
  or _50089_ (_17620_, _17619_, _17615_);
  and _50090_ (_25318_, _17620_, _27355_);
  nor _50091_ (_17621_, _01660_, _26489_);
  and _50092_ (_17622_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _50093_ (_17623_, _17622_, _17621_);
  and _50094_ (_25319_, _17623_, _27355_);
  and _50095_ (_17624_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _50096_ (_17625_, _17415_, _26482_);
  or _50097_ (_17626_, _17625_, _17624_);
  and _50098_ (_25320_, _17626_, _27355_);
  and _50099_ (_17627_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _50100_ (_17628_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _50101_ (_17629_, _17628_, _17604_);
  nor _50102_ (_17630_, _01660_, _26475_);
  or _50103_ (_17631_, _17630_, _17629_);
  or _50104_ (_17632_, _17631_, _17627_);
  and _50105_ (_25322_, _17632_, _27355_);
  not _50106_ (_17633_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _50107_ (_17634_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _50108_ (_17635_, _17634_, _17633_);
  and _50109_ (_17636_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _27355_);
  and _50110_ (_25387_, _17636_, _17635_);
  nor _50111_ (_17637_, _17635_, rst);
  nand _50112_ (_17638_, _17634_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _50113_ (_17639_, _17634_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _50114_ (_17640_, _17639_, _17638_);
  and _50115_ (_25388_, _17640_, _17637_);
  nor _50116_ (_17641_, _02004_, _02053_);
  and _50117_ (_17642_, _01811_, _02142_);
  and _50118_ (_17643_, _17642_, _01907_);
  and _50119_ (_17644_, _17643_, _17641_);
  and _50120_ (_17645_, _17644_, _27034_);
  nor _50121_ (_17646_, _17645_, _15901_);
  not _50122_ (_17647_, _01854_);
  and _50123_ (_17648_, _01952_, _17647_);
  and _50124_ (_17649_, _17648_, _27840_);
  or _50125_ (_17650_, _17649_, _02129_);
  nor _50126_ (_17651_, _01952_, _01854_);
  and _50127_ (_17652_, _17651_, _17402_);
  and _50128_ (_17653_, _01952_, _01854_);
  and _50129_ (_17654_, _17653_, _27829_);
  not _50130_ (_17655_, _01952_);
  and _50131_ (_17656_, _17655_, _01854_);
  and _50132_ (_17657_, _17656_, _27852_);
  or _50133_ (_17658_, _17657_, _17654_);
  or _50134_ (_17659_, _17658_, _17652_);
  or _50135_ (_17660_, _17659_, _17650_);
  not _50136_ (_17661_, _02129_);
  and _50137_ (_17662_, _17648_, _17554_);
  or _50138_ (_17663_, _17662_, _17661_);
  and _50139_ (_17664_, _17651_, _27827_);
  and _50140_ (_17665_, _17653_, _26522_);
  and _50141_ (_17666_, _17656_, _27805_);
  or _50142_ (_17667_, _17666_, _17665_);
  or _50143_ (_17668_, _17667_, _17664_);
  or _50144_ (_17669_, _17668_, _17663_);
  nand _50145_ (_17670_, _17669_, _17660_);
  nor _50146_ (_17671_, _17670_, _17646_);
  not _50147_ (_17672_, _02053_);
  and _50148_ (_17673_, _02004_, _17672_);
  not _50149_ (_17674_, _01907_);
  and _50150_ (_17675_, _17642_, _17674_);
  and _50151_ (_17676_, _17675_, _17673_);
  or _50152_ (_17677_, _27115_, _27100_);
  nand _50153_ (_17678_, _27115_, _27100_);
  nand _50154_ (_17679_, _17678_, _17677_);
  nand _50155_ (_17680_, _27071_, _27070_);
  nand _50156_ (_17681_, _27088_, _17680_);
  or _50157_ (_17682_, _27088_, _17680_);
  and _50158_ (_17683_, _17682_, _17681_);
  nand _50159_ (_17684_, _17683_, _17679_);
  or _50160_ (_17685_, _17683_, _17679_);
  nand _50161_ (_17686_, _17685_, _17684_);
  or _50162_ (_17687_, _27135_, _27125_);
  nand _50163_ (_17688_, _27135_, _27125_);
  nand _50164_ (_17689_, _17688_, _17687_);
  nand _50165_ (_17690_, _27146_, _27060_);
  or _50166_ (_17691_, _27146_, _27060_);
  and _50167_ (_17692_, _17691_, _17690_);
  nand _50168_ (_17693_, _17692_, _17689_);
  or _50169_ (_17694_, _17692_, _17689_);
  nand _50170_ (_17695_, _17694_, _17693_);
  nand _50171_ (_17696_, _17695_, _17686_);
  or _50172_ (_17697_, _17695_, _17686_);
  nand _50173_ (_17698_, _17697_, _17696_);
  nand _50174_ (_17699_, _17698_, _02129_);
  or _50175_ (_17700_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _50176_ (_17701_, _17700_, _17653_);
  and _50177_ (_17702_, _17701_, _17699_);
  and _50178_ (_17703_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _50179_ (_17704_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _50180_ (_17705_, _17704_, _17703_);
  and _50181_ (_17706_, _17705_, _17661_);
  and _50182_ (_17707_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _50183_ (_17708_, _02129_, _26928_);
  or _50184_ (_17709_, _17708_, _17707_);
  and _50185_ (_17710_, _17709_, _17651_);
  and _50186_ (_17711_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _50187_ (_17712_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _50188_ (_17713_, _17712_, _17711_);
  and _50189_ (_17714_, _17713_, _02129_);
  or _50190_ (_17715_, _17714_, _17710_);
  or _50191_ (_17716_, _17715_, _17706_);
  or _50192_ (_17717_, _17716_, _17702_);
  and _50193_ (_17718_, _17717_, _17676_);
  not _50194_ (_17719_, _17642_);
  and _50195_ (_17720_, _17673_, _01907_);
  or _50196_ (_17721_, _17720_, _17719_);
  nor _50197_ (_17722_, _01811_, _01748_);
  and _50198_ (_17723_, _17722_, _01907_);
  and _50199_ (_17724_, _17723_, _17673_);
  not _50200_ (_17725_, _01811_);
  and _50201_ (_17726_, _02053_, _02142_);
  nand _50202_ (_17727_, _17726_, _17725_);
  nand _50203_ (_17728_, _17727_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _50204_ (_17729_, _17728_, _17724_);
  and _50205_ (_17730_, _17729_, _17721_);
  and _50206_ (_17731_, _17675_, _17641_);
  and _50207_ (_17732_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _50208_ (_17733_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _50209_ (_17734_, _17733_, _17732_);
  and _50210_ (_17735_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _50211_ (_17736_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _50212_ (_17737_, _17736_, _17735_);
  or _50213_ (_17738_, _17737_, _17734_);
  and _50214_ (_17739_, _17738_, _17731_);
  and _50215_ (_17740_, _17722_, _17674_);
  nor _50216_ (_17741_, _02004_, _17672_);
  and _50217_ (_17742_, _17741_, _17740_);
  and _50218_ (_17743_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _50219_ (_17744_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _50220_ (_17745_, _17744_, _17743_);
  and _50221_ (_17746_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _50222_ (_17747_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _50223_ (_17748_, _17747_, _17746_);
  or _50224_ (_17749_, _17748_, _17745_);
  and _50225_ (_17750_, _17749_, _17742_);
  or _50226_ (_17751_, _17750_, _17739_);
  and _50227_ (_17752_, _17751_, _02129_);
  or _50228_ (_17753_, _17752_, _17730_);
  and _50229_ (_17754_, _15895_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nor _50230_ (_17755_, _15349_, _26307_);
  and _50231_ (_17756_, _17755_, _15420_);
  nor _50232_ (_17757_, _15418_, _26402_);
  and _50233_ (_17758_, _26327_, _26374_);
  not _50234_ (_17759_, _17758_);
  and _50235_ (_17760_, _17759_, _17757_);
  and _50236_ (_17761_, _26281_, _26322_);
  nor _50237_ (_17762_, _17761_, _26347_);
  not _50238_ (_17763_, _15351_);
  and _50239_ (_17764_, _17763_, _26321_);
  and _50240_ (_17765_, _17764_, _17762_);
  and _50241_ (_17766_, _17765_, _17760_);
  and _50242_ (_17767_, _17766_, _15673_);
  and _50243_ (_17768_, _17767_, _17756_);
  and _50244_ (_17769_, _17768_, _26305_);
  nor _50245_ (_17770_, _17769_, _26393_);
  or _50246_ (_17771_, _17770_, p2_in[4]);
  not _50247_ (_17772_, _17770_);
  or _50248_ (_17773_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _50249_ (_17774_, _17773_, _17771_);
  and _50250_ (_17775_, _17774_, _17653_);
  or _50251_ (_17776_, _17775_, _02129_);
  or _50252_ (_17777_, _17770_, p2_in[7]);
  or _50253_ (_17778_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _50254_ (_17779_, _17778_, _17777_);
  and _50255_ (_17780_, _17779_, _17651_);
  or _50256_ (_17781_, _17770_, p2_in[5]);
  or _50257_ (_17782_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _50258_ (_17783_, _17782_, _17781_);
  and _50259_ (_17784_, _17783_, _17648_);
  or _50260_ (_17785_, _17770_, p2_in[6]);
  or _50261_ (_17786_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _50262_ (_17787_, _17786_, _17785_);
  and _50263_ (_17788_, _17787_, _17656_);
  or _50264_ (_17789_, _17788_, _17784_);
  or _50265_ (_17790_, _17789_, _17780_);
  or _50266_ (_17791_, _17790_, _17776_);
  and _50267_ (_17792_, _17741_, _17643_);
  nor _50268_ (_17793_, _17770_, p2_in[0]);
  and _50269_ (_17794_, _17770_, _27415_);
  nor _50270_ (_17795_, _17794_, _17793_);
  and _50271_ (_17796_, _17795_, _17653_);
  or _50272_ (_17797_, _17796_, _17661_);
  or _50273_ (_17798_, _17770_, p2_in[2]);
  or _50274_ (_17799_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _50275_ (_17800_, _17799_, _17798_);
  and _50276_ (_17801_, _17800_, _17656_);
  or _50277_ (_17802_, _17770_, p2_in[1]);
  or _50278_ (_17803_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _50279_ (_17804_, _17803_, _17802_);
  and _50280_ (_17805_, _17804_, _17648_);
  or _50281_ (_17806_, _17770_, p2_in[3]);
  or _50282_ (_17807_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _50283_ (_17808_, _17807_, _17806_);
  and _50284_ (_17809_, _17808_, _17651_);
  or _50285_ (_17810_, _17809_, _17805_);
  or _50286_ (_17811_, _17810_, _17801_);
  or _50287_ (_17812_, _17811_, _17797_);
  and _50288_ (_17813_, _17812_, _17792_);
  and _50289_ (_17814_, _17813_, _17791_);
  or _50290_ (_17815_, _17814_, _17754_);
  and _50291_ (_17816_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _50292_ (_17817_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _50293_ (_17818_, _17817_, _17816_);
  and _50294_ (_17819_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _50295_ (_17820_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _50296_ (_17821_, _17820_, _17819_);
  or _50297_ (_17822_, _17821_, _17818_);
  and _50298_ (_17823_, _17822_, _17742_);
  and _50299_ (_17825_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _50300_ (_17826_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _50301_ (_17827_, _17826_, _17825_);
  and _50302_ (_17828_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _50303_ (_17829_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _50304_ (_17830_, _17829_, _17828_);
  or _50305_ (_17831_, _17830_, _17827_);
  and _50306_ (_17832_, _17831_, _17731_);
  or _50307_ (_17833_, _17832_, _17823_);
  and _50308_ (_17834_, _17833_, _17661_);
  and _50309_ (_17835_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _50310_ (_17836_, _17835_, _02129_);
  and _50311_ (_17837_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _50312_ (_17838_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _50313_ (_17839_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _50314_ (_17840_, _17839_, _17838_);
  or _50315_ (_17841_, _17840_, _17837_);
  or _50316_ (_17842_, _17841_, _17836_);
  and _50317_ (_17843_, _02004_, _02053_);
  and _50318_ (_17844_, _17740_, _17843_);
  and _50319_ (_17845_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _50320_ (_17846_, _17845_, _17661_);
  and _50321_ (_17847_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _50322_ (_17848_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _50323_ (_17849_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _50324_ (_17850_, _17849_, _17848_);
  or _50325_ (_17851_, _17850_, _17847_);
  or _50326_ (_17852_, _17851_, _17846_);
  and _50327_ (_17853_, _17852_, _17844_);
  and _50328_ (_17854_, _17853_, _17842_);
  or _50329_ (_17855_, _17854_, _17834_);
  or _50330_ (_17856_, _17855_, _17815_);
  or _50331_ (_17857_, _17856_, _17753_);
  or _50332_ (_17858_, _17770_, p0_in[2]);
  or _50333_ (_17859_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _50334_ (_17860_, _17859_, _17858_);
  and _50335_ (_17861_, _17860_, _17656_);
  nor _50336_ (_17862_, _17770_, p0_in[0]);
  and _50337_ (_17863_, _17770_, _27220_);
  nor _50338_ (_17864_, _17863_, _17862_);
  and _50339_ (_17865_, _17864_, _17653_);
  or _50340_ (_17866_, _17865_, _17861_);
  or _50341_ (_17867_, _17770_, p0_in[3]);
  or _50342_ (_17868_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _50343_ (_17869_, _17868_, _17867_);
  and _50344_ (_17870_, _17869_, _17651_);
  or _50345_ (_17871_, _17770_, p0_in[1]);
  or _50346_ (_17872_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _50347_ (_17873_, _17872_, _17871_);
  and _50348_ (_17874_, _17873_, _17648_);
  or _50349_ (_17875_, _17874_, _17870_);
  or _50350_ (_17876_, _17875_, _17866_);
  and _50351_ (_17877_, _17876_, _17643_);
  or _50352_ (_17878_, _17770_, p1_in[3]);
  or _50353_ (_17879_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _50354_ (_17880_, _17879_, _17878_);
  and _50355_ (_17881_, _17880_, _17651_);
  or _50356_ (_17882_, _17770_, p1_in[1]);
  or _50357_ (_17883_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _50358_ (_17884_, _17883_, _17882_);
  and _50359_ (_17885_, _17884_, _17648_);
  or _50360_ (_17886_, _17885_, _17881_);
  or _50361_ (_17887_, _17770_, p1_in[2]);
  or _50362_ (_17888_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _50363_ (_17889_, _17888_, _17887_);
  and _50364_ (_17890_, _17889_, _17656_);
  nor _50365_ (_17891_, _17770_, p1_in[0]);
  and _50366_ (_17892_, _17770_, _27321_);
  nor _50367_ (_17893_, _17892_, _17891_);
  and _50368_ (_17894_, _17893_, _17653_);
  or _50369_ (_17895_, _17894_, _17890_);
  or _50370_ (_17896_, _17895_, _17886_);
  and _50371_ (_17897_, _17896_, _17675_);
  or _50372_ (_17898_, _17897_, _17877_);
  and _50373_ (_17899_, _17898_, _02129_);
  or _50374_ (_17900_, _17770_, p1_in[6]);
  or _50375_ (_17901_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _50376_ (_17902_, _17901_, _17900_);
  and _50377_ (_17903_, _17902_, _17656_);
  or _50378_ (_17904_, _17770_, p1_in[4]);
  or _50379_ (_17905_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _50380_ (_17906_, _17905_, _17904_);
  and _50381_ (_17907_, _17906_, _17653_);
  or _50382_ (_17908_, _17907_, _17903_);
  or _50383_ (_17909_, _17770_, p1_in[7]);
  or _50384_ (_17910_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _50385_ (_17911_, _17910_, _17909_);
  and _50386_ (_17912_, _17911_, _17651_);
  or _50387_ (_17913_, _17770_, p1_in[5]);
  or _50388_ (_17914_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _50389_ (_17915_, _17914_, _17913_);
  and _50390_ (_17916_, _17915_, _17648_);
  or _50391_ (_17917_, _17916_, _17912_);
  or _50392_ (_17918_, _17917_, _17908_);
  and _50393_ (_17919_, _17918_, _17675_);
  or _50394_ (_17920_, _17770_, p0_in[6]);
  or _50395_ (_17921_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _50396_ (_17922_, _17921_, _17920_);
  and _50397_ (_17923_, _17922_, _17656_);
  or _50398_ (_17924_, _17770_, p0_in[4]);
  or _50399_ (_17925_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _50400_ (_17926_, _17925_, _17924_);
  and _50401_ (_17927_, _17926_, _17653_);
  or _50402_ (_17928_, _17927_, _17923_);
  or _50403_ (_17929_, _17770_, p0_in[7]);
  or _50404_ (_17930_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _50405_ (_17931_, _17930_, _17929_);
  and _50406_ (_17932_, _17931_, _17651_);
  or _50407_ (_17933_, _17770_, p0_in[5]);
  or _50408_ (_17934_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _50409_ (_17935_, _17934_, _17933_);
  and _50410_ (_17936_, _17935_, _17648_);
  or _50411_ (_17937_, _17936_, _17932_);
  or _50412_ (_17938_, _17937_, _17928_);
  and _50413_ (_17939_, _17938_, _17643_);
  or _50414_ (_17940_, _17939_, _17919_);
  and _50415_ (_17941_, _17940_, _17661_);
  or _50416_ (_17942_, _17941_, _17899_);
  and _50417_ (_17943_, _17942_, _17843_);
  and _50418_ (_17944_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _50419_ (_17945_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _50420_ (_17946_, _17945_, _17944_);
  and _50421_ (_17947_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _50422_ (_17948_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _50423_ (_17949_, _17948_, _17947_);
  or _50424_ (_17950_, _17949_, _17946_);
  and _50425_ (_17951_, _17950_, _17741_);
  and _50426_ (_17952_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _50427_ (_17953_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _50428_ (_17954_, _17953_, _17952_);
  and _50429_ (_17955_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _50430_ (_17956_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _50431_ (_17957_, _17956_, _17955_);
  or _50432_ (_17958_, _17957_, _17954_);
  and _50433_ (_17959_, _17958_, _17843_);
  or _50434_ (_17960_, _17959_, _17951_);
  and _50435_ (_17961_, _17960_, _02129_);
  and _50436_ (_17962_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _50437_ (_17963_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _50438_ (_17964_, _17963_, _17962_);
  and _50439_ (_17965_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _50440_ (_17966_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _50441_ (_17967_, _17966_, _17965_);
  or _50442_ (_17968_, _17967_, _17964_);
  and _50443_ (_17969_, _17968_, _17843_);
  and _50444_ (_17970_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _50445_ (_17971_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _50446_ (_17972_, _17971_, _17970_);
  and _50447_ (_17973_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _50448_ (_17974_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _50449_ (_17975_, _17974_, _17973_);
  or _50450_ (_17976_, _17975_, _17972_);
  and _50451_ (_17977_, _17976_, _17741_);
  or _50452_ (_17978_, _17977_, _17969_);
  and _50453_ (_17979_, _17978_, _17661_);
  or _50454_ (_17980_, _17979_, _17961_);
  and _50455_ (_17981_, _17980_, _17723_);
  nor _50456_ (_17982_, _17770_, p3_in[0]);
  and _50457_ (_17983_, _17770_, _27499_);
  nor _50458_ (_17984_, _17983_, _17982_);
  and _50459_ (_17985_, _17984_, _17653_);
  or _50460_ (_17986_, _17985_, _17661_);
  or _50461_ (_17987_, _17770_, p3_in[2]);
  or _50462_ (_17988_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _50463_ (_17989_, _17988_, _17987_);
  and _50464_ (_17990_, _17989_, _17656_);
  or _50465_ (_17991_, _17770_, p3_in[3]);
  or _50466_ (_17992_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _50467_ (_17993_, _17992_, _17991_);
  and _50468_ (_17994_, _17993_, _17651_);
  or _50469_ (_17995_, _17770_, p3_in[1]);
  or _50470_ (_17996_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _50471_ (_17997_, _17996_, _17995_);
  and _50472_ (_17998_, _17997_, _17648_);
  or _50473_ (_17999_, _17998_, _17994_);
  or _50474_ (_18000_, _17999_, _17990_);
  or _50475_ (_18001_, _18000_, _17986_);
  and _50476_ (_18002_, _17741_, _17675_);
  or _50477_ (_18003_, _17770_, p3_in[4]);
  or _50478_ (_18004_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _50479_ (_18005_, _18004_, _18003_);
  and _50480_ (_18006_, _18005_, _17653_);
  or _50481_ (_18007_, _18006_, _02129_);
  or _50482_ (_18008_, _17770_, p3_in[6]);
  or _50483_ (_18009_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _50484_ (_18010_, _18009_, _18008_);
  and _50485_ (_18011_, _18010_, _17656_);
  or _50486_ (_18012_, _17770_, p3_in[7]);
  or _50487_ (_18013_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _50488_ (_18014_, _18013_, _18012_);
  and _50489_ (_18015_, _18014_, _17651_);
  or _50490_ (_18016_, _17770_, p3_in[5]);
  or _50491_ (_18017_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _50492_ (_18018_, _18017_, _18016_);
  and _50493_ (_18019_, _18018_, _17648_);
  or _50494_ (_18020_, _18019_, _18015_);
  or _50495_ (_18021_, _18020_, _18011_);
  or _50496_ (_18022_, _18021_, _18007_);
  and _50497_ (_18023_, _18022_, _18002_);
  and _50498_ (_18024_, _18023_, _18001_);
  and _50499_ (_18025_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _50500_ (_18026_, _18025_, _02129_);
  and _50501_ (_18027_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _50502_ (_18028_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _50503_ (_18029_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _50504_ (_18030_, _18029_, _18028_);
  or _50505_ (_18031_, _18030_, _18027_);
  or _50506_ (_18032_, _18031_, _18026_);
  and _50507_ (_18033_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _50508_ (_18034_, _18033_, _17661_);
  and _50509_ (_18035_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _50510_ (_18036_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _50511_ (_18037_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _50512_ (_18038_, _18037_, _18036_);
  or _50513_ (_18039_, _18038_, _18035_);
  or _50514_ (_18040_, _18039_, _18034_);
  and _50515_ (_18041_, _18040_, _17724_);
  and _50516_ (_18042_, _18041_, _18032_);
  and _50517_ (_18043_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _50518_ (_18044_, _18043_, _02129_);
  and _50519_ (_18045_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _50520_ (_18046_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _50521_ (_18047_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _50522_ (_18048_, _18047_, _18046_);
  or _50523_ (_18049_, _18048_, _18045_);
  or _50524_ (_18050_, _18049_, _18044_);
  and _50525_ (_18051_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _50526_ (_18052_, _18051_, _17661_);
  and _50527_ (_18053_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _50528_ (_18054_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _50529_ (_18055_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _50530_ (_18056_, _18055_, _18054_);
  or _50531_ (_18057_, _18056_, _18053_);
  or _50532_ (_18058_, _18057_, _18052_);
  and _50533_ (_18059_, _18058_, _17644_);
  and _50534_ (_18060_, _18059_, _18050_);
  or _50535_ (_18061_, _18060_, _18042_);
  or _50536_ (_18062_, _18061_, _18024_);
  or _50537_ (_18063_, _18062_, _17981_);
  or _50538_ (_18064_, _18063_, _17943_);
  or _50539_ (_18065_, _18064_, _17857_);
  or _50540_ (_18066_, _18065_, _17718_);
  nand _50541_ (_18067_, _17754_, _25514_);
  and _50542_ (_18068_, _18067_, _17646_);
  and _50543_ (_18069_, _18068_, _18066_);
  or _50544_ (_18070_, _18069_, _17671_);
  and _50545_ (_25389_, _18070_, _27355_);
  and _50546_ (_18071_, _02129_, _01811_);
  and _50547_ (_18072_, _18071_, _17653_);
  and _50548_ (_18073_, _01907_, _02142_);
  and _50549_ (_18074_, _18073_, _17641_);
  and _50550_ (_18075_, _18074_, _18072_);
  and _50551_ (_18076_, _18075_, _27034_);
  and _50552_ (_18077_, _17651_, _17661_);
  not _50553_ (_18078_, _18077_);
  and _50554_ (_18079_, _18078_, _27048_);
  and _50555_ (_18080_, _18079_, _15882_);
  nor _50556_ (_18081_, _18080_, _18076_);
  and _50557_ (_18082_, _18081_, _15898_);
  and _50558_ (_18083_, _17843_, _18073_);
  and _50559_ (_18084_, _18071_, _17651_);
  and _50560_ (_18085_, _18084_, _18083_);
  and _50561_ (_18086_, _18085_, _26591_);
  and _50562_ (_18087_, _17674_, _02004_);
  and _50563_ (_18088_, _18072_, _02142_);
  and _50564_ (_18089_, _18088_, _17672_);
  and _50565_ (_18090_, _18089_, _18087_);
  and _50566_ (_18091_, _18090_, _26933_);
  and _50567_ (_18092_, _18075_, _27044_);
  or _50568_ (_18093_, _18092_, _18091_);
  nor _50569_ (_18094_, _18093_, _18086_);
  nor _50570_ (_18095_, _18094_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _50571_ (_18096_, _18095_);
  and _50572_ (_18097_, _18096_, _18082_);
  and _50573_ (_18098_, _18071_, _17656_);
  and _50574_ (_18099_, _18098_, _18083_);
  and _50575_ (_18100_, _18099_, _26591_);
  or _50576_ (_18101_, _18100_, rst);
  nor _50577_ (_25391_, _18101_, _18097_);
  not _50578_ (_18102_, _18100_);
  not _50579_ (_18103_, _18090_);
  and _50580_ (_18104_, _02129_, _17725_);
  and _50581_ (_18105_, _18104_, _17651_);
  and _50582_ (_18106_, _18105_, _18083_);
  and _50583_ (_18107_, _18104_, _17653_);
  and _50584_ (_18108_, _18087_, _17726_);
  and _50585_ (_18109_, _18108_, _18107_);
  nor _50586_ (_18110_, _18109_, _18106_);
  and _50587_ (_18111_, _18107_, _18083_);
  nor _50588_ (_18112_, _02129_, _01811_);
  and _50589_ (_18113_, _18112_, _17653_);
  and _50590_ (_18114_, _18113_, _18083_);
  nor _50591_ (_18115_, _18114_, _18111_);
  and _50592_ (_18116_, _18115_, _18110_);
  and _50593_ (_18117_, _17741_, _18073_);
  and _50594_ (_18118_, _18117_, _18107_);
  and _50595_ (_18119_, _18112_, _17648_);
  and _50596_ (_18120_, _18119_, _18083_);
  nor _50597_ (_18121_, _18120_, _18118_);
  and _50598_ (_18122_, _18104_, _17656_);
  and _50599_ (_18123_, _18122_, _18083_);
  and _50600_ (_18124_, _18104_, _17648_);
  and _50601_ (_18125_, _18124_, _18108_);
  nor _50602_ (_18126_, _18125_, _18123_);
  and _50603_ (_18127_, _18126_, _18121_);
  and _50604_ (_18128_, _18127_, _18116_);
  and _50605_ (_18129_, _18128_, _18103_);
  and _50606_ (_18130_, _17673_, _18073_);
  and _50607_ (_18131_, _18130_, _18113_);
  and _50608_ (_18132_, _18130_, _18105_);
  and _50609_ (_18133_, _18077_, _01811_);
  and _50610_ (_18134_, _18133_, _18083_);
  or _50611_ (_18135_, _18134_, _18132_);
  nor _50612_ (_18136_, _18135_, _18131_);
  and _50613_ (_18137_, _18130_, _18119_);
  and _50614_ (_18138_, _18130_, _18122_);
  nor _50615_ (_18139_, _18138_, _18137_);
  nor _50616_ (_18140_, _01907_, _02004_);
  and _50617_ (_18141_, _18140_, _17726_);
  nand _50618_ (_18142_, _18141_, _18133_);
  not _50619_ (_18143_, _18071_);
  nand _50620_ (_18144_, _18083_, _17648_);
  or _50621_ (_18145_, _18144_, _18143_);
  and _50622_ (_18146_, _18145_, _18142_);
  and _50623_ (_18147_, _18146_, _18139_);
  not _50624_ (_18148_, _18104_);
  or _50625_ (_18149_, _18144_, _18148_);
  nor _50626_ (_18150_, _18099_, _18085_);
  and _50627_ (_18151_, _18150_, _18149_);
  and _50628_ (_18152_, _18130_, _18107_);
  not _50629_ (_18153_, _17673_);
  and _50630_ (_18154_, _18088_, _18153_);
  nor _50631_ (_18155_, _18154_, _18152_);
  and _50632_ (_18156_, _18155_, _18151_);
  and _50633_ (_18157_, _18156_, _18147_);
  and _50634_ (_18158_, _18157_, _18136_);
  and _50635_ (_18159_, _18158_, _18129_);
  not _50636_ (_18160_, _18159_);
  nand _50637_ (_18161_, _18160_, _18097_);
  and _50638_ (_18162_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _50639_ (_18163_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _50640_ (_18164_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _50641_ (_18165_, _18164_, _18163_);
  and _50642_ (_18166_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _50643_ (_18167_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _50644_ (_18168_, _18167_, _18166_);
  or _50645_ (_18169_, _18168_, _18165_);
  and _50646_ (_18170_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _50647_ (_18171_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _50648_ (_18172_, _18171_, _18170_);
  and _50649_ (_18173_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _50650_ (_18174_, _18141_, _18133_);
  and _50651_ (_18175_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _50652_ (_18176_, _18175_, _18173_);
  or _50653_ (_18177_, _18176_, _18172_);
  or _50654_ (_18178_, _18177_, _18169_);
  and _50655_ (_18179_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _50656_ (_18180_, _18124_, _18083_);
  and _50657_ (_18181_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _50658_ (_18182_, _18181_, _18179_);
  and _50659_ (_18183_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _50660_ (_18184_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _50661_ (_18185_, _18184_, _18183_);
  or _50662_ (_18186_, _18185_, _18182_);
  and _50663_ (_18187_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _50664_ (_18188_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _50665_ (_18189_, _18188_, _18187_);
  and _50666_ (_18190_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _50667_ (_18191_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _50668_ (_18192_, _18191_, _18190_);
  or _50669_ (_18193_, _18192_, _18189_);
  or _50670_ (_18194_, _18193_, _18186_);
  or _50671_ (_18195_, _18194_, _18178_);
  and _50672_ (_18196_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _50673_ (_18197_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or _50674_ (_18198_, _18197_, _18196_);
  and _50675_ (_18199_, _18140_, _18089_);
  and _50676_ (_18200_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _50677_ (_18201_, _18071_, _17648_);
  and _50678_ (_18202_, _18201_, _18083_);
  and _50679_ (_18203_, _18202_, _26545_);
  or _50680_ (_18204_, _18203_, _18200_);
  or _50681_ (_18205_, _18204_, _18198_);
  and _50682_ (_18206_, _18083_, _18072_);
  and _50683_ (_18207_, _18206_, _17931_);
  and _50684_ (_18208_, _18108_, _18072_);
  and _50685_ (_18209_, _18208_, _17911_);
  or _50686_ (_18210_, _18209_, _18207_);
  and _50687_ (_18211_, _18141_, _18072_);
  and _50688_ (_18212_, _18211_, _18014_);
  and _50689_ (_18213_, _18117_, _18072_);
  and _50690_ (_18214_, _18213_, _17779_);
  or _50691_ (_18215_, _18214_, _18212_);
  or _50692_ (_18216_, _18215_, _18210_);
  or _50693_ (_18217_, _18216_, _18205_);
  and _50694_ (_18218_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _50695_ (_18219_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _50696_ (_18220_, _18219_, _18218_);
  or _50697_ (_18221_, _18220_, _18217_);
  or _50698_ (_18222_, _18221_, _18195_);
  and _50699_ (_18223_, _18222_, _18097_);
  or _50700_ (_18224_, _18223_, _18162_);
  and _50701_ (_18225_, _18224_, _18102_);
  and _50702_ (_18226_, _18100_, _25441_);
  or _50703_ (_18227_, _18226_, _18225_);
  and _50704_ (_25392_, _18227_, _27355_);
  nor _50705_ (_25485_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _50706_ (_18228_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _50707_ (_18229_, _17634_, rst);
  and _50708_ (_25486_, _18229_, _18228_);
  nor _50709_ (_18230_, _17634_, _17633_);
  or _50710_ (_18231_, _18230_, _17635_);
  and _50711_ (_18232_, _17638_, _27355_);
  and _50712_ (_25487_, _18232_, _18231_);
  or _50713_ (_18233_, _18103_, _17698_);
  nand _50714_ (_18234_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _50715_ (_18235_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _50716_ (_18236_, _18235_, _18234_);
  nand _50717_ (_18237_, _18206_, _17864_);
  nand _50718_ (_18238_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _50719_ (_18239_, _18238_, _18237_);
  and _50720_ (_18240_, _18239_, _18236_);
  nand _50721_ (_18241_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand _50722_ (_18242_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _50723_ (_18243_, _18242_, _18241_);
  nand _50724_ (_18244_, _18211_, _17984_);
  nand _50725_ (_18245_, _18213_, _17795_);
  and _50726_ (_18246_, _18245_, _18244_);
  and _50727_ (_18247_, _18246_, _18243_);
  and _50728_ (_18248_, _18247_, _18240_);
  nand _50729_ (_18249_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _50730_ (_18250_, _18208_, _17893_);
  nand _50731_ (_18251_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _50732_ (_18252_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _50733_ (_18253_, _18252_, _18251_);
  and _50734_ (_18254_, _18253_, _18250_);
  and _50735_ (_18255_, _18254_, _18249_);
  and _50736_ (_18256_, _18255_, _18248_);
  nand _50737_ (_18257_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand _50738_ (_18258_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _50739_ (_18259_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _50740_ (_18260_, _18259_, _18258_);
  and _50741_ (_18261_, _18260_, _18257_);
  nand _50742_ (_18262_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _50743_ (_18263_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _50744_ (_18264_, _18263_, _18262_);
  nand _50745_ (_18265_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _50746_ (_18266_, _18145_, _26553_);
  and _50747_ (_18267_, _18266_, _18265_);
  and _50748_ (_18268_, _18267_, _18264_);
  nand _50749_ (_18269_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _50750_ (_18270_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _50751_ (_18271_, _18270_, _18269_);
  nand _50752_ (_18272_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _50753_ (_18273_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _50754_ (_18274_, _18273_, _18272_);
  and _50755_ (_18275_, _18274_, _18271_);
  nand _50756_ (_18276_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _50757_ (_18277_, _18149_, _27720_);
  and _50758_ (_18278_, _18277_, _18276_);
  and _50759_ (_18279_, _18278_, _18275_);
  and _50760_ (_18280_, _18279_, _18268_);
  and _50761_ (_18281_, _18280_, _18261_);
  and _50762_ (_18282_, _18281_, _18256_);
  nand _50763_ (_18283_, _18282_, _18233_);
  and _50764_ (_18284_, _18283_, _18097_);
  and _50765_ (_18285_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _50766_ (_18286_, _18285_, _18100_);
  or _50767_ (_18287_, _18286_, _18284_);
  nand _50768_ (_18288_, _18100_, _25562_);
  and _50769_ (_18289_, _18288_, _27355_);
  and _50770_ (_25488_, _18289_, _18287_);
  and _50771_ (_18290_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _50772_ (_18291_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _50773_ (_18292_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _50774_ (_18293_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _50775_ (_18294_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _50776_ (_18295_, _18294_, _18293_);
  or _50777_ (_18296_, _18295_, _18292_);
  or _50778_ (_18297_, _18296_, _18291_);
  or _50779_ (_18298_, _18297_, _18290_);
  and _50780_ (_18299_, _18213_, _17804_);
  and _50781_ (_18300_, _18211_, _17997_);
  or _50782_ (_18301_, _18300_, _18299_);
  and _50783_ (_18302_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _50784_ (_18303_, _18208_, _17884_);
  or _50785_ (_18304_, _18303_, _18302_);
  or _50786_ (_18305_, _18304_, _18301_);
  and _50787_ (_18306_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _50788_ (_18307_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _50789_ (_18308_, _18307_, _18306_);
  or _50790_ (_18309_, _18308_, _18305_);
  and _50791_ (_18310_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _50792_ (_18311_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _50793_ (_18312_, _18311_, _18310_);
  and _50794_ (_18313_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _50795_ (_18314_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or _50796_ (_18315_, _18314_, _18313_);
  or _50797_ (_18316_, _18315_, _18312_);
  and _50798_ (_18317_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _50799_ (_18318_, _18206_, _17873_);
  or _50800_ (_18319_, _18318_, _18317_);
  and _50801_ (_18320_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _50802_ (_18321_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _50803_ (_18322_, _18321_, _18320_);
  or _50804_ (_18323_, _18322_, _18319_);
  or _50805_ (_18324_, _18323_, _18316_);
  or _50806_ (_18325_, _18324_, _18309_);
  and _50807_ (_18326_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _50808_ (_18327_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _50809_ (_18328_, _18149_, _27701_);
  or _50810_ (_18329_, _18328_, _18327_);
  or _50811_ (_18330_, _18329_, _18326_);
  and _50812_ (_18331_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _50813_ (_18332_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _50814_ (_18333_, _18332_, _18331_);
  and _50815_ (_18334_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _50816_ (_18335_, _18145_, _26559_);
  or _50817_ (_18336_, _18335_, _18334_);
  or _50818_ (_18337_, _18336_, _18333_);
  or _50819_ (_18338_, _18337_, _18330_);
  or _50820_ (_18339_, _18338_, _18325_);
  or _50821_ (_18340_, _18339_, _18298_);
  and _50822_ (_18341_, _18340_, _18097_);
  and _50823_ (_18342_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _50824_ (_18343_, _18342_, _18341_);
  or _50825_ (_18344_, _18343_, _18100_);
  or _50826_ (_18345_, _18102_, _25639_);
  and _50827_ (_18346_, _18345_, _27355_);
  and _50828_ (_25489_, _18346_, _18344_);
  and _50829_ (_18347_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _50830_ (_18348_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _50831_ (_18349_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _50832_ (_18350_, _18349_, _18348_);
  and _50833_ (_18351_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _50834_ (_18352_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _50835_ (_18353_, _18352_, _18351_);
  or _50836_ (_18354_, _18353_, _18350_);
  and _50837_ (_18355_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _50838_ (_18356_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _50839_ (_18357_, _18356_, _18355_);
  and _50840_ (_18358_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _50841_ (_18359_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _50842_ (_18360_, _18359_, _18358_);
  or _50843_ (_18361_, _18360_, _18357_);
  or _50844_ (_18362_, _18361_, _18354_);
  and _50845_ (_18363_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _50846_ (_18364_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _50847_ (_18365_, _18364_, _18363_);
  and _50848_ (_18366_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _50849_ (_18367_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _50850_ (_18368_, _18367_, _18366_);
  or _50851_ (_18369_, _18368_, _18365_);
  and _50852_ (_18370_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _50853_ (_18371_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _50854_ (_18372_, _18371_, _18370_);
  and _50855_ (_18373_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _50856_ (_18374_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _50857_ (_18375_, _18374_, _18373_);
  or _50858_ (_18376_, _18375_, _18372_);
  or _50859_ (_18377_, _18376_, _18369_);
  or _50860_ (_18378_, _18377_, _18362_);
  and _50861_ (_18379_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _50862_ (_18380_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _50863_ (_18381_, _18380_, _18379_);
  and _50864_ (_18382_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _50865_ (_18383_, _18202_, _02108_);
  or _50866_ (_18384_, _18383_, _18382_);
  or _50867_ (_18385_, _18384_, _18381_);
  and _50868_ (_18386_, _18211_, _17989_);
  and _50869_ (_18387_, _18213_, _17800_);
  or _50870_ (_18388_, _18387_, _18386_);
  and _50871_ (_18389_, _18206_, _17860_);
  and _50872_ (_18390_, _18208_, _17889_);
  or _50873_ (_18391_, _18390_, _18389_);
  or _50874_ (_18392_, _18391_, _18388_);
  or _50875_ (_18393_, _18392_, _18385_);
  and _50876_ (_18394_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _50877_ (_18395_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _50878_ (_18396_, _18395_, _18394_);
  or _50879_ (_18397_, _18396_, _18393_);
  or _50880_ (_18398_, _18397_, _18378_);
  and _50881_ (_18399_, _18398_, _18097_);
  or _50882_ (_18400_, _18399_, _18100_);
  or _50883_ (_18401_, _18400_, _18347_);
  nand _50884_ (_18402_, _18100_, _25704_);
  and _50885_ (_18403_, _18402_, _27355_);
  and _50886_ (_25490_, _18403_, _18401_);
  and _50887_ (_18404_, _18208_, _17880_);
  and _50888_ (_18405_, _18206_, _17869_);
  and _50889_ (_18406_, _18213_, _17808_);
  or _50890_ (_18407_, _18406_, _18405_);
  or _50891_ (_18408_, _18407_, _18404_);
  and _50892_ (_18409_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _50893_ (_18410_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _50894_ (_18411_, _18410_, _18409_);
  and _50895_ (_18412_, _18211_, _17993_);
  nor _50896_ (_18413_, _18145_, _26571_);
  or _50897_ (_18414_, _18413_, _18412_);
  or _50898_ (_18415_, _18414_, _18411_);
  or _50899_ (_18416_, _18415_, _18408_);
  and _50900_ (_18417_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _50901_ (_18418_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _50902_ (_18419_, _18418_, _18417_);
  and _50903_ (_18420_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _50904_ (_18421_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _50905_ (_18422_, _18421_, _18420_);
  or _50906_ (_18423_, _18422_, _18419_);
  and _50907_ (_18424_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _50908_ (_18425_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _50909_ (_18426_, _18425_, _18424_);
  and _50910_ (_18427_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _50911_ (_18428_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _50912_ (_18429_, _18428_, _18427_);
  or _50913_ (_18430_, _18429_, _18426_);
  or _50914_ (_18431_, _18430_, _18423_);
  and _50915_ (_18432_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _50916_ (_18433_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _50917_ (_18434_, _18433_, _18432_);
  and _50918_ (_18435_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _50919_ (_18436_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _50920_ (_18437_, _18436_, _18435_);
  or _50921_ (_18438_, _18437_, _18434_);
  and _50922_ (_18439_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _50923_ (_18440_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _50924_ (_18441_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _50925_ (_18442_, _18441_, _18440_);
  or _50926_ (_18443_, _18442_, _18439_);
  and _50927_ (_18444_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _50928_ (_18445_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _50929_ (_18446_, _18445_, _18444_);
  and _50930_ (_18447_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _50931_ (_18448_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _50932_ (_18449_, _18448_, _18447_);
  or _50933_ (_18450_, _18449_, _18446_);
  or _50934_ (_18451_, _18450_, _18443_);
  or _50935_ (_18452_, _18451_, _18438_);
  or _50936_ (_18453_, _18452_, _18431_);
  or _50937_ (_18454_, _18453_, _18416_);
  and _50938_ (_18455_, _18454_, _18097_);
  and _50939_ (_18456_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or _50940_ (_18457_, _18456_, _18455_);
  or _50941_ (_18458_, _18457_, _18100_);
  nand _50942_ (_18459_, _18100_, _25769_);
  and _50943_ (_18460_, _18459_, _27355_);
  and _50944_ (_25492_, _18460_, _18458_);
  and _50945_ (_18461_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _50946_ (_18462_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _50947_ (_18463_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _50948_ (_18464_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _50949_ (_18465_, _18464_, _18463_);
  and _50950_ (_18466_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _50951_ (_18467_, _18466_, _18465_);
  or _50952_ (_18468_, _18467_, _18462_);
  or _50953_ (_18469_, _18468_, _18461_);
  and _50954_ (_18470_, _18208_, _17906_);
  and _50955_ (_18471_, _18206_, _17926_);
  or _50956_ (_18472_, _18471_, _18470_);
  and _50957_ (_18473_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _50958_ (_18474_, _18213_, _17774_);
  or _50959_ (_18475_, _18474_, _18473_);
  or _50960_ (_18476_, _18475_, _18472_);
  and _50961_ (_18477_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _50962_ (_18478_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _50963_ (_18479_, _18478_, _18477_);
  or _50964_ (_18480_, _18479_, _18476_);
  and _50965_ (_18481_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _50966_ (_18482_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _50967_ (_18483_, _18482_, _18481_);
  and _50968_ (_18484_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _50969_ (_18485_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _50970_ (_18486_, _18485_, _18484_);
  or _50971_ (_18487_, _18486_, _18483_);
  and _50972_ (_18488_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _50973_ (_18489_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or _50974_ (_18490_, _18489_, _18488_);
  and _50975_ (_18491_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _50976_ (_18492_, _18211_, _18005_);
  or _50977_ (_18493_, _18492_, _18491_);
  or _50978_ (_18494_, _18493_, _18490_);
  or _50979_ (_18495_, _18494_, _18487_);
  or _50980_ (_18496_, _18495_, _18480_);
  nor _50981_ (_18497_, _18149_, _27580_);
  and _50982_ (_18498_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _50983_ (_18499_, _18145_, _26577_);
  or _50984_ (_18500_, _18499_, _18498_);
  or _50985_ (_18501_, _18500_, _18497_);
  and _50986_ (_18502_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _50987_ (_18503_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _50988_ (_18504_, _18503_, _18502_);
  and _50989_ (_18505_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _50990_ (_18506_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _50991_ (_18507_, _18506_, _18505_);
  or _50992_ (_18508_, _18507_, _18504_);
  or _50993_ (_18509_, _18508_, _18501_);
  or _50994_ (_18510_, _18509_, _18496_);
  or _50995_ (_18511_, _18510_, _18469_);
  and _50996_ (_18512_, _18511_, _18097_);
  and _50997_ (_18513_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _50998_ (_18514_, _18513_, _18512_);
  or _50999_ (_18515_, _18514_, _18100_);
  or _51000_ (_18516_, _18102_, _25830_);
  and _51001_ (_18517_, _18516_, _27355_);
  and _51002_ (_25493_, _18517_, _18515_);
  and _51003_ (_18518_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _51004_ (_18519_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _51005_ (_18520_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _51006_ (_18521_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _51007_ (_18522_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _51008_ (_18523_, _18522_, _18521_);
  or _51009_ (_18524_, _18523_, _18520_);
  or _51010_ (_18525_, _18524_, _18519_);
  or _51011_ (_18526_, _18525_, _18518_);
  and _51012_ (_18527_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _51013_ (_18528_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _51014_ (_18529_, _18528_, _18527_);
  and _51015_ (_18530_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _51016_ (_18531_, _18208_, _17915_);
  or _51017_ (_18532_, _18531_, _18530_);
  or _51018_ (_18533_, _18532_, _18529_);
  and _51019_ (_18534_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _51020_ (_18535_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _51021_ (_18536_, _18535_, _18534_);
  or _51022_ (_18537_, _18536_, _18533_);
  and _51023_ (_18538_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _51024_ (_18539_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _51025_ (_18540_, _18539_, _18538_);
  and _51026_ (_18541_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _51027_ (_18542_, _18211_, _18018_);
  or _51028_ (_18543_, _18542_, _18541_);
  or _51029_ (_18544_, _18543_, _18540_);
  and _51030_ (_18545_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _51031_ (_18546_, _18213_, _17783_);
  or _51032_ (_18547_, _18546_, _18545_);
  and _51033_ (_18548_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _51034_ (_18549_, _18206_, _17935_);
  or _51035_ (_18550_, _18549_, _18548_);
  or _51036_ (_18551_, _18550_, _18547_);
  or _51037_ (_18552_, _18551_, _18544_);
  or _51038_ (_18553_, _18552_, _18537_);
  and _51039_ (_18554_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _51040_ (_18555_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _51041_ (_18556_, _18145_, _26583_);
  or _51042_ (_18557_, _18556_, _18555_);
  or _51043_ (_18558_, _18557_, _18554_);
  and _51044_ (_18559_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _51045_ (_18560_, _18149_, _27582_);
  or _51046_ (_18561_, _18560_, _18559_);
  and _51047_ (_18562_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _51048_ (_18563_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _51049_ (_18564_, _18563_, _18562_);
  or _51050_ (_18565_, _18564_, _18561_);
  or _51051_ (_18566_, _18565_, _18558_);
  or _51052_ (_18567_, _18566_, _18553_);
  or _51053_ (_18568_, _18567_, _18526_);
  and _51054_ (_18569_, _18568_, _18097_);
  and _51055_ (_18570_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _51056_ (_18571_, _18570_, _18569_);
  or _51057_ (_18572_, _18571_, _18100_);
  or _51058_ (_18573_, _18102_, _25898_);
  and _51059_ (_18574_, _18573_, _27355_);
  and _51060_ (_25494_, _18574_, _18572_);
  nand _51061_ (_18575_, _18100_, _25963_);
  and _51062_ (_18576_, _18575_, _27355_);
  and _51063_ (_18577_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _51064_ (_18578_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _51065_ (_18579_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _51066_ (_18580_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _51067_ (_18581_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _51068_ (_18582_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or _51069_ (_18583_, _18582_, _18581_);
  or _51070_ (_18584_, _18583_, _18580_);
  or _51071_ (_18585_, _18584_, _18579_);
  or _51072_ (_18586_, _18585_, _18578_);
  and _51073_ (_18587_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _51074_ (_18588_, _18211_, _18010_);
  or _51075_ (_18589_, _18588_, _18587_);
  and _51076_ (_18590_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _51077_ (_18591_, _18208_, _17902_);
  or _51078_ (_18592_, _18591_, _18590_);
  or _51079_ (_18593_, _18592_, _18589_);
  and _51080_ (_18594_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _51081_ (_18595_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _51082_ (_18596_, _18595_, _18594_);
  or _51083_ (_18597_, _18596_, _18593_);
  and _51084_ (_18598_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _51085_ (_18599_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _51086_ (_18600_, _18599_, _18598_);
  and _51087_ (_18601_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _51088_ (_18602_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _51089_ (_18603_, _18602_, _18601_);
  or _51090_ (_18604_, _18603_, _18600_);
  and _51091_ (_18605_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _51092_ (_18606_, _18213_, _17787_);
  or _51093_ (_18607_, _18606_, _18605_);
  and _51094_ (_18608_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _51095_ (_18609_, _18206_, _17922_);
  or _51096_ (_18610_, _18609_, _18608_);
  or _51097_ (_18611_, _18610_, _18607_);
  or _51098_ (_18612_, _18611_, _18604_);
  or _51099_ (_18613_, _18612_, _18597_);
  and _51100_ (_18614_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _51101_ (_18615_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _51102_ (_18616_, _18145_, _26589_);
  or _51103_ (_18617_, _18616_, _18615_);
  or _51104_ (_18618_, _18617_, _18614_);
  and _51105_ (_18619_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _51106_ (_18620_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _51107_ (_18621_, _18620_, _18619_);
  and _51108_ (_18622_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _51109_ (_18623_, _18149_, _27591_);
  or _51110_ (_18624_, _18623_, _18622_);
  or _51111_ (_18625_, _18624_, _18621_);
  or _51112_ (_18626_, _18625_, _18618_);
  or _51113_ (_18627_, _18626_, _18613_);
  or _51114_ (_18628_, _18627_, _18586_);
  and _51115_ (_18629_, _18628_, _18097_);
  or _51116_ (_18630_, _18629_, _18577_);
  or _51117_ (_18631_, _18630_, _18100_);
  and _51118_ (_25495_, _18631_, _18576_);
  and _51119_ (_25567_, _02141_, _27355_);
  and _51120_ (_25568_, _03058_, _27355_);
  nor _51121_ (_25571_, _02129_, rst);
  and _51122_ (_25586_, _02983_, _27355_);
  and _51123_ (_25587_, _02997_, _27355_);
  and _51124_ (_25588_, _03007_, _27355_);
  and _51125_ (_25589_, _03016_, _27355_);
  and _51126_ (_25590_, _03026_, _27355_);
  and _51127_ (_25591_, _03036_, _27355_);
  and _51128_ (_25592_, _03047_, _27355_);
  nor _51129_ (_25593_, _01854_, rst);
  nor _51130_ (_25594_, _01952_, rst);
  nor _51131_ (_18632_, _16708_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _51132_ (_18633_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _51133_ (_18634_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _18633_);
  nor _51134_ (_18635_, _18634_, _18632_);
  not _51135_ (_18636_, _18635_);
  nor _51136_ (_18637_, _16726_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _51137_ (_18638_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _18633_);
  nor _51138_ (_18639_, _18638_, _18637_);
  nor _51139_ (_18640_, _18639_, _18636_);
  and _51140_ (_18641_, _18640_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _51141_ (_18642_, _18639_, _18635_);
  and _51142_ (_18643_, _18642_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _51143_ (_18644_, _18643_, _18641_);
  and _51144_ (_18645_, _18639_, _18636_);
  and _51145_ (_18646_, _18645_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _51146_ (_18647_, _18639_, _18635_);
  and _51147_ (_18648_, _18647_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _51148_ (_18649_, _18648_, _18646_);
  and _51149_ (_18650_, _18649_, _18644_);
  nor _51150_ (_18651_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _51151_ (_18652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _18633_);
  nor _51152_ (_18653_, _18652_, _18651_);
  nor _51153_ (_18654_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _51154_ (_18655_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _18633_);
  nor _51155_ (_18656_, _18655_, _18654_);
  nor _51156_ (_18657_, _18656_, _18653_);
  not _51157_ (_18658_, _18657_);
  nor _51158_ (_18659_, _18658_, _18650_);
  and _51159_ (_18660_, _18642_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _51160_ (_18661_, _18647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _51161_ (_18662_, _18661_, _18660_);
  and _51162_ (_18663_, _18645_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51163_ (_18664_, _18640_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _51164_ (_18665_, _18664_, _18663_);
  and _51165_ (_18666_, _18665_, _18662_);
  and _51166_ (_18667_, _18656_, _18653_);
  not _51167_ (_18668_, _18667_);
  nor _51168_ (_18669_, _18668_, _18666_);
  nor _51169_ (_18670_, _18669_, _18659_);
  and _51170_ (_18671_, _18642_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _51171_ (_18672_, _18647_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _51172_ (_18673_, _18672_, _18671_);
  and _51173_ (_18674_, _18645_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _51174_ (_18675_, _18640_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _51175_ (_18676_, _18675_, _18674_);
  and _51176_ (_18677_, _18676_, _18673_);
  not _51177_ (_18678_, _18653_);
  and _51178_ (_18679_, _18656_, _18678_);
  not _51179_ (_18680_, _18679_);
  nor _51180_ (_18681_, _18680_, _18677_);
  and _51181_ (_18682_, _18640_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _51182_ (_18683_, _18647_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _51183_ (_18684_, _18683_, _18682_);
  and _51184_ (_18685_, _18645_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _51185_ (_18686_, _18642_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _51186_ (_18687_, _18686_, _18685_);
  and _51187_ (_18688_, _18687_, _18684_);
  not _51188_ (_18689_, _18656_);
  and _51189_ (_18690_, _18689_, _18653_);
  not _51190_ (_18691_, _18690_);
  nor _51191_ (_18692_, _18691_, _18688_);
  nor _51192_ (_18693_, _18692_, _18681_);
  and _51193_ (_18694_, _18693_, _18670_);
  not _51194_ (_18695_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _51195_ (_18696_, _18653_, _18695_);
  or _51196_ (_18697_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _51197_ (_18698_, _18697_, _18696_);
  not _51198_ (_18699_, _18639_);
  and _51199_ (_18700_, _18656_, _18635_);
  and _51200_ (_18701_, _18700_, _18699_);
  and _51201_ (_18702_, _18701_, _18698_);
  not _51202_ (_18703_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _51203_ (_18704_, _18653_, _18703_);
  or _51204_ (_18705_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _51205_ (_18706_, _18705_, _18704_);
  and _51206_ (_18707_, _18700_, _18639_);
  and _51207_ (_18708_, _18707_, _18706_);
  or _51208_ (_18709_, _18708_, _18702_);
  and _51209_ (_18710_, _18689_, _18635_);
  not _51210_ (_18711_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _51211_ (_18712_, _18653_, _18711_);
  or _51212_ (_18713_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _51213_ (_18714_, _18713_, _18712_);
  and _51214_ (_18715_, _18714_, _18639_);
  not _51215_ (_18716_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _51216_ (_18717_, _18653_, _18716_);
  or _51217_ (_18718_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _51218_ (_18719_, _18718_, _18717_);
  and _51219_ (_18720_, _18719_, _18699_);
  or _51220_ (_18721_, _18720_, _18715_);
  and _51221_ (_18722_, _18721_, _18710_);
  not _51222_ (_18723_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _51223_ (_18724_, _18653_, _18723_);
  or _51224_ (_18725_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _51225_ (_18726_, _18725_, _18724_);
  and _51226_ (_18727_, _18726_, _18656_);
  not _51227_ (_18728_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _51228_ (_18729_, _18653_, _18728_);
  or _51229_ (_18730_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _51230_ (_18731_, _18730_, _18729_);
  and _51231_ (_18732_, _18731_, _18689_);
  or _51232_ (_18733_, _18732_, _18727_);
  and _51233_ (_18734_, _18733_, _18639_);
  not _51234_ (_18735_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _51235_ (_18736_, _18653_, _18735_);
  or _51236_ (_18737_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _51237_ (_18738_, _18737_, _18736_);
  and _51238_ (_18739_, _18738_, _18656_);
  not _51239_ (_18740_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _51240_ (_18741_, _18653_, _18740_);
  or _51241_ (_18742_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _51242_ (_18743_, _18742_, _18741_);
  and _51243_ (_18744_, _18743_, _18689_);
  nor _51244_ (_18745_, _18744_, _18739_);
  nor _51245_ (_18746_, _18745_, _18639_);
  or _51246_ (_18747_, _18746_, _18734_);
  and _51247_ (_18748_, _18747_, _18636_);
  or _51248_ (_18749_, _18748_, _18722_);
  nor _51249_ (_18750_, _18749_, _18709_);
  nor _51250_ (_18751_, _18750_, _18694_);
  and _51251_ (_18752_, _18694_, word_in[7]);
  or _51252_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _18752_, _18751_);
  and _51253_ (_18753_, _18667_, _18635_);
  nor _51254_ (_18754_, _18753_, _18699_);
  and _51255_ (_18755_, _18667_, _18640_);
  nor _51256_ (_18756_, _18755_, _18754_);
  nor _51257_ (_18757_, _18667_, _18635_);
  nor _51258_ (_18758_, _18757_, _18753_);
  not _51259_ (_18759_, _18758_);
  and _51260_ (_18760_, _18759_, _18756_);
  and _51261_ (_18761_, _18760_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _51262_ (_18762_, _18761_);
  not _51263_ (_18763_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _51264_ (_18764_, _18756_, _18763_);
  nor _51265_ (_18765_, _18756_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _51266_ (_18766_, _18765_, _18759_);
  and _51267_ (_18767_, _18766_, _18764_);
  nor _51268_ (_18768_, _18758_, _18756_);
  and _51269_ (_18769_, _18768_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _51270_ (_18770_, _18769_, _18767_);
  and _51271_ (_18771_, _18770_, _18762_);
  nor _51272_ (_18772_, _18771_, _18658_);
  and _51273_ (_18773_, _18760_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _51274_ (_18774_, _18773_);
  not _51275_ (_18775_, _18756_);
  or _51276_ (_18776_, _18775_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _51277_ (_18777_, _18756_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _51278_ (_18778_, _18777_, _18759_);
  and _51279_ (_18779_, _18778_, _18776_);
  and _51280_ (_18780_, _18768_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _51281_ (_18781_, _18780_, _18779_);
  and _51282_ (_18782_, _18781_, _18774_);
  nor _51283_ (_18783_, _18782_, _18680_);
  nor _51284_ (_18784_, _18783_, _18772_);
  and _51285_ (_18785_, _18760_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _51286_ (_18786_, _18785_);
  not _51287_ (_18787_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _51288_ (_18788_, _18756_, _18787_);
  nor _51289_ (_18789_, _18756_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _51290_ (_18790_, _18789_, _18759_);
  and _51291_ (_18791_, _18790_, _18788_);
  and _51292_ (_18792_, _18768_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _51293_ (_18793_, _18792_, _18791_);
  and _51294_ (_18794_, _18793_, _18786_);
  nor _51295_ (_18795_, _18794_, _18668_);
  and _51296_ (_18796_, _18760_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _51297_ (_18797_, _18796_);
  not _51298_ (_18798_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _51299_ (_18799_, _18756_, _18798_);
  nor _51300_ (_18800_, _18756_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _51301_ (_18801_, _18800_, _18759_);
  and _51302_ (_18802_, _18801_, _18799_);
  and _51303_ (_18803_, _18768_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _51304_ (_18804_, _18803_, _18802_);
  and _51305_ (_18805_, _18804_, _18797_);
  nor _51306_ (_18806_, _18805_, _18691_);
  nor _51307_ (_18807_, _18806_, _18795_);
  and _51308_ (_18808_, _18807_, _18784_);
  or _51309_ (_18809_, _18667_, _18657_);
  not _51310_ (_18810_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _51311_ (_18811_, _18653_, _18810_);
  or _51312_ (_18812_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _51313_ (_18813_, _18812_, _18811_);
  and _51314_ (_18814_, _18813_, _18809_);
  not _51315_ (_18815_, _18809_);
  and _51316_ (_18816_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor _51317_ (_18817_, _18653_, _18735_);
  or _51318_ (_18818_, _18817_, _18816_);
  and _51319_ (_18819_, _18818_, _18815_);
  or _51320_ (_18820_, _18819_, _18814_);
  or _51321_ (_18821_, _18820_, _18758_);
  not _51322_ (_18822_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _51323_ (_18823_, _18653_, _18822_);
  or _51324_ (_18824_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _51325_ (_18825_, _18824_, _18823_);
  and _51326_ (_18826_, _18825_, _18809_);
  not _51327_ (_18827_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _51328_ (_18828_, _18653_, _18827_);
  or _51329_ (_18829_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _51330_ (_18830_, _18829_, _18828_);
  and _51331_ (_18831_, _18830_, _18815_);
  nor _51332_ (_18832_, _18831_, _18826_);
  nand _51333_ (_18833_, _18832_, _18758_);
  and _51334_ (_18834_, _18833_, _18756_);
  and _51335_ (_18835_, _18834_, _18821_);
  not _51336_ (_18836_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _51337_ (_18837_, _18653_, _18836_);
  or _51338_ (_18838_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _51339_ (_18839_, _18838_, _18837_);
  and _51340_ (_18840_, _18839_, _18809_);
  not _51341_ (_18841_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _51342_ (_18842_, _18653_, _18841_);
  or _51343_ (_18843_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _51344_ (_18844_, _18843_, _18842_);
  and _51345_ (_18845_, _18844_, _18815_);
  or _51346_ (_18846_, _18845_, _18840_);
  or _51347_ (_18847_, _18846_, _18758_);
  not _51348_ (_18848_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _51349_ (_18849_, _18653_, _18848_);
  or _51350_ (_18850_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _51351_ (_18851_, _18850_, _18849_);
  and _51352_ (_18852_, _18851_, _18809_);
  not _51353_ (_18853_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _51354_ (_18854_, _18653_, _18853_);
  or _51355_ (_18855_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _51356_ (_18856_, _18855_, _18854_);
  and _51357_ (_18857_, _18856_, _18815_);
  nor _51358_ (_18858_, _18857_, _18852_);
  nand _51359_ (_18859_, _18858_, _18758_);
  nand _51360_ (_18860_, _18859_, _18847_);
  nor _51361_ (_18861_, _18860_, _18756_);
  nor _51362_ (_18862_, _18861_, _18835_);
  nor _51363_ (_18863_, _18862_, _18808_);
  and _51364_ (_18864_, _18808_, word_in[15]);
  or _51365_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _18864_, _18863_);
  not _51366_ (_18865_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _51367_ (_18866_, _18701_);
  or _51368_ (_18867_, _18700_, _18699_);
  and _51369_ (_18868_, _18867_, _18866_);
  and _51370_ (_18869_, _18868_, _18865_);
  and _51371_ (_18870_, _18689_, _18642_);
  nor _51372_ (_18871_, _18707_, _18870_);
  not _51373_ (_18872_, _18871_);
  nor _51374_ (_18873_, _18689_, _18635_);
  nor _51375_ (_18874_, _18873_, _18710_);
  and _51376_ (_18875_, _18874_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _51377_ (_18876_, _18875_, _18872_);
  nor _51378_ (_18877_, _18876_, _18869_);
  and _51379_ (_18878_, _18868_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _51380_ (_18879_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _51381_ (_18880_, _18868_, _18879_);
  nor _51382_ (_18881_, _18880_, _18878_);
  nor _51383_ (_18882_, _18881_, _18636_);
  nor _51384_ (_18883_, _18882_, _18877_);
  nor _51385_ (_18884_, _18883_, _18656_);
  and _51386_ (_18885_, _18868_, _18763_);
  not _51387_ (_18886_, _18873_);
  not _51388_ (_18887_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _51389_ (_18888_, _18639_, _18887_);
  nor _51390_ (_18889_, _18888_, _18886_);
  not _51391_ (_18891_, _18889_);
  nor _51392_ (_18892_, _18891_, _18885_);
  not _51393_ (_18894_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _51394_ (_18895_, _18868_, _18894_);
  and _51395_ (_18897_, _18700_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _51396_ (_18898_, _18897_, _18707_);
  nor _51397_ (_18900_, _18898_, _18895_);
  or _51398_ (_18901_, _18900_, _18678_);
  or _51399_ (_18903_, _18901_, _18892_);
  nor _51400_ (_18904_, _18903_, _18884_);
  not _51401_ (_18906_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _51402_ (_18907_, _18868_, _18906_);
  and _51403_ (_18909_, _18874_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _51404_ (_18910_, _18909_, _18872_);
  nor _51405_ (_18912_, _18910_, _18907_);
  and _51406_ (_18913_, _18868_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not _51407_ (_18915_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _51408_ (_18916_, _18868_, _18915_);
  nor _51409_ (_18918_, _18916_, _18913_);
  nor _51410_ (_18919_, _18918_, _18636_);
  nor _51411_ (_18921_, _18919_, _18912_);
  nor _51412_ (_18922_, _18921_, _18656_);
  and _51413_ (_18924_, _18868_, _18787_);
  not _51414_ (_18925_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _51415_ (_18927_, _18639_, _18925_);
  nor _51416_ (_18928_, _18927_, _18886_);
  not _51417_ (_18929_, _18928_);
  nor _51418_ (_18930_, _18929_, _18924_);
  not _51419_ (_18931_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _51420_ (_18932_, _18868_, _18931_);
  and _51421_ (_18933_, _18700_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _51422_ (_18934_, _18933_, _18707_);
  nor _51423_ (_18935_, _18934_, _18932_);
  or _51424_ (_18936_, _18935_, _18653_);
  or _51425_ (_18937_, _18936_, _18930_);
  nor _51426_ (_18938_, _18937_, _18922_);
  nor _51427_ (_18939_, _18938_, _18904_);
  or _51428_ (_18940_, _18738_, _18656_);
  or _51429_ (_18941_, _18743_, _18689_);
  and _51430_ (_18942_, _18941_, _18940_);
  and _51431_ (_18943_, _18942_, _18874_);
  and _51432_ (_18944_, _18710_, _18698_);
  and _51433_ (_18945_, _18719_, _18873_);
  or _51434_ (_18946_, _18945_, _18944_);
  or _51435_ (_18947_, _18946_, _18943_);
  and _51436_ (_18948_, _18947_, _18868_);
  or _51437_ (_18949_, _18726_, _18656_);
  or _51438_ (_18950_, _18731_, _18689_);
  and _51439_ (_18951_, _18950_, _18949_);
  and _51440_ (_18952_, _18951_, _18874_);
  and _51441_ (_18953_, _18710_, _18706_);
  and _51442_ (_18954_, _18714_, _18873_);
  or _51443_ (_18955_, _18954_, _18953_);
  nor _51444_ (_18956_, _18955_, _18952_);
  nor _51445_ (_18957_, _18956_, _18868_);
  or _51446_ (_18958_, _18957_, _18948_);
  and _51447_ (_18959_, _18958_, _18939_);
  not _51448_ (_18960_, _18939_);
  and _51449_ (_18961_, _18960_, word_in[23]);
  or _51450_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _18961_, _18959_);
  and _51451_ (_18962_, _18658_, _18635_);
  nor _51452_ (_18963_, _18658_, _18635_);
  nor _51453_ (_18964_, _18963_, _18962_);
  and _51454_ (_18965_, _18962_, _18639_);
  nor _51455_ (_18966_, _18962_, _18639_);
  nor _51456_ (_18967_, _18966_, _18965_);
  nor _51457_ (_18968_, _18967_, _18865_);
  and _51458_ (_18969_, _18967_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _51459_ (_18970_, _18969_, _18968_);
  nor _51460_ (_18971_, _18970_, _18964_);
  nand _51461_ (_18972_, _18967_, _18879_);
  not _51462_ (_18973_, _18964_);
  nor _51463_ (_18974_, _18967_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _51464_ (_18975_, _18974_, _18973_);
  and _51465_ (_18976_, _18975_, _18972_);
  nor _51466_ (_18977_, _18976_, _18971_);
  nor _51467_ (_18978_, _18977_, _18658_);
  nor _51468_ (_18979_, _18967_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not _51469_ (_18980_, _18979_);
  nor _51470_ (_18981_, _18973_, _18888_);
  and _51471_ (_18982_, _18981_, _18980_);
  nor _51472_ (_18983_, _18967_, _18894_);
  and _51473_ (_18985_, _18967_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _51474_ (_18987_, _18985_, _18983_);
  nor _51475_ (_18988_, _18987_, _18964_);
  nor _51476_ (_18990_, _18988_, _18982_);
  nor _51477_ (_18991_, _18990_, _18680_);
  nor _51478_ (_18993_, _18991_, _18978_);
  nor _51479_ (_18994_, _18967_, _18906_);
  and _51480_ (_18996_, _18967_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _51481_ (_18997_, _18996_, _18994_);
  nor _51482_ (_18999_, _18997_, _18964_);
  nand _51483_ (_19000_, _18967_, _18915_);
  nor _51484_ (_19002_, _18967_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _51485_ (_19003_, _19002_, _18973_);
  and _51486_ (_19005_, _19003_, _19000_);
  nor _51487_ (_19006_, _19005_, _18999_);
  nor _51488_ (_19008_, _19006_, _18668_);
  nor _51489_ (_19009_, _18967_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not _51490_ (_19011_, _19009_);
  nor _51491_ (_19012_, _18973_, _18927_);
  and _51492_ (_19014_, _19012_, _19011_);
  nor _51493_ (_19015_, _18967_, _18931_);
  and _51494_ (_19017_, _18967_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _51495_ (_19018_, _19017_, _19015_);
  nor _51496_ (_19020_, _19018_, _18964_);
  nor _51497_ (_19021_, _19020_, _19014_);
  nor _51498_ (_19022_, _19021_, _18691_);
  nor _51499_ (_19023_, _19022_, _19008_);
  and _51500_ (_19024_, _19023_, _18993_);
  and _51501_ (_19025_, _18844_, _18809_);
  and _51502_ (_19026_, _18839_, _18815_);
  or _51503_ (_19027_, _19026_, _19025_);
  or _51504_ (_19028_, _19027_, _18964_);
  and _51505_ (_19029_, _18856_, _18809_);
  and _51506_ (_19030_, _18851_, _18815_);
  nor _51507_ (_19031_, _19030_, _19029_);
  nand _51508_ (_19032_, _19031_, _18964_);
  and _51509_ (_19033_, _19032_, _19028_);
  and _51510_ (_19034_, _19033_, _18967_);
  not _51511_ (_19035_, _18967_);
  and _51512_ (_19036_, _18818_, _18809_);
  and _51513_ (_19037_, _18813_, _18815_);
  nor _51514_ (_19038_, _19037_, _19036_);
  nor _51515_ (_19039_, _19038_, _18964_);
  and _51516_ (_19040_, _18830_, _18809_);
  and _51517_ (_19041_, _18825_, _18815_);
  or _51518_ (_19042_, _19041_, _19040_);
  and _51519_ (_19043_, _19042_, _18964_);
  or _51520_ (_19044_, _19043_, _19039_);
  and _51521_ (_19045_, _19044_, _19035_);
  nor _51522_ (_19046_, _19045_, _19034_);
  nor _51523_ (_19047_, _19046_, _19024_);
  and _51524_ (_19048_, _19024_, word_in[31]);
  or _51525_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _19048_, _19047_);
  or _51526_ (_19049_, _18647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _51527_ (_25618_, _19049_, _27355_);
  and _51528_ (_19050_, _19024_, _27355_);
  and _51529_ (_19051_, _19050_, _18967_);
  and _51530_ (_19052_, _19051_, _18964_);
  and _51531_ (_19053_, _19052_, _18657_);
  not _51532_ (_19054_, _19053_);
  and _51533_ (_19055_, _18904_, _27355_);
  and _51534_ (_19056_, _19055_, _18689_);
  nor _51535_ (_19057_, _18939_, rst);
  nor _51536_ (_19058_, _18874_, _18699_);
  and _51537_ (_19059_, _19058_, _19057_);
  and _51538_ (_19060_, _19059_, _19056_);
  not _51539_ (_19061_, _19060_);
  and _51540_ (_19062_, _18808_, _27355_);
  and _51541_ (_19063_, _19062_, _18758_);
  and _51542_ (_19064_, _19063_, _18775_);
  and _51543_ (_19065_, _19064_, _18679_);
  and _51544_ (_19066_, _18753_, _18639_);
  and _51545_ (_19067_, _18694_, _27355_);
  and _51546_ (_19068_, _19067_, word_in[7]);
  and _51547_ (_19069_, _19068_, _19066_);
  nand _51548_ (_19070_, _19067_, _19066_);
  and _51549_ (_19071_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _51550_ (_19072_, _19071_, _19069_);
  nor _51551_ (_19073_, _19072_, _19065_);
  and _51552_ (_19074_, _19062_, word_in[15]);
  and _51553_ (_19075_, _19074_, _19065_);
  or _51554_ (_19076_, _19075_, _19073_);
  and _51555_ (_19077_, _19076_, _19061_);
  and _51556_ (_19078_, _19060_, word_in[23]);
  or _51557_ (_19079_, _19078_, _19077_);
  and _51558_ (_19080_, _19079_, _19054_);
  and _51559_ (_19081_, _19050_, word_in[31]);
  and _51560_ (_19082_, _19081_, _19053_);
  or _51561_ (_25622_, _19082_, _19080_);
  and _51562_ (_19083_, _18657_, _18642_);
  or _51563_ (_19084_, _18965_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _51564_ (_19085_, _19084_, _19083_);
  and _51565_ (_25625_, _19085_, _27355_);
  or _51566_ (_19086_, _19066_, _18870_);
  and _51567_ (_19087_, _18679_, _18647_);
  or _51568_ (_19088_, _19087_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _51569_ (_19089_, _19088_, _19086_);
  and _51570_ (_25629_, _19089_, _27355_);
  and _51571_ (_19090_, _18679_, _18642_);
  or _51572_ (_19091_, _19090_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _51573_ (_19092_, _19091_, _19086_);
  and _51574_ (_25634_, _19092_, _27355_);
  or _51575_ (_19093_, _18642_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _51576_ (_25640_, _19093_, _27355_);
  and _51577_ (_19094_, _18667_, _18642_);
  and _51578_ (_19095_, _18668_, _18642_);
  and _51579_ (_19096_, _19095_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _51580_ (_19097_, _19096_, _19094_);
  not _51581_ (_19098_, _18642_);
  and _51582_ (_19099_, _18657_, _18640_);
  nand _51583_ (_19100_, _18966_, _18668_);
  and _51584_ (_19101_, _19100_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _51585_ (_19102_, _19101_, _19099_);
  and _51586_ (_19103_, _19102_, _19098_);
  nor _51587_ (_19104_, _19103_, _19097_);
  nor _51588_ (_19105_, _19104_, _18760_);
  or _51589_ (_19106_, _19102_, _19096_);
  and _51590_ (_19107_, _19106_, _19066_);
  and _51591_ (_19108_, _18815_, _18642_);
  and _51592_ (_19109_, _18870_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _51593_ (_19110_, _19109_, _19108_);
  or _51594_ (_19111_, _19110_, _19107_);
  or _51595_ (_19112_, _19111_, _19105_);
  and _51596_ (_25647_, _19112_, _27355_);
  and _51597_ (_19113_, _18690_, _18640_);
  or _51598_ (_19114_, _19113_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _51599_ (_19115_, _18966_, _19066_);
  and _51600_ (_19116_, _19115_, _19114_);
  or _51601_ (_19117_, _19116_, _19099_);
  and _51602_ (_19118_, _18690_, _18642_);
  and _51603_ (_19119_, _19118_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _51604_ (_19120_, _19119_, _19090_);
  and _51605_ (_19121_, _19083_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _51606_ (_19122_, _19114_, _19066_);
  or _51607_ (_19123_, _19122_, _19121_);
  or _51608_ (_19124_, _19123_, _19120_);
  or _51609_ (_19125_, _19124_, _19094_);
  or _51610_ (_19126_, _19125_, _19117_);
  and _51611_ (_25655_, _19126_, _27355_);
  or _51612_ (_19127_, _19094_, _19099_);
  or _51613_ (_19128_, _19127_, _19113_);
  and _51614_ (_19129_, _19095_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _51615_ (_19130_, _18700_, _18639_);
  and _51616_ (_19131_, _18679_, _18640_);
  or _51617_ (_19132_, _18653_, _18639_);
  nor _51618_ (_19133_, _18642_, _18798_);
  and _51619_ (_19134_, _19133_, _19132_);
  or _51620_ (_19135_, _19134_, _19131_);
  and _51621_ (_19136_, _19135_, _19130_);
  or _51622_ (_19137_, _19136_, _19129_);
  or _51623_ (_19138_, _19137_, _19128_);
  and _51624_ (_25663_, _19138_, _27355_);
  or _51625_ (_19139_, _18874_, _18639_);
  not _51626_ (_19140_, _19139_);
  nor _51627_ (_19141_, _19140_, _19086_);
  and _51628_ (_19142_, _18664_, _18689_);
  nand _51629_ (_19143_, _18680_, _18640_);
  and _51630_ (_19144_, _19143_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _51631_ (_19145_, _19144_, _19142_);
  or _51632_ (_19146_, _19145_, _18755_);
  and _51633_ (_19147_, _19146_, _18775_);
  and _51634_ (_19148_, _19094_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _51635_ (_19149_, _19148_, _19131_);
  or _51636_ (_19150_, _19149_, _19142_);
  or _51637_ (_19151_, _19150_, _19147_);
  and _51638_ (_19152_, _19151_, _19141_);
  and _51639_ (_19153_, _19145_, _19066_);
  or _51640_ (_19154_, _19148_, _19099_);
  and _51641_ (_19155_, _18870_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _51642_ (_19156_, _19090_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _51643_ (_19157_, _19156_, _19155_);
  or _51644_ (_19158_, _19157_, _19154_);
  or _51645_ (_19159_, _19158_, _19153_);
  or _51646_ (_19160_, _19159_, _19113_);
  or _51647_ (_19161_, _19160_, _19152_);
  and _51648_ (_25673_, _19161_, _27355_);
  and _51649_ (_19162_, _18815_, _18640_);
  and _51650_ (_19163_, _18963_, _18639_);
  or _51651_ (_19164_, _19163_, _18755_);
  or _51652_ (_19165_, _19164_, _19162_);
  or _51653_ (_19166_, _19165_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _51654_ (_25683_, _19166_, _27355_);
  not _51655_ (_19167_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _51656_ (_19168_, _19130_, _19167_);
  and _51657_ (_19169_, _18690_, _18645_);
  or _51658_ (_19170_, _19169_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _51659_ (_19171_, _19170_, _19130_);
  or _51660_ (_19172_, _19171_, _18963_);
  and _51661_ (_19173_, _19172_, _18639_);
  or _51662_ (_19174_, _19173_, _18755_);
  or _51663_ (_19175_, _19174_, _19131_);
  or _51664_ (_19176_, _19175_, _19168_);
  and _51665_ (_28201_[9], _19176_, _27355_);
  or _51666_ (_19177_, _19058_, _19087_);
  or _51667_ (_19178_, _19177_, _19066_);
  and _51668_ (_19179_, _19083_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _51669_ (_19180_, _18679_, _18645_);
  and _51670_ (_19181_, _19108_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _51671_ (_19182_, _19181_, _19180_);
  or _51672_ (_19183_, _19182_, _19179_);
  or _51673_ (_19184_, _19127_, _19162_);
  and _51674_ (_19185_, _19184_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _51675_ (_19186_, _19164_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _51676_ (_19187_, _18757_);
  and _51677_ (_19188_, _19187_, _18639_);
  or _51678_ (_19189_, _19188_, _19169_);
  and _51679_ (_19190_, _19189_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _51680_ (_19191_, _19190_, _19186_);
  or _51681_ (_19192_, _19191_, _19185_);
  or _51682_ (_19193_, _19192_, _19183_);
  and _51683_ (_19194_, _19193_, _19178_);
  not _51684_ (_19195_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _51685_ (_19196_, _19139_, _19195_);
  and _51686_ (_19197_, _19131_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _51687_ (_19198_, _18870_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _51688_ (_19199_, _19198_, _18755_);
  or _51689_ (_19200_, _19199_, _19197_);
  or _51690_ (_19201_, _19200_, _19196_);
  or _51691_ (_19202_, _19201_, _19169_);
  or _51692_ (_19203_, _19202_, _19163_);
  or _51693_ (_19204_, _19203_, _19194_);
  and _51694_ (_28201_[10], _19204_, _27355_);
  and _51695_ (_19205_, _18667_, _18645_);
  or _51696_ (_19206_, _19205_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51697_ (_19207_, _19187_, _18754_);
  and _51698_ (_19208_, _19207_, _19206_);
  and _51699_ (_19209_, _18663_, _18689_);
  and _51700_ (_19210_, _18755_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _51701_ (_19211_, _19210_, _19180_);
  or _51702_ (_19212_, _19211_, _19209_);
  or _51703_ (_19213_, _19099_, _19113_);
  and _51704_ (_19214_, _19213_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51705_ (_19215_, _19131_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51706_ (_19216_, _19094_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51707_ (_19217_, _19108_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _51708_ (_19218_, _19217_, _19216_);
  or _51709_ (_19219_, _19218_, _19215_);
  or _51710_ (_19220_, _19219_, _19214_);
  or _51711_ (_19221_, _19220_, _19212_);
  or _51712_ (_19222_, _19221_, _19208_);
  and _51713_ (_19223_, _19222_, _19177_);
  and _51714_ (_19224_, _19066_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _51715_ (_19225_, _19083_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _51716_ (_19226_, _19225_, _19163_);
  or _51717_ (_19227_, _19226_, _19210_);
  or _51718_ (_19228_, _19227_, _19220_);
  or _51719_ (_19229_, _19228_, _19169_);
  or _51720_ (_19230_, _19229_, _19224_);
  or _51721_ (_19231_, _19230_, _19223_);
  and _51722_ (_28201_[11], _19231_, _27355_);
  and _51723_ (_19232_, _18965_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _51724_ (_19233_, _18690_, _18647_);
  not _51725_ (_19234_, _19233_);
  and _51726_ (_19235_, _19058_, _19234_);
  and _51727_ (_19236_, _19108_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _51728_ (_19237_, _19162_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _51729_ (_19238_, _19237_, _19236_);
  or _51730_ (_19239_, _19238_, _19235_);
  and _51731_ (_19240_, _19099_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _51732_ (_19241_, _18963_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _51733_ (_19242_, _19241_, _19169_);
  or _51734_ (_19243_, _19242_, _19240_);
  and _51735_ (_19244_, _19094_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _51736_ (_19245_, _18755_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _51737_ (_19246_, _19245_, _19244_);
  or _51738_ (_19247_, _19246_, _19243_);
  or _51739_ (_19248_, _19247_, _19239_);
  or _51740_ (_19249_, _19248_, _19232_);
  and _51741_ (_28201_[12], _19249_, _27355_);
  or _51742_ (_19250_, _19058_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _51743_ (_28201_[13], _19250_, _27355_);
  or _51744_ (_19251_, _19207_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _51745_ (_28201_[14], _19251_, _27355_);
  and _51746_ (_19252_, _19050_, word_in[24]);
  and _51747_ (_19253_, _19050_, _18964_);
  nor _51748_ (_19254_, _19051_, _19253_);
  and _51749_ (_19255_, _19254_, _18690_);
  and _51750_ (_19256_, _19255_, _19252_);
  and _51751_ (_19257_, _19057_, _18689_);
  nor _51752_ (_19258_, _19257_, _19055_);
  and _51753_ (_19259_, _19258_, _19057_);
  and _51754_ (_19260_, _19259_, _18872_);
  not _51755_ (_19261_, _19260_);
  or _51756_ (_19262_, _19261_, word_in[16]);
  and _51757_ (_19263_, _19255_, _19050_);
  not _51758_ (_19264_, _19263_);
  and _51759_ (_19265_, _19062_, _19066_);
  and _51760_ (_19266_, _19067_, word_in[0]);
  and _51761_ (_19267_, _19266_, _19083_);
  not _51762_ (_19268_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _51763_ (_19269_, _19067_, _19083_);
  nor _51764_ (_19270_, _19269_, _19268_);
  or _51765_ (_19271_, _19270_, _19267_);
  or _51766_ (_19272_, _19271_, _19265_);
  not _51767_ (_19273_, _19265_);
  or _51768_ (_19274_, _19273_, word_in[8]);
  and _51769_ (_19275_, _19274_, _19272_);
  or _51770_ (_19276_, _19275_, _19260_);
  and _51771_ (_19277_, _19276_, _19264_);
  and _51772_ (_19278_, _19277_, _19262_);
  or _51773_ (_28202_[0], _19278_, _19256_);
  and _51774_ (_19279_, _19050_, word_in[25]);
  and _51775_ (_19280_, _19279_, _19255_);
  or _51776_ (_19281_, _19261_, word_in[17]);
  and _51777_ (_19282_, _19062_, word_in[9]);
  and _51778_ (_19283_, _19282_, _19066_);
  not _51779_ (_19284_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or _51780_ (_19285_, _19269_, _19284_);
  and _51781_ (_19286_, _19067_, word_in[1]);
  nand _51782_ (_19287_, _19286_, _19269_);
  and _51783_ (_19288_, _19287_, _19285_);
  nor _51784_ (_19289_, _19288_, _19265_);
  or _51785_ (_19290_, _19289_, _19283_);
  or _51786_ (_19291_, _19290_, _19260_);
  and _51787_ (_19292_, _19291_, _19264_);
  and _51788_ (_19293_, _19292_, _19281_);
  or _51789_ (_28202_[1], _19293_, _19280_);
  and _51790_ (_19294_, _19050_, word_in[26]);
  and _51791_ (_19295_, _19294_, _19255_);
  or _51792_ (_19296_, _19261_, word_in[18]);
  not _51793_ (_19297_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _51794_ (_19298_, _19269_, _19297_);
  and _51795_ (_19299_, _19067_, word_in[2]);
  and _51796_ (_19300_, _19299_, _19269_);
  or _51797_ (_19301_, _19300_, _19298_);
  or _51798_ (_19302_, _19301_, _19265_);
  or _51799_ (_19303_, _19273_, word_in[10]);
  and _51800_ (_19304_, _19303_, _19302_);
  or _51801_ (_19305_, _19304_, _19260_);
  and _51802_ (_19306_, _19305_, _19264_);
  and _51803_ (_19307_, _19306_, _19296_);
  or _51804_ (_28202_[2], _19307_, _19295_);
  and _51805_ (_19308_, _19050_, word_in[27]);
  and _51806_ (_19309_, _19308_, _19255_);
  or _51807_ (_19310_, _19261_, word_in[19]);
  not _51808_ (_19311_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _51809_ (_19312_, _19269_, _19311_);
  and _51810_ (_19313_, _19067_, word_in[3]);
  and _51811_ (_19314_, _19313_, _19269_);
  or _51812_ (_19315_, _19314_, _19312_);
  or _51813_ (_19316_, _19315_, _19265_);
  or _51814_ (_19317_, _19273_, word_in[11]);
  and _51815_ (_19318_, _19317_, _19316_);
  or _51816_ (_19319_, _19318_, _19260_);
  and _51817_ (_19320_, _19319_, _19264_);
  and _51818_ (_19321_, _19320_, _19310_);
  or _51819_ (_28202_[3], _19321_, _19309_);
  and _51820_ (_19322_, _19050_, word_in[28]);
  and _51821_ (_19323_, _19322_, _19255_);
  or _51822_ (_19324_, _19261_, word_in[20]);
  not _51823_ (_19325_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _51824_ (_19326_, _19269_, _19325_);
  and _51825_ (_19327_, _19067_, word_in[4]);
  and _51826_ (_19328_, _19327_, _19083_);
  or _51827_ (_19329_, _19328_, _19326_);
  or _51828_ (_19330_, _19329_, _19265_);
  or _51829_ (_19331_, _19273_, word_in[12]);
  and _51830_ (_19332_, _19331_, _19330_);
  or _51831_ (_19333_, _19332_, _19260_);
  and _51832_ (_19334_, _19333_, _19264_);
  and _51833_ (_19335_, _19334_, _19324_);
  or _51834_ (_28202_[4], _19335_, _19323_);
  or _51835_ (_19336_, _19261_, word_in[21]);
  not _51836_ (_19337_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _51837_ (_19338_, _19269_, _19337_);
  and _51838_ (_19339_, _19067_, word_in[5]);
  and _51839_ (_19340_, _19339_, _19269_);
  or _51840_ (_19341_, _19340_, _19338_);
  or _51841_ (_19342_, _19341_, _19265_);
  or _51842_ (_19343_, _19273_, word_in[13]);
  and _51843_ (_19344_, _19343_, _19342_);
  or _51844_ (_19345_, _19344_, _19260_);
  and _51845_ (_19346_, _19345_, _19264_);
  and _51846_ (_19347_, _19346_, _19336_);
  and _51847_ (_19348_, _19050_, word_in[29]);
  and _51848_ (_19349_, _19348_, _19263_);
  or _51849_ (_28202_[5], _19349_, _19347_);
  and _51850_ (_19350_, _19050_, word_in[30]);
  and _51851_ (_19351_, _19350_, _19255_);
  or _51852_ (_19352_, _19261_, word_in[22]);
  not _51853_ (_19353_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _51854_ (_19354_, _19269_, _19353_);
  and _51855_ (_19355_, _19067_, word_in[6]);
  and _51856_ (_19356_, _19355_, _19269_);
  or _51857_ (_19357_, _19356_, _19354_);
  or _51858_ (_19358_, _19357_, _19265_);
  or _51859_ (_19359_, _19273_, word_in[14]);
  and _51860_ (_19360_, _19359_, _19358_);
  or _51861_ (_19361_, _19360_, _19260_);
  and _51862_ (_19362_, _19361_, _19264_);
  and _51863_ (_19363_, _19362_, _19352_);
  or _51864_ (_28202_[6], _19363_, _19351_);
  and _51865_ (_19364_, _19255_, _19081_);
  or _51866_ (_19365_, _19261_, word_in[23]);
  nor _51867_ (_19366_, _19269_, _18810_);
  and _51868_ (_19367_, _19269_, _19068_);
  or _51869_ (_19368_, _19367_, _19366_);
  or _51870_ (_19369_, _19368_, _19265_);
  or _51871_ (_19370_, _19273_, word_in[15]);
  and _51872_ (_19371_, _19370_, _19369_);
  or _51873_ (_19372_, _19371_, _19260_);
  and _51874_ (_19373_, _19372_, _19264_);
  and _51875_ (_19374_, _19373_, _19365_);
  or _51876_ (_28202_[7], _19374_, _19364_);
  and _51877_ (_19375_, _19050_, _18679_);
  and _51878_ (_19376_, _19375_, _19254_);
  and _51879_ (_19377_, _19376_, _19252_);
  and _51880_ (_19378_, _19057_, _18871_);
  and _51881_ (_19379_, _19055_, _18656_);
  not _51882_ (_19380_, _19379_);
  nor _51883_ (_19381_, _19380_, _19378_);
  and _51884_ (_19382_, _19062_, _19083_);
  and _51885_ (_19383_, _19266_, _19118_);
  nand _51886_ (_19384_, _19067_, _19118_);
  and _51887_ (_19385_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or _51888_ (_19386_, _19385_, _19383_);
  or _51889_ (_19387_, _19386_, _19382_);
  not _51890_ (_19388_, _19382_);
  or _51891_ (_19389_, _19388_, word_in[8]);
  and _51892_ (_19390_, _19389_, _19387_);
  or _51893_ (_19391_, _19390_, _19381_);
  not _51894_ (_19392_, _19376_);
  and _51895_ (_19393_, _19057_, word_in[16]);
  not _51896_ (_19394_, _19381_);
  or _51897_ (_19395_, _19394_, _19393_);
  and _51898_ (_19396_, _19395_, _19392_);
  and _51899_ (_19397_, _19396_, _19391_);
  or _51900_ (_28209_[0], _19397_, _19377_);
  and _51901_ (_19398_, _19286_, _19118_);
  and _51902_ (_19399_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _51903_ (_19400_, _19399_, _19398_);
  nor _51904_ (_19401_, _19400_, _19382_);
  and _51905_ (_19402_, _19382_, word_in[9]);
  nor _51906_ (_19403_, _19402_, _19401_);
  nor _51907_ (_19404_, _19403_, _19381_);
  and _51908_ (_19405_, _19057_, word_in[17]);
  and _51909_ (_19406_, _19381_, _19405_);
  or _51910_ (_19407_, _19406_, _19376_);
  or _51911_ (_19408_, _19407_, _19404_);
  or _51912_ (_19409_, _19392_, _19279_);
  and _51913_ (_28209_[1], _19409_, _19408_);
  and _51914_ (_19410_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _51915_ (_19411_, _19299_, _19118_);
  nor _51916_ (_19412_, _19411_, _19410_);
  nor _51917_ (_19413_, _19412_, _19382_);
  and _51918_ (_19414_, _19382_, word_in[10]);
  nor _51919_ (_19415_, _19414_, _19413_);
  nor _51920_ (_19416_, _19415_, _19381_);
  and _51921_ (_19417_, _19057_, word_in[18]);
  and _51922_ (_19418_, _19381_, _19417_);
  or _51923_ (_19419_, _19418_, _19376_);
  or _51924_ (_19420_, _19419_, _19416_);
  or _51925_ (_19421_, _19392_, _19294_);
  and _51926_ (_28209_[2], _19421_, _19420_);
  and _51927_ (_19422_, _19313_, _19118_);
  and _51928_ (_19423_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _51929_ (_19424_, _19423_, _19422_);
  nor _51930_ (_19425_, _19424_, _19382_);
  and _51931_ (_19426_, _19382_, word_in[11]);
  nor _51932_ (_19427_, _19426_, _19425_);
  nor _51933_ (_19428_, _19427_, _19381_);
  and _51934_ (_19429_, _19057_, word_in[19]);
  and _51935_ (_19430_, _19381_, _19429_);
  or _51936_ (_19431_, _19430_, _19376_);
  or _51937_ (_19432_, _19431_, _19428_);
  or _51938_ (_19433_, _19392_, _19308_);
  and _51939_ (_28209_[3], _19433_, _19432_);
  and _51940_ (_19434_, _19327_, _19118_);
  and _51941_ (_19435_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or _51942_ (_19436_, _19435_, _19434_);
  or _51943_ (_19437_, _19436_, _19382_);
  or _51944_ (_19438_, _19388_, word_in[12]);
  nand _51945_ (_19439_, _19438_, _19437_);
  nor _51946_ (_19440_, _19439_, _19381_);
  and _51947_ (_19441_, _19057_, word_in[20]);
  and _51948_ (_19442_, _19381_, _19441_);
  or _51949_ (_19443_, _19442_, _19376_);
  or _51950_ (_19444_, _19443_, _19440_);
  or _51951_ (_19445_, _19392_, word_in[28]);
  and _51952_ (_28209_[4], _19445_, _19444_);
  and _51953_ (_19446_, _19339_, _19118_);
  and _51954_ (_19447_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or _51955_ (_19448_, _19447_, _19446_);
  or _51956_ (_19449_, _19448_, _19382_);
  or _51957_ (_19450_, _19388_, word_in[13]);
  nand _51958_ (_19451_, _19450_, _19449_);
  nor _51959_ (_19452_, _19451_, _19381_);
  and _51960_ (_19453_, _19057_, word_in[21]);
  and _51961_ (_19454_, _19381_, _19453_);
  or _51962_ (_19455_, _19454_, _19376_);
  or _51963_ (_19456_, _19455_, _19452_);
  or _51964_ (_19457_, _19392_, word_in[29]);
  and _51965_ (_28209_[5], _19457_, _19456_);
  and _51966_ (_19458_, _19355_, _19118_);
  and _51967_ (_19459_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _51968_ (_19460_, _19459_, _19458_);
  nor _51969_ (_19461_, _19460_, _19382_);
  and _51970_ (_19462_, _19382_, word_in[14]);
  nor _51971_ (_19463_, _19462_, _19461_);
  nor _51972_ (_19464_, _19463_, _19381_);
  and _51973_ (_19465_, _19057_, word_in[22]);
  and _51974_ (_19466_, _19381_, _19465_);
  or _51975_ (_19467_, _19466_, _19376_);
  or _51976_ (_19468_, _19467_, _19464_);
  or _51977_ (_19469_, _19392_, _19350_);
  and _51978_ (_28209_[6], _19469_, _19468_);
  and _51979_ (_19470_, _19068_, _19118_);
  and _51980_ (_19471_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _51981_ (_19472_, _19471_, _19470_);
  nor _51982_ (_19473_, _19472_, _19382_);
  and _51983_ (_19474_, _19382_, word_in[15]);
  nor _51984_ (_19475_, _19474_, _19473_);
  nor _51985_ (_19476_, _19475_, _19381_);
  and _51986_ (_19477_, _19057_, word_in[23]);
  and _51987_ (_19478_, _19381_, _19477_);
  or _51988_ (_19479_, _19478_, _19376_);
  or _51989_ (_19480_, _19479_, _19476_);
  or _51990_ (_19481_, _19392_, _19081_);
  and _51991_ (_28209_[7], _19481_, _19480_);
  and _51992_ (_19482_, _19050_, _18667_);
  and _51993_ (_19483_, _19482_, _19254_);
  not _51994_ (_19484_, _19483_);
  not _51995_ (_19485_, _19055_);
  and _51996_ (_19486_, _19257_, _19485_);
  and _51997_ (_19487_, _19486_, _18872_);
  and _51998_ (_19488_, _19062_, _19118_);
  nand _51999_ (_19489_, _19067_, _19090_);
  and _52000_ (_19490_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _52001_ (_19491_, _19266_, _19090_);
  nor _52002_ (_19492_, _19491_, _19490_);
  nor _52003_ (_19493_, _19492_, _19488_);
  and _52004_ (_19494_, _19488_, word_in[8]);
  nor _52005_ (_19495_, _19494_, _19493_);
  nor _52006_ (_19496_, _19495_, _19487_);
  and _52007_ (_19497_, _19487_, _19393_);
  or _52008_ (_19499_, _19497_, _19496_);
  and _52009_ (_19500_, _19499_, _19484_);
  and _52010_ (_19501_, _19483_, word_in[24]);
  or _52011_ (_28210_[0], _19501_, _19500_);
  and _52012_ (_19502_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _52013_ (_19503_, _19286_, _19090_);
  or _52014_ (_19504_, _19503_, _19502_);
  or _52015_ (_19505_, _19504_, _19488_);
  not _52016_ (_19506_, _19488_);
  or _52017_ (_19507_, _19506_, word_in[9]);
  nand _52018_ (_19509_, _19507_, _19505_);
  nor _52019_ (_19510_, _19509_, _19487_);
  and _52020_ (_19511_, _19487_, _19405_);
  or _52021_ (_19512_, _19511_, _19483_);
  or _52022_ (_19513_, _19512_, _19510_);
  or _52023_ (_19514_, _19484_, word_in[25]);
  and _52024_ (_28210_[1], _19514_, _19513_);
  and _52025_ (_19515_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _52026_ (_19516_, _19299_, _19090_);
  nor _52027_ (_19517_, _19516_, _19515_);
  nor _52028_ (_19519_, _19517_, _19488_);
  and _52029_ (_19520_, _19488_, word_in[10]);
  nor _52030_ (_19521_, _19520_, _19519_);
  nor _52031_ (_19522_, _19521_, _19487_);
  and _52032_ (_19523_, _19487_, _19417_);
  or _52033_ (_19524_, _19523_, _19522_);
  and _52034_ (_19525_, _19524_, _19484_);
  and _52035_ (_19526_, _19483_, word_in[26]);
  or _52036_ (_28210_[2], _19526_, _19525_);
  and _52037_ (_19527_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _52038_ (_19529_, _19313_, _19090_);
  nor _52039_ (_19530_, _19529_, _19527_);
  nor _52040_ (_19531_, _19530_, _19488_);
  and _52041_ (_19532_, _19488_, word_in[11]);
  nor _52042_ (_19533_, _19532_, _19531_);
  nor _52043_ (_19534_, _19533_, _19487_);
  and _52044_ (_19535_, _19487_, _19429_);
  or _52045_ (_19536_, _19535_, _19534_);
  and _52046_ (_19537_, _19536_, _19484_);
  and _52047_ (_19538_, _19483_, word_in[27]);
  or _52048_ (_28210_[3], _19538_, _19537_);
  and _52049_ (_19540_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _52050_ (_19541_, _19327_, _19090_);
  nor _52051_ (_19542_, _19541_, _19540_);
  nor _52052_ (_19543_, _19542_, _19488_);
  and _52053_ (_19544_, _19488_, word_in[12]);
  nor _52054_ (_19545_, _19544_, _19543_);
  nor _52055_ (_19546_, _19545_, _19487_);
  and _52056_ (_19547_, _19487_, _19441_);
  or _52057_ (_19548_, _19547_, _19546_);
  and _52058_ (_19550_, _19548_, _19484_);
  and _52059_ (_19551_, _19483_, word_in[28]);
  or _52060_ (_28210_[4], _19551_, _19550_);
  and _52061_ (_19552_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _52062_ (_19553_, _19339_, _19090_);
  or _52063_ (_19554_, _19553_, _19552_);
  or _52064_ (_19555_, _19554_, _19488_);
  or _52065_ (_19556_, _19506_, word_in[13]);
  nand _52066_ (_19557_, _19556_, _19555_);
  nor _52067_ (_19558_, _19557_, _19487_);
  and _52068_ (_19560_, _19487_, _19453_);
  or _52069_ (_19561_, _19560_, _19483_);
  or _52070_ (_19562_, _19561_, _19558_);
  or _52071_ (_19563_, _19484_, word_in[29]);
  and _52072_ (_28210_[5], _19563_, _19562_);
  and _52073_ (_19564_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _52074_ (_19565_, _19355_, _19090_);
  nor _52075_ (_19566_, _19565_, _19564_);
  nor _52076_ (_19567_, _19566_, _19488_);
  and _52077_ (_19568_, _19488_, word_in[14]);
  nor _52078_ (_19569_, _19568_, _19567_);
  nor _52079_ (_19570_, _19569_, _19487_);
  and _52080_ (_19571_, _19487_, _19465_);
  or _52081_ (_19572_, _19571_, _19570_);
  and _52082_ (_19573_, _19572_, _19484_);
  and _52083_ (_19574_, _19483_, word_in[30]);
  or _52084_ (_28210_[6], _19574_, _19573_);
  and _52085_ (_19575_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _52086_ (_19576_, _19068_, _19090_);
  nor _52087_ (_19577_, _19576_, _19575_);
  nor _52088_ (_19578_, _19577_, _19488_);
  and _52089_ (_19579_, _19488_, word_in[15]);
  nor _52090_ (_19580_, _19579_, _19578_);
  nor _52091_ (_19581_, _19580_, _19487_);
  and _52092_ (_19582_, _19487_, _19477_);
  or _52093_ (_19583_, _19582_, _19581_);
  and _52094_ (_19584_, _19583_, _19484_);
  and _52095_ (_19585_, _19483_, word_in[31]);
  or _52096_ (_28210_[7], _19585_, _19584_);
  not _52097_ (_19586_, _19056_);
  nor _52098_ (_19587_, _19378_, _19586_);
  and _52099_ (_19588_, _19062_, _19090_);
  nand _52100_ (_19589_, _19067_, _19094_);
  and _52101_ (_19590_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _52102_ (_19591_, _19266_, _19094_);
  or _52103_ (_19592_, _19591_, _19590_);
  or _52104_ (_19593_, _19592_, _19588_);
  not _52105_ (_19594_, _19588_);
  or _52106_ (_19595_, _19594_, word_in[8]);
  and _52107_ (_19596_, _19595_, _19593_);
  or _52108_ (_19597_, _19596_, _19587_);
  and _52109_ (_19598_, _19050_, _19083_);
  not _52110_ (_19599_, _19598_);
  not _52111_ (_19600_, _19587_);
  or _52112_ (_19601_, _19600_, _19393_);
  and _52113_ (_19602_, _19601_, _19599_);
  and _52114_ (_19603_, _19602_, _19597_);
  and _52115_ (_19604_, _19598_, word_in[24]);
  or _52116_ (_28211_[0], _19604_, _19603_);
  and _52117_ (_19605_, _19587_, _19405_);
  and _52118_ (_19606_, _19286_, _19094_);
  and _52119_ (_19607_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _52120_ (_19608_, _19607_, _19606_);
  nor _52121_ (_19609_, _19608_, _19588_);
  and _52122_ (_19610_, _19588_, word_in[9]);
  nor _52123_ (_19611_, _19610_, _19609_);
  nor _52124_ (_19612_, _19611_, _19587_);
  or _52125_ (_19613_, _19612_, _19605_);
  and _52126_ (_19614_, _19613_, _19599_);
  and _52127_ (_19615_, _19598_, word_in[25]);
  or _52128_ (_28211_[1], _19615_, _19614_);
  and _52129_ (_19616_, _19587_, _19417_);
  and _52130_ (_19617_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _52131_ (_19618_, _19299_, _19094_);
  nor _52132_ (_19619_, _19618_, _19617_);
  nor _52133_ (_19620_, _19619_, _19588_);
  and _52134_ (_19621_, _19588_, word_in[10]);
  nor _52135_ (_19622_, _19621_, _19620_);
  nor _52136_ (_19623_, _19622_, _19587_);
  or _52137_ (_19624_, _19623_, _19616_);
  and _52138_ (_19625_, _19624_, _19599_);
  and _52139_ (_19626_, _19598_, word_in[26]);
  or _52140_ (_28211_[2], _19626_, _19625_);
  and _52141_ (_19627_, _19598_, _19308_);
  and _52142_ (_19628_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _52143_ (_19629_, _19313_, _19094_);
  or _52144_ (_19630_, _19629_, _19628_);
  or _52145_ (_19631_, _19630_, _19588_);
  or _52146_ (_19632_, _19594_, word_in[11]);
  and _52147_ (_19633_, _19632_, _19631_);
  or _52148_ (_19634_, _19633_, _19587_);
  or _52149_ (_19635_, _19600_, _19429_);
  and _52150_ (_19636_, _19635_, _19599_);
  and _52151_ (_19637_, _19636_, _19634_);
  or _52152_ (_28211_[3], _19637_, _19627_);
  and _52153_ (_19638_, _19587_, _19441_);
  and _52154_ (_19639_, _19327_, _19094_);
  and _52155_ (_19640_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _52156_ (_19641_, _19640_, _19639_);
  nor _52157_ (_19642_, _19641_, _19588_);
  and _52158_ (_19643_, _19588_, word_in[12]);
  nor _52159_ (_19644_, _19643_, _19642_);
  nor _52160_ (_19645_, _19644_, _19587_);
  or _52161_ (_19646_, _19645_, _19638_);
  and _52162_ (_19647_, _19646_, _19599_);
  and _52163_ (_19648_, _19598_, word_in[28]);
  or _52164_ (_28211_[4], _19648_, _19647_);
  and _52165_ (_19649_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _52166_ (_19650_, _19339_, _19094_);
  or _52167_ (_19651_, _19650_, _19649_);
  or _52168_ (_19652_, _19651_, _19588_);
  or _52169_ (_19653_, _19594_, word_in[13]);
  and _52170_ (_19654_, _19653_, _19652_);
  or _52171_ (_19655_, _19654_, _19587_);
  or _52172_ (_19656_, _19600_, _19453_);
  and _52173_ (_19657_, _19656_, _19599_);
  and _52174_ (_19658_, _19657_, _19655_);
  and _52175_ (_19659_, _19598_, word_in[29]);
  or _52176_ (_28211_[5], _19659_, _19658_);
  and _52177_ (_19660_, _19587_, _19465_);
  and _52178_ (_19661_, _19355_, _19094_);
  and _52179_ (_19662_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _52180_ (_19663_, _19662_, _19661_);
  nor _52181_ (_19664_, _19663_, _19588_);
  and _52182_ (_19665_, _19588_, word_in[14]);
  nor _52183_ (_19666_, _19665_, _19664_);
  nor _52184_ (_19667_, _19666_, _19587_);
  or _52185_ (_19668_, _19667_, _19660_);
  and _52186_ (_19669_, _19668_, _19599_);
  and _52187_ (_19670_, _19598_, word_in[30]);
  or _52188_ (_28211_[6], _19670_, _19669_);
  and _52189_ (_19671_, _19587_, _19477_);
  and _52190_ (_19672_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _52191_ (_19673_, _19068_, _19094_);
  nor _52192_ (_19674_, _19673_, _19672_);
  nor _52193_ (_19675_, _19674_, _19588_);
  and _52194_ (_19676_, _19588_, word_in[15]);
  nor _52195_ (_19677_, _19676_, _19675_);
  nor _52196_ (_19678_, _19677_, _19587_);
  or _52197_ (_19679_, _19678_, _19671_);
  and _52198_ (_19680_, _19679_, _19599_);
  and _52199_ (_19681_, _19598_, word_in[31]);
  or _52200_ (_28211_[7], _19681_, _19680_);
  and _52201_ (_19682_, _19253_, _18699_);
  and _52202_ (_19683_, _19682_, _18690_);
  not _52203_ (_19684_, _19683_);
  and _52204_ (_19685_, _19140_, _19057_);
  and _52205_ (_19686_, _19685_, _19258_);
  and _52206_ (_19687_, _19062_, _19094_);
  not _52207_ (_19688_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _52208_ (_19689_, _19067_, _19099_);
  nor _52209_ (_19690_, _19689_, _19688_);
  and _52210_ (_19691_, _19266_, _19099_);
  nor _52211_ (_19692_, _19691_, _19690_);
  nor _52212_ (_19693_, _19692_, _19687_);
  and _52213_ (_19694_, _19687_, word_in[8]);
  nor _52214_ (_19695_, _19694_, _19693_);
  nor _52215_ (_19696_, _19695_, _19686_);
  and _52216_ (_19697_, _19686_, _19393_);
  or _52217_ (_19698_, _19697_, _19696_);
  and _52218_ (_19699_, _19698_, _19684_);
  and _52219_ (_19700_, _19683_, _19252_);
  or _52220_ (_28212_[0], _19700_, _19699_);
  not _52221_ (_19701_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _52222_ (_19702_, _19689_, _19701_);
  and _52223_ (_19703_, _19286_, _19099_);
  or _52224_ (_19704_, _19703_, _19702_);
  or _52225_ (_19705_, _19704_, _19687_);
  not _52226_ (_19706_, _19687_);
  or _52227_ (_19707_, _19706_, word_in[9]);
  and _52228_ (_19708_, _19707_, _19705_);
  or _52229_ (_19709_, _19708_, _19686_);
  not _52230_ (_19710_, _19686_);
  or _52231_ (_19711_, _19710_, _19405_);
  and _52232_ (_19712_, _19711_, _19709_);
  or _52233_ (_19713_, _19712_, _19683_);
  or _52234_ (_19714_, _19684_, _19279_);
  and _52235_ (_28212_[1], _19714_, _19713_);
  not _52236_ (_19715_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _52237_ (_19716_, _19689_, _19715_);
  and _52238_ (_19717_, _19299_, _19099_);
  nor _52239_ (_19718_, _19717_, _19716_);
  nor _52240_ (_19719_, _19718_, _19687_);
  and _52241_ (_19720_, _19687_, word_in[10]);
  nor _52242_ (_19721_, _19720_, _19719_);
  nor _52243_ (_19722_, _19721_, _19686_);
  and _52244_ (_19723_, _19686_, _19417_);
  or _52245_ (_19724_, _19723_, _19722_);
  and _52246_ (_19725_, _19724_, _19684_);
  and _52247_ (_19726_, _19683_, _19294_);
  or _52248_ (_28212_[2], _19726_, _19725_);
  not _52249_ (_19727_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _52250_ (_19728_, _19689_, _19727_);
  and _52251_ (_19729_, _19313_, _19099_);
  nor _52252_ (_19730_, _19729_, _19728_);
  nor _52253_ (_19731_, _19730_, _19687_);
  and _52254_ (_19732_, _19687_, word_in[11]);
  nor _52255_ (_19733_, _19732_, _19731_);
  nor _52256_ (_19734_, _19733_, _19686_);
  and _52257_ (_19735_, _19686_, _19429_);
  or _52258_ (_19736_, _19735_, _19734_);
  and _52259_ (_19737_, _19736_, _19684_);
  and _52260_ (_19738_, _19683_, _19308_);
  or _52261_ (_28212_[3], _19738_, _19737_);
  not _52262_ (_19739_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _52263_ (_19740_, _19689_, _19739_);
  and _52264_ (_19741_, _19327_, _19099_);
  nor _52265_ (_19742_, _19741_, _19740_);
  nor _52266_ (_19743_, _19742_, _19687_);
  and _52267_ (_19744_, _19687_, word_in[12]);
  nor _52268_ (_19745_, _19744_, _19743_);
  nor _52269_ (_19746_, _19745_, _19686_);
  and _52270_ (_19747_, _19686_, _19441_);
  or _52271_ (_19748_, _19747_, _19746_);
  and _52272_ (_19749_, _19748_, _19684_);
  and _52273_ (_19750_, _19683_, _19322_);
  or _52274_ (_28212_[4], _19750_, _19749_);
  not _52275_ (_19751_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _52276_ (_19752_, _19689_, _19751_);
  and _52277_ (_19753_, _19339_, _19099_);
  or _52278_ (_19754_, _19753_, _19752_);
  or _52279_ (_19755_, _19754_, _19687_);
  or _52280_ (_19756_, _19706_, word_in[13]);
  and _52281_ (_19757_, _19756_, _19755_);
  or _52282_ (_19758_, _19757_, _19686_);
  or _52283_ (_19759_, _19710_, _19453_);
  and _52284_ (_19760_, _19759_, _19758_);
  or _52285_ (_19761_, _19760_, _19683_);
  or _52286_ (_19762_, _19684_, _19348_);
  and _52287_ (_28212_[5], _19762_, _19761_);
  not _52288_ (_19763_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _52289_ (_19764_, _19689_, _19763_);
  and _52290_ (_19765_, _19355_, _19099_);
  or _52291_ (_19766_, _19765_, _19764_);
  or _52292_ (_19767_, _19766_, _19687_);
  or _52293_ (_19768_, _19706_, word_in[14]);
  and _52294_ (_19769_, _19768_, _19767_);
  or _52295_ (_19770_, _19769_, _19686_);
  or _52296_ (_19771_, _19710_, _19465_);
  and _52297_ (_19772_, _19771_, _19770_);
  or _52298_ (_19773_, _19772_, _19683_);
  or _52299_ (_19774_, _19684_, _19350_);
  and _52300_ (_28212_[6], _19774_, _19773_);
  nor _52301_ (_19775_, _19689_, _18822_);
  and _52302_ (_19776_, _19689_, _19068_);
  or _52303_ (_19777_, _19776_, _19775_);
  or _52304_ (_19778_, _19777_, _19687_);
  or _52305_ (_19779_, _19706_, word_in[15]);
  and _52306_ (_19780_, _19779_, _19778_);
  or _52307_ (_19781_, _19780_, _19686_);
  or _52308_ (_19782_, _19710_, _19477_);
  and _52309_ (_19783_, _19782_, _19781_);
  or _52310_ (_19784_, _19783_, _19683_);
  or _52311_ (_19785_, _19684_, _19081_);
  and _52312_ (_28212_[7], _19785_, _19784_);
  and _52313_ (_19786_, _19685_, _19379_);
  not _52314_ (_19787_, _19786_);
  and _52315_ (_19788_, _19063_, _18756_);
  and _52316_ (_19789_, _19788_, _18657_);
  not _52317_ (_19790_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _52318_ (_19791_, _19067_, _19113_);
  nor _52319_ (_19792_, _19791_, _19790_);
  and _52320_ (_19793_, _19266_, _19113_);
  nor _52321_ (_19794_, _19793_, _19792_);
  nor _52322_ (_19795_, _19794_, _19789_);
  and _52323_ (_19796_, _19062_, word_in[8]);
  and _52324_ (_19797_, _19789_, _19796_);
  or _52325_ (_19798_, _19797_, _19795_);
  and _52326_ (_19799_, _19798_, _19787_);
  and _52327_ (_19800_, _19682_, _18679_);
  and _52328_ (_19801_, _19786_, _19393_);
  or _52329_ (_19802_, _19801_, _19800_);
  or _52330_ (_19803_, _19802_, _19799_);
  not _52331_ (_19804_, _19800_);
  or _52332_ (_19805_, _19804_, _19252_);
  and _52333_ (_28213_[0], _19805_, _19803_);
  not _52334_ (_19806_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _52335_ (_19807_, _19791_, _19806_);
  and _52336_ (_19808_, _19286_, _19113_);
  nor _52337_ (_19809_, _19808_, _19807_);
  nor _52338_ (_19810_, _19809_, _19789_);
  and _52339_ (_19811_, _19789_, _19282_);
  or _52340_ (_19812_, _19811_, _19810_);
  or _52341_ (_19813_, _19812_, _19786_);
  or _52342_ (_19814_, _19787_, _19405_);
  and _52343_ (_19815_, _19814_, _19804_);
  and _52344_ (_19816_, _19815_, _19813_);
  and _52345_ (_19817_, _19800_, _19279_);
  or _52346_ (_28213_[1], _19817_, _19816_);
  not _52347_ (_19818_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _52348_ (_19819_, _19791_, _19818_);
  and _52349_ (_19820_, _19299_, _19113_);
  nor _52350_ (_19821_, _19820_, _19819_);
  nor _52351_ (_19822_, _19821_, _19789_);
  and _52352_ (_19823_, _19062_, word_in[10]);
  and _52353_ (_19824_, _19789_, _19823_);
  or _52354_ (_19825_, _19824_, _19822_);
  and _52355_ (_19826_, _19825_, _19787_);
  and _52356_ (_19827_, _19786_, _19417_);
  or _52357_ (_19828_, _19827_, _19800_);
  or _52358_ (_19829_, _19828_, _19826_);
  or _52359_ (_19830_, _19804_, _19294_);
  and _52360_ (_28213_[2], _19830_, _19829_);
  not _52361_ (_19831_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _52362_ (_19832_, _19791_, _19831_);
  and _52363_ (_19833_, _19313_, _19113_);
  nor _52364_ (_19834_, _19833_, _19832_);
  nor _52365_ (_19835_, _19834_, _19789_);
  and _52366_ (_19836_, _19062_, word_in[11]);
  and _52367_ (_19837_, _19789_, _19836_);
  or _52368_ (_19838_, _19837_, _19835_);
  and _52369_ (_19839_, _19838_, _19787_);
  and _52370_ (_19840_, _19786_, _19429_);
  or _52371_ (_19841_, _19840_, _19800_);
  or _52372_ (_19842_, _19841_, _19839_);
  or _52373_ (_19843_, _19804_, _19308_);
  and _52374_ (_28213_[3], _19843_, _19842_);
  not _52375_ (_19844_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _52376_ (_19845_, _19791_, _19844_);
  and _52377_ (_19846_, _19327_, _19113_);
  or _52378_ (_19847_, _19846_, _19845_);
  or _52379_ (_19848_, _19847_, _19789_);
  and _52380_ (_19849_, _19062_, word_in[12]);
  not _52381_ (_19850_, _19789_);
  or _52382_ (_19851_, _19850_, _19849_);
  and _52383_ (_19852_, _19851_, _19848_);
  or _52384_ (_19853_, _19852_, _19786_);
  or _52385_ (_19854_, _19787_, _19441_);
  and _52386_ (_19855_, _19854_, _19804_);
  and _52387_ (_19856_, _19855_, _19853_);
  and _52388_ (_19857_, _19800_, _19322_);
  or _52389_ (_28213_[4], _19857_, _19856_);
  and _52390_ (_19858_, _19786_, _19453_);
  not _52391_ (_19859_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _52392_ (_19860_, _19791_, _19859_);
  and _52393_ (_19861_, _19339_, _19113_);
  nor _52394_ (_19862_, _19861_, _19860_);
  nor _52395_ (_19863_, _19862_, _19789_);
  and _52396_ (_19864_, _19062_, word_in[13]);
  and _52397_ (_19865_, _19789_, _19864_);
  or _52398_ (_19866_, _19865_, _19863_);
  and _52399_ (_19867_, _19866_, _19787_);
  or _52400_ (_19868_, _19867_, _19858_);
  and _52401_ (_19869_, _19868_, _19804_);
  and _52402_ (_19870_, _19800_, _19348_);
  or _52403_ (_28213_[5], _19870_, _19869_);
  not _52404_ (_19871_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _52405_ (_19872_, _19791_, _19871_);
  and _52406_ (_19873_, _19355_, _19113_);
  nor _52407_ (_19874_, _19873_, _19872_);
  nor _52408_ (_19875_, _19874_, _19789_);
  and _52409_ (_19876_, _19062_, word_in[14]);
  and _52410_ (_19877_, _19789_, _19876_);
  or _52411_ (_19878_, _19877_, _19875_);
  and _52412_ (_19879_, _19878_, _19787_);
  and _52413_ (_19880_, _19786_, _19465_);
  or _52414_ (_19881_, _19880_, _19800_);
  or _52415_ (_19882_, _19881_, _19879_);
  or _52416_ (_19883_, _19804_, _19350_);
  and _52417_ (_28213_[6], _19883_, _19882_);
  and _52418_ (_19884_, _19791_, word_in[7]);
  nor _52419_ (_19885_, _19791_, _18716_);
  nor _52420_ (_19886_, _19885_, _19884_);
  nor _52421_ (_19887_, _19886_, _19789_);
  and _52422_ (_19888_, _19789_, _19074_);
  or _52423_ (_19889_, _19888_, _19887_);
  and _52424_ (_19890_, _19889_, _19787_);
  and _52425_ (_19891_, _19786_, _19477_);
  or _52426_ (_19892_, _19891_, _19800_);
  or _52427_ (_19893_, _19892_, _19890_);
  or _52428_ (_19894_, _19804_, _19081_);
  and _52429_ (_28213_[7], _19894_, _19893_);
  and _52430_ (_19895_, _19685_, _19486_);
  and _52431_ (_19896_, _19788_, _18690_);
  and _52432_ (_19897_, _19067_, _19131_);
  and _52433_ (_19898_, _19897_, word_in[0]);
  not _52434_ (_19899_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _52435_ (_19900_, _19897_, _19899_);
  nor _52436_ (_19901_, _19900_, _19898_);
  nor _52437_ (_19902_, _19901_, _19896_);
  and _52438_ (_19903_, _19896_, _19796_);
  or _52439_ (_19904_, _19903_, _19902_);
  or _52440_ (_19905_, _19904_, _19895_);
  and _52441_ (_19906_, _19682_, _18667_);
  not _52442_ (_19907_, _19906_);
  not _52443_ (_19908_, _19895_);
  or _52444_ (_19909_, _19908_, _19393_);
  and _52445_ (_19910_, _19909_, _19907_);
  and _52446_ (_19911_, _19910_, _19905_);
  and _52447_ (_19912_, _19906_, _19252_);
  or _52448_ (_28214_[0], _19912_, _19911_);
  not _52449_ (_19913_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _52450_ (_19914_, _19897_, _19913_);
  and _52451_ (_19915_, _19897_, _19286_);
  or _52452_ (_19916_, _19915_, _19914_);
  or _52453_ (_19917_, _19916_, _19896_);
  not _52454_ (_19918_, _19896_);
  or _52455_ (_19919_, _19918_, _19282_);
  and _52456_ (_19920_, _19919_, _19917_);
  or _52457_ (_19921_, _19920_, _19895_);
  or _52458_ (_19922_, _19908_, _19405_);
  and _52459_ (_19923_, _19922_, _19907_);
  and _52460_ (_19924_, _19923_, _19921_);
  and _52461_ (_19925_, _19906_, _19279_);
  or _52462_ (_28214_[1], _19925_, _19924_);
  not _52463_ (_19926_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _52464_ (_19927_, _19897_, _19926_);
  and _52465_ (_19928_, _19897_, _19299_);
  or _52466_ (_19929_, _19928_, _19927_);
  or _52467_ (_19930_, _19929_, _19896_);
  or _52468_ (_19931_, _19918_, _19823_);
  and _52469_ (_19932_, _19931_, _19930_);
  or _52470_ (_19933_, _19932_, _19895_);
  or _52471_ (_19934_, _19908_, _19417_);
  and _52472_ (_19935_, _19934_, _19933_);
  or _52473_ (_19936_, _19935_, _19906_);
  or _52474_ (_19937_, _19907_, _19294_);
  and _52475_ (_28214_[2], _19937_, _19936_);
  or _52476_ (_19938_, _19908_, _19429_);
  not _52477_ (_19939_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _52478_ (_19940_, _19897_, _19939_);
  and _52479_ (_19941_, _19897_, _19313_);
  or _52480_ (_19942_, _19941_, _19940_);
  or _52481_ (_19943_, _19942_, _19896_);
  or _52482_ (_19944_, _19918_, _19836_);
  and _52483_ (_19945_, _19944_, _19943_);
  or _52484_ (_19946_, _19945_, _19895_);
  and _52485_ (_19947_, _19946_, _19938_);
  or _52486_ (_19948_, _19947_, _19906_);
  or _52487_ (_19949_, _19907_, _19308_);
  and _52488_ (_28214_[3], _19949_, _19948_);
  not _52489_ (_19950_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _52490_ (_19951_, _19897_, _19950_);
  and _52491_ (_19952_, _19897_, _19327_);
  or _52492_ (_19953_, _19952_, _19951_);
  or _52493_ (_19954_, _19953_, _19896_);
  or _52494_ (_19955_, _19918_, _19849_);
  and _52495_ (_19956_, _19955_, _19954_);
  or _52496_ (_19957_, _19956_, _19895_);
  or _52497_ (_19958_, _19908_, _19441_);
  and _52498_ (_19959_, _19958_, _19907_);
  and _52499_ (_19960_, _19959_, _19957_);
  and _52500_ (_19961_, _19906_, _19322_);
  or _52501_ (_28214_[4], _19961_, _19960_);
  not _52502_ (_19962_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _52503_ (_19963_, _19897_, _19962_);
  and _52504_ (_19964_, _19897_, _19339_);
  or _52505_ (_19965_, _19964_, _19963_);
  or _52506_ (_19966_, _19965_, _19896_);
  or _52507_ (_19967_, _19918_, _19864_);
  and _52508_ (_19968_, _19967_, _19966_);
  or _52509_ (_19969_, _19968_, _19895_);
  or _52510_ (_19970_, _19908_, _19453_);
  and _52511_ (_19971_, _19970_, _19907_);
  and _52512_ (_19972_, _19971_, _19969_);
  and _52513_ (_19973_, _19906_, _19348_);
  or _52514_ (_28214_[5], _19973_, _19972_);
  or _52515_ (_19974_, _19908_, _19465_);
  not _52516_ (_19975_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _52517_ (_19976_, _19897_, _19975_);
  and _52518_ (_19977_, _19897_, _19355_);
  or _52519_ (_19978_, _19977_, _19976_);
  or _52520_ (_19979_, _19978_, _19896_);
  or _52521_ (_19980_, _19918_, _19876_);
  and _52522_ (_19981_, _19980_, _19979_);
  or _52523_ (_19982_, _19981_, _19895_);
  and _52524_ (_19983_, _19982_, _19974_);
  or _52525_ (_19984_, _19983_, _19906_);
  or _52526_ (_19985_, _19907_, _19350_);
  and _52527_ (_28214_[6], _19985_, _19984_);
  nor _52528_ (_19986_, _19897_, _18827_);
  and _52529_ (_19987_, _19897_, _19068_);
  or _52530_ (_19988_, _19987_, _19986_);
  or _52531_ (_19989_, _19988_, _19896_);
  or _52532_ (_19990_, _19918_, _19074_);
  and _52533_ (_19991_, _19990_, _19989_);
  or _52534_ (_19992_, _19991_, _19895_);
  or _52535_ (_19993_, _19908_, _19477_);
  and _52536_ (_19994_, _19993_, _19907_);
  and _52537_ (_19995_, _19994_, _19992_);
  and _52538_ (_19996_, _19906_, _19081_);
  or _52539_ (_28214_[7], _19996_, _19995_);
  and _52540_ (_19997_, _19252_, _19099_);
  and _52541_ (_19998_, _19685_, _19056_);
  and _52542_ (_19999_, _19788_, _18679_);
  and _52543_ (_20000_, _19067_, _18755_);
  and _52544_ (_20001_, _20000_, word_in[0]);
  not _52545_ (_20002_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _52546_ (_20003_, _20000_, _20002_);
  nor _52547_ (_20004_, _20003_, _20001_);
  nor _52548_ (_20005_, _20004_, _19999_);
  and _52549_ (_20006_, _19999_, _19796_);
  or _52550_ (_20007_, _20006_, _20005_);
  or _52551_ (_20008_, _20007_, _19998_);
  and _52552_ (_20009_, _19050_, _19099_);
  not _52553_ (_20010_, _20009_);
  not _52554_ (_20011_, _19998_);
  or _52555_ (_20012_, _20011_, _19393_);
  and _52556_ (_20013_, _20012_, _20010_);
  and _52557_ (_20014_, _20013_, _20008_);
  or _52558_ (_28215_[0], _20014_, _19997_);
  and _52559_ (_20015_, _19279_, _19099_);
  not _52560_ (_20016_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _52561_ (_20017_, _20000_, _20016_);
  and _52562_ (_20018_, _20000_, _19286_);
  or _52563_ (_20019_, _20018_, _20017_);
  or _52564_ (_20020_, _20019_, _19999_);
  not _52565_ (_20021_, _19999_);
  or _52566_ (_20022_, _20021_, _19282_);
  and _52567_ (_20023_, _20022_, _20020_);
  or _52568_ (_20024_, _20023_, _19998_);
  or _52569_ (_20025_, _20011_, _19405_);
  and _52570_ (_20026_, _20025_, _20010_);
  and _52571_ (_20027_, _20026_, _20024_);
  or _52572_ (_28215_[1], _20027_, _20015_);
  and _52573_ (_20028_, _19294_, _19099_);
  and _52574_ (_20029_, _20000_, word_in[2]);
  not _52575_ (_20030_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _52576_ (_20031_, _20000_, _20030_);
  nor _52577_ (_20032_, _20031_, _20029_);
  nor _52578_ (_20033_, _20032_, _19999_);
  and _52579_ (_20034_, _19999_, _19823_);
  or _52580_ (_20035_, _20034_, _20033_);
  or _52581_ (_20036_, _20035_, _19998_);
  or _52582_ (_20037_, _20011_, _19417_);
  and _52583_ (_20038_, _20037_, _20010_);
  and _52584_ (_20039_, _20038_, _20036_);
  or _52585_ (_28215_[2], _20039_, _20028_);
  and _52586_ (_20040_, _19308_, _19099_);
  and _52587_ (_20041_, _20000_, word_in[3]);
  not _52588_ (_20042_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _52589_ (_20043_, _20000_, _20042_);
  nor _52590_ (_20044_, _20043_, _20041_);
  nor _52591_ (_20045_, _20044_, _19999_);
  and _52592_ (_20046_, _19999_, _19836_);
  or _52593_ (_20047_, _20046_, _20045_);
  or _52594_ (_20048_, _20047_, _19998_);
  or _52595_ (_20049_, _20011_, _19429_);
  and _52596_ (_20050_, _20049_, _20010_);
  and _52597_ (_20051_, _20050_, _20048_);
  or _52598_ (_28215_[3], _20051_, _20040_);
  and _52599_ (_20052_, _20000_, word_in[4]);
  not _52600_ (_20053_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _52601_ (_20054_, _20000_, _20053_);
  nor _52602_ (_20055_, _20054_, _20052_);
  nor _52603_ (_20056_, _20055_, _19999_);
  and _52604_ (_20057_, _19999_, _19849_);
  or _52605_ (_20058_, _20057_, _20056_);
  and _52606_ (_20059_, _20058_, _20011_);
  and _52607_ (_20060_, _19998_, _19441_);
  or _52608_ (_20061_, _20060_, _20059_);
  and _52609_ (_20062_, _20061_, _20010_);
  and _52610_ (_20063_, _20009_, word_in[28]);
  or _52611_ (_28215_[4], _20063_, _20062_);
  and _52612_ (_20064_, _20009_, word_in[29]);
  and _52613_ (_20065_, _20000_, word_in[5]);
  not _52614_ (_20066_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _52615_ (_20067_, _20000_, _20066_);
  nor _52616_ (_20068_, _20067_, _20065_);
  nor _52617_ (_20069_, _20068_, _19999_);
  and _52618_ (_20070_, _19999_, _19864_);
  or _52619_ (_20071_, _20070_, _20069_);
  or _52620_ (_20072_, _20071_, _19998_);
  or _52621_ (_20073_, _20011_, _19453_);
  and _52622_ (_20074_, _20073_, _20010_);
  and _52623_ (_20075_, _20074_, _20072_);
  or _52624_ (_28215_[5], _20075_, _20064_);
  not _52625_ (_20076_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _52626_ (_20077_, _20000_, _20076_);
  and _52627_ (_20078_, _20000_, _19355_);
  or _52628_ (_20079_, _20078_, _20077_);
  or _52629_ (_20080_, _20079_, _19999_);
  or _52630_ (_20081_, _20021_, _19876_);
  and _52631_ (_20082_, _20081_, _20080_);
  or _52632_ (_20083_, _20082_, _19998_);
  or _52633_ (_20084_, _20011_, _19465_);
  and _52634_ (_20085_, _20084_, _20083_);
  or _52635_ (_20086_, _20085_, _20009_);
  or _52636_ (_20087_, _20010_, word_in[30]);
  and _52637_ (_28215_[6], _20087_, _20086_);
  and _52638_ (_20088_, _20009_, word_in[31]);
  and _52639_ (_20089_, _20000_, word_in[7]);
  nor _52640_ (_20090_, _20000_, _18695_);
  nor _52641_ (_20091_, _20090_, _20089_);
  nor _52642_ (_20092_, _20091_, _19999_);
  and _52643_ (_20093_, _19999_, _19074_);
  or _52644_ (_20094_, _20093_, _20092_);
  or _52645_ (_20095_, _20094_, _19998_);
  or _52646_ (_20096_, _20011_, _19477_);
  and _52647_ (_20097_, _20096_, _20010_);
  and _52648_ (_20098_, _20097_, _20095_);
  or _52649_ (_28215_[7], _20098_, _20088_);
  and _52650_ (_20099_, _19051_, _18973_);
  and _52651_ (_20100_, _20099_, _18690_);
  not _52652_ (_20101_, _20100_);
  and _52653_ (_20102_, _18689_, _18645_);
  or _52654_ (_20103_, _20102_, _18701_);
  and _52655_ (_20104_, _20103_, _19057_);
  and _52656_ (_20105_, _20104_, _19258_);
  and _52657_ (_20106_, _19062_, _18755_);
  and _52658_ (_20107_, _19067_, _19163_);
  and _52659_ (_20108_, _20107_, word_in[0]);
  not _52660_ (_20109_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _52661_ (_20110_, _20107_, _20109_);
  nor _52662_ (_20111_, _20110_, _20108_);
  nor _52663_ (_20112_, _20111_, _20106_);
  and _52664_ (_20113_, _20106_, word_in[8]);
  nor _52665_ (_20114_, _20113_, _20112_);
  nor _52666_ (_20115_, _20114_, _20105_);
  and _52667_ (_20116_, _20105_, word_in[16]);
  or _52668_ (_20117_, _20116_, _20115_);
  and _52669_ (_20118_, _20117_, _20101_);
  and _52670_ (_20119_, _20100_, _19252_);
  or _52671_ (_28216_[0], _20119_, _20118_);
  not _52672_ (_20120_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _52673_ (_20121_, _20107_, _20120_);
  and _52674_ (_20122_, _20107_, _19286_);
  or _52675_ (_20123_, _20122_, _20121_);
  or _52676_ (_20124_, _20123_, _20106_);
  not _52677_ (_20125_, _20106_);
  or _52678_ (_20126_, _20125_, word_in[9]);
  and _52679_ (_20127_, _20126_, _20124_);
  or _52680_ (_20128_, _20127_, _20105_);
  not _52681_ (_20129_, _20105_);
  or _52682_ (_20130_, _20129_, word_in[17]);
  and _52683_ (_20131_, _20130_, _20128_);
  or _52684_ (_20132_, _20131_, _20100_);
  or _52685_ (_20133_, _20101_, _19279_);
  and _52686_ (_28216_[1], _20133_, _20132_);
  and _52687_ (_20134_, _20107_, word_in[2]);
  not _52688_ (_20135_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _52689_ (_20136_, _20107_, _20135_);
  nor _52690_ (_20137_, _20136_, _20134_);
  nor _52691_ (_20138_, _20137_, _20106_);
  and _52692_ (_20139_, _20106_, word_in[10]);
  nor _52693_ (_20140_, _20139_, _20138_);
  nor _52694_ (_20141_, _20140_, _20105_);
  and _52695_ (_20142_, _20105_, word_in[18]);
  or _52696_ (_20143_, _20142_, _20141_);
  and _52697_ (_20144_, _20143_, _20101_);
  and _52698_ (_20145_, _20100_, _19294_);
  or _52699_ (_28216_[2], _20145_, _20144_);
  and _52700_ (_20146_, _20107_, word_in[3]);
  not _52701_ (_20147_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _52702_ (_20148_, _20107_, _20147_);
  nor _52703_ (_20149_, _20148_, _20146_);
  nor _52704_ (_20150_, _20149_, _20106_);
  and _52705_ (_20151_, _20106_, word_in[11]);
  nor _52706_ (_20152_, _20151_, _20150_);
  nor _52707_ (_20153_, _20152_, _20105_);
  and _52708_ (_20154_, _20105_, word_in[19]);
  or _52709_ (_20155_, _20154_, _20153_);
  and _52710_ (_20156_, _20155_, _20101_);
  and _52711_ (_20157_, _20100_, _19308_);
  or _52712_ (_28216_[3], _20157_, _20156_);
  not _52713_ (_20158_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _52714_ (_20159_, _20107_, _20158_);
  and _52715_ (_20160_, _20107_, _19327_);
  or _52716_ (_20161_, _20160_, _20159_);
  or _52717_ (_20162_, _20161_, _20106_);
  or _52718_ (_20163_, _20125_, word_in[12]);
  and _52719_ (_20164_, _20163_, _20162_);
  or _52720_ (_20165_, _20164_, _20105_);
  or _52721_ (_20166_, _20129_, word_in[20]);
  and _52722_ (_20167_, _20166_, _20165_);
  or _52723_ (_20168_, _20167_, _20100_);
  or _52724_ (_20169_, _20101_, _19322_);
  and _52725_ (_28216_[4], _20169_, _20168_);
  not _52726_ (_20170_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _52727_ (_20171_, _20107_, _20170_);
  and _52728_ (_20172_, _20107_, _19339_);
  or _52729_ (_20173_, _20172_, _20171_);
  or _52730_ (_20174_, _20173_, _20106_);
  or _52731_ (_20175_, _20125_, word_in[13]);
  and _52732_ (_20176_, _20175_, _20174_);
  or _52733_ (_20177_, _20176_, _20105_);
  or _52734_ (_20178_, _20129_, word_in[21]);
  and _52735_ (_20179_, _20178_, _20177_);
  or _52736_ (_20180_, _20179_, _20100_);
  or _52737_ (_20181_, _20101_, _19348_);
  and _52738_ (_28216_[5], _20181_, _20180_);
  not _52739_ (_20182_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _52740_ (_20183_, _20107_, _20182_);
  and _52741_ (_20184_, _20107_, _19355_);
  or _52742_ (_20185_, _20184_, _20183_);
  or _52743_ (_20186_, _20185_, _20106_);
  or _52744_ (_20187_, _20125_, word_in[14]);
  and _52745_ (_20188_, _20187_, _20186_);
  or _52746_ (_20189_, _20188_, _20105_);
  or _52747_ (_20190_, _20129_, word_in[22]);
  and _52748_ (_20191_, _20190_, _20189_);
  or _52749_ (_20192_, _20191_, _20100_);
  or _52750_ (_20193_, _20101_, _19350_);
  and _52751_ (_28216_[6], _20193_, _20192_);
  and _52752_ (_20194_, _20107_, word_in[7]);
  nor _52753_ (_20195_, _20107_, _18836_);
  nor _52754_ (_20196_, _20195_, _20194_);
  nor _52755_ (_20197_, _20196_, _20106_);
  and _52756_ (_20198_, _20106_, word_in[15]);
  nor _52757_ (_20199_, _20198_, _20197_);
  nor _52758_ (_20200_, _20199_, _20105_);
  and _52759_ (_20201_, _20105_, word_in[23]);
  or _52760_ (_20202_, _20201_, _20200_);
  and _52761_ (_20203_, _20202_, _20101_);
  and _52762_ (_20204_, _20100_, _19081_);
  or _52763_ (_28216_[7], _20204_, _20203_);
  and _52764_ (_20205_, _20104_, _19379_);
  and _52765_ (_20206_, _19062_, _18768_);
  and _52766_ (_20207_, _20206_, _18657_);
  and _52767_ (_20208_, _19266_, _19169_);
  not _52768_ (_20209_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _52769_ (_20210_, _19067_, _19169_);
  nor _52770_ (_20211_, _20210_, _20209_);
  nor _52771_ (_20212_, _20211_, _20208_);
  nor _52772_ (_20213_, _20212_, _20207_);
  and _52773_ (_20214_, _20207_, word_in[8]);
  nor _52774_ (_20215_, _20214_, _20213_);
  nor _52775_ (_20216_, _20215_, _20205_);
  and _52776_ (_20217_, _20099_, _18679_);
  and _52777_ (_20218_, _20205_, _19393_);
  or _52778_ (_20219_, _20218_, _20217_);
  or _52779_ (_20220_, _20219_, _20216_);
  not _52780_ (_20221_, _20217_);
  or _52781_ (_20222_, _20221_, _19252_);
  and _52782_ (_28217_[0], _20222_, _20220_);
  not _52783_ (_20223_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _52784_ (_20224_, _20210_, _20223_);
  and _52785_ (_20225_, _19286_, _19169_);
  or _52786_ (_20226_, _20225_, _20224_);
  or _52787_ (_20227_, _20226_, _20207_);
  not _52788_ (_20228_, _20207_);
  or _52789_ (_20229_, _20228_, word_in[9]);
  and _52790_ (_20230_, _20229_, _20227_);
  or _52791_ (_20231_, _20230_, _20205_);
  not _52792_ (_20232_, _20205_);
  or _52793_ (_20233_, _20232_, _19405_);
  and _52794_ (_20234_, _20233_, _20231_);
  or _52795_ (_20235_, _20234_, _20217_);
  or _52796_ (_20236_, _20221_, _19279_);
  and _52797_ (_28217_[1], _20236_, _20235_);
  not _52798_ (_20237_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _52799_ (_20238_, _20210_, _20237_);
  and _52800_ (_20239_, _19299_, _19169_);
  or _52801_ (_20240_, _20239_, _20238_);
  or _52802_ (_20241_, _20240_, _20207_);
  or _52803_ (_20242_, _20228_, word_in[10]);
  and _52804_ (_20243_, _20242_, _20241_);
  or _52805_ (_20244_, _20243_, _20205_);
  or _52806_ (_20245_, _20232_, _19417_);
  and _52807_ (_20246_, _20245_, _20244_);
  or _52808_ (_20247_, _20246_, _20217_);
  or _52809_ (_20248_, _20221_, _19294_);
  and _52810_ (_28217_[2], _20248_, _20247_);
  not _52811_ (_20249_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _52812_ (_20250_, _20210_, _20249_);
  and _52813_ (_20251_, _19313_, _19169_);
  nor _52814_ (_20252_, _20251_, _20250_);
  nor _52815_ (_20253_, _20252_, _20207_);
  and _52816_ (_20254_, _20207_, word_in[11]);
  nor _52817_ (_20255_, _20254_, _20253_);
  nor _52818_ (_20256_, _20255_, _20205_);
  and _52819_ (_20257_, _20205_, _19429_);
  or _52820_ (_20258_, _20257_, _20256_);
  and _52821_ (_20259_, _20258_, _20221_);
  and _52822_ (_20260_, _20217_, _19308_);
  or _52823_ (_28217_[3], _20260_, _20259_);
  not _52824_ (_20261_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _52825_ (_20262_, _20210_, _20261_);
  and _52826_ (_20263_, _19327_, _19169_);
  or _52827_ (_20264_, _20263_, _20262_);
  or _52828_ (_20265_, _20264_, _20207_);
  or _52829_ (_20266_, _20228_, word_in[12]);
  and _52830_ (_20267_, _20266_, _20265_);
  or _52831_ (_20268_, _20267_, _20205_);
  or _52832_ (_20269_, _20232_, _19441_);
  and _52833_ (_20270_, _20269_, _20268_);
  or _52834_ (_20271_, _20270_, _20217_);
  or _52835_ (_20272_, _20221_, _19322_);
  and _52836_ (_28217_[4], _20272_, _20271_);
  not _52837_ (_20273_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _52838_ (_20274_, _20210_, _20273_);
  and _52839_ (_20275_, _20210_, _19339_);
  or _52840_ (_20276_, _20275_, _20274_);
  or _52841_ (_20277_, _20276_, _20207_);
  or _52842_ (_20278_, _20228_, word_in[13]);
  and _52843_ (_20279_, _20278_, _20277_);
  or _52844_ (_20280_, _20279_, _20205_);
  or _52845_ (_20281_, _20232_, _19453_);
  and _52846_ (_20282_, _20281_, _20221_);
  and _52847_ (_20283_, _20282_, _20280_);
  and _52848_ (_20284_, _20217_, _19348_);
  or _52849_ (_28217_[5], _20284_, _20283_);
  and _52850_ (_20285_, _20210_, word_in[6]);
  not _52851_ (_20286_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _52852_ (_20287_, _20210_, _20286_);
  nor _52853_ (_20288_, _20287_, _20285_);
  nor _52854_ (_20289_, _20288_, _20207_);
  and _52855_ (_20290_, _20207_, word_in[14]);
  or _52856_ (_20291_, _20290_, _20289_);
  or _52857_ (_20292_, _20291_, _20205_);
  or _52858_ (_20293_, _20232_, _19465_);
  and _52859_ (_20294_, _20293_, _20221_);
  and _52860_ (_20295_, _20294_, _20292_);
  and _52861_ (_20296_, _20217_, _19350_);
  or _52862_ (_28217_[6], _20296_, _20295_);
  and _52863_ (_20297_, _20210_, word_in[7]);
  nor _52864_ (_20298_, _20210_, _18728_);
  nor _52865_ (_20299_, _20298_, _20297_);
  nor _52866_ (_20300_, _20299_, _20207_);
  and _52867_ (_20301_, _20207_, word_in[15]);
  nor _52868_ (_20302_, _20301_, _20300_);
  nor _52869_ (_20303_, _20302_, _20205_);
  and _52870_ (_20304_, _20205_, _19477_);
  or _52871_ (_20305_, _20304_, _20303_);
  and _52872_ (_20306_, _20305_, _20221_);
  and _52873_ (_20307_, _20217_, _19081_);
  or _52874_ (_28217_[7], _20307_, _20306_);
  and _52875_ (_20308_, _19051_, _18753_);
  not _52876_ (_20309_, _20308_);
  and _52877_ (_20310_, _20104_, _19486_);
  and _52878_ (_20311_, _20206_, _18690_);
  not _52879_ (_20312_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _52880_ (_20313_, _19067_, _19180_);
  nor _52881_ (_20314_, _20313_, _20312_);
  and _52882_ (_20315_, _20313_, _19266_);
  nor _52883_ (_20316_, _20315_, _20314_);
  nor _52884_ (_20317_, _20316_, _20311_);
  and _52885_ (_20318_, _20311_, word_in[8]);
  nor _52886_ (_20319_, _20318_, _20317_);
  nor _52887_ (_20320_, _20319_, _20310_);
  and _52888_ (_20321_, _20310_, _19393_);
  or _52889_ (_20322_, _20321_, _20320_);
  and _52890_ (_20323_, _20322_, _20309_);
  and _52891_ (_20324_, _20308_, _19252_);
  or _52892_ (_28203_[0], _20324_, _20323_);
  not _52893_ (_20325_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _52894_ (_20326_, _20313_, _20325_);
  and _52895_ (_20327_, _20313_, _19286_);
  or _52896_ (_20328_, _20327_, _20326_);
  or _52897_ (_20329_, _20328_, _20311_);
  not _52898_ (_20330_, _20311_);
  or _52899_ (_20331_, _20330_, word_in[9]);
  and _52900_ (_20332_, _20331_, _20329_);
  or _52901_ (_20333_, _20332_, _20310_);
  not _52902_ (_20334_, _20310_);
  or _52903_ (_20335_, _20334_, _19405_);
  and _52904_ (_20336_, _20335_, _20309_);
  and _52905_ (_20337_, _20336_, _20333_);
  and _52906_ (_20338_, _20308_, _19279_);
  or _52907_ (_28203_[1], _20338_, _20337_);
  not _52908_ (_20339_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _52909_ (_20340_, _20313_, _20339_);
  and _52910_ (_20341_, _20313_, _19299_);
  or _52911_ (_20342_, _20341_, _20340_);
  or _52912_ (_20343_, _20342_, _20311_);
  or _52913_ (_20344_, _20330_, word_in[10]);
  and _52914_ (_20345_, _20344_, _20343_);
  or _52915_ (_20346_, _20345_, _20310_);
  or _52916_ (_20347_, _20334_, _19417_);
  and _52917_ (_20348_, _20347_, _20309_);
  and _52918_ (_20349_, _20348_, _20346_);
  and _52919_ (_20350_, _20308_, _19294_);
  or _52920_ (_28203_[2], _20350_, _20349_);
  and _52921_ (_20351_, _20310_, _19429_);
  and _52922_ (_20352_, _20313_, word_in[3]);
  not _52923_ (_20353_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _52924_ (_20354_, _20313_, _20353_);
  nor _52925_ (_20355_, _20354_, _20352_);
  nor _52926_ (_20356_, _20355_, _20311_);
  and _52927_ (_20357_, _20311_, word_in[11]);
  nor _52928_ (_20358_, _20357_, _20356_);
  nor _52929_ (_20359_, _20358_, _20310_);
  or _52930_ (_20360_, _20359_, _20351_);
  and _52931_ (_20361_, _20360_, _20309_);
  and _52932_ (_20362_, _20308_, _19308_);
  or _52933_ (_28203_[3], _20362_, _20361_);
  not _52934_ (_20363_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _52935_ (_20364_, _20313_, _20363_);
  and _52936_ (_20365_, _20313_, _19327_);
  or _52937_ (_20366_, _20365_, _20364_);
  or _52938_ (_20367_, _20366_, _20311_);
  or _52939_ (_20368_, _20330_, word_in[12]);
  nand _52940_ (_20369_, _20368_, _20367_);
  nor _52941_ (_20370_, _20369_, _20310_);
  and _52942_ (_20371_, _20310_, _19441_);
  or _52943_ (_20372_, _20371_, _20308_);
  or _52944_ (_20373_, _20372_, _20370_);
  or _52945_ (_20374_, _20309_, _19322_);
  and _52946_ (_28203_[4], _20374_, _20373_);
  not _52947_ (_20375_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _52948_ (_20376_, _20313_, _20375_);
  and _52949_ (_20377_, _20313_, _19339_);
  or _52950_ (_20378_, _20377_, _20376_);
  or _52951_ (_20379_, _20378_, _20311_);
  or _52952_ (_20380_, _20330_, word_in[13]);
  and _52953_ (_20381_, _20380_, _20379_);
  or _52954_ (_20382_, _20381_, _20310_);
  or _52955_ (_20383_, _20334_, _19453_);
  and _52956_ (_20384_, _20383_, _20309_);
  and _52957_ (_20385_, _20384_, _20382_);
  and _52958_ (_20386_, _20308_, _19348_);
  or _52959_ (_28203_[5], _20386_, _20385_);
  and _52960_ (_20387_, _20313_, word_in[6]);
  not _52961_ (_20388_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _52962_ (_20389_, _20313_, _20388_);
  nor _52963_ (_20390_, _20389_, _20387_);
  nor _52964_ (_20391_, _20390_, _20311_);
  and _52965_ (_20392_, _20311_, word_in[14]);
  or _52966_ (_20393_, _20392_, _20391_);
  or _52967_ (_20394_, _20393_, _20310_);
  or _52968_ (_20395_, _20334_, _19465_);
  and _52969_ (_20396_, _20395_, _20309_);
  and _52970_ (_20397_, _20396_, _20394_);
  and _52971_ (_20398_, _20308_, _19350_);
  or _52972_ (_28203_[6], _20398_, _20397_);
  nor _52973_ (_20399_, _20313_, _18841_);
  and _52974_ (_20400_, _20313_, _19068_);
  or _52975_ (_20401_, _20400_, _20399_);
  or _52976_ (_20402_, _20401_, _20311_);
  or _52977_ (_20403_, _20330_, word_in[15]);
  and _52978_ (_20404_, _20403_, _20402_);
  or _52979_ (_20405_, _20404_, _20310_);
  or _52980_ (_20406_, _20334_, _19477_);
  and _52981_ (_20407_, _20406_, _20309_);
  and _52982_ (_20408_, _20407_, _20405_);
  and _52983_ (_20409_, _20308_, _19081_);
  or _52984_ (_28203_[7], _20409_, _20408_);
  and _52985_ (_20410_, _20104_, _19056_);
  and _52986_ (_20411_, _20206_, _18679_);
  not _52987_ (_20412_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _52988_ (_20413_, _19067_, _19205_);
  nor _52989_ (_20414_, _20413_, _20412_);
  and _52990_ (_20415_, _20413_, _19266_);
  or _52991_ (_20416_, _20415_, _20414_);
  or _52992_ (_20417_, _20416_, _20411_);
  not _52993_ (_20418_, _20411_);
  or _52994_ (_20419_, _20418_, word_in[8]);
  and _52995_ (_20420_, _20419_, _20417_);
  or _52996_ (_20421_, _20420_, _20410_);
  and _52997_ (_20422_, _19050_, _19163_);
  not _52998_ (_20423_, _20422_);
  not _52999_ (_20424_, _20410_);
  or _53000_ (_20425_, _20424_, word_in[16]);
  and _53001_ (_20426_, _20425_, _20423_);
  and _53002_ (_20427_, _20426_, _20421_);
  and _53003_ (_20428_, _20422_, word_in[24]);
  or _53004_ (_28204_[0], _20428_, _20427_);
  not _53005_ (_20429_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _53006_ (_20430_, _20413_, _20429_);
  and _53007_ (_20431_, _20413_, _19286_);
  or _53008_ (_20432_, _20431_, _20430_);
  or _53009_ (_20433_, _20432_, _20411_);
  or _53010_ (_20434_, _20418_, word_in[9]);
  and _53011_ (_20435_, _20434_, _20433_);
  or _53012_ (_20436_, _20435_, _20410_);
  or _53013_ (_20437_, _20424_, word_in[17]);
  and _53014_ (_20438_, _20437_, _20423_);
  and _53015_ (_20439_, _20438_, _20436_);
  and _53016_ (_20440_, _20422_, word_in[25]);
  or _53017_ (_28204_[1], _20440_, _20439_);
  and _53018_ (_20441_, _20413_, word_in[2]);
  not _53019_ (_20442_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _53020_ (_20443_, _20413_, _20442_);
  nor _53021_ (_20444_, _20443_, _20441_);
  nor _53022_ (_20445_, _20444_, _20411_);
  and _53023_ (_20446_, _20411_, word_in[10]);
  nor _53024_ (_20447_, _20446_, _20445_);
  nor _53025_ (_20448_, _20447_, _20410_);
  and _53026_ (_20449_, _20410_, word_in[18]);
  or _53027_ (_20450_, _20449_, _20448_);
  and _53028_ (_20451_, _20450_, _20423_);
  and _53029_ (_20452_, _20422_, word_in[26]);
  or _53030_ (_28204_[2], _20452_, _20451_);
  not _53031_ (_20453_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _53032_ (_20454_, _20413_, _20453_);
  and _53033_ (_20455_, _20413_, _19313_);
  or _53034_ (_20456_, _20455_, _20454_);
  or _53035_ (_20457_, _20456_, _20411_);
  or _53036_ (_20458_, _20418_, word_in[11]);
  and _53037_ (_20459_, _20458_, _20457_);
  or _53038_ (_20460_, _20459_, _20410_);
  or _53039_ (_20461_, _20424_, word_in[19]);
  and _53040_ (_20462_, _20461_, _20423_);
  and _53041_ (_20463_, _20462_, _20460_);
  and _53042_ (_20464_, _20422_, word_in[27]);
  or _53043_ (_28204_[3], _20464_, _20463_);
  not _53044_ (_20465_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _53045_ (_20466_, _20413_, _20465_);
  and _53046_ (_20467_, _20413_, _19327_);
  or _53047_ (_20468_, _20467_, _20466_);
  or _53048_ (_20469_, _20468_, _20411_);
  or _53049_ (_20470_, _20418_, word_in[12]);
  and _53050_ (_20471_, _20470_, _20469_);
  or _53051_ (_20472_, _20471_, _20410_);
  or _53052_ (_20473_, _20424_, word_in[20]);
  and _53053_ (_20474_, _20473_, _20423_);
  and _53054_ (_20475_, _20474_, _20472_);
  and _53055_ (_20476_, _20422_, word_in[28]);
  or _53056_ (_28204_[4], _20476_, _20475_);
  not _53057_ (_20477_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _53058_ (_20478_, _20413_, _20477_);
  and _53059_ (_20479_, _20413_, _19339_);
  or _53060_ (_20480_, _20479_, _20478_);
  or _53061_ (_20481_, _20480_, _20411_);
  or _53062_ (_20482_, _20418_, word_in[13]);
  and _53063_ (_20483_, _20482_, _20481_);
  or _53064_ (_20484_, _20483_, _20410_);
  or _53065_ (_20485_, _20424_, _19453_);
  and _53066_ (_20486_, _20485_, _20423_);
  and _53067_ (_20487_, _20486_, _20484_);
  and _53068_ (_20488_, _20422_, word_in[29]);
  or _53069_ (_28204_[5], _20488_, _20487_);
  and _53070_ (_20489_, _20413_, word_in[6]);
  not _53071_ (_20490_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _53072_ (_20491_, _20413_, _20490_);
  nor _53073_ (_20492_, _20491_, _20489_);
  nor _53074_ (_20493_, _20492_, _20411_);
  and _53075_ (_20494_, _20411_, word_in[14]);
  nor _53076_ (_20495_, _20494_, _20493_);
  nor _53077_ (_20496_, _20495_, _20410_);
  and _53078_ (_20497_, _20410_, word_in[22]);
  or _53079_ (_20498_, _20497_, _20496_);
  and _53080_ (_20499_, _20498_, _20423_);
  and _53081_ (_20500_, _20422_, word_in[30]);
  or _53082_ (_28204_[6], _20500_, _20499_);
  nor _53083_ (_20501_, _20413_, _18723_);
  and _53084_ (_20502_, _20413_, _19068_);
  or _53085_ (_20503_, _20502_, _20501_);
  or _53086_ (_20504_, _20503_, _20411_);
  or _53087_ (_20505_, _20418_, word_in[15]);
  and _53088_ (_20506_, _20505_, _20504_);
  or _53089_ (_20507_, _20506_, _20410_);
  or _53090_ (_20508_, _20424_, word_in[23]);
  and _53091_ (_20509_, _20508_, _20423_);
  and _53092_ (_20510_, _20509_, _20507_);
  and _53093_ (_20511_, _20422_, word_in[31]);
  or _53094_ (_28204_[7], _20511_, _20510_);
  and _53095_ (_20512_, _19052_, _18690_);
  and _53096_ (_20513_, _19258_, _19059_);
  and _53097_ (_20514_, _19062_, _19205_);
  and _53098_ (_20515_, _18657_, _18647_);
  and _53099_ (_20516_, _19067_, _20515_);
  and _53100_ (_20517_, _20516_, _19266_);
  not _53101_ (_20518_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _53102_ (_20519_, _20516_, _20518_);
  or _53103_ (_20520_, _20519_, _20517_);
  or _53104_ (_20521_, _20520_, _20514_);
  not _53105_ (_20522_, _20514_);
  or _53106_ (_20523_, _20522_, word_in[8]);
  and _53107_ (_20524_, _20523_, _20521_);
  or _53108_ (_20525_, _20524_, _20513_);
  not _53109_ (_20526_, _20513_);
  or _53110_ (_20527_, _20526_, word_in[16]);
  and _53111_ (_20528_, _20527_, _20525_);
  or _53112_ (_20529_, _20528_, _20512_);
  not _53113_ (_20530_, _20512_);
  or _53114_ (_20531_, _20530_, _19252_);
  and _53115_ (_28205_[0], _20531_, _20529_);
  not _53116_ (_20532_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _53117_ (_20533_, _20516_, _20532_);
  and _53118_ (_20534_, _20516_, _19286_);
  nor _53119_ (_20535_, _20534_, _20533_);
  nor _53120_ (_20536_, _20535_, _20514_);
  and _53121_ (_20537_, _20514_, word_in[9]);
  nor _53122_ (_20538_, _20537_, _20536_);
  nor _53123_ (_20539_, _20538_, _20513_);
  and _53124_ (_20540_, _20513_, word_in[17]);
  or _53125_ (_20541_, _20540_, _20539_);
  and _53126_ (_20542_, _20541_, _20530_);
  and _53127_ (_20543_, _20512_, _19279_);
  or _53128_ (_28205_[1], _20543_, _20542_);
  not _53129_ (_20544_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _53130_ (_20545_, _20516_, _20544_);
  and _53131_ (_20546_, _20516_, _19299_);
  or _53132_ (_20547_, _20546_, _20545_);
  or _53133_ (_20548_, _20547_, _20514_);
  or _53134_ (_20549_, _20522_, word_in[10]);
  and _53135_ (_20550_, _20549_, _20548_);
  or _53136_ (_20551_, _20550_, _20513_);
  or _53137_ (_20552_, _20526_, word_in[18]);
  and _53138_ (_20553_, _20552_, _20551_);
  or _53139_ (_20554_, _20553_, _20512_);
  or _53140_ (_20555_, _20530_, _19294_);
  and _53141_ (_28205_[2], _20555_, _20554_);
  and _53142_ (_20556_, _20516_, word_in[3]);
  not _53143_ (_20557_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _53144_ (_20558_, _20516_, _20557_);
  nor _53145_ (_20559_, _20558_, _20556_);
  nor _53146_ (_20560_, _20559_, _20514_);
  and _53147_ (_20561_, _20514_, word_in[11]);
  nor _53148_ (_20562_, _20561_, _20560_);
  nor _53149_ (_20563_, _20562_, _20513_);
  and _53150_ (_20564_, _20513_, word_in[19]);
  or _53151_ (_20565_, _20564_, _20563_);
  and _53152_ (_20566_, _20565_, _20530_);
  and _53153_ (_20567_, _20512_, _19308_);
  or _53154_ (_28205_[3], _20567_, _20566_);
  not _53155_ (_20568_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _53156_ (_20569_, _20516_, _20568_);
  and _53157_ (_20570_, _20516_, _19327_);
  or _53158_ (_20571_, _20570_, _20569_);
  or _53159_ (_20572_, _20571_, _20514_);
  or _53160_ (_20573_, _20522_, word_in[12]);
  and _53161_ (_20574_, _20573_, _20572_);
  or _53162_ (_20575_, _20574_, _20513_);
  or _53163_ (_20576_, _20526_, word_in[20]);
  and _53164_ (_20577_, _20576_, _20575_);
  or _53165_ (_20578_, _20577_, _20512_);
  or _53166_ (_20579_, _20530_, _19322_);
  and _53167_ (_28205_[4], _20579_, _20578_);
  not _53168_ (_20580_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _53169_ (_20581_, _20516_, _20580_);
  and _53170_ (_20582_, _20516_, word_in[5]);
  nor _53171_ (_20583_, _20582_, _20581_);
  nor _53172_ (_20584_, _20583_, _20514_);
  and _53173_ (_20585_, _20514_, word_in[13]);
  nor _53174_ (_20586_, _20585_, _20584_);
  nor _53175_ (_20587_, _20586_, _20513_);
  and _53176_ (_20588_, _20513_, word_in[21]);
  or _53177_ (_20589_, _20588_, _20587_);
  and _53178_ (_20590_, _20589_, _20530_);
  and _53179_ (_20591_, _20512_, _19348_);
  or _53180_ (_28205_[5], _20591_, _20590_);
  and _53181_ (_20592_, _20516_, word_in[6]);
  not _53182_ (_20593_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _53183_ (_20594_, _20516_, _20593_);
  nor _53184_ (_20595_, _20594_, _20592_);
  nor _53185_ (_20596_, _20595_, _20514_);
  and _53186_ (_20597_, _20514_, word_in[14]);
  nor _53187_ (_20598_, _20597_, _20596_);
  nor _53188_ (_20599_, _20598_, _20513_);
  and _53189_ (_20600_, _20513_, word_in[22]);
  or _53190_ (_20601_, _20600_, _20599_);
  and _53191_ (_20602_, _20601_, _20530_);
  and _53192_ (_20603_, _20512_, _19350_);
  or _53193_ (_28205_[6], _20603_, _20602_);
  nor _53194_ (_20604_, _20516_, _18848_);
  and _53195_ (_20605_, _20516_, _19068_);
  or _53196_ (_20606_, _20605_, _20604_);
  or _53197_ (_20607_, _20606_, _20514_);
  or _53198_ (_20608_, _20522_, word_in[15]);
  and _53199_ (_20609_, _20608_, _20607_);
  or _53200_ (_20610_, _20609_, _20513_);
  or _53201_ (_20611_, _20526_, word_in[23]);
  and _53202_ (_20612_, _20611_, _20610_);
  or _53203_ (_20613_, _20612_, _20512_);
  or _53204_ (_20614_, _20530_, _19081_);
  and _53205_ (_28205_[7], _20614_, _20613_);
  and _53206_ (_20615_, _19052_, _18679_);
  not _53207_ (_20616_, _20615_);
  and _53208_ (_20617_, _19379_, _19059_);
  not _53209_ (_20618_, _20617_);
  and _53210_ (_20619_, _19064_, _18657_);
  not _53211_ (_20620_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _53212_ (_20621_, _19067_, _19233_);
  nor _53213_ (_20622_, _20621_, _20620_);
  and _53214_ (_20623_, _19266_, _19233_);
  nor _53215_ (_20624_, _20623_, _20622_);
  nor _53216_ (_20625_, _20624_, _20619_);
  and _53217_ (_20626_, _20619_, _19796_);
  or _53218_ (_20627_, _20626_, _20625_);
  and _53219_ (_20628_, _20627_, _20618_);
  and _53220_ (_20629_, _20617_, _19393_);
  or _53221_ (_20630_, _20629_, _20628_);
  and _53222_ (_20631_, _20630_, _20616_);
  and _53223_ (_20632_, _20615_, _19252_);
  or _53224_ (_28206_[0], _20632_, _20631_);
  not _53225_ (_20633_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _53226_ (_20634_, _20621_, _20633_);
  and _53227_ (_20635_, _19286_, _19233_);
  nor _53228_ (_20636_, _20635_, _20634_);
  nor _53229_ (_20637_, _20636_, _20619_);
  and _53230_ (_20638_, _20619_, _19282_);
  or _53231_ (_20639_, _20638_, _20637_);
  or _53232_ (_20640_, _20639_, _20617_);
  or _53233_ (_20641_, _20618_, _19405_);
  and _53234_ (_20642_, _20641_, _20616_);
  and _53235_ (_20643_, _20642_, _20640_);
  and _53236_ (_20644_, _20615_, _19279_);
  or _53237_ (_28206_[1], _20644_, _20643_);
  not _53238_ (_20645_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _53239_ (_20646_, _20621_, _20645_);
  and _53240_ (_20647_, _20621_, _19299_);
  or _53241_ (_20648_, _20647_, _20646_);
  or _53242_ (_20649_, _20648_, _20619_);
  not _53243_ (_20650_, _20619_);
  or _53244_ (_20651_, _20650_, _19823_);
  and _53245_ (_20652_, _20651_, _20649_);
  or _53246_ (_20653_, _20652_, _20617_);
  or _53247_ (_20654_, _20618_, _19417_);
  and _53248_ (_20655_, _20654_, _20616_);
  and _53249_ (_20656_, _20655_, _20653_);
  and _53250_ (_20657_, _20615_, _19294_);
  or _53251_ (_28206_[2], _20657_, _20656_);
  and _53252_ (_20658_, _20621_, word_in[3]);
  not _53253_ (_20659_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _53254_ (_20660_, _20621_, _20659_);
  nor _53255_ (_20661_, _20660_, _20658_);
  nor _53256_ (_20662_, _20661_, _20619_);
  and _53257_ (_20663_, _20619_, _19836_);
  or _53258_ (_20664_, _20663_, _20662_);
  and _53259_ (_20665_, _20664_, _20618_);
  and _53260_ (_20666_, _20617_, _19429_);
  or _53261_ (_20667_, _20666_, _20615_);
  or _53262_ (_20668_, _20667_, _20665_);
  or _53263_ (_20669_, _20616_, _19308_);
  and _53264_ (_28206_[3], _20669_, _20668_);
  not _53265_ (_20670_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _53266_ (_20671_, _20621_, _20670_);
  and _53267_ (_20672_, _19327_, _19233_);
  nor _53268_ (_20673_, _20672_, _20671_);
  nor _53269_ (_20674_, _20673_, _20619_);
  and _53270_ (_20675_, _20619_, _19849_);
  or _53271_ (_20676_, _20675_, _20674_);
  and _53272_ (_20677_, _20676_, _20618_);
  and _53273_ (_20678_, _20617_, _19441_);
  or _53274_ (_20679_, _20678_, _20677_);
  and _53275_ (_20680_, _20679_, _20616_);
  and _53276_ (_20681_, _20615_, _19322_);
  or _53277_ (_28206_[4], _20681_, _20680_);
  not _53278_ (_20682_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _53279_ (_20683_, _20621_, _20682_);
  and _53280_ (_20684_, _20621_, _19339_);
  or _53281_ (_20685_, _20684_, _20683_);
  or _53282_ (_20686_, _20685_, _20619_);
  or _53283_ (_20687_, _20650_, _19864_);
  and _53284_ (_20688_, _20687_, _20686_);
  or _53285_ (_20689_, _20688_, _20617_);
  or _53286_ (_20690_, _20618_, _19453_);
  and _53287_ (_20691_, _20690_, _20616_);
  and _53288_ (_20692_, _20691_, _20689_);
  and _53289_ (_20693_, _20615_, _19348_);
  or _53290_ (_28206_[5], _20693_, _20692_);
  not _53291_ (_20694_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _53292_ (_20695_, _20621_, _20694_);
  and _53293_ (_20696_, _20621_, _19355_);
  or _53294_ (_20697_, _20696_, _20695_);
  or _53295_ (_20698_, _20697_, _20619_);
  or _53296_ (_20699_, _20650_, _19876_);
  and _53297_ (_20700_, _20699_, _20698_);
  or _53298_ (_20701_, _20700_, _20617_);
  or _53299_ (_20702_, _20618_, _19465_);
  and _53300_ (_20703_, _20702_, _20701_);
  or _53301_ (_20704_, _20703_, _20615_);
  or _53302_ (_20705_, _20616_, _19350_);
  and _53303_ (_28206_[6], _20705_, _20704_);
  nor _53304_ (_20706_, _20621_, _18711_);
  and _53305_ (_20707_, _20621_, _19068_);
  or _53306_ (_20708_, _20707_, _20706_);
  or _53307_ (_20709_, _20708_, _20619_);
  or _53308_ (_20710_, _20650_, _19074_);
  and _53309_ (_20711_, _20710_, _20709_);
  or _53310_ (_20712_, _20711_, _20617_);
  or _53311_ (_20713_, _20618_, _19477_);
  and _53312_ (_20714_, _20713_, _20616_);
  and _53313_ (_20715_, _20714_, _20712_);
  and _53314_ (_20716_, _20615_, _19081_);
  or _53315_ (_28206_[7], _20716_, _20715_);
  and _53316_ (_20717_, _19486_, _19058_);
  and _53317_ (_20718_, _19064_, _18690_);
  not _53318_ (_20719_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _53319_ (_20720_, _19067_, _19087_);
  nor _53320_ (_20721_, _20720_, _20719_);
  and _53321_ (_20722_, _20720_, _19266_);
  nor _53322_ (_20723_, _20722_, _20721_);
  nor _53323_ (_20724_, _20723_, _20718_);
  and _53324_ (_20725_, _20718_, _19796_);
  nor _53325_ (_20726_, _20725_, _20724_);
  nor _53326_ (_20727_, _20726_, _20717_);
  and _53327_ (_20728_, _19052_, _18667_);
  and _53328_ (_20729_, _20717_, _19393_);
  or _53329_ (_20730_, _20729_, _20728_);
  or _53330_ (_20731_, _20730_, _20727_);
  not _53331_ (_20732_, _20728_);
  or _53332_ (_20733_, _20732_, _19252_);
  and _53333_ (_28207_[0], _20733_, _20731_);
  not _53334_ (_20734_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _53335_ (_20735_, _20720_, _20734_);
  and _53336_ (_20736_, _20720_, _19286_);
  or _53337_ (_20737_, _20736_, _20735_);
  or _53338_ (_20738_, _20737_, _20718_);
  not _53339_ (_20739_, _20718_);
  or _53340_ (_20740_, _20739_, _19282_);
  and _53341_ (_20741_, _20740_, _20738_);
  or _53342_ (_20742_, _20741_, _20717_);
  not _53343_ (_20743_, _20717_);
  or _53344_ (_20744_, _20743_, _19405_);
  and _53345_ (_20745_, _20744_, _20732_);
  and _53346_ (_20746_, _20745_, _20742_);
  and _53347_ (_20747_, _20728_, _19279_);
  or _53348_ (_28207_[1], _20747_, _20746_);
  not _53349_ (_20748_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _53350_ (_20749_, _20720_, _20748_);
  and _53351_ (_20750_, _20720_, _19299_);
  or _53352_ (_20751_, _20750_, _20749_);
  or _53353_ (_20752_, _20751_, _20718_);
  or _53354_ (_20753_, _20739_, _19823_);
  and _53355_ (_20754_, _20753_, _20752_);
  or _53356_ (_20755_, _20754_, _20717_);
  or _53357_ (_20756_, _20743_, _19417_);
  and _53358_ (_20757_, _20756_, _20755_);
  or _53359_ (_20758_, _20757_, _20728_);
  or _53360_ (_20759_, _20732_, _19294_);
  and _53361_ (_28207_[2], _20759_, _20758_);
  not _53362_ (_20760_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _53363_ (_20761_, _20720_, _20760_);
  and _53364_ (_20762_, _20720_, _19313_);
  or _53365_ (_20763_, _20762_, _20761_);
  or _53366_ (_20764_, _20763_, _20718_);
  or _53367_ (_20765_, _20739_, _19836_);
  and _53368_ (_20766_, _20765_, _20764_);
  or _53369_ (_20767_, _20766_, _20717_);
  or _53370_ (_20768_, _20743_, _19429_);
  and _53371_ (_20769_, _20768_, _20767_);
  or _53372_ (_20770_, _20769_, _20728_);
  or _53373_ (_20771_, _20732_, _19308_);
  and _53374_ (_28207_[3], _20771_, _20770_);
  not _53375_ (_20772_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _53376_ (_20773_, _20720_, _20772_);
  and _53377_ (_20774_, _20720_, _19327_);
  or _53378_ (_20775_, _20774_, _20773_);
  or _53379_ (_20776_, _20775_, _20718_);
  or _53380_ (_20777_, _20739_, _19849_);
  and _53381_ (_20778_, _20777_, _20776_);
  or _53382_ (_20779_, _20778_, _20717_);
  or _53383_ (_20780_, _20743_, _19441_);
  and _53384_ (_20781_, _20780_, _20779_);
  or _53385_ (_20782_, _20781_, _20728_);
  or _53386_ (_20783_, _20732_, _19322_);
  and _53387_ (_28207_[4], _20783_, _20782_);
  and _53388_ (_20784_, _20720_, word_in[5]);
  not _53389_ (_20785_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _53390_ (_20786_, _20720_, _20785_);
  nor _53391_ (_20787_, _20786_, _20784_);
  nor _53392_ (_20788_, _20787_, _20718_);
  and _53393_ (_20789_, _20718_, _19864_);
  or _53394_ (_20790_, _20789_, _20788_);
  or _53395_ (_20791_, _20790_, _20717_);
  or _53396_ (_20792_, _20743_, _19453_);
  and _53397_ (_20793_, _20792_, _20732_);
  and _53398_ (_20794_, _20793_, _20791_);
  and _53399_ (_20795_, _20728_, _19348_);
  or _53400_ (_28207_[5], _20795_, _20794_);
  not _53401_ (_20796_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _53402_ (_20797_, _20720_, _20796_);
  and _53403_ (_20798_, _20720_, _19355_);
  or _53404_ (_20799_, _20798_, _20797_);
  or _53405_ (_20800_, _20799_, _20718_);
  or _53406_ (_20801_, _20739_, _19876_);
  and _53407_ (_20802_, _20801_, _20800_);
  or _53408_ (_20803_, _20802_, _20717_);
  or _53409_ (_20804_, _20743_, _19465_);
  and _53410_ (_20805_, _20804_, _20803_);
  or _53411_ (_20806_, _20805_, _20728_);
  or _53412_ (_20807_, _20732_, _19350_);
  and _53413_ (_28207_[6], _20807_, _20806_);
  nor _53414_ (_20808_, _20720_, _18853_);
  and _53415_ (_20809_, _20720_, _19068_);
  or _53416_ (_20810_, _20809_, _20808_);
  or _53417_ (_20811_, _20810_, _20718_);
  or _53418_ (_20812_, _20739_, _19074_);
  and _53419_ (_20813_, _20812_, _20811_);
  or _53420_ (_20814_, _20813_, _20717_);
  or _53421_ (_20815_, _20743_, _19477_);
  and _53422_ (_20816_, _20815_, _20732_);
  and _53423_ (_20817_, _20816_, _20814_);
  and _53424_ (_20818_, _20728_, _19081_);
  or _53425_ (_28207_[7], _20818_, _20817_);
  and _53426_ (_20819_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _53427_ (_20820_, _19266_, _19066_);
  nor _53428_ (_20821_, _20820_, _20819_);
  nor _53429_ (_20822_, _20821_, _19065_);
  and _53430_ (_20823_, _19796_, _19065_);
  or _53431_ (_20824_, _20823_, _20822_);
  and _53432_ (_20825_, _20824_, _19061_);
  and _53433_ (_20826_, _19060_, word_in[16]);
  or _53434_ (_20827_, _20826_, _20825_);
  and _53435_ (_20828_, _20827_, _19054_);
  and _53436_ (_20829_, _19252_, _19053_);
  or _53437_ (_28208_[0], _20829_, _20828_);
  and _53438_ (_20830_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _53439_ (_20831_, _19286_, _19066_);
  nor _53440_ (_20832_, _20831_, _20830_);
  nor _53441_ (_20833_, _20832_, _19065_);
  and _53442_ (_20834_, _19282_, _19065_);
  or _53443_ (_20835_, _20834_, _20833_);
  and _53444_ (_20836_, _20835_, _19061_);
  and _53445_ (_20837_, _19060_, word_in[17]);
  or _53446_ (_20838_, _20837_, _20836_);
  and _53447_ (_20839_, _20838_, _19054_);
  and _53448_ (_20840_, _19279_, _19053_);
  or _53449_ (_28208_[1], _20840_, _20839_);
  and _53450_ (_20841_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _53451_ (_20842_, _19299_, _19066_);
  nor _53452_ (_20843_, _20842_, _20841_);
  nor _53453_ (_20844_, _20843_, _19065_);
  and _53454_ (_20845_, _19823_, _19065_);
  or _53455_ (_20846_, _20845_, _20844_);
  and _53456_ (_20847_, _20846_, _19061_);
  and _53457_ (_20848_, _19060_, word_in[18]);
  or _53458_ (_20849_, _20848_, _20847_);
  and _53459_ (_20850_, _20849_, _19054_);
  and _53460_ (_20851_, _19294_, _19053_);
  or _53461_ (_28208_[2], _20851_, _20850_);
  and _53462_ (_20852_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _53463_ (_20853_, _19313_, _19066_);
  nor _53464_ (_20854_, _20853_, _20852_);
  nor _53465_ (_20855_, _20854_, _19065_);
  and _53466_ (_20856_, _19836_, _19065_);
  or _53467_ (_20857_, _20856_, _20855_);
  and _53468_ (_20858_, _20857_, _19061_);
  and _53469_ (_20859_, _19060_, word_in[19]);
  or _53470_ (_20860_, _20859_, _20858_);
  and _53471_ (_20861_, _20860_, _19054_);
  and _53472_ (_20862_, _19308_, _19053_);
  or _53473_ (_28208_[3], _20862_, _20861_);
  and _53474_ (_20863_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _53475_ (_20864_, _19327_, _19066_);
  nor _53476_ (_20865_, _20864_, _20863_);
  nor _53477_ (_20866_, _20865_, _19065_);
  and _53478_ (_20867_, _19849_, _19065_);
  or _53479_ (_20868_, _20867_, _20866_);
  and _53480_ (_20869_, _20868_, _19061_);
  and _53481_ (_20870_, _19060_, word_in[20]);
  or _53482_ (_20871_, _20870_, _20869_);
  and _53483_ (_20872_, _20871_, _19054_);
  and _53484_ (_20873_, _19322_, _19053_);
  or _53485_ (_28208_[4], _20873_, _20872_);
  and _53486_ (_20874_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _53487_ (_20875_, _19339_, _19066_);
  nor _53488_ (_20876_, _20875_, _20874_);
  nor _53489_ (_20877_, _20876_, _19065_);
  and _53490_ (_20878_, _19864_, _19065_);
  or _53491_ (_20879_, _20878_, _20877_);
  and _53492_ (_20880_, _20879_, _19061_);
  and _53493_ (_20881_, _19060_, word_in[21]);
  or _53494_ (_20882_, _20881_, _20880_);
  and _53495_ (_20883_, _20882_, _19054_);
  and _53496_ (_20884_, _19348_, _19053_);
  or _53497_ (_28208_[5], _20884_, _20883_);
  and _53498_ (_20885_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _53499_ (_20886_, _19355_, _19066_);
  nor _53500_ (_20887_, _20886_, _20885_);
  nor _53501_ (_20888_, _20887_, _19065_);
  and _53502_ (_20889_, _19876_, _19065_);
  or _53503_ (_20890_, _20889_, _20888_);
  and _53504_ (_20891_, _20890_, _19061_);
  and _53505_ (_20892_, _19060_, word_in[22]);
  or _53506_ (_20893_, _20892_, _20891_);
  and _53507_ (_20894_, _20893_, _19054_);
  and _53508_ (_20895_, _19350_, _19053_);
  or _53509_ (_28208_[6], _20895_, _20894_);
  and _53510_ (_20896_, _18694_, word_in[0]);
  nand _53511_ (_20897_, _18653_, _20412_);
  or _53512_ (_20898_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _53513_ (_20899_, _20898_, _20897_);
  and _53514_ (_20900_, _20899_, _18873_);
  nand _53515_ (_20901_, _18653_, _20620_);
  or _53516_ (_20902_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _53517_ (_20903_, _20902_, _20901_);
  and _53518_ (_20904_, _20903_, _18710_);
  nor _53519_ (_20905_, _18656_, _18635_);
  nand _53520_ (_20906_, _18653_, _20209_);
  or _53521_ (_20907_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _53522_ (_20908_, _20907_, _20906_);
  and _53523_ (_20909_, _20908_, _20905_);
  or _53524_ (_20910_, _20909_, _20904_);
  or _53525_ (_20911_, _20910_, _20900_);
  and _53526_ (_20912_, _20911_, _18639_);
  nand _53527_ (_20913_, _18653_, _19790_);
  or _53528_ (_20914_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _53529_ (_20915_, _20914_, _20913_);
  and _53530_ (_20916_, _20915_, _18710_);
  not _53531_ (_20917_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _53532_ (_20918_, _18653_, _20917_);
  or _53533_ (_20919_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _53534_ (_20920_, _20919_, _20918_);
  and _53535_ (_20921_, _20920_, _20905_);
  or _53536_ (_20922_, _20921_, _20916_);
  nand _53537_ (_20923_, _18653_, _20002_);
  or _53538_ (_20924_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _53539_ (_20925_, _20924_, _20923_);
  and _53540_ (_20926_, _20925_, _18700_);
  not _53541_ (_20927_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _53542_ (_20928_, _18653_, _20927_);
  or _53543_ (_20929_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _53544_ (_20930_, _20929_, _20928_);
  and _53545_ (_20931_, _20930_, _18873_);
  or _53546_ (_20932_, _20931_, _20926_);
  or _53547_ (_20933_, _20932_, _20922_);
  and _53548_ (_20934_, _20933_, _18699_);
  not _53549_ (_20935_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand _53550_ (_20936_, _18653_, _20935_);
  or _53551_ (_20937_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _53552_ (_20938_, _20937_, _20936_);
  and _53553_ (_20939_, _20938_, _18707_);
  or _53554_ (_20940_, _20939_, _20934_);
  nor _53555_ (_20941_, _20940_, _20912_);
  nor _53556_ (_20942_, _20941_, _18694_);
  or _53557_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _20942_, _20896_);
  and _53558_ (_20943_, _18694_, word_in[1]);
  nand _53559_ (_20944_, _18653_, _20223_);
  or _53560_ (_20945_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _53561_ (_20946_, _20945_, _20944_);
  and _53562_ (_20947_, _20946_, _20905_);
  nand _53563_ (_20948_, _18653_, _20429_);
  or _53564_ (_20949_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _53565_ (_20950_, _20949_, _20948_);
  and _53566_ (_20951_, _20950_, _18873_);
  or _53567_ (_20952_, _20951_, _20947_);
  nand _53568_ (_20953_, _18653_, _20633_);
  or _53569_ (_20954_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _53570_ (_20955_, _20954_, _20953_);
  and _53571_ (_20956_, _20955_, _18710_);
  or _53572_ (_20957_, _20956_, _20952_);
  and _53573_ (_20958_, _20957_, _18639_);
  nand _53574_ (_20959_, _18653_, _19806_);
  or _53575_ (_20960_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _53576_ (_20961_, _20960_, _20959_);
  and _53577_ (_20962_, _20961_, _18710_);
  not _53578_ (_20963_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand _53579_ (_20964_, _18653_, _20963_);
  or _53580_ (_20965_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _53581_ (_20966_, _20965_, _20964_);
  and _53582_ (_20967_, _20966_, _18873_);
  or _53583_ (_20968_, _20967_, _20962_);
  nand _53584_ (_20969_, _18653_, _20016_);
  or _53585_ (_20970_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _53586_ (_20971_, _20970_, _20969_);
  and _53587_ (_20972_, _20971_, _18700_);
  not _53588_ (_20973_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand _53589_ (_20974_, _18653_, _20973_);
  or _53590_ (_20975_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _53591_ (_20976_, _20975_, _20974_);
  and _53592_ (_20977_, _20976_, _20905_);
  or _53593_ (_20978_, _20977_, _20972_);
  or _53594_ (_20979_, _20978_, _20968_);
  and _53595_ (_20980_, _20979_, _18699_);
  not _53596_ (_20981_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nand _53597_ (_20982_, _18653_, _20981_);
  or _53598_ (_20983_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _53599_ (_20984_, _20983_, _20982_);
  and _53600_ (_20985_, _20984_, _18707_);
  or _53601_ (_20986_, _20985_, _20980_);
  nor _53602_ (_20987_, _20986_, _20958_);
  nor _53603_ (_20988_, _20987_, _18694_);
  or _53604_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _20988_, _20943_);
  and _53605_ (_20989_, _18694_, word_in[2]);
  nand _53606_ (_20990_, _18653_, _20442_);
  or _53607_ (_20991_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _53608_ (_20992_, _20991_, _20990_);
  and _53609_ (_20993_, _20992_, _18873_);
  nand _53610_ (_20994_, _18653_, _20645_);
  or _53611_ (_20995_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _53612_ (_20996_, _20995_, _20994_);
  and _53613_ (_20997_, _20996_, _18710_);
  nand _53614_ (_20998_, _18653_, _20237_);
  or _53615_ (_20999_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _53616_ (_21000_, _20999_, _20998_);
  and _53617_ (_21001_, _21000_, _20905_);
  or _53618_ (_21002_, _21001_, _20997_);
  or _53619_ (_21003_, _21002_, _20993_);
  and _53620_ (_21004_, _21003_, _18639_);
  nand _53621_ (_21005_, _18653_, _19818_);
  or _53622_ (_21006_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _53623_ (_21007_, _21006_, _21005_);
  and _53624_ (_21008_, _21007_, _18710_);
  not _53625_ (_21009_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _53626_ (_21010_, _18653_, _21009_);
  or _53627_ (_21011_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _53628_ (_21012_, _21011_, _21010_);
  and _53629_ (_21013_, _21012_, _20905_);
  or _53630_ (_21014_, _21013_, _21008_);
  nand _53631_ (_21015_, _18653_, _20030_);
  or _53632_ (_21016_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _53633_ (_21017_, _21016_, _21015_);
  and _53634_ (_21018_, _21017_, _18700_);
  not _53635_ (_21019_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _53636_ (_21020_, _18653_, _21019_);
  or _53637_ (_21021_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _53638_ (_21022_, _21021_, _21020_);
  and _53639_ (_21023_, _21022_, _18873_);
  or _53640_ (_21024_, _21023_, _21018_);
  or _53641_ (_21025_, _21024_, _21014_);
  and _53642_ (_21026_, _21025_, _18699_);
  not _53643_ (_21027_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nand _53644_ (_21028_, _18653_, _21027_);
  or _53645_ (_21029_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _53646_ (_21030_, _21029_, _21028_);
  and _53647_ (_21031_, _21030_, _18707_);
  or _53648_ (_21032_, _21031_, _21026_);
  nor _53649_ (_21033_, _21032_, _21004_);
  nor _53650_ (_21034_, _21033_, _18694_);
  or _53651_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _21034_, _20989_);
  and _53652_ (_21035_, _18694_, word_in[3]);
  nand _53653_ (_21036_, _18653_, _19831_);
  or _53654_ (_21037_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _53655_ (_21038_, _21037_, _21036_);
  and _53656_ (_21039_, _21038_, _18710_);
  not _53657_ (_21040_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand _53658_ (_21041_, _18653_, _21040_);
  or _53659_ (_21042_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _53660_ (_21043_, _21042_, _21041_);
  and _53661_ (_21044_, _21043_, _18873_);
  or _53662_ (_21045_, _21044_, _21039_);
  nand _53663_ (_21046_, _18653_, _20042_);
  or _53664_ (_21047_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _53665_ (_21048_, _21047_, _21046_);
  and _53666_ (_21049_, _21048_, _18700_);
  not _53667_ (_21050_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nand _53668_ (_21051_, _18653_, _21050_);
  or _53669_ (_21052_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _53670_ (_21053_, _21052_, _21051_);
  and _53671_ (_21054_, _21053_, _20905_);
  or _53672_ (_21055_, _21054_, _21049_);
  or _53673_ (_21056_, _21055_, _21045_);
  and _53674_ (_21057_, _21056_, _18699_);
  nand _53675_ (_21058_, _18653_, _20249_);
  or _53676_ (_21059_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _53677_ (_21060_, _21059_, _21058_);
  and _53678_ (_21061_, _21060_, _20905_);
  nand _53679_ (_21062_, _18653_, _20453_);
  or _53680_ (_21063_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _53681_ (_21064_, _21063_, _21062_);
  and _53682_ (_21065_, _21064_, _18873_);
  or _53683_ (_21066_, _21065_, _21061_);
  nand _53684_ (_21067_, _18653_, _20659_);
  or _53685_ (_21068_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _53686_ (_21069_, _21068_, _21067_);
  and _53687_ (_21070_, _21069_, _18710_);
  or _53688_ (_21071_, _21070_, _21066_);
  and _53689_ (_21072_, _21071_, _18639_);
  not _53690_ (_21073_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nand _53691_ (_21074_, _18653_, _21073_);
  or _53692_ (_21075_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _53693_ (_21076_, _21075_, _21074_);
  and _53694_ (_21077_, _21076_, _18707_);
  or _53695_ (_21078_, _21077_, _21072_);
  nor _53696_ (_21079_, _21078_, _21057_);
  nor _53697_ (_21080_, _21079_, _18694_);
  or _53698_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _21080_, _21035_);
  and _53699_ (_21081_, _18694_, word_in[4]);
  nand _53700_ (_21082_, _18653_, _19844_);
  or _53701_ (_21083_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _53702_ (_21084_, _21083_, _21082_);
  and _53703_ (_21085_, _21084_, _18710_);
  not _53704_ (_21086_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand _53705_ (_21087_, _18653_, _21086_);
  or _53706_ (_21088_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _53707_ (_21089_, _21088_, _21087_);
  and _53708_ (_21090_, _21089_, _20905_);
  or _53709_ (_21091_, _21090_, _21085_);
  nand _53710_ (_21092_, _18653_, _20053_);
  or _53711_ (_21093_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _53712_ (_21094_, _21093_, _21092_);
  and _53713_ (_21095_, _21094_, _18700_);
  not _53714_ (_21096_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand _53715_ (_21097_, _18653_, _21096_);
  or _53716_ (_21098_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _53717_ (_21099_, _21098_, _21097_);
  and _53718_ (_21100_, _21099_, _18873_);
  or _53719_ (_21101_, _21100_, _21095_);
  or _53720_ (_21102_, _21101_, _21091_);
  and _53721_ (_21103_, _21102_, _18699_);
  nand _53722_ (_21104_, _18653_, _20465_);
  or _53723_ (_21105_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _53724_ (_21106_, _21105_, _21104_);
  and _53725_ (_21107_, _21106_, _18873_);
  nand _53726_ (_21108_, _18653_, _20670_);
  or _53727_ (_21109_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _53728_ (_21110_, _21109_, _21108_);
  and _53729_ (_21111_, _21110_, _18710_);
  nand _53730_ (_21112_, _18653_, _20261_);
  or _53731_ (_21113_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _53732_ (_21114_, _21113_, _21112_);
  and _53733_ (_21115_, _21114_, _20905_);
  or _53734_ (_21116_, _21115_, _21111_);
  or _53735_ (_21117_, _21116_, _21107_);
  and _53736_ (_21118_, _21117_, _18639_);
  not _53737_ (_21119_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand _53738_ (_21120_, _18653_, _21119_);
  or _53739_ (_21121_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _53740_ (_21122_, _21121_, _21120_);
  and _53741_ (_21123_, _21122_, _18707_);
  or _53742_ (_21124_, _21123_, _21118_);
  nor _53743_ (_21125_, _21124_, _21103_);
  nor _53744_ (_21126_, _21125_, _18694_);
  or _53745_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _21126_, _21081_);
  and _53746_ (_21127_, _18694_, word_in[5]);
  nand _53747_ (_21128_, _18653_, _20477_);
  or _53748_ (_21129_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _53749_ (_21130_, _21129_, _21128_);
  and _53750_ (_21131_, _21130_, _18873_);
  nand _53751_ (_21132_, _18653_, _20682_);
  or _53752_ (_21133_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _53753_ (_21134_, _21133_, _21132_);
  and _53754_ (_21135_, _21134_, _18710_);
  nand _53755_ (_21136_, _18653_, _20273_);
  or _53756_ (_21137_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _53757_ (_21138_, _21137_, _21136_);
  and _53758_ (_21139_, _21138_, _20905_);
  or _53759_ (_21140_, _21139_, _21135_);
  or _53760_ (_21141_, _21140_, _21131_);
  and _53761_ (_21142_, _21141_, _18639_);
  nand _53762_ (_21143_, _18653_, _19859_);
  or _53763_ (_21144_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _53764_ (_21145_, _21144_, _21143_);
  and _53765_ (_21146_, _21145_, _18710_);
  not _53766_ (_21147_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nand _53767_ (_21148_, _18653_, _21147_);
  or _53768_ (_21149_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _53769_ (_21150_, _21149_, _21148_);
  and _53770_ (_21151_, _21150_, _20905_);
  or _53771_ (_21152_, _21151_, _21146_);
  nand _53772_ (_21153_, _18653_, _20066_);
  or _53773_ (_21154_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _53774_ (_21155_, _21154_, _21153_);
  and _53775_ (_21156_, _21155_, _18700_);
  not _53776_ (_21157_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand _53777_ (_21158_, _18653_, _21157_);
  or _53778_ (_21159_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _53779_ (_21160_, _21159_, _21158_);
  and _53780_ (_21161_, _21160_, _18873_);
  or _53781_ (_21162_, _21161_, _21156_);
  or _53782_ (_21163_, _21162_, _21152_);
  and _53783_ (_21164_, _21163_, _18699_);
  not _53784_ (_21165_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand _53785_ (_21166_, _18653_, _21165_);
  or _53786_ (_21167_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _53787_ (_21168_, _21167_, _21166_);
  and _53788_ (_21169_, _21168_, _18707_);
  or _53789_ (_21170_, _21169_, _21164_);
  nor _53790_ (_21171_, _21170_, _21142_);
  nor _53791_ (_21172_, _21171_, _18694_);
  or _53792_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _21172_, _21127_);
  and _53793_ (_21173_, _18694_, word_in[6]);
  nand _53794_ (_21174_, _18653_, _20490_);
  or _53795_ (_21175_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _53796_ (_21176_, _21175_, _21174_);
  and _53797_ (_21177_, _21176_, _18873_);
  nand _53798_ (_21178_, _18653_, _20694_);
  or _53799_ (_21179_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _53800_ (_21180_, _21179_, _21178_);
  and _53801_ (_21181_, _21180_, _18710_);
  nand _53802_ (_21182_, _18653_, _20286_);
  or _53803_ (_21183_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _53804_ (_21184_, _21183_, _21182_);
  and _53805_ (_21185_, _21184_, _20905_);
  or _53806_ (_21186_, _21185_, _21181_);
  or _53807_ (_21187_, _21186_, _21177_);
  and _53808_ (_21188_, _21187_, _18639_);
  nand _53809_ (_21189_, _18653_, _19871_);
  or _53810_ (_21190_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _53811_ (_21191_, _21190_, _21189_);
  and _53812_ (_21192_, _21191_, _18710_);
  not _53813_ (_21193_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nand _53814_ (_21194_, _18653_, _21193_);
  or _53815_ (_21195_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _53816_ (_21196_, _21195_, _21194_);
  and _53817_ (_21197_, _21196_, _18873_);
  or _53818_ (_21198_, _21197_, _21192_);
  nand _53819_ (_21199_, _18653_, _20076_);
  or _53820_ (_21200_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _53821_ (_21201_, _21200_, _21199_);
  and _53822_ (_21202_, _21201_, _18700_);
  not _53823_ (_21203_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nand _53824_ (_21204_, _18653_, _21203_);
  or _53825_ (_21205_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _53826_ (_21206_, _21205_, _21204_);
  and _53827_ (_21207_, _21206_, _20905_);
  or _53828_ (_21208_, _21207_, _21202_);
  or _53829_ (_21209_, _21208_, _21198_);
  and _53830_ (_21210_, _21209_, _18699_);
  not _53831_ (_21211_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nand _53832_ (_21212_, _18653_, _21211_);
  or _53833_ (_21213_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _53834_ (_21214_, _21213_, _21212_);
  and _53835_ (_21215_, _21214_, _18707_);
  or _53836_ (_21216_, _21215_, _21210_);
  nor _53837_ (_21217_, _21216_, _21188_);
  nor _53838_ (_21218_, _21217_, _18694_);
  or _53839_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _21218_, _21173_);
  and _53840_ (_21219_, _18808_, word_in[8]);
  nand _53841_ (_21220_, _18653_, _19268_);
  or _53842_ (_21221_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _53843_ (_21222_, _21221_, _21220_);
  and _53844_ (_21223_, _21222_, _18809_);
  and _53845_ (_21224_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _53846_ (_21225_, _18653_, _20927_);
  or _53847_ (_21226_, _21225_, _21224_);
  and _53848_ (_21227_, _21226_, _18815_);
  nor _53849_ (_21228_, _21227_, _21223_);
  nor _53850_ (_21229_, _21228_, _18758_);
  nand _53851_ (_21230_, _18653_, _19688_);
  or _53852_ (_21231_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _53853_ (_21232_, _21231_, _21230_);
  and _53854_ (_21233_, _21232_, _18809_);
  nand _53855_ (_21234_, _18653_, _19899_);
  or _53856_ (_21235_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _53857_ (_21236_, _21235_, _21234_);
  and _53858_ (_21237_, _21236_, _18815_);
  or _53859_ (_21238_, _21237_, _21233_);
  and _53860_ (_21239_, _21238_, _18758_);
  or _53861_ (_21240_, _21239_, _21229_);
  and _53862_ (_21241_, _21240_, _18756_);
  nand _53863_ (_21242_, _18653_, _20109_);
  or _53864_ (_21243_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _53865_ (_21244_, _21243_, _21242_);
  and _53866_ (_21245_, _21244_, _18809_);
  nand _53867_ (_21246_, _18653_, _20312_);
  or _53868_ (_21247_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _53869_ (_21248_, _21247_, _21246_);
  and _53870_ (_21249_, _21248_, _18815_);
  nor _53871_ (_21250_, _21249_, _21245_);
  nor _53872_ (_21251_, _21250_, _18758_);
  nand _53873_ (_21252_, _18653_, _20518_);
  or _53874_ (_21253_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _53875_ (_21254_, _21253_, _21252_);
  and _53876_ (_21255_, _21254_, _18809_);
  nand _53877_ (_21256_, _18653_, _20719_);
  or _53878_ (_21257_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _53879_ (_21258_, _21257_, _21256_);
  and _53880_ (_21259_, _21258_, _18815_);
  or _53881_ (_21260_, _21259_, _21255_);
  and _53882_ (_21261_, _21260_, _18758_);
  nor _53883_ (_21262_, _21261_, _21251_);
  nor _53884_ (_21263_, _21262_, _18756_);
  nor _53885_ (_21264_, _21263_, _21241_);
  nor _53886_ (_21265_, _21264_, _18808_);
  or _53887_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _21265_, _21219_);
  and _53888_ (_21266_, _18808_, word_in[9]);
  nand _53889_ (_21267_, _18653_, _19284_);
  or _53890_ (_21268_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _53891_ (_21269_, _21268_, _21267_);
  and _53892_ (_21270_, _21269_, _18809_);
  and _53893_ (_21271_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _53894_ (_21272_, _18653_, _20963_);
  or _53895_ (_21273_, _21272_, _21271_);
  and _53896_ (_21274_, _21273_, _18815_);
  nor _53897_ (_21275_, _21274_, _21270_);
  nor _53898_ (_21276_, _21275_, _18758_);
  nand _53899_ (_21277_, _18653_, _19701_);
  or _53900_ (_21278_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _53901_ (_21279_, _21278_, _21277_);
  and _53902_ (_21280_, _21279_, _18809_);
  nand _53903_ (_21281_, _18653_, _19913_);
  or _53904_ (_21282_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _53905_ (_21283_, _21282_, _21281_);
  and _53906_ (_21284_, _21283_, _18815_);
  or _53907_ (_21285_, _21284_, _21280_);
  and _53908_ (_21286_, _21285_, _18758_);
  or _53909_ (_21287_, _21286_, _21276_);
  and _53910_ (_21288_, _21287_, _18756_);
  nand _53911_ (_21289_, _18653_, _20120_);
  or _53912_ (_21290_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _53913_ (_21291_, _21290_, _21289_);
  and _53914_ (_21292_, _21291_, _18809_);
  nand _53915_ (_21293_, _18653_, _20325_);
  or _53916_ (_21294_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _53917_ (_21295_, _21294_, _21293_);
  and _53918_ (_21296_, _21295_, _18815_);
  nor _53919_ (_21297_, _21296_, _21292_);
  nor _53920_ (_21298_, _21297_, _18758_);
  nand _53921_ (_21299_, _18653_, _20532_);
  or _53922_ (_21300_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _53923_ (_21301_, _21300_, _21299_);
  and _53924_ (_21302_, _21301_, _18809_);
  nand _53925_ (_21303_, _18653_, _20734_);
  or _53926_ (_21304_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _53927_ (_21305_, _21304_, _21303_);
  and _53928_ (_21306_, _21305_, _18815_);
  or _53929_ (_21307_, _21306_, _21302_);
  and _53930_ (_21308_, _21307_, _18758_);
  nor _53931_ (_21309_, _21308_, _21298_);
  nor _53932_ (_21310_, _21309_, _18756_);
  nor _53933_ (_21311_, _21310_, _21288_);
  nor _53934_ (_21312_, _21311_, _18808_);
  or _53935_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _21312_, _21266_);
  and _53936_ (_21313_, _18808_, word_in[10]);
  nand _53937_ (_21314_, _18653_, _19297_);
  or _53938_ (_21315_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _53939_ (_21316_, _21315_, _21314_);
  and _53940_ (_21317_, _21316_, _18809_);
  and _53941_ (_21318_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _53942_ (_21319_, _18653_, _21019_);
  or _53943_ (_21320_, _21319_, _21318_);
  and _53944_ (_21321_, _21320_, _18815_);
  nor _53945_ (_21322_, _21321_, _21317_);
  nor _53946_ (_21323_, _21322_, _18758_);
  nand _53947_ (_21324_, _18653_, _19715_);
  or _53948_ (_21325_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _53949_ (_21326_, _21325_, _21324_);
  and _53950_ (_21327_, _21326_, _18809_);
  nand _53951_ (_21328_, _18653_, _19926_);
  or _53952_ (_21329_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _53953_ (_21330_, _21329_, _21328_);
  and _53954_ (_21331_, _21330_, _18815_);
  or _53955_ (_21332_, _21331_, _21327_);
  and _53956_ (_21333_, _21332_, _18758_);
  or _53957_ (_21334_, _21333_, _21323_);
  and _53958_ (_21335_, _21334_, _18756_);
  nand _53959_ (_21336_, _18653_, _20135_);
  or _53960_ (_21337_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _53961_ (_21338_, _21337_, _21336_);
  and _53962_ (_21339_, _21338_, _18809_);
  nand _53963_ (_21340_, _18653_, _20339_);
  or _53964_ (_21341_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _53965_ (_21342_, _21341_, _21340_);
  and _53966_ (_21343_, _21342_, _18815_);
  nor _53967_ (_21344_, _21343_, _21339_);
  nor _53968_ (_21345_, _21344_, _18758_);
  nand _53969_ (_21346_, _18653_, _20544_);
  or _53970_ (_21347_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _53971_ (_21348_, _21347_, _21346_);
  and _53972_ (_21349_, _21348_, _18809_);
  nand _53973_ (_21350_, _18653_, _20748_);
  or _53974_ (_21351_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _53975_ (_21352_, _21351_, _21350_);
  and _53976_ (_21353_, _21352_, _18815_);
  or _53977_ (_21354_, _21353_, _21349_);
  and _53978_ (_21355_, _21354_, _18758_);
  nor _53979_ (_21356_, _21355_, _21345_);
  nor _53980_ (_21357_, _21356_, _18756_);
  nor _53981_ (_21358_, _21357_, _21335_);
  nor _53982_ (_21359_, _21358_, _18808_);
  or _53983_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _21359_, _21313_);
  and _53984_ (_21360_, _18808_, word_in[11]);
  nand _53985_ (_21361_, _18653_, _19311_);
  or _53986_ (_21362_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _53987_ (_21363_, _21362_, _21361_);
  and _53988_ (_21364_, _21363_, _18809_);
  and _53989_ (_21365_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _53990_ (_21366_, _18653_, _21040_);
  or _53991_ (_21367_, _21366_, _21365_);
  and _53992_ (_21368_, _21367_, _18815_);
  nor _53993_ (_21369_, _21368_, _21364_);
  nor _53994_ (_21370_, _21369_, _18758_);
  nand _53995_ (_21371_, _18653_, _19727_);
  or _53996_ (_21372_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _53997_ (_21373_, _21372_, _21371_);
  and _53998_ (_21374_, _21373_, _18809_);
  nand _53999_ (_21375_, _18653_, _19939_);
  or _54000_ (_21376_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _54001_ (_21377_, _21376_, _21375_);
  and _54002_ (_21378_, _21377_, _18815_);
  or _54003_ (_21379_, _21378_, _21374_);
  and _54004_ (_21380_, _21379_, _18758_);
  or _54005_ (_21381_, _21380_, _21370_);
  and _54006_ (_21382_, _21381_, _18756_);
  nand _54007_ (_21383_, _18653_, _20147_);
  or _54008_ (_21384_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _54009_ (_21385_, _21384_, _21383_);
  and _54010_ (_21386_, _21385_, _18809_);
  nand _54011_ (_21387_, _18653_, _20353_);
  or _54012_ (_21388_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _54013_ (_21389_, _21388_, _21387_);
  and _54014_ (_21390_, _21389_, _18815_);
  nor _54015_ (_21391_, _21390_, _21386_);
  nor _54016_ (_21392_, _21391_, _18758_);
  nand _54017_ (_21393_, _18653_, _20557_);
  or _54018_ (_21394_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _54019_ (_21395_, _21394_, _21393_);
  and _54020_ (_21396_, _21395_, _18809_);
  nand _54021_ (_21397_, _18653_, _20760_);
  or _54022_ (_21398_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _54023_ (_21399_, _21398_, _21397_);
  and _54024_ (_21400_, _21399_, _18815_);
  or _54025_ (_21401_, _21400_, _21396_);
  and _54026_ (_21402_, _21401_, _18758_);
  nor _54027_ (_21403_, _21402_, _21392_);
  nor _54028_ (_21404_, _21403_, _18756_);
  nor _54029_ (_21405_, _21404_, _21382_);
  nor _54030_ (_21406_, _21405_, _18808_);
  or _54031_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _21406_, _21360_);
  and _54032_ (_21407_, _18808_, word_in[12]);
  nand _54033_ (_21408_, _18653_, _19325_);
  or _54034_ (_21409_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _54035_ (_21410_, _21409_, _21408_);
  and _54036_ (_21411_, _21410_, _18809_);
  and _54037_ (_21412_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _54038_ (_21413_, _18653_, _21096_);
  or _54039_ (_21414_, _21413_, _21412_);
  and _54040_ (_21415_, _21414_, _18815_);
  nor _54041_ (_21416_, _21415_, _21411_);
  nor _54042_ (_21417_, _21416_, _18758_);
  nand _54043_ (_21418_, _18653_, _19739_);
  or _54044_ (_21419_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _54045_ (_21420_, _21419_, _21418_);
  and _54046_ (_21421_, _21420_, _18809_);
  nand _54047_ (_21422_, _18653_, _19950_);
  or _54048_ (_21423_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _54049_ (_21424_, _21423_, _21422_);
  and _54050_ (_21425_, _21424_, _18815_);
  or _54051_ (_21426_, _21425_, _21421_);
  and _54052_ (_21427_, _21426_, _18758_);
  or _54053_ (_21428_, _21427_, _21417_);
  and _54054_ (_21429_, _21428_, _18756_);
  nand _54055_ (_21430_, _18653_, _20158_);
  or _54056_ (_21431_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _54057_ (_21432_, _21431_, _21430_);
  and _54058_ (_21433_, _21432_, _18809_);
  nand _54059_ (_21434_, _18653_, _20363_);
  or _54060_ (_21435_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _54061_ (_21436_, _21435_, _21434_);
  and _54062_ (_21437_, _21436_, _18815_);
  nor _54063_ (_21438_, _21437_, _21433_);
  nor _54064_ (_21439_, _21438_, _18758_);
  nand _54065_ (_21440_, _18653_, _20568_);
  or _54066_ (_21441_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _54067_ (_21442_, _21441_, _21440_);
  and _54068_ (_21443_, _21442_, _18809_);
  nand _54069_ (_21444_, _18653_, _20772_);
  or _54070_ (_21445_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _54071_ (_21446_, _21445_, _21444_);
  and _54072_ (_21447_, _21446_, _18815_);
  or _54073_ (_21448_, _21447_, _21443_);
  and _54074_ (_21449_, _21448_, _18758_);
  nor _54075_ (_21450_, _21449_, _21439_);
  nor _54076_ (_21451_, _21450_, _18756_);
  nor _54077_ (_21452_, _21451_, _21429_);
  nor _54078_ (_21453_, _21452_, _18808_);
  or _54079_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _21453_, _21407_);
  and _54080_ (_21454_, _18808_, word_in[13]);
  nand _54081_ (_21455_, _18653_, _19337_);
  or _54082_ (_21456_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _54083_ (_21457_, _21456_, _21455_);
  and _54084_ (_21458_, _21457_, _18809_);
  and _54085_ (_21459_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _54086_ (_21460_, _18653_, _21157_);
  or _54087_ (_21461_, _21460_, _21459_);
  and _54088_ (_21462_, _21461_, _18815_);
  nor _54089_ (_21463_, _21462_, _21458_);
  nor _54090_ (_21464_, _21463_, _18758_);
  nand _54091_ (_21465_, _18653_, _19751_);
  or _54092_ (_21466_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _54093_ (_21467_, _21466_, _21465_);
  and _54094_ (_21468_, _21467_, _18809_);
  nand _54095_ (_21469_, _18653_, _19962_);
  or _54096_ (_21470_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _54097_ (_21471_, _21470_, _21469_);
  and _54098_ (_21472_, _21471_, _18815_);
  or _54099_ (_21473_, _21472_, _21468_);
  and _54100_ (_21474_, _21473_, _18758_);
  or _54101_ (_21475_, _21474_, _21464_);
  and _54102_ (_21476_, _21475_, _18756_);
  nand _54103_ (_21477_, _18653_, _20170_);
  or _54104_ (_21478_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _54105_ (_21479_, _21478_, _21477_);
  and _54106_ (_21480_, _21479_, _18809_);
  nand _54107_ (_21481_, _18653_, _20375_);
  or _54108_ (_21482_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _54109_ (_21483_, _21482_, _21481_);
  and _54110_ (_21484_, _21483_, _18815_);
  nor _54111_ (_21485_, _21484_, _21480_);
  nor _54112_ (_21486_, _21485_, _18758_);
  nand _54113_ (_21487_, _18653_, _20580_);
  or _54114_ (_21488_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _54115_ (_21489_, _21488_, _21487_);
  and _54116_ (_21490_, _21489_, _18809_);
  nand _54117_ (_21491_, _18653_, _20785_);
  or _54118_ (_21492_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _54119_ (_21493_, _21492_, _21491_);
  and _54120_ (_21494_, _21493_, _18815_);
  or _54121_ (_21495_, _21494_, _21490_);
  and _54122_ (_21496_, _21495_, _18758_);
  nor _54123_ (_21497_, _21496_, _21486_);
  nor _54124_ (_21498_, _21497_, _18756_);
  nor _54125_ (_21499_, _21498_, _21476_);
  nor _54126_ (_21500_, _21499_, _18808_);
  or _54127_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _21500_, _21454_);
  and _54128_ (_21501_, _18808_, word_in[14]);
  nand _54129_ (_21502_, _18653_, _19353_);
  or _54130_ (_21503_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _54131_ (_21504_, _21503_, _21502_);
  and _54132_ (_21505_, _21504_, _18809_);
  and _54133_ (_21506_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _54134_ (_21507_, _18653_, _21193_);
  or _54135_ (_21508_, _21507_, _21506_);
  and _54136_ (_21509_, _21508_, _18815_);
  nor _54137_ (_21510_, _21509_, _21505_);
  nor _54138_ (_21511_, _21510_, _18758_);
  nand _54139_ (_21512_, _18653_, _19763_);
  or _54140_ (_21513_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _54141_ (_21514_, _21513_, _21512_);
  and _54142_ (_21515_, _21514_, _18809_);
  nand _54143_ (_21516_, _18653_, _19975_);
  or _54144_ (_21517_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _54145_ (_21518_, _21517_, _21516_);
  and _54146_ (_21519_, _21518_, _18815_);
  or _54147_ (_21520_, _21519_, _21515_);
  and _54148_ (_21521_, _21520_, _18758_);
  or _54149_ (_21522_, _21521_, _21511_);
  and _54150_ (_21523_, _21522_, _18756_);
  nand _54151_ (_21524_, _18653_, _20182_);
  or _54152_ (_21525_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _54153_ (_21526_, _21525_, _21524_);
  and _54154_ (_21527_, _21526_, _18809_);
  nand _54155_ (_21528_, _18653_, _20388_);
  or _54156_ (_21529_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _54157_ (_21530_, _21529_, _21528_);
  and _54158_ (_21531_, _21530_, _18815_);
  nor _54159_ (_21532_, _21531_, _21527_);
  nor _54160_ (_21533_, _21532_, _18758_);
  nand _54161_ (_21534_, _18653_, _20593_);
  or _54162_ (_21535_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _54163_ (_21536_, _21535_, _21534_);
  and _54164_ (_21537_, _21536_, _18809_);
  nand _54165_ (_21538_, _18653_, _20796_);
  or _54166_ (_21539_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _54167_ (_21540_, _21539_, _21538_);
  and _54168_ (_21541_, _21540_, _18815_);
  or _54169_ (_21542_, _21541_, _21537_);
  and _54170_ (_21543_, _21542_, _18758_);
  nor _54171_ (_21544_, _21543_, _21533_);
  nor _54172_ (_21545_, _21544_, _18756_);
  nor _54173_ (_21546_, _21545_, _21523_);
  nor _54174_ (_21547_, _21546_, _18808_);
  or _54175_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _21547_, _21501_);
  and _54176_ (_21548_, _18960_, word_in[16]);
  and _54177_ (_21549_, _20903_, _18873_);
  and _54178_ (_21550_, _20899_, _20905_);
  or _54179_ (_21551_, _21550_, _21549_);
  and _54180_ (_21552_, _20938_, _18710_);
  and _54181_ (_21553_, _20908_, _18700_);
  or _54182_ (_21554_, _21553_, _21552_);
  or _54183_ (_21555_, _21554_, _21551_);
  or _54184_ (_21556_, _21555_, _18868_);
  and _54185_ (_21557_, _20925_, _18710_);
  and _54186_ (_21558_, _20930_, _20905_);
  or _54187_ (_21559_, _21558_, _21557_);
  and _54188_ (_21560_, _20915_, _18873_);
  and _54189_ (_21561_, _20920_, _18700_);
  or _54190_ (_21562_, _21561_, _21560_);
  nor _54191_ (_21563_, _21562_, _21559_);
  nand _54192_ (_21564_, _21563_, _18868_);
  and _54193_ (_21565_, _21564_, _21556_);
  and _54194_ (_21566_, _21565_, _18939_);
  or _54195_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _21566_, _21548_);
  and _54196_ (_21567_, _18960_, word_in[17]);
  and _54197_ (_21568_, _20946_, _18700_);
  and _54198_ (_21569_, _20950_, _20905_);
  or _54199_ (_21570_, _21569_, _21568_);
  and _54200_ (_21571_, _20984_, _18710_);
  and _54201_ (_21572_, _20955_, _18873_);
  or _54202_ (_21573_, _21572_, _21571_);
  or _54203_ (_21574_, _21573_, _21570_);
  or _54204_ (_21575_, _21574_, _18868_);
  and _54205_ (_21576_, _20961_, _18873_);
  and _54206_ (_21577_, _20966_, _20905_);
  or _54207_ (_21578_, _21577_, _21576_);
  and _54208_ (_21579_, _20971_, _18710_);
  and _54209_ (_21580_, _20976_, _18700_);
  or _54210_ (_21581_, _21580_, _21579_);
  nor _54211_ (_21582_, _21581_, _21578_);
  nand _54212_ (_21583_, _21582_, _18868_);
  and _54213_ (_21584_, _21583_, _21575_);
  and _54214_ (_21585_, _21584_, _18939_);
  or _54215_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _21585_, _21567_);
  and _54216_ (_21586_, _18960_, word_in[18]);
  and _54217_ (_21587_, _21030_, _18710_);
  and _54218_ (_21588_, _20996_, _18873_);
  or _54219_ (_21589_, _21588_, _21587_);
  and _54220_ (_21590_, _21000_, _18700_);
  and _54221_ (_21591_, _20992_, _20905_);
  or _54222_ (_21592_, _21591_, _21590_);
  or _54223_ (_21593_, _21592_, _21589_);
  or _54224_ (_21594_, _21593_, _18868_);
  and _54225_ (_21595_, _21007_, _18873_);
  and _54226_ (_21596_, _21022_, _20905_);
  or _54227_ (_21597_, _21596_, _21595_);
  and _54228_ (_21598_, _21017_, _18710_);
  and _54229_ (_21599_, _21012_, _18700_);
  or _54230_ (_21600_, _21599_, _21598_);
  nor _54231_ (_21601_, _21600_, _21597_);
  nand _54232_ (_21602_, _21601_, _18868_);
  and _54233_ (_21603_, _21602_, _21594_);
  and _54234_ (_21604_, _21603_, _18939_);
  or _54235_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _21604_, _21586_);
  and _54236_ (_21605_, _18960_, word_in[19]);
  and _54237_ (_21606_, _21076_, _18710_);
  and _54238_ (_21607_, _21069_, _18873_);
  or _54239_ (_21608_, _21607_, _21606_);
  and _54240_ (_21609_, _21060_, _18700_);
  and _54241_ (_21610_, _21064_, _20905_);
  or _54242_ (_21611_, _21610_, _21609_);
  or _54243_ (_21612_, _21611_, _21608_);
  or _54244_ (_21613_, _21612_, _18868_);
  and _54245_ (_21614_, _21038_, _18873_);
  and _54246_ (_21615_, _21043_, _20905_);
  or _54247_ (_21616_, _21615_, _21614_);
  and _54248_ (_21617_, _21048_, _18710_);
  and _54249_ (_21618_, _21053_, _18700_);
  or _54250_ (_21619_, _21618_, _21617_);
  nor _54251_ (_21620_, _21619_, _21616_);
  nand _54252_ (_21621_, _21620_, _18868_);
  and _54253_ (_21622_, _21621_, _21613_);
  and _54254_ (_21623_, _21622_, _18939_);
  or _54255_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _21623_, _21605_);
  and _54256_ (_21624_, _18960_, word_in[20]);
  and _54257_ (_21625_, _21094_, _18710_);
  and _54258_ (_21626_, _21084_, _18873_);
  or _54259_ (_21627_, _21626_, _21625_);
  and _54260_ (_21628_, _21089_, _18700_);
  and _54261_ (_21629_, _21099_, _20905_);
  or _54262_ (_21630_, _21629_, _21628_);
  nor _54263_ (_21631_, _21630_, _21627_);
  nand _54264_ (_21632_, _21631_, _18868_);
  and _54265_ (_21633_, _21110_, _18873_);
  and _54266_ (_21634_, _21106_, _20905_);
  or _54267_ (_21635_, _21634_, _21633_);
  and _54268_ (_21636_, _21122_, _18710_);
  and _54269_ (_21637_, _21114_, _18700_);
  or _54270_ (_21638_, _21637_, _21636_);
  or _54271_ (_21639_, _21638_, _21635_);
  or _54272_ (_21640_, _21639_, _18868_);
  and _54273_ (_21641_, _21640_, _21632_);
  and _54274_ (_21642_, _21641_, _18939_);
  or _54275_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _21642_, _21624_);
  and _54276_ (_21643_, _18960_, word_in[21]);
  and _54277_ (_21644_, _21168_, _18710_);
  and _54278_ (_21645_, _21134_, _18873_);
  or _54279_ (_21646_, _21645_, _21644_);
  and _54280_ (_21647_, _21138_, _18700_);
  and _54281_ (_21648_, _21130_, _20905_);
  or _54282_ (_21649_, _21648_, _21647_);
  or _54283_ (_21650_, _21649_, _21646_);
  or _54284_ (_21651_, _21650_, _18868_);
  and _54285_ (_21652_, _21155_, _18710_);
  and _54286_ (_21653_, _21145_, _18873_);
  or _54287_ (_21654_, _21653_, _21652_);
  and _54288_ (_21655_, _21150_, _18700_);
  and _54289_ (_21656_, _21160_, _20905_);
  or _54290_ (_21657_, _21656_, _21655_);
  nor _54291_ (_21658_, _21657_, _21654_);
  nand _54292_ (_21659_, _21658_, _18868_);
  and _54293_ (_21660_, _21659_, _21651_);
  and _54294_ (_21661_, _21660_, _18939_);
  or _54295_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _21661_, _21643_);
  and _54296_ (_21662_, _18960_, word_in[22]);
  and _54297_ (_21663_, _21180_, _18873_);
  and _54298_ (_21664_, _21176_, _20905_);
  or _54299_ (_21665_, _21664_, _21663_);
  and _54300_ (_21666_, _21214_, _18710_);
  and _54301_ (_21667_, _21184_, _18700_);
  or _54302_ (_21668_, _21667_, _21666_);
  or _54303_ (_21669_, _21668_, _21665_);
  or _54304_ (_21670_, _21669_, _18868_);
  and _54305_ (_21671_, _21191_, _18873_);
  and _54306_ (_21672_, _21196_, _20905_);
  or _54307_ (_21673_, _21672_, _21671_);
  and _54308_ (_21674_, _21201_, _18710_);
  and _54309_ (_21675_, _21206_, _18700_);
  or _54310_ (_21676_, _21675_, _21674_);
  nor _54311_ (_21677_, _21676_, _21673_);
  nand _54312_ (_21678_, _21677_, _18868_);
  and _54313_ (_21679_, _21678_, _21670_);
  and _54314_ (_21680_, _21679_, _18939_);
  or _54315_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _21680_, _21662_);
  and _54316_ (_21681_, _19024_, word_in[24]);
  and _54317_ (_21682_, _21226_, _18809_);
  and _54318_ (_21683_, _21222_, _18815_);
  or _54319_ (_21684_, _21683_, _21682_);
  or _54320_ (_21685_, _21684_, _18964_);
  and _54321_ (_21686_, _21236_, _18809_);
  and _54322_ (_21687_, _21232_, _18815_);
  nor _54323_ (_21688_, _21687_, _21686_);
  and _54324_ (_21689_, _21688_, _18964_);
  nor _54325_ (_21690_, _21689_, _18967_);
  and _54326_ (_21691_, _21690_, _21685_);
  and _54327_ (_21692_, _21248_, _18809_);
  and _54328_ (_21693_, _21244_, _18815_);
  or _54329_ (_21694_, _21693_, _21692_);
  or _54330_ (_21695_, _21694_, _18964_);
  and _54331_ (_21696_, _21258_, _18809_);
  and _54332_ (_21697_, _21254_, _18815_);
  nor _54333_ (_21698_, _21697_, _21696_);
  nand _54334_ (_21699_, _21698_, _18964_);
  and _54335_ (_21700_, _21699_, _18967_);
  and _54336_ (_21701_, _21700_, _21695_);
  nor _54337_ (_21702_, _21701_, _21691_);
  nor _54338_ (_21703_, _21702_, _19024_);
  or _54339_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _21703_, _21681_);
  and _54340_ (_21704_, _19024_, word_in[25]);
  or _54341_ (_21705_, _21269_, _18809_);
  or _54342_ (_21706_, _21273_, _18815_);
  and _54343_ (_21707_, _21706_, _21705_);
  or _54344_ (_21708_, _21707_, _18964_);
  or _54345_ (_21709_, _21279_, _18809_);
  or _54346_ (_21710_, _21283_, _18815_);
  nand _54347_ (_21711_, _21710_, _21709_);
  nand _54348_ (_21712_, _21711_, _18964_);
  and _54349_ (_21713_, _21712_, _21708_);
  and _54350_ (_21714_, _21713_, _19035_);
  and _54351_ (_21715_, _21291_, _18815_);
  and _54352_ (_21716_, _21295_, _18809_);
  or _54353_ (_21717_, _21716_, _21715_);
  or _54354_ (_21718_, _21717_, _18964_);
  and _54355_ (_21719_, _21305_, _18809_);
  and _54356_ (_21720_, _21301_, _18815_);
  nor _54357_ (_21721_, _21720_, _21719_);
  nand _54358_ (_21722_, _21721_, _18964_);
  and _54359_ (_21723_, _21722_, _21718_);
  and _54360_ (_21724_, _21723_, _18967_);
  nor _54361_ (_21725_, _21724_, _21714_);
  nor _54362_ (_21726_, _21725_, _19024_);
  or _54363_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _21726_, _21704_);
  and _54364_ (_21727_, _19024_, word_in[26]);
  or _54365_ (_21728_, _21326_, _18809_);
  or _54366_ (_21729_, _21330_, _18815_);
  nand _54367_ (_21730_, _21729_, _21728_);
  nand _54368_ (_21731_, _21730_, _18964_);
  or _54369_ (_21732_, _21316_, _18809_);
  or _54370_ (_21733_, _21320_, _18815_);
  and _54371_ (_21734_, _21733_, _21732_);
  or _54372_ (_21735_, _21734_, _18964_);
  and _54373_ (_21736_, _21735_, _21731_);
  and _54374_ (_21737_, _21736_, _19035_);
  and _54375_ (_21738_, _21338_, _18815_);
  and _54376_ (_21739_, _21342_, _18809_);
  or _54377_ (_21740_, _21739_, _21738_);
  or _54378_ (_21741_, _21740_, _18964_);
  and _54379_ (_21742_, _21352_, _18809_);
  and _54380_ (_21743_, _21348_, _18815_);
  nor _54381_ (_21744_, _21743_, _21742_);
  nand _54382_ (_21745_, _21744_, _18964_);
  and _54383_ (_21746_, _21745_, _21741_);
  and _54384_ (_21747_, _21746_, _18967_);
  nor _54385_ (_21748_, _21747_, _21737_);
  nor _54386_ (_21749_, _21748_, _19024_);
  or _54387_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _21749_, _21727_);
  and _54388_ (_21750_, _19024_, word_in[27]);
  and _54389_ (_21751_, _21367_, _18809_);
  and _54390_ (_21752_, _21363_, _18815_);
  or _54391_ (_21753_, _21752_, _21751_);
  or _54392_ (_21754_, _21753_, _18964_);
  and _54393_ (_21755_, _21377_, _18809_);
  and _54394_ (_21756_, _21373_, _18815_);
  nor _54395_ (_21757_, _21756_, _21755_);
  and _54396_ (_21758_, _21757_, _18964_);
  nor _54397_ (_21759_, _21758_, _18967_);
  and _54398_ (_21760_, _21759_, _21754_);
  and _54399_ (_21761_, _21389_, _18809_);
  and _54400_ (_21762_, _21385_, _18815_);
  or _54401_ (_21763_, _21762_, _21761_);
  or _54402_ (_21764_, _21763_, _18964_);
  and _54403_ (_21765_, _21399_, _18809_);
  and _54404_ (_21766_, _21395_, _18815_);
  nor _54405_ (_21767_, _21766_, _21765_);
  nand _54406_ (_21768_, _21767_, _18964_);
  and _54407_ (_21769_, _21768_, _18967_);
  and _54408_ (_21770_, _21769_, _21764_);
  nor _54409_ (_21771_, _21770_, _21760_);
  nor _54410_ (_21772_, _21771_, _19024_);
  or _54411_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _21772_, _21750_);
  and _54412_ (_21773_, _19024_, word_in[28]);
  or _54413_ (_21774_, _21410_, _18809_);
  or _54414_ (_21775_, _21414_, _18815_);
  and _54415_ (_21776_, _21775_, _21774_);
  or _54416_ (_21777_, _21776_, _18964_);
  or _54417_ (_21778_, _21420_, _18809_);
  or _54418_ (_21779_, _21424_, _18815_);
  nand _54419_ (_21780_, _21779_, _21778_);
  nand _54420_ (_21781_, _21780_, _18964_);
  and _54421_ (_21782_, _21781_, _21777_);
  and _54422_ (_21783_, _21782_, _19035_);
  and _54423_ (_21784_, _21432_, _18815_);
  and _54424_ (_21785_, _21436_, _18809_);
  or _54425_ (_21786_, _21785_, _21784_);
  or _54426_ (_21787_, _21786_, _18964_);
  and _54427_ (_21788_, _21446_, _18809_);
  and _54428_ (_21789_, _21442_, _18815_);
  nor _54429_ (_21790_, _21789_, _21788_);
  nand _54430_ (_21791_, _21790_, _18964_);
  and _54431_ (_21792_, _21791_, _21787_);
  and _54432_ (_21793_, _21792_, _18967_);
  nor _54433_ (_21794_, _21793_, _21783_);
  nor _54434_ (_21795_, _21794_, _19024_);
  or _54435_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _21795_, _21773_);
  and _54436_ (_21796_, _19024_, word_in[29]);
  and _54437_ (_21797_, _21461_, _18809_);
  and _54438_ (_21798_, _21457_, _18815_);
  or _54439_ (_21799_, _21798_, _21797_);
  or _54440_ (_21800_, _21799_, _18964_);
  and _54441_ (_21801_, _21471_, _18809_);
  and _54442_ (_21802_, _21467_, _18815_);
  nor _54443_ (_21803_, _21802_, _21801_);
  and _54444_ (_21804_, _21803_, _18964_);
  nor _54445_ (_21805_, _21804_, _18967_);
  and _54446_ (_21806_, _21805_, _21800_);
  and _54447_ (_21807_, _21483_, _18809_);
  and _54448_ (_21808_, _21479_, _18815_);
  or _54449_ (_21809_, _21808_, _21807_);
  or _54450_ (_21810_, _21809_, _18964_);
  and _54451_ (_21811_, _21493_, _18809_);
  and _54452_ (_21812_, _21489_, _18815_);
  nor _54453_ (_21813_, _21812_, _21811_);
  nand _54454_ (_21814_, _21813_, _18964_);
  and _54455_ (_21815_, _21814_, _18967_);
  and _54456_ (_21816_, _21815_, _21810_);
  nor _54457_ (_21817_, _21816_, _21806_);
  nor _54458_ (_21818_, _21817_, _19024_);
  or _54459_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _21818_, _21796_);
  and _54460_ (_21819_, _19024_, word_in[30]);
  or _54461_ (_21820_, _21504_, _18809_);
  or _54462_ (_21821_, _21508_, _18815_);
  and _54463_ (_21822_, _21821_, _21820_);
  or _54464_ (_21823_, _21822_, _18964_);
  or _54465_ (_21824_, _21514_, _18809_);
  or _54466_ (_21825_, _21518_, _18815_);
  nand _54467_ (_21826_, _21825_, _21824_);
  nand _54468_ (_21827_, _21826_, _18964_);
  and _54469_ (_21828_, _21827_, _21823_);
  and _54470_ (_21829_, _21828_, _19035_);
  and _54471_ (_21830_, _21526_, _18815_);
  and _54472_ (_21831_, _21530_, _18809_);
  or _54473_ (_21832_, _21831_, _21830_);
  or _54474_ (_21833_, _21832_, _18964_);
  and _54475_ (_21834_, _21540_, _18809_);
  and _54476_ (_21835_, _21536_, _18815_);
  nor _54477_ (_21836_, _21835_, _21834_);
  nand _54478_ (_21837_, _21836_, _18964_);
  and _54479_ (_21838_, _21837_, _21833_);
  and _54480_ (_21839_, _21838_, _18967_);
  nor _54481_ (_21840_, _21839_, _21829_);
  nor _54482_ (_21841_, _21840_, _19024_);
  or _54483_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _21841_, _21819_);
  not _54484_ (_21842_, first_instr);
  nor _54485_ (_21843_, pc_log_change, _21842_);
  or _54486_ (_00001_, _21843_, rst);
  or _54487_ (_21844_, pc_log_change_r, cy_reg);
  nand _54488_ (_21845_, pc_log_change_r, _26928_);
  and _54489_ (_00000_, _21845_, _21844_);
  and _54490_ (_21846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _54491_ (_21847_, _21846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _54492_ (_21848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _54493_ (_21849_, _21848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _54494_ (_21850_, _21849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _54495_ (_21851_, _21850_, _21847_);
  and _54496_ (_21852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _54497_ (_21853_, _21852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _54498_ (_21854_, _21853_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _54499_ (_21855_, _21854_, _21851_);
  and _54500_ (_21856_, _21855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _54501_ (_21857_, _21856_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _54502_ (_21858_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _54503_ (_21859_, _21858_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _54504_ (_21860_, _21858_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _54505_ (_21861_, _21860_, _21859_);
  and _54506_ (_21862_, _21861_, cy_reg);
  nor _54507_ (_21863_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _54508_ (_21864_, _21863_);
  and _54509_ (_21865_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _16515_);
  and _54510_ (_21866_, _21846_, _16527_);
  nor _54511_ (_21867_, _21846_, _16527_);
  nor _54512_ (_21868_, _21867_, _21866_);
  nor _54513_ (_21869_, _21868_, _16515_);
  nor _54514_ (_21870_, _21869_, _21865_);
  not _54515_ (_21871_, _21870_);
  and _54516_ (_21872_, _16523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _54517_ (_21873_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _16519_);
  nor _54518_ (_21874_, _21873_, _21872_);
  and _54519_ (_21875_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54520_ (_21876_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54521_ (_21877_, _21876_, _21875_);
  nor _54522_ (_21878_, _21877_, _18894_);
  and _54523_ (_21879_, _21877_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _54524_ (_21880_, _21879_, _21878_);
  nor _54525_ (_21881_, _21880_, _21871_);
  nor _54526_ (_21882_, _21877_, _19167_);
  and _54527_ (_21883_, _21877_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _54528_ (_21884_, _21883_, _21882_);
  nor _54529_ (_21885_, _21884_, _21870_);
  nor _54530_ (_21886_, _21885_, _21881_);
  nor _54531_ (_21887_, _21886_, _21864_);
  and _54532_ (_21888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _16515_);
  not _54533_ (_21889_, _21888_);
  nor _54534_ (_21890_, _21877_, _18865_);
  and _54535_ (_21891_, _21877_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _54536_ (_21892_, _21891_, _21890_);
  nor _54537_ (_21893_, _21892_, _21871_);
  not _54538_ (_21894_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _54539_ (_21895_, _21877_, _21894_);
  and _54540_ (_21896_, _21877_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _54541_ (_21897_, _21896_, _21895_);
  nor _54542_ (_21898_, _21897_, _21870_);
  nor _54543_ (_21899_, _21898_, _21893_);
  nor _54544_ (_21900_, _21899_, _21889_);
  nor _54545_ (_21901_, _21900_, _21887_);
  and _54546_ (_21902_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _54547_ (_21903_, _21902_);
  nor _54548_ (_21904_, _21877_, _18931_);
  and _54549_ (_21905_, _21877_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _54550_ (_21906_, _21905_, _21904_);
  nor _54551_ (_21907_, _21906_, _21871_);
  not _54552_ (_21908_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _54553_ (_21909_, _21877_, _21908_);
  and _54554_ (_21910_, _21877_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _54555_ (_21911_, _21910_, _21909_);
  nor _54556_ (_21912_, _21911_, _21870_);
  nor _54557_ (_21913_, _21912_, _21907_);
  nor _54558_ (_21914_, _21913_, _21903_);
  and _54559_ (_21915_, _16519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _54560_ (_21916_, _21915_);
  nor _54561_ (_21917_, _21877_, _18906_);
  and _54562_ (_21918_, _21877_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _54563_ (_21919_, _21918_, _21917_);
  nor _54564_ (_21920_, _21919_, _21871_);
  nor _54565_ (_21921_, _21877_, _19195_);
  and _54566_ (_21922_, _21877_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _54567_ (_21923_, _21922_, _21921_);
  nor _54568_ (_21924_, _21923_, _21870_);
  nor _54569_ (_21925_, _21924_, _21920_);
  nor _54570_ (_21926_, _21925_, _21916_);
  nor _54571_ (_21927_, _21926_, _21914_);
  and _54572_ (_21928_, _21927_, _21901_);
  not _54573_ (_21929_, _21877_);
  and _54574_ (_21930_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _54575_ (_21931_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _54576_ (_21932_, _21931_, _21930_);
  and _54577_ (_21933_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _54578_ (_21934_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _54579_ (_21935_, _21934_, _21933_);
  and _54580_ (_21936_, _21935_, _21932_);
  and _54581_ (_21937_, _21936_, _21929_);
  and _54582_ (_21938_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _54583_ (_21939_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _54584_ (_21940_, _21939_, _21938_);
  and _54585_ (_21941_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _54586_ (_21942_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _54587_ (_21943_, _21942_, _21941_);
  and _54588_ (_21944_, _21943_, _21940_);
  and _54589_ (_21945_, _21944_, _21877_);
  or _54590_ (_21946_, _21945_, _21871_);
  nor _54591_ (_21947_, _21946_, _21937_);
  and _54592_ (_21948_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _54593_ (_21949_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _54594_ (_21950_, _21949_, _21948_);
  and _54595_ (_21951_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _54596_ (_21952_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _54597_ (_21953_, _21952_, _21951_);
  and _54598_ (_21954_, _21953_, _21950_);
  nor _54599_ (_21955_, _21954_, _21877_);
  and _54600_ (_21956_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _54601_ (_21957_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _54602_ (_21958_, _21957_, _21956_);
  and _54603_ (_21959_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _54604_ (_21960_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _54605_ (_21961_, _21960_, _21959_);
  and _54606_ (_21962_, _21961_, _21958_);
  nor _54607_ (_21963_, _21962_, _21929_);
  or _54608_ (_21964_, _21963_, _21955_);
  and _54609_ (_21965_, _21964_, _21871_);
  nor _54610_ (_21966_, _21965_, _21947_);
  nor _54611_ (_21967_, _21966_, _21928_);
  nor _54612_ (_21968_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _54613_ (_21969_, _21968_, _21858_);
  and _54614_ (_21970_, _21969_, _21967_);
  nor _54615_ (_21971_, _21969_, _21967_);
  nor _54616_ (_21972_, _21971_, _21970_);
  not _54617_ (_21973_, _21972_);
  nor _54618_ (_21974_, _21856_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _54619_ (_21975_, _21974_, _21857_);
  nor _54620_ (_21976_, _21975_, _21967_);
  and _54621_ (_21977_, _21975_, _21967_);
  not _54622_ (_21978_, _21977_);
  nor _54623_ (_21979_, _21855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _54624_ (_21980_, _21979_, _21856_);
  and _54625_ (_21981_, _21980_, _21967_);
  and _54626_ (_21982_, _21853_, _21851_);
  nor _54627_ (_21983_, _21982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _54628_ (_21984_, _21982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _54629_ (_21985_, _21984_, _21983_);
  and _54630_ (_21986_, _21985_, _21967_);
  nor _54631_ (_21987_, _21985_, _21967_);
  and _54632_ (_21988_, _21851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _54633_ (_21989_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _54634_ (_21990_, _21989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _54635_ (_21991_, _21990_, _21982_);
  and _54636_ (_21992_, _21991_, _21967_);
  nor _54637_ (_21993_, _21991_, _21967_);
  nor _54638_ (_21994_, _21993_, _21992_);
  not _54639_ (_21995_, _21994_);
  nor _54640_ (_21996_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _54641_ (_21997_, _21996_, _21989_);
  and _54642_ (_21998_, _21997_, _21967_);
  nor _54643_ (_21999_, _21851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _54644_ (_22000_, _21999_, _21988_);
  and _54645_ (_22001_, _22000_, _21967_);
  nor _54646_ (_22002_, _21997_, _21967_);
  nor _54647_ (_22003_, _22002_, _21998_);
  and _54648_ (_22004_, _21849_, _21847_);
  nor _54649_ (_22005_, _22004_, _16540_);
  and _54650_ (_22006_, _22004_, _16540_);
  nor _54651_ (_22007_, _22006_, _22005_);
  not _54652_ (_22008_, _22007_);
  and _54653_ (_22009_, _22008_, _21967_);
  nor _54654_ (_22010_, _22008_, _21967_);
  and _54655_ (_22011_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _54656_ (_22012_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _54657_ (_22013_, _22012_, _22011_);
  and _54658_ (_22014_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _54659_ (_22015_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _54660_ (_22016_, _22015_, _22014_);
  and _54661_ (_22017_, _22016_, _22013_);
  and _54662_ (_22018_, _22017_, _21929_);
  and _54663_ (_22019_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _54664_ (_22020_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _54665_ (_22021_, _22020_, _22019_);
  and _54666_ (_22022_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _54667_ (_22023_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _54668_ (_22024_, _22023_, _22022_);
  and _54669_ (_22025_, _22024_, _22021_);
  and _54670_ (_22026_, _22025_, _21877_);
  or _54671_ (_22027_, _22026_, _21871_);
  nor _54672_ (_22028_, _22027_, _22018_);
  and _54673_ (_22029_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _54674_ (_22030_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _54675_ (_22031_, _22030_, _22029_);
  and _54676_ (_22032_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _54677_ (_22033_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _54678_ (_22034_, _22033_, _22032_);
  and _54679_ (_22035_, _22034_, _22031_);
  nor _54680_ (_22036_, _22035_, _21877_);
  and _54681_ (_22037_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _54682_ (_22038_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _54683_ (_22039_, _22038_, _22037_);
  and _54684_ (_22040_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _54685_ (_22041_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _54686_ (_22042_, _22041_, _22040_);
  and _54687_ (_22043_, _22042_, _22039_);
  nor _54688_ (_22044_, _22043_, _21929_);
  or _54689_ (_22045_, _22044_, _22036_);
  and _54690_ (_22046_, _22045_, _21871_);
  nor _54691_ (_22047_, _22046_, _22028_);
  nor _54692_ (_22048_, _22047_, _21928_);
  and _54693_ (_22049_, _21848_, _21847_);
  nor _54694_ (_22050_, _22049_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _54695_ (_22051_, _22050_, _22004_);
  and _54696_ (_22052_, _22051_, _22048_);
  nor _54697_ (_22053_, _22051_, _22048_);
  nor _54698_ (_22054_, _22053_, _22052_);
  not _54699_ (_22055_, _22054_);
  and _54700_ (_22056_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _54701_ (_22057_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _54702_ (_22058_, _22057_, _22056_);
  and _54703_ (_22059_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _54704_ (_22060_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _54705_ (_22061_, _22060_, _22059_);
  and _54706_ (_22062_, _22061_, _22058_);
  and _54707_ (_22063_, _22062_, _21929_);
  and _54708_ (_22064_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _54709_ (_22065_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _54710_ (_22066_, _22065_, _22064_);
  and _54711_ (_22067_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _54712_ (_22068_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _54713_ (_22069_, _22068_, _22067_);
  and _54714_ (_22070_, _22069_, _22066_);
  and _54715_ (_22071_, _22070_, _21877_);
  or _54716_ (_22072_, _22071_, _21871_);
  nor _54717_ (_22073_, _22072_, _22063_);
  and _54718_ (_22074_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _54719_ (_22075_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _54720_ (_22076_, _22075_, _22074_);
  and _54721_ (_22077_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _54722_ (_22078_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _54723_ (_22079_, _22078_, _22077_);
  and _54724_ (_22080_, _22079_, _22076_);
  nor _54725_ (_22081_, _22080_, _21877_);
  and _54726_ (_22082_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _54727_ (_22083_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _54728_ (_22084_, _22083_, _22082_);
  and _54729_ (_22085_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _54730_ (_22086_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _54731_ (_22087_, _22086_, _22085_);
  and _54732_ (_22088_, _22087_, _22084_);
  nor _54733_ (_22089_, _22088_, _21929_);
  or _54734_ (_22090_, _22089_, _22081_);
  and _54735_ (_22091_, _22090_, _21871_);
  nor _54736_ (_22092_, _22091_, _22073_);
  nor _54737_ (_22093_, _22092_, _21928_);
  and _54738_ (_22094_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _54739_ (_22095_, _22094_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _54740_ (_22096_, _22095_, _22049_);
  and _54741_ (_22097_, _22096_, _22093_);
  nor _54742_ (_22098_, _22096_, _22093_);
  nor _54743_ (_22099_, _22098_, _22097_);
  not _54744_ (_22100_, _22099_);
  and _54745_ (_22101_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _54746_ (_22102_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _54747_ (_22103_, _22102_, _22101_);
  and _54748_ (_22104_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _54749_ (_22105_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _54750_ (_22106_, _22105_, _22104_);
  and _54751_ (_22107_, _22106_, _22103_);
  and _54752_ (_22108_, _22107_, _21929_);
  and _54753_ (_22109_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _54754_ (_22110_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _54755_ (_22111_, _22110_, _22109_);
  and _54756_ (_22112_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _54757_ (_22113_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _54758_ (_22114_, _22113_, _22112_);
  and _54759_ (_22115_, _22114_, _22111_);
  and _54760_ (_22116_, _22115_, _21877_);
  or _54761_ (_22117_, _22116_, _21871_);
  nor _54762_ (_22118_, _22117_, _22108_);
  and _54763_ (_22119_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _54764_ (_22120_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _54765_ (_22121_, _22120_, _22119_);
  and _54766_ (_22122_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _54767_ (_22123_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _54768_ (_22124_, _22123_, _22122_);
  and _54769_ (_22125_, _22124_, _22121_);
  nor _54770_ (_22126_, _22125_, _21877_);
  and _54771_ (_22127_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _54772_ (_22128_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _54773_ (_22129_, _22128_, _22127_);
  and _54774_ (_22130_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _54775_ (_22131_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _54776_ (_22132_, _22131_, _22130_);
  and _54777_ (_22133_, _22132_, _22129_);
  nor _54778_ (_22134_, _22133_, _21929_);
  or _54779_ (_22135_, _22134_, _22126_);
  and _54780_ (_22136_, _22135_, _21871_);
  nor _54781_ (_22137_, _22136_, _22118_);
  nor _54782_ (_22138_, _22137_, _21928_);
  nor _54783_ (_22139_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _54784_ (_22140_, _22139_, _22094_);
  and _54785_ (_22141_, _22140_, _22138_);
  not _54786_ (_22142_, _21868_);
  and _54787_ (_22143_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _54788_ (_22144_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _54789_ (_22145_, _22144_, _22143_);
  and _54790_ (_22146_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _54791_ (_22147_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _54792_ (_22148_, _22147_, _22146_);
  and _54793_ (_22149_, _22148_, _22145_);
  and _54794_ (_22150_, _22149_, _21929_);
  and _54795_ (_22151_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _54796_ (_22152_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _54797_ (_22153_, _22152_, _22151_);
  and _54798_ (_22154_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _54799_ (_22155_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _54800_ (_22156_, _22155_, _22154_);
  and _54801_ (_22157_, _22156_, _22153_);
  and _54802_ (_22158_, _22157_, _21877_);
  or _54803_ (_22159_, _22158_, _21871_);
  nor _54804_ (_22160_, _22159_, _22150_);
  and _54805_ (_22161_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _54806_ (_22162_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _54807_ (_22163_, _22162_, _22161_);
  and _54808_ (_22164_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _54809_ (_22165_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _54810_ (_22166_, _22165_, _22164_);
  and _54811_ (_22167_, _22166_, _22163_);
  nor _54812_ (_22168_, _22167_, _21877_);
  and _54813_ (_22169_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _54814_ (_22170_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _54815_ (_22171_, _22170_, _22169_);
  and _54816_ (_22172_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _54817_ (_22173_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _54818_ (_22174_, _22173_, _22172_);
  and _54819_ (_22175_, _22174_, _22171_);
  nor _54820_ (_22176_, _22175_, _21929_);
  or _54821_ (_22177_, _22176_, _22168_);
  and _54822_ (_22178_, _22177_, _21871_);
  nor _54823_ (_22179_, _22178_, _22160_);
  nor _54824_ (_22180_, _22179_, _21928_);
  and _54825_ (_22181_, _22180_, _22142_);
  nor _54826_ (_22182_, _22180_, _22142_);
  nor _54827_ (_22183_, _22182_, _22181_);
  not _54828_ (_22184_, _22183_);
  not _54829_ (_22185_, _21874_);
  and _54830_ (_22186_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _54831_ (_22187_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _54832_ (_22188_, _22187_, _22186_);
  and _54833_ (_22189_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _54834_ (_22190_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _54835_ (_22191_, _22190_, _22189_);
  and _54836_ (_22192_, _22191_, _22188_);
  and _54837_ (_22193_, _22192_, _21929_);
  and _54838_ (_22194_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _54839_ (_22195_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _54840_ (_22196_, _22195_, _22194_);
  and _54841_ (_22197_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _54842_ (_22198_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _54843_ (_22199_, _22198_, _22197_);
  and _54844_ (_22200_, _22199_, _22196_);
  and _54845_ (_22201_, _22200_, _21877_);
  or _54846_ (_22202_, _22201_, _21871_);
  nor _54847_ (_22203_, _22202_, _22193_);
  and _54848_ (_22204_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _54849_ (_22205_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _54850_ (_22206_, _22205_, _22204_);
  and _54851_ (_22207_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _54852_ (_22208_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _54853_ (_22209_, _22208_, _22207_);
  and _54854_ (_22210_, _22209_, _22206_);
  nor _54855_ (_22211_, _22210_, _21877_);
  and _54856_ (_22212_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _54857_ (_22213_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _54858_ (_22214_, _22213_, _22212_);
  and _54859_ (_22215_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _54860_ (_22216_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _54861_ (_22217_, _22216_, _22215_);
  and _54862_ (_22218_, _22217_, _22214_);
  nor _54863_ (_22219_, _22218_, _21929_);
  or _54864_ (_22220_, _22219_, _22211_);
  and _54865_ (_22221_, _22220_, _21871_);
  nor _54866_ (_22222_, _22221_, _22203_);
  nor _54867_ (_22223_, _22222_, _21928_);
  and _54868_ (_22224_, _22223_, _22185_);
  and _54869_ (_22225_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _54870_ (_22226_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _54871_ (_22227_, _22226_, _22225_);
  and _54872_ (_22228_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _54873_ (_22229_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _54874_ (_22230_, _22229_, _22228_);
  and _54875_ (_22231_, _22230_, _22227_);
  and _54876_ (_22232_, _22231_, _21929_);
  and _54877_ (_22233_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _54878_ (_22234_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _54879_ (_22235_, _22234_, _22233_);
  and _54880_ (_22236_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _54881_ (_22237_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _54882_ (_22238_, _22237_, _22236_);
  and _54883_ (_22239_, _22238_, _22235_);
  and _54884_ (_22240_, _22239_, _21877_);
  or _54885_ (_22241_, _22240_, _21871_);
  nor _54886_ (_22242_, _22241_, _22232_);
  and _54887_ (_22243_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _54888_ (_22244_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _54889_ (_22245_, _22244_, _22243_);
  and _54890_ (_22246_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _54891_ (_22247_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _54892_ (_22248_, _22247_, _22246_);
  and _54893_ (_22249_, _22248_, _22245_);
  nor _54894_ (_22250_, _22249_, _21877_);
  and _54895_ (_22251_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _54896_ (_22252_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _54897_ (_22253_, _22252_, _22251_);
  and _54898_ (_22254_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _54899_ (_22255_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _54900_ (_22256_, _22255_, _22254_);
  and _54901_ (_22257_, _22256_, _22253_);
  nor _54902_ (_22258_, _22257_, _21929_);
  or _54903_ (_22259_, _22258_, _22250_);
  and _54904_ (_22260_, _22259_, _21871_);
  nor _54905_ (_22261_, _22260_, _22242_);
  nor _54906_ (_22262_, _22261_, _21928_);
  and _54907_ (_22263_, _22262_, _16519_);
  and _54908_ (_22264_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _54909_ (_22265_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _54910_ (_22266_, _22265_, _22264_);
  and _54911_ (_22267_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _54912_ (_22268_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _54913_ (_22269_, _22268_, _22267_);
  and _54914_ (_22270_, _22269_, _22266_);
  and _54915_ (_22271_, _22270_, _21929_);
  and _54916_ (_22272_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _54917_ (_22273_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _54918_ (_22274_, _22273_, _22272_);
  and _54919_ (_22275_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _54920_ (_22276_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _54921_ (_22277_, _22276_, _22275_);
  and _54922_ (_22278_, _22277_, _22274_);
  and _54923_ (_22279_, _22278_, _21877_);
  or _54924_ (_22280_, _22279_, _21871_);
  nor _54925_ (_22281_, _22280_, _22271_);
  and _54926_ (_22282_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _54927_ (_22283_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _54928_ (_22284_, _22283_, _22282_);
  and _54929_ (_22285_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _54930_ (_22286_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _54931_ (_22287_, _22286_, _22285_);
  and _54932_ (_22288_, _22287_, _22284_);
  nor _54933_ (_22289_, _22288_, _21877_);
  and _54934_ (_22290_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _54935_ (_22291_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _54936_ (_22292_, _22291_, _22290_);
  and _54937_ (_22293_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _54938_ (_22294_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _54939_ (_22295_, _22294_, _22293_);
  and _54940_ (_22296_, _22295_, _22292_);
  nor _54941_ (_22297_, _22296_, _21929_);
  or _54942_ (_22298_, _22297_, _22289_);
  and _54943_ (_22299_, _22298_, _21871_);
  nor _54944_ (_22300_, _22299_, _22281_);
  nor _54945_ (_22301_, _22300_, _21928_);
  and _54946_ (_22302_, _22301_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54947_ (_22303_, _22262_, _16519_);
  nor _54948_ (_22304_, _22303_, _22263_);
  and _54949_ (_22305_, _22304_, _22302_);
  nor _54950_ (_22306_, _22305_, _22263_);
  nor _54951_ (_22307_, _22223_, _22185_);
  nor _54952_ (_22308_, _22307_, _22224_);
  not _54953_ (_22309_, _22308_);
  nor _54954_ (_22310_, _22309_, _22306_);
  nor _54955_ (_22311_, _22310_, _22224_);
  nor _54956_ (_22312_, _22311_, _22184_);
  nor _54957_ (_22313_, _22312_, _22181_);
  nor _54958_ (_22314_, _22140_, _22138_);
  nor _54959_ (_22315_, _22314_, _22141_);
  not _54960_ (_22316_, _22315_);
  nor _54961_ (_22317_, _22316_, _22313_);
  nor _54962_ (_22318_, _22317_, _22141_);
  nor _54963_ (_22319_, _22318_, _22100_);
  nor _54964_ (_22320_, _22319_, _22097_);
  nor _54965_ (_22321_, _22320_, _22055_);
  nor _54966_ (_22322_, _22321_, _22052_);
  nor _54967_ (_22323_, _22322_, _22010_);
  or _54968_ (_22324_, _22323_, _22009_);
  nor _54969_ (_22325_, _22000_, _21967_);
  nor _54970_ (_22326_, _22325_, _22001_);
  and _54971_ (_22327_, _22326_, _22324_);
  and _54972_ (_22328_, _22327_, _22003_);
  or _54973_ (_22329_, _22328_, _22001_);
  nor _54974_ (_22330_, _22329_, _21998_);
  nor _54975_ (_22331_, _22330_, _21995_);
  nor _54976_ (_22332_, _22331_, _21992_);
  nor _54977_ (_22333_, _22332_, _21987_);
  or _54978_ (_22334_, _22333_, _21986_);
  nor _54979_ (_22335_, _21980_, _21967_);
  nor _54980_ (_22336_, _22335_, _21981_);
  and _54981_ (_22337_, _22336_, _22334_);
  nor _54982_ (_22338_, _22337_, _21981_);
  and _54983_ (_22339_, _22338_, _21978_);
  or _54984_ (_22340_, _22339_, _21976_);
  nor _54985_ (_22341_, _22340_, _21973_);
  nor _54986_ (_22342_, _22341_, _21970_);
  and _54987_ (_22343_, _21967_, _21861_);
  nor _54988_ (_22344_, _21967_, _21861_);
  or _54989_ (_22345_, _22344_, _22343_);
  and _54990_ (_22346_, _22345_, _22342_);
  nor _54991_ (_22347_, _22345_, _22342_);
  or _54992_ (_22348_, _22347_, _22346_);
  nor _54993_ (_22349_, _22348_, cy_reg);
  nor _54994_ (_22350_, _22349_, _21862_);
  nor _54995_ (_22351_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _54996_ (_22352_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _54997_ (_22353_, _21969_, cy_reg);
  not _54998_ (_22354_, cy_reg);
  and _54999_ (_22355_, _22340_, _21973_);
  nor _55000_ (_22356_, _22355_, _22341_);
  and _55001_ (_22357_, _22356_, _22354_);
  nor _55002_ (_22358_, _22357_, _22353_);
  nor _55003_ (_22359_, _22358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _55004_ (_22360_, _22358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _55005_ (_22361_, _21976_, _21977_);
  nor _55006_ (_22362_, _22361_, _22338_);
  and _55007_ (_22363_, _22361_, _22338_);
  nor _55008_ (_22364_, _22363_, _22362_);
  nor _55009_ (_22365_, _22364_, cy_reg);
  and _55010_ (_22366_, _21975_, cy_reg);
  nor _55011_ (_22367_, _22366_, _22365_);
  and _55012_ (_22368_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _55013_ (_22369_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _55014_ (_22370_, _22336_, _22334_);
  nor _55015_ (_22371_, _22370_, _22337_);
  nor _55016_ (_22372_, _22371_, cy_reg);
  nor _55017_ (_22373_, _21980_, _22354_);
  nor _55018_ (_22374_, _22373_, _22372_);
  nor _55019_ (_22375_, _22374_, _16503_);
  and _55020_ (_22376_, _22374_, _16503_);
  and _55021_ (_22377_, _21985_, cy_reg);
  nor _55022_ (_22378_, _21986_, _21987_);
  nor _55023_ (_22379_, _22378_, _22332_);
  and _55024_ (_22380_, _22378_, _22332_);
  nor _55025_ (_22381_, _22380_, _22379_);
  nor _55026_ (_22382_, _22381_, cy_reg);
  nor _55027_ (_22383_, _22382_, _22377_);
  and _55028_ (_22384_, _22383_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _55029_ (_22385_, _22383_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _55030_ (_22386_, _22327_, _22001_);
  and _55031_ (_22387_, _22386_, _22003_);
  nor _55032_ (_22388_, _22386_, _22003_);
  nor _55033_ (_22389_, _22388_, _22387_);
  nor _55034_ (_22390_, _22389_, cy_reg);
  and _55035_ (_22391_, _21997_, cy_reg);
  nor _55036_ (_22392_, _22391_, _22390_);
  nand _55037_ (_22393_, _22392_, _16491_);
  or _55038_ (_22394_, _22392_, _16491_);
  and _55039_ (_22395_, _22394_, _22393_);
  nor _55040_ (_22396_, _22000_, _16487_);
  and _55041_ (_22397_, _22000_, _16487_);
  or _55042_ (_22398_, _22397_, _22396_);
  or _55043_ (_22399_, _22007_, _16483_);
  nand _55044_ (_22400_, _22007_, _16483_);
  and _55045_ (_22401_, _22400_, _22399_);
  or _55046_ (_22402_, _22401_, _22354_);
  or _55047_ (_22403_, _22402_, _22398_);
  nor _55048_ (_22404_, _22326_, _22324_);
  nor _55049_ (_22405_, _22404_, _22327_);
  or _55050_ (_22406_, _22405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _55051_ (_22407_, _22405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _55052_ (_22408_, _22407_, _22406_);
  nor _55053_ (_22409_, _22009_, _22010_);
  nor _55054_ (_22410_, _22409_, _22322_);
  and _55055_ (_22411_, _22409_, _22322_);
  nor _55056_ (_22412_, _22411_, _22410_);
  nor _55057_ (_22413_, _22412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _55058_ (_22414_, _22412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _55059_ (_22415_, _22414_, _22413_);
  or _55060_ (_22416_, _22415_, cy_reg);
  or _55061_ (_22417_, _22416_, _22408_);
  and _55062_ (_22418_, _22417_, _22403_);
  and _55063_ (_22419_, _22051_, cy_reg);
  and _55064_ (_22420_, _22320_, _22055_);
  nor _55065_ (_22421_, _22420_, _22321_);
  and _55066_ (_22422_, _22421_, _22354_);
  nor _55067_ (_22423_, _22422_, _22419_);
  nor _55068_ (_22424_, _22423_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _55069_ (_22425_, _22423_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _55070_ (_22426_, _22318_, _22100_);
  nor _55071_ (_22427_, _22426_, _22319_);
  and _55072_ (_22428_, _22427_, _22354_);
  and _55073_ (_22429_, _22096_, cy_reg);
  nor _55074_ (_22430_, _22429_, _22428_);
  and _55075_ (_22431_, _22430_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _55076_ (_22432_, _22430_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _55077_ (_22433_, _22140_, cy_reg);
  and _55078_ (_22434_, _22316_, _22313_);
  nor _55079_ (_22435_, _22434_, _22317_);
  and _55080_ (_22436_, _22435_, _22354_);
  nor _55081_ (_22437_, _22436_, _22433_);
  and _55082_ (_22438_, _22437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _55083_ (_22439_, _22437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _55084_ (_22440_, _22311_, _22184_);
  nor _55085_ (_22441_, _22440_, _22312_);
  and _55086_ (_22442_, _22441_, _22354_);
  nor _55087_ (_22443_, _21868_, _22354_);
  nor _55088_ (_22444_, _22443_, _22442_);
  nor _55089_ (_22445_, _22444_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55090_ (_22446_, _22444_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55091_ (_22447_, cy_reg, _16519_);
  nor _55092_ (_22448_, _22304_, _22302_);
  nor _55093_ (_22449_, _22448_, _22305_);
  and _55094_ (_22450_, _22449_, _22354_);
  nor _55095_ (_22451_, _22450_, _22447_);
  and _55096_ (_22452_, _22451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _55097_ (_22453_, _22301_, _22354_);
  and _55098_ (_22454_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _55099_ (_22455_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _55100_ (_22456_, _22455_, _22454_);
  nor _55101_ (_22457_, _22456_, _22453_);
  and _55102_ (_22458_, _22456_, _22301_);
  and _55103_ (_22459_, _22458_, _22354_);
  or _55104_ (_22460_, _22459_, _22457_);
  nor _55105_ (_22461_, _22451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _55106_ (_22462_, _22461_, _22460_);
  or _55107_ (_22463_, _22462_, _22452_);
  and _55108_ (_22464_, _22309_, _22306_);
  nor _55109_ (_22465_, _22464_, _22310_);
  and _55110_ (_22466_, _22465_, _22354_);
  nor _55111_ (_22467_, _21874_, _22354_);
  nor _55112_ (_22468_, _22467_, _22466_);
  nor _55113_ (_22469_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _55114_ (_22470_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _55115_ (_22471_, _22470_, _22469_);
  or _55116_ (_22472_, _22471_, _22463_);
  or _55117_ (_22473_, _22472_, _22446_);
  or _55118_ (_22474_, _22473_, _22445_);
  or _55119_ (_22475_, _22474_, _22439_);
  or _55120_ (_22476_, _22475_, _22438_);
  or _55121_ (_22477_, _22476_, _22432_);
  or _55122_ (_22478_, _22477_, _22431_);
  or _55123_ (_22479_, _22478_, _22425_);
  or _55124_ (_22480_, _22479_, _22424_);
  or _55125_ (_22481_, _22480_, _22418_);
  or _55126_ (_22482_, _22481_, _22395_);
  and _55127_ (_22483_, _21991_, cy_reg);
  and _55128_ (_22484_, _22330_, _21995_);
  nor _55129_ (_22485_, _22484_, _22331_);
  and _55130_ (_22486_, _22485_, _22354_);
  nor _55131_ (_22487_, _22486_, _22483_);
  and _55132_ (_22488_, _22487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _55133_ (_22489_, _22487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or _55134_ (_22490_, _22489_, _22488_);
  or _55135_ (_22491_, _22490_, _22482_);
  or _55136_ (_22492_, _22491_, _22385_);
  or _55137_ (_22493_, _22492_, _22384_);
  or _55138_ (_22494_, _22493_, _22376_);
  or _55139_ (_22495_, _22494_, _22375_);
  or _55140_ (_22496_, _22495_, _22369_);
  or _55141_ (_22497_, _22496_, _22368_);
  or _55142_ (_22498_, _22497_, _22360_);
  or _55143_ (_22499_, _22498_, _22359_);
  or _55144_ (_22500_, _22499_, _22352_);
  or _55145_ (_22501_, _22500_, _22351_);
  and _55146_ (_22502_, _18925_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55147_ (_22503_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55148_ (_22504_, _22503_, _22502_);
  and _55149_ (_22505_, _22504_, _21873_);
  nor _55150_ (_22506_, _22505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55151_ (_22507_, _18915_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _55152_ (_22508_, _22507_);
  nor _55153_ (_22509_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55154_ (_22510_, _22509_, _16523_);
  and _55155_ (_22511_, _22510_, _22508_);
  and _55156_ (_22512_, _19195_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55157_ (_22513_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55158_ (_22514_, _22513_, _22512_);
  and _55159_ (_22515_, _22514_, _16523_);
  nor _55160_ (_22516_, _22515_, _22511_);
  nor _55161_ (_22517_, _22516_, _16519_);
  nor _55162_ (_22518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _55163_ (_22519_, _21908_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55164_ (_22520_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55165_ (_22521_, _22520_, _22519_);
  and _55166_ (_22522_, _22521_, _22518_);
  nor _55167_ (_22523_, _22522_, _22517_);
  and _55168_ (_22524_, _22523_, _22506_);
  nor _55169_ (_22525_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _55170_ (_22526_, _22525_);
  and _55171_ (_22527_, _18879_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55172_ (_22528_, _22527_, _16523_);
  and _55173_ (_22529_, _22528_, _22526_);
  and _55174_ (_22530_, _21894_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55175_ (_22531_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55176_ (_22532_, _22531_, _22530_);
  and _55177_ (_22533_, _22532_, _16523_);
  nor _55178_ (_22534_, _22533_, _22529_);
  nor _55179_ (_22535_, _22534_, _16519_);
  nor _55180_ (_22536_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _55181_ (_22537_, _19167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55182_ (_22538_, _22537_, _22536_);
  and _55183_ (_22539_, _22538_, _22518_);
  nor _55184_ (_22540_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _55185_ (_22541_, _18887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55186_ (_22542_, _22541_, _22540_);
  and _55187_ (_22543_, _22542_, _21873_);
  or _55188_ (_22544_, _22543_, _16515_);
  or _55189_ (_22545_, _22544_, _22539_);
  nor _55190_ (_22546_, _22545_, _22535_);
  nor _55191_ (_22547_, _22546_, _22524_);
  nor _55192_ (_22548_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55193_ (_22549_, _21040_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55194_ (_22550_, _22549_, _22548_);
  and _55195_ (_22551_, _22550_, _21872_);
  nor _55196_ (_22552_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55197_ (_22553_, _19831_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55198_ (_22554_, _22553_, _22552_);
  and _55199_ (_22555_, _22554_, _21873_);
  nor _55200_ (_22556_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55201_ (_22557_, _21050_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55202_ (_22558_, _22557_, _22556_);
  and _55203_ (_22559_, _22558_, _22518_);
  nor _55204_ (_22560_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55205_ (_22561_, _20042_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55206_ (_22562_, _22561_, _22560_);
  and _55207_ (_22563_, _22562_, _21846_);
  or _55208_ (_22564_, _22563_, _22559_);
  or _55209_ (_22565_, _22564_, _22555_);
  or _55210_ (_22566_, _22565_, _22551_);
  and _55211_ (_22567_, _22566_, _16527_);
  nor _55212_ (_22568_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55213_ (_22569_, _20453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55214_ (_22570_, _22569_, _22568_);
  and _55215_ (_22571_, _22570_, _21872_);
  nor _55216_ (_22572_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55217_ (_22573_, _20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55218_ (_22574_, _22573_, _22572_);
  and _55219_ (_22575_, _22574_, _21873_);
  nor _55220_ (_22576_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55221_ (_22577_, _20249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55222_ (_22578_, _22577_, _22576_);
  and _55223_ (_22579_, _22578_, _22518_);
  nor _55224_ (_22580_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55225_ (_22581_, _21073_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55226_ (_22582_, _22581_, _22580_);
  and _55227_ (_22583_, _22582_, _21846_);
  or _55228_ (_22584_, _22583_, _22579_);
  or _55229_ (_22585_, _22584_, _22575_);
  or _55230_ (_22586_, _22585_, _22571_);
  and _55231_ (_22587_, _22586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55232_ (_22588_, _22587_, _22567_);
  and _55233_ (_22589_, _22588_, _22547_);
  nor _55234_ (_22590_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55235_ (_22591_, _21019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55236_ (_22592_, _22591_, _22590_);
  and _55237_ (_22593_, _22592_, _21872_);
  nor _55238_ (_22594_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55239_ (_22595_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55240_ (_22596_, _22595_, _22594_);
  and _55241_ (_22597_, _22596_, _21873_);
  nor _55242_ (_22598_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55243_ (_22599_, _21009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55244_ (_22600_, _22599_, _22598_);
  and _55245_ (_22601_, _22600_, _22518_);
  nor _55246_ (_22602_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55247_ (_22603_, _20030_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55248_ (_22604_, _22603_, _22602_);
  and _55249_ (_22605_, _22604_, _21846_);
  or _55250_ (_22606_, _22605_, _22601_);
  or _55251_ (_22607_, _22606_, _22597_);
  or _55252_ (_22608_, _22607_, _22593_);
  and _55253_ (_22609_, _22608_, _16527_);
  nor _55254_ (_22610_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55255_ (_22611_, _20442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55256_ (_22612_, _22611_, _22610_);
  and _55257_ (_22613_, _22612_, _21872_);
  nor _55258_ (_22614_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55259_ (_22615_, _20645_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55260_ (_22616_, _22615_, _22614_);
  and _55261_ (_22617_, _22616_, _21873_);
  nor _55262_ (_22618_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55263_ (_22619_, _20237_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55264_ (_22620_, _22619_, _22618_);
  and _55265_ (_22621_, _22620_, _22518_);
  nor _55266_ (_22622_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55267_ (_22623_, _21027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55268_ (_22624_, _22623_, _22622_);
  and _55269_ (_22625_, _22624_, _21846_);
  or _55270_ (_22626_, _22625_, _22621_);
  or _55271_ (_22627_, _22626_, _22617_);
  or _55272_ (_22628_, _22627_, _22613_);
  and _55273_ (_22629_, _22628_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55274_ (_22630_, _22629_, _22609_);
  and _55275_ (_22631_, _22630_, _22547_);
  nor _55276_ (_22632_, _22631_, _22589_);
  nor _55277_ (_22633_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55278_ (_22634_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55279_ (_22635_, _22634_, _22633_);
  and _55280_ (_22636_, _22635_, _21872_);
  nor _55281_ (_22637_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55282_ (_22638_, _19806_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55283_ (_22639_, _22638_, _22637_);
  and _55284_ (_22640_, _22639_, _21873_);
  nor _55285_ (_22641_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55286_ (_22642_, _20973_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55287_ (_22643_, _22642_, _22641_);
  and _55288_ (_22644_, _22643_, _22518_);
  nor _55289_ (_22645_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55290_ (_22646_, _20016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55291_ (_22647_, _22646_, _22645_);
  and _55292_ (_22648_, _22647_, _21846_);
  or _55293_ (_22649_, _22648_, _22644_);
  or _55294_ (_22650_, _22649_, _22640_);
  or _55295_ (_22651_, _22650_, _22636_);
  and _55296_ (_22652_, _22651_, _16527_);
  nor _55297_ (_22653_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55298_ (_22654_, _20429_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55299_ (_22655_, _22654_, _22653_);
  and _55300_ (_22656_, _22655_, _21872_);
  nor _55301_ (_22657_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55302_ (_22658_, _20633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55303_ (_22659_, _22658_, _22657_);
  and _55304_ (_22660_, _22659_, _21873_);
  nor _55305_ (_22661_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55306_ (_22662_, _20223_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55307_ (_22663_, _22662_, _22661_);
  and _55308_ (_22664_, _22663_, _22518_);
  nor _55309_ (_22665_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55310_ (_22666_, _20981_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55311_ (_22667_, _22666_, _22665_);
  and _55312_ (_22668_, _22667_, _21846_);
  or _55313_ (_22669_, _22668_, _22664_);
  or _55314_ (_22670_, _22669_, _22660_);
  or _55315_ (_22671_, _22670_, _22656_);
  and _55316_ (_22672_, _22671_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55317_ (_22673_, _22672_, _22652_);
  and _55318_ (_22674_, _22673_, _22547_);
  nor _55319_ (_22675_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55320_ (_22676_, _20620_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55321_ (_22677_, _22676_, _22675_);
  and _55322_ (_22678_, _22677_, _21873_);
  nor _55323_ (_22679_, _22678_, _16527_);
  nor _55324_ (_22680_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55325_ (_22681_, _20209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55326_ (_22682_, _22681_, _22680_);
  and _55327_ (_22683_, _22682_, _22518_);
  nor _55328_ (_22684_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55329_ (_22685_, _20412_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55330_ (_22686_, _22685_, _22684_);
  and _55331_ (_22687_, _22686_, _21872_);
  nor _55332_ (_22688_, _22687_, _22683_);
  nor _55333_ (_22689_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55334_ (_22690_, _20935_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55335_ (_22691_, _22690_, _22689_);
  and _55336_ (_22692_, _22691_, _21846_);
  not _55337_ (_22693_, _22692_);
  and _55338_ (_22694_, _22693_, _22688_);
  and _55339_ (_22695_, _22694_, _22679_);
  nor _55340_ (_22696_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55341_ (_22697_, _19790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55342_ (_22698_, _22697_, _22696_);
  and _55343_ (_22699_, _22698_, _21873_);
  nor _55344_ (_22700_, _22699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55345_ (_22701_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55346_ (_22702_, _20917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55347_ (_22703_, _22702_, _22701_);
  and _55348_ (_22704_, _22703_, _22518_);
  nor _55349_ (_22705_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55350_ (_22706_, _20927_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55351_ (_22707_, _22706_, _22705_);
  and _55352_ (_22708_, _22707_, _21872_);
  nor _55353_ (_22709_, _22708_, _22704_);
  nor _55354_ (_22710_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55355_ (_22711_, _20002_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55356_ (_22712_, _22711_, _22710_);
  and _55357_ (_22713_, _22712_, _21846_);
  not _55358_ (_22714_, _22713_);
  and _55359_ (_22715_, _22714_, _22709_);
  and _55360_ (_22716_, _22715_, _22700_);
  nor _55361_ (_22717_, _22716_, _22695_);
  and _55362_ (_22718_, _22717_, _22547_);
  nor _55363_ (_22719_, _22718_, _22674_);
  and _55364_ (_22720_, _22719_, _22632_);
  nor _55365_ (_22721_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55366_ (_22722_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55367_ (_22723_, _22722_, _22721_);
  and _55368_ (_22724_, _22723_, _21872_);
  nor _55369_ (_22725_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55370_ (_22726_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55371_ (_22727_, _22726_, _22725_);
  and _55372_ (_22728_, _22727_, _21873_);
  nor _55373_ (_22729_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55374_ (_22730_, _21086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55375_ (_22731_, _22730_, _22729_);
  and _55376_ (_22732_, _22731_, _22518_);
  nor _55377_ (_22733_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55378_ (_22734_, _20053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55379_ (_22735_, _22734_, _22733_);
  and _55380_ (_22736_, _22735_, _21846_);
  or _55381_ (_22737_, _22736_, _22732_);
  or _55382_ (_22738_, _22737_, _22728_);
  or _55383_ (_22739_, _22738_, _22724_);
  and _55384_ (_22740_, _22739_, _16527_);
  nor _55385_ (_22741_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55386_ (_22742_, _20465_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55387_ (_22743_, _22742_, _22741_);
  and _55388_ (_22744_, _22743_, _21872_);
  nor _55389_ (_22745_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55390_ (_22746_, _20670_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55391_ (_22747_, _22746_, _22745_);
  and _55392_ (_22748_, _22747_, _21873_);
  nor _55393_ (_22749_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55394_ (_22750_, _20261_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55395_ (_22751_, _22750_, _22749_);
  and _55396_ (_22752_, _22751_, _22518_);
  nor _55397_ (_22753_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55398_ (_22754_, _21119_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55399_ (_22755_, _22754_, _22753_);
  and _55400_ (_22756_, _22755_, _21846_);
  or _55401_ (_22757_, _22756_, _22752_);
  or _55402_ (_22758_, _22757_, _22748_);
  or _55403_ (_22759_, _22758_, _22744_);
  and _55404_ (_22760_, _22759_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55405_ (_22761_, _22760_, _22740_);
  and _55406_ (_22762_, _22761_, _22547_);
  nor _55407_ (_22763_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55408_ (_22764_, _21157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55409_ (_22765_, _22764_, _22763_);
  and _55410_ (_22766_, _22765_, _21872_);
  nor _55411_ (_22767_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55412_ (_22768_, _19859_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55413_ (_22769_, _22768_, _22767_);
  and _55414_ (_22770_, _22769_, _21873_);
  nor _55415_ (_22771_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55416_ (_22772_, _21147_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55417_ (_22773_, _22772_, _22771_);
  and _55418_ (_22774_, _22773_, _22518_);
  nor _55419_ (_22775_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55420_ (_22776_, _20066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55421_ (_22777_, _22776_, _22775_);
  and _55422_ (_22778_, _22777_, _21846_);
  or _55423_ (_22779_, _22778_, _22774_);
  or _55424_ (_22780_, _22779_, _22770_);
  or _55425_ (_22781_, _22780_, _22766_);
  and _55426_ (_22782_, _22781_, _16527_);
  nor _55427_ (_22783_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55428_ (_22784_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55429_ (_22785_, _22784_, _22783_);
  and _55430_ (_22786_, _22785_, _21872_);
  nor _55431_ (_22787_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55432_ (_22788_, _20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55433_ (_22789_, _22788_, _22787_);
  and _55434_ (_22790_, _22789_, _21873_);
  nor _55435_ (_22791_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55436_ (_22792_, _20273_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55437_ (_22793_, _22792_, _22791_);
  and _55438_ (_22794_, _22793_, _22518_);
  nor _55439_ (_22795_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55440_ (_22796_, _21165_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55441_ (_22797_, _22796_, _22795_);
  and _55442_ (_22798_, _22797_, _21846_);
  or _55443_ (_22799_, _22798_, _22794_);
  or _55444_ (_22800_, _22799_, _22790_);
  or _55445_ (_22801_, _22800_, _22786_);
  and _55446_ (_22802_, _22801_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55447_ (_22803_, _22802_, _22782_);
  and _55448_ (_22804_, _22803_, _22547_);
  not _55449_ (_22805_, _22804_);
  and _55450_ (_22806_, _22805_, _22762_);
  and _55451_ (_22807_, _22806_, _22720_);
  or _55452_ (_22808_, \oc8051_symbolic_cxrom1.regvalid [1], _16467_);
  and _55453_ (_22809_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _55454_ (_22810_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55455_ (_22811_, _22810_, _22809_);
  and _55456_ (_22812_, _22811_, _22808_);
  or _55457_ (_22813_, \oc8051_symbolic_cxrom1.regvalid [13], _16467_);
  or _55458_ (_22814_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55459_ (_22815_, _22814_, _22813_);
  and _55460_ (_22816_, _16463_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _55461_ (_22817_, _22816_, _22815_);
  or _55462_ (_22818_, _22817_, _22812_);
  nor _55463_ (_22819_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _55464_ (_22820_, _22819_, _16463_);
  nor _55465_ (_22821_, _22820_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55466_ (_22822_, _22820_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _55467_ (_22823_, _22822_, _22821_);
  and _55468_ (_22824_, _22823_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _55469_ (_22825_, _22819_, _16463_);
  nor _55470_ (_22826_, _22825_, _22820_);
  nand _55471_ (_22827_, \oc8051_symbolic_cxrom1.regvalid [7], _16467_);
  nand _55472_ (_22828_, _22827_, _22826_);
  or _55473_ (_22829_, _22828_, _22824_);
  and _55474_ (_22830_, _22829_, _16459_);
  nand _55475_ (_22831_, _22823_, _21894_);
  or _55476_ (_22832_, _22823_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _55477_ (_22833_, _22832_, _22831_);
  or _55478_ (_22834_, _22826_, _22833_);
  and _55479_ (_22835_, _22834_, _22830_);
  or _55480_ (_22836_, _22835_, _22818_);
  and _55481_ (_22837_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55482_ (_22838_, \oc8051_symbolic_cxrom1.regvalid [0], _16467_);
  or _55483_ (_22839_, _22838_, _22837_);
  and _55484_ (_22840_, _22839_, _16463_);
  and _55485_ (_22841_, \oc8051_symbolic_cxrom1.regvalid [4], _16467_);
  and _55486_ (_22842_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _55487_ (_22843_, _22842_, _22841_);
  and _55488_ (_22844_, _22843_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _55489_ (_22845_, _22844_, _22840_);
  and _55490_ (_22846_, _22845_, _16459_);
  and _55491_ (_22847_, _22809_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _55492_ (_22848_, _22847_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55493_ (_22849_, _22847_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _55494_ (_22850_, _22849_, _22848_);
  or _55495_ (_22851_, _22850_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _55496_ (_22852_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _55497_ (_22853_, _22852_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _55498_ (_22854_, _22853_, _22847_);
  and _55499_ (_22855_, _22854_, _22813_);
  and _55500_ (_22856_, _22855_, _22851_);
  or _55501_ (_22857_, _22850_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _55502_ (_22858_, _22854_);
  nand _55503_ (_22859_, _22850_, _19167_);
  and _55504_ (_22860_, _22859_, _22858_);
  and _55505_ (_22861_, _22860_, _22857_);
  or _55506_ (_22862_, _22861_, _22856_);
  and _55507_ (_22863_, _22862_, _22846_);
  or _55508_ (_22864_, _22850_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _55509_ (_22865_, \oc8051_symbolic_cxrom1.regvalid [15], _16467_);
  and _55510_ (_22866_, _22865_, _22854_);
  and _55511_ (_22867_, _22866_, _22864_);
  or _55512_ (_22868_, _22850_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _55513_ (_22869_, _22850_, _21894_);
  and _55514_ (_22870_, _22869_, _22858_);
  and _55515_ (_22871_, _22870_, _22868_);
  or _55516_ (_22872_, _22871_, _22867_);
  and _55517_ (_22873_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55518_ (_22874_, \oc8051_symbolic_cxrom1.regvalid [6], _16467_);
  or _55519_ (_22875_, _22874_, _16463_);
  or _55520_ (_22876_, _22875_, _22873_);
  or _55521_ (_22877_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _55522_ (_22878_, \oc8051_symbolic_cxrom1.regvalid [10], _16467_);
  and _55523_ (_22879_, _22878_, _22877_);
  or _55524_ (_22880_, _22879_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _55525_ (_22881_, _22880_, _22876_);
  and _55526_ (_22882_, _22881_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _55527_ (_22883_, _22843_, _22816_);
  or _55528_ (_22884_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _55529_ (_22885_, \oc8051_symbolic_cxrom1.regvalid [0], _16467_);
  and _55530_ (_22886_, _22885_, _22809_);
  and _55531_ (_22887_, _22886_, _22884_);
  or _55532_ (_22888_, _22887_, _22883_);
  and _55533_ (_22889_, _22888_, _22882_);
  and _55534_ (_22890_, _22889_, _22872_);
  or _55535_ (_22891_, _22890_, _22863_);
  or _55536_ (_22892_, _22888_, _22881_);
  and _55537_ (_22893_, _22892_, _16455_);
  and _55538_ (_22894_, _22893_, _22891_);
  and _55539_ (_22895_, _22894_, _22836_);
  or _55540_ (_22896_, \oc8051_symbolic_cxrom1.regvalid [2], _16459_);
  or _55541_ (_22897_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _55542_ (_22898_, _22897_, _22896_);
  or _55543_ (_22899_, _22898_, _22823_);
  or _55544_ (_22900_, \oc8051_symbolic_cxrom1.regvalid [10], _16459_);
  or _55545_ (_22901_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _55546_ (_22902_, _22901_, _22900_);
  and _55547_ (_22903_, _22902_, _22823_);
  nor _55548_ (_22904_, _22903_, _22826_);
  and _55549_ (_22905_, _22904_, _22899_);
  and _55550_ (_22906_, _22823_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _55551_ (_22907_, _22841_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _55552_ (_22908_, _22907_, _22906_);
  and _55553_ (_22909_, _22823_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _55554_ (_22910_, _22874_, _16459_);
  or _55555_ (_22911_, _22910_, _22909_);
  and _55556_ (_22912_, _22911_, _22826_);
  and _55557_ (_22913_, _22912_, _22908_);
  or _55558_ (_22914_, _22913_, _22905_);
  or _55559_ (_22915_, _22850_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _55560_ (_22916_, \oc8051_symbolic_cxrom1.regvalid [14], _16467_);
  and _55561_ (_22917_, _22916_, _22915_);
  or _55562_ (_22918_, _22917_, _22858_);
  nand _55563_ (_22919_, _22850_, _19195_);
  or _55564_ (_22920_, _22850_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _55565_ (_22921_, _22920_, _22919_);
  or _55566_ (_22922_, _22921_, _22854_);
  and _55567_ (_22923_, _22922_, _22918_);
  or _55568_ (_22924_, _22923_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _55569_ (_22925_, _22850_, _18931_);
  and _55570_ (_22926_, _22850_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _55571_ (_22927_, _22926_, _22925_);
  and _55572_ (_22928_, _22927_, _22858_);
  or _55573_ (_22929_, _22850_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _55574_ (_22930_, \oc8051_symbolic_cxrom1.regvalid [12], _16467_);
  and _55575_ (_22931_, _22930_, _22854_);
  and _55576_ (_22932_, _22931_, _22929_);
  or _55577_ (_22933_, _22932_, _16459_);
  or _55578_ (_22934_, _22933_, _22928_);
  or _55579_ (_22935_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55580_ (_22936_, _22935_, _22865_);
  or _55581_ (_22937_, _22936_, _16463_);
  or _55582_ (_22938_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _55583_ (_22939_, \oc8051_symbolic_cxrom1.regvalid [11], _16467_);
  and _55584_ (_22940_, _22939_, _22938_);
  or _55585_ (_22941_, _22940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _55586_ (_22942_, _22941_, _22937_);
  and _55587_ (_22943_, _22942_, _22852_);
  and _55588_ (_22944_, _16459_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _55589_ (_22945_, _22815_, _16463_);
  or _55590_ (_22946_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _55591_ (_22947_, \oc8051_symbolic_cxrom1.regvalid [9], _16467_);
  and _55592_ (_22948_, _22947_, _22946_);
  or _55593_ (_22949_, _22948_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _55594_ (_22950_, _22949_, _22945_);
  and _55595_ (_22951_, _22950_, _22944_);
  or _55596_ (_22952_, _22951_, _22943_);
  and _55597_ (_22953_, _22942_, _16459_);
  or _55598_ (_22954_, _22953_, _22818_);
  and _55599_ (_22955_, _22954_, _22952_);
  and _55600_ (_22956_, _22955_, _22934_);
  and _55601_ (_22957_, _22956_, _22924_);
  and _55602_ (_22958_, _22957_, _22914_);
  or _55603_ (_22959_, _22958_, _22895_);
  nor _55604_ (_22960_, _21863_, _16523_);
  and _55605_ (_22961_, _22960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55606_ (_22962_, _22960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55607_ (_22963_, _22962_, _22961_);
  nand _55608_ (_22964_, _22963_, _18879_);
  and _55609_ (_22965_, _21876_, _16519_);
  nor _55610_ (_22966_, _22965_, _22960_);
  and _55611_ (_22967_, _22966_, _22526_);
  and _55612_ (_22968_, _22967_, _22964_);
  not _55613_ (_22969_, _22966_);
  and _55614_ (_22970_, _22963_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _55615_ (_22971_, _22963_, _18865_);
  or _55616_ (_22972_, _22971_, _22970_);
  and _55617_ (_22973_, _22972_, _22969_);
  or _55618_ (_22974_, _22973_, _22968_);
  and _55619_ (_22975_, _22974_, _21863_);
  nand _55620_ (_22976_, _22963_, _18887_);
  nor _55621_ (_22977_, _22969_, _22540_);
  and _55622_ (_22978_, _22977_, _22976_);
  and _55623_ (_22979_, _22963_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _55624_ (_22980_, _22963_, _18894_);
  or _55625_ (_22981_, _22980_, _22979_);
  and _55626_ (_22982_, _22981_, _22969_);
  or _55627_ (_22983_, _22982_, _22978_);
  and _55628_ (_22984_, _22983_, _21888_);
  or _55629_ (_22985_, _22984_, _22975_);
  or _55630_ (_22986_, _22963_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _55631_ (_22987_, _22966_, _22508_);
  and _55632_ (_22988_, _22987_, _22986_);
  and _55633_ (_22989_, _22963_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _55634_ (_22990_, _22963_, _18906_);
  or _55635_ (_22991_, _22990_, _22989_);
  and _55636_ (_22992_, _22991_, _22969_);
  or _55637_ (_22993_, _22992_, _22988_);
  and _55638_ (_22994_, _22993_, _21902_);
  or _55639_ (_22995_, _22963_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _55640_ (_22996_, _22969_, _22502_);
  and _55641_ (_22997_, _22996_, _22995_);
  and _55642_ (_22998_, _22963_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _55643_ (_22999_, _22963_, _18931_);
  or _55644_ (_23000_, _22999_, _22998_);
  and _55645_ (_23001_, _23000_, _22969_);
  or _55646_ (_23002_, _23001_, _22997_);
  and _55647_ (_23003_, _23002_, _21915_);
  or _55648_ (_23004_, _23003_, _22994_);
  or _55649_ (_23005_, _23004_, _22985_);
  nor _55650_ (_23006_, _22516_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _55651_ (_23007_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55652_ (_23008_, \oc8051_symbolic_cxrom1.regvalid [0], _16527_);
  and _55653_ (_23009_, _23008_, _21846_);
  and _55654_ (_23010_, _23009_, _23007_);
  and _55655_ (_23011_, _22504_, _21872_);
  or _55656_ (_23012_, _23011_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _55657_ (_23013_, _23012_, _23010_);
  or _55658_ (_23014_, _23013_, _23006_);
  nor _55659_ (_23015_, _22534_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _55660_ (_23016_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55661_ (_23017_, \oc8051_symbolic_cxrom1.regvalid [1], _16527_);
  and _55662_ (_23018_, _23017_, _21846_);
  and _55663_ (_23019_, _23018_, _23016_);
  and _55664_ (_23020_, _22542_, _21872_);
  or _55665_ (_23021_, _23020_, _16515_);
  or _55666_ (_23022_, _23021_, _23019_);
  or _55667_ (_23023_, _23022_, _23015_);
  and _55668_ (_23024_, _23023_, _23014_);
  and _55669_ (_23025_, pc_log_change, _21842_);
  and _55670_ (_23026_, _23025_, _22547_);
  nand _55671_ (_23027_, _23026_, _23024_);
  nor _55672_ (_23028_, _23027_, _21928_);
  and _55673_ (_23029_, _23028_, _23005_);
  and _55674_ (_23030_, _23029_, _22959_);
  nor _55675_ (_23031_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55676_ (_23032_, _21193_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55677_ (_23033_, _23032_, _23031_);
  and _55678_ (_23034_, _23033_, _21872_);
  nor _55679_ (_23035_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55680_ (_23036_, _19871_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55681_ (_23037_, _23036_, _23035_);
  and _55682_ (_23038_, _23037_, _21873_);
  nor _55683_ (_23039_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55684_ (_23040_, _21203_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55685_ (_23041_, _23040_, _23039_);
  and _55686_ (_23042_, _23041_, _22518_);
  nor _55687_ (_23043_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55688_ (_23044_, _20076_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55689_ (_23045_, _23044_, _23043_);
  and _55690_ (_23046_, _23045_, _21846_);
  or _55691_ (_23047_, _23046_, _23042_);
  or _55692_ (_23048_, _23047_, _23038_);
  or _55693_ (_23049_, _23048_, _23034_);
  and _55694_ (_23050_, _23049_, _16527_);
  nor _55695_ (_23051_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55696_ (_23052_, _20490_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55697_ (_23053_, _23052_, _23051_);
  and _55698_ (_23054_, _23053_, _21872_);
  nor _55699_ (_23055_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55700_ (_23056_, _20694_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55701_ (_23057_, _23056_, _23055_);
  and _55702_ (_23058_, _23057_, _21873_);
  nor _55703_ (_23059_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55704_ (_23060_, _20286_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55705_ (_23061_, _23060_, _23059_);
  and _55706_ (_23062_, _23061_, _22518_);
  nor _55707_ (_23063_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55708_ (_23064_, _21211_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55709_ (_23065_, _23064_, _23063_);
  and _55710_ (_23066_, _23065_, _21846_);
  or _55711_ (_23067_, _23066_, _23062_);
  or _55712_ (_23068_, _23067_, _23058_);
  or _55713_ (_23069_, _23068_, _23054_);
  and _55714_ (_23070_, _23069_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55715_ (_23071_, _23070_, _23050_);
  and _55716_ (_23072_, _23071_, _22547_);
  nor _55717_ (_23073_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55718_ (_23074_, _18740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55719_ (_23075_, _23074_, _23073_);
  and _55720_ (_23076_, _23075_, _22518_);
  nor _55721_ (_23077_, _23076_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _55722_ (_23078_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55723_ (_23079_, _18716_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55724_ (_23080_, _23079_, _23078_);
  and _55725_ (_23081_, _23080_, _21873_);
  not _55726_ (_23082_, _23081_);
  nor _55727_ (_23083_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55728_ (_23084_, _18735_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55729_ (_23085_, _23084_, _23083_);
  and _55730_ (_23086_, _23085_, _21872_);
  nor _55731_ (_23087_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55732_ (_23088_, _18695_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55733_ (_23089_, _23088_, _23087_);
  and _55734_ (_23090_, _23089_, _21846_);
  nor _55735_ (_23091_, _23090_, _23086_);
  and _55736_ (_23092_, _23091_, _23082_);
  and _55737_ (_23093_, _23092_, _23077_);
  nor _55738_ (_23094_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55739_ (_23095_, _18728_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55740_ (_23096_, _23095_, _23094_);
  and _55741_ (_23097_, _23096_, _22518_);
  nor _55742_ (_23098_, _23097_, _16527_);
  nor _55743_ (_23099_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55744_ (_23100_, _18711_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55745_ (_23101_, _23100_, _23099_);
  and _55746_ (_23102_, _23101_, _21873_);
  not _55747_ (_23103_, _23102_);
  nor _55748_ (_23104_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55749_ (_23105_, _18723_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55750_ (_23106_, _23105_, _23104_);
  and _55751_ (_23107_, _23106_, _21872_);
  nor _55752_ (_23108_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _55753_ (_23109_, _18703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _55754_ (_23110_, _23109_, _23108_);
  and _55755_ (_23111_, _23110_, _21846_);
  nor _55756_ (_23112_, _23111_, _23107_);
  and _55757_ (_23113_, _23112_, _23103_);
  and _55758_ (_23114_, _23113_, _23098_);
  nor _55759_ (_23115_, _23114_, _23093_);
  not _55760_ (_23116_, _23115_);
  and _55761_ (_23117_, _23116_, _23072_);
  and _55762_ (_23118_, _23117_, _23030_);
  and _55763_ (_23119_, _23118_, _22807_);
  and _55764_ (property_invalid_jnc, _23119_, _22501_);
  and _55765_ (_23120_, _21861_, _22354_);
  nor _55766_ (_23121_, _22348_, _22354_);
  nor _55767_ (_23122_, _23121_, _23120_);
  nor _55768_ (_23123_, _23122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _55769_ (_23124_, _23122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _55770_ (_23125_, _21969_, _22354_);
  and _55771_ (_23126_, _22356_, cy_reg);
  nor _55772_ (_23127_, _23126_, _23125_);
  nor _55773_ (_23128_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _55774_ (_23129_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _55775_ (_23130_, _21975_, _22354_);
  nor _55776_ (_23131_, _22364_, _22354_);
  nor _55777_ (_23132_, _23131_, _23130_);
  and _55778_ (_23133_, _23132_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _55779_ (_23134_, _23132_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _55780_ (_23135_, _21980_, cy_reg);
  nor _55781_ (_23136_, _22371_, _22354_);
  nor _55782_ (_23137_, _23136_, _23135_);
  nor _55783_ (_23138_, _23137_, _16503_);
  and _55784_ (_23139_, _23137_, _16503_);
  and _55785_ (_23140_, _21985_, _22354_);
  nor _55786_ (_23141_, _22381_, _22354_);
  nor _55787_ (_23142_, _23141_, _23140_);
  and _55788_ (_23143_, _23142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _55789_ (_23144_, _23142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _55790_ (_23145_, _21997_, _22354_);
  nor _55791_ (_23146_, _22389_, _22354_);
  nor _55792_ (_23147_, _23146_, _23145_);
  nor _55793_ (_23148_, _23147_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _55794_ (_23149_, _23147_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _55795_ (_23150_, _22000_, _22354_);
  and _55796_ (_23151_, _22405_, cy_reg);
  nor _55797_ (_23152_, _23151_, _23150_);
  and _55798_ (_23153_, _23152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _55799_ (_23154_, _23152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _55800_ (_23155_, _22007_, cy_reg);
  nor _55801_ (_23156_, _22412_, _22354_);
  nor _55802_ (_23157_, _23156_, _23155_);
  nor _55803_ (_23158_, _23157_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _55804_ (_23159_, _23157_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _55805_ (_23160_, _22051_, _22354_);
  and _55806_ (_23161_, _22421_, cy_reg);
  nor _55807_ (_23162_, _23161_, _23160_);
  nor _55808_ (_23163_, _23162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _55809_ (_23164_, _23162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _55810_ (_23165_, _22096_, _22354_);
  and _55811_ (_23166_, _22427_, cy_reg);
  nor _55812_ (_23167_, _23166_, _23165_);
  nor _55813_ (_23168_, _23167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _55814_ (_23169_, _23167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _55815_ (_23170_, _22140_, _22354_);
  and _55816_ (_23171_, _22435_, cy_reg);
  nor _55817_ (_23172_, _23171_, _23170_);
  nor _55818_ (_23173_, _23172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _55819_ (_23174_, _23172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _55820_ (_23175_, _21868_, cy_reg);
  and _55821_ (_23176_, _22441_, cy_reg);
  nor _55822_ (_23177_, _23176_, _23175_);
  nor _55823_ (_23178_, _23177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55824_ (_23179_, _23177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55825_ (_23180_, _22465_, cy_reg);
  nor _55826_ (_23181_, _21874_, cy_reg);
  nor _55827_ (_23182_, _23181_, _23180_);
  nor _55828_ (_23183_, _23182_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _55829_ (_23184_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _55830_ (_23185_, _22449_, cy_reg);
  nor _55831_ (_23186_, _23185_, _23184_);
  and _55832_ (_23187_, _23186_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _55833_ (_23188_, _22456_, _22301_);
  or _55834_ (_23189_, _23188_, _22458_);
  or _55835_ (_23190_, _23189_, _22354_);
  nand _55836_ (_23191_, _22456_, _22354_);
  and _55837_ (_23192_, _23191_, _23190_);
  nor _55838_ (_23193_, _23186_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _55839_ (_23194_, _23193_, _23192_);
  or _55840_ (_23195_, _23194_, _23187_);
  and _55841_ (_23196_, _23182_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _55842_ (_23197_, _23196_, _23195_);
  or _55843_ (_23198_, _23197_, _23183_);
  or _55844_ (_23199_, _23198_, _23179_);
  or _55845_ (_23200_, _23199_, _23178_);
  or _55846_ (_23201_, _23200_, _23174_);
  or _55847_ (_23202_, _23201_, _23173_);
  or _55848_ (_23203_, _23202_, _23169_);
  or _55849_ (_23204_, _23203_, _23168_);
  or _55850_ (_23205_, _23204_, _23164_);
  or _55851_ (_23206_, _23205_, _23163_);
  or _55852_ (_23207_, _23206_, _23159_);
  or _55853_ (_23208_, _23207_, _23158_);
  or _55854_ (_23209_, _23208_, _23154_);
  or _55855_ (_23210_, _23209_, _23153_);
  or _55856_ (_23211_, _23210_, _23149_);
  or _55857_ (_23212_, _23211_, _23148_);
  and _55858_ (_23213_, _21991_, _22354_);
  and _55859_ (_23214_, _22485_, cy_reg);
  nor _55860_ (_23215_, _23214_, _23213_);
  and _55861_ (_23216_, _23215_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _55862_ (_23217_, _23215_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or _55863_ (_23218_, _23217_, _23216_);
  or _55864_ (_23219_, _23218_, _23212_);
  or _55865_ (_23220_, _23219_, _23144_);
  or _55866_ (_23221_, _23220_, _23143_);
  or _55867_ (_23222_, _23221_, _23139_);
  or _55868_ (_23223_, _23222_, _23138_);
  or _55869_ (_23224_, _23223_, _23134_);
  or _55870_ (_23225_, _23224_, _23133_);
  or _55871_ (_23226_, _23225_, _23129_);
  or _55872_ (_23227_, _23226_, _23128_);
  or _55873_ (_23228_, _23227_, _23124_);
  or _55874_ (_23229_, _23228_, _23123_);
  nor _55875_ (_23230_, _22804_, _22762_);
  and _55876_ (_23231_, _23230_, _22720_);
  and _55877_ (_23232_, _23231_, _23118_);
  and _55878_ (property_invalid_jc, _23232_, _23229_);
  or _55879_ (_23233_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _55880_ (_23234_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _55881_ (_23235_, _23234_, _23233_);
  or _55882_ (_23236_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _55883_ (_23237_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _55884_ (_23238_, _23237_, _23236_);
  or _55885_ (_23239_, _23238_, _23235_);
  nor _55886_ (_23240_, _22301_, _16455_);
  or _55887_ (_23241_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _55888_ (_23242_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _55889_ (_23243_, _23242_, _23241_);
  nor _55890_ (_23244_, _21975_, _16507_);
  and _55891_ (_23245_, _21975_, _16507_);
  or _55892_ (_23246_, _23245_, _23244_);
  or _55893_ (_23247_, _21980_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _55894_ (_23248_, _21980_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _55895_ (_23249_, _23248_, _23247_);
  or _55896_ (_23250_, _23249_, _23246_);
  or _55897_ (_23251_, _21969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _55898_ (_23252_, _21969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _55899_ (_23253_, _23252_, _23251_);
  or _55900_ (_23254_, _23253_, _23250_);
  or _55901_ (_23255_, _23254_, _23243_);
  or _55902_ (_23256_, _23255_, _23240_);
  and _55903_ (_23257_, _22301_, _16455_);
  nor _55904_ (_23258_, _22223_, _16463_);
  or _55905_ (_23259_, _23258_, _23257_);
  or _55906_ (_23260_, _23259_, _23256_);
  or _55907_ (_23261_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _55908_ (_23262_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _55909_ (_23263_, _23262_, _23261_);
  and _55910_ (_23264_, _22804_, _16487_);
  nor _55911_ (_23265_, _22804_, _16487_);
  or _55912_ (_23266_, _23265_, _23264_);
  and _55913_ (_23267_, _23072_, _16491_);
  nor _55914_ (_23268_, _23072_, _16491_);
  or _55915_ (_23269_, _23268_, _23267_);
  or _55916_ (_23270_, _23269_, _23266_);
  nor _55917_ (_23271_, _21985_, _16499_);
  and _55918_ (_23272_, _21985_, _16499_);
  or _55919_ (_23273_, _23272_, _23271_);
  and _55920_ (_23274_, _23115_, _22547_);
  nor _55921_ (_23275_, _23274_, _16495_);
  and _55922_ (_23276_, _23274_, _16495_);
  or _55923_ (_23277_, _23276_, _23275_);
  or _55924_ (_23278_, _23277_, _23273_);
  or _55925_ (_23279_, _23278_, _23270_);
  or _55926_ (_23280_, _23279_, _23263_);
  or _55927_ (_23281_, _23280_, _23260_);
  and _55928_ (_23282_, _22048_, _16479_);
  and _55929_ (_23283_, _21967_, _16483_);
  nor _55930_ (_23284_, _21967_, _16483_);
  or _55931_ (_23285_, _23284_, _23283_);
  or _55932_ (_23286_, _23285_, _23282_);
  and _55933_ (_23287_, _22138_, _16471_);
  nor _55934_ (_23288_, _22048_, _16479_);
  or _55935_ (_23289_, _23288_, _23287_);
  and _55936_ (_23290_, _22223_, _16463_);
  nor _55937_ (_23291_, _22138_, _16471_);
  or _55938_ (_23292_, _23291_, _23290_);
  or _55939_ (_23293_, _23292_, _23289_);
  or _55940_ (_23294_, _23293_, _23286_);
  or _55941_ (_23295_, _23294_, _23281_);
  or _55942_ (_23296_, _23295_, _23239_);
  not _55943_ (_23297_, _22673_);
  and _55944_ (_23298_, _22718_, _22632_);
  and _55945_ (_23299_, _23298_, _23297_);
  and _55946_ (_23300_, _23299_, _23030_);
  and _55947_ (property_invalid_ajmp, _23300_, _23296_);
  and _55948_ (_23301_, _22691_, _21873_);
  and _55949_ (_23302_, _22677_, _21872_);
  or _55950_ (_23303_, _23302_, _23301_);
  and _55951_ (_23304_, _22686_, _22518_);
  and _55952_ (_23305_, _22682_, _21846_);
  or _55953_ (_23306_, _23305_, _23304_);
  or _55954_ (_23307_, _23306_, _23303_);
  and _55955_ (_23308_, _23307_, _22142_);
  and _55956_ (_23309_, _22712_, _21873_);
  and _55957_ (_23310_, _22698_, _21872_);
  or _55958_ (_23311_, _23310_, _23309_);
  and _55959_ (_23312_, _22707_, _22518_);
  and _55960_ (_23313_, _22703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _55961_ (_23314_, _23313_, _23312_);
  or _55962_ (_23315_, _23314_, _23311_);
  and _55963_ (_23316_, _23315_, _21868_);
  or _55964_ (_23317_, _23316_, _23308_);
  and _55965_ (_23318_, _23317_, _23024_);
  and _55966_ (_23319_, _23318_, _16455_);
  nor _55967_ (_23320_, _23318_, _16455_);
  or _55968_ (_23321_, _23320_, _23319_);
  and _55969_ (_23322_, _22647_, _21873_);
  or _55970_ (_23323_, _23322_, _22142_);
  and _55971_ (_23324_, _22643_, _21846_);
  and _55972_ (_23325_, _22635_, _22518_);
  and _55973_ (_23326_, _22639_, _21872_);
  or _55974_ (_23327_, _23326_, _23325_);
  or _55975_ (_23328_, _23327_, _23324_);
  or _55976_ (_23329_, _23328_, _23323_);
  and _55977_ (_23330_, _22663_, _21846_);
  or _55978_ (_23331_, _23330_, _21868_);
  and _55979_ (_23332_, _22659_, _21872_);
  and _55980_ (_23333_, _22655_, _22518_);
  and _55981_ (_23334_, _22667_, _21873_);
  or _55982_ (_23335_, _23334_, _23333_);
  or _55983_ (_23336_, _23335_, _23332_);
  or _55984_ (_23337_, _23336_, _23331_);
  and _55985_ (_23338_, _23337_, _23329_);
  and _55986_ (_23339_, _23338_, _23024_);
  nor _55987_ (_23340_, _23339_, _16459_);
  and _55988_ (_23341_, _23339_, _16459_);
  or _55989_ (_23342_, _23341_, _23340_);
  or _55990_ (_23343_, _23342_, _23321_);
  and _55991_ (_23344_, _22562_, _21873_);
  or _55992_ (_23345_, _23344_, _22142_);
  and _55993_ (_23346_, _22558_, _21846_);
  and _55994_ (_23347_, _22550_, _22518_);
  and _55995_ (_23348_, _22554_, _21872_);
  or _55996_ (_23349_, _23348_, _23347_);
  or _55997_ (_23350_, _23349_, _23346_);
  or _55998_ (_23351_, _23350_, _23345_);
  and _55999_ (_23352_, _22578_, _21846_);
  or _56000_ (_23353_, _23352_, _21868_);
  and _56001_ (_23354_, _22574_, _21872_);
  and _56002_ (_23355_, _22570_, _22518_);
  and _56003_ (_23356_, _22582_, _21873_);
  or _56004_ (_23357_, _23356_, _23355_);
  or _56005_ (_23358_, _23357_, _23354_);
  or _56006_ (_23359_, _23358_, _23353_);
  and _56007_ (_23360_, _23359_, _23351_);
  and _56008_ (_23361_, _23360_, _23024_);
  nand _56009_ (_23362_, _23361_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _56010_ (_23363_, _23361_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _56011_ (_23364_, _23363_, _23362_);
  and _56012_ (_23365_, _22604_, _21873_);
  or _56013_ (_23366_, _23365_, _22142_);
  and _56014_ (_23367_, _22600_, _21846_);
  and _56015_ (_23368_, _22592_, _22518_);
  and _56016_ (_23369_, _22596_, _21872_);
  or _56017_ (_23370_, _23369_, _23368_);
  or _56018_ (_23371_, _23370_, _23367_);
  or _56019_ (_23372_, _23371_, _23366_);
  and _56020_ (_23373_, _22620_, _21846_);
  or _56021_ (_23374_, _23373_, _21868_);
  and _56022_ (_23375_, _22616_, _21872_);
  and _56023_ (_23376_, _22612_, _22518_);
  and _56024_ (_23377_, _22624_, _21873_);
  or _56025_ (_23378_, _23377_, _23376_);
  or _56026_ (_23379_, _23378_, _23375_);
  or _56027_ (_23380_, _23379_, _23374_);
  and _56028_ (_23381_, _23380_, _23372_);
  and _56029_ (_23382_, _23381_, _23024_);
  nand _56030_ (_23383_, _23382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _56031_ (_23384_, _23382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _56032_ (_23385_, _23384_, _23383_);
  or _56033_ (_23386_, _23385_, _23364_);
  or _56034_ (_23387_, _23386_, _23343_);
  and _56035_ (_23388_, _22727_, _21872_);
  or _56036_ (_23389_, _23388_, _22142_);
  and _56037_ (_23390_, _22723_, _22518_);
  and _56038_ (_23391_, _22731_, _21846_);
  or _56039_ (_23392_, _23391_, _23390_);
  and _56040_ (_23393_, _22735_, _21873_);
  or _56041_ (_23394_, _23393_, _23392_);
  or _56042_ (_23395_, _23394_, _23389_);
  and _56043_ (_23396_, _22751_, _21846_);
  or _56044_ (_23397_, _23396_, _21868_);
  and _56045_ (_23398_, _22747_, _21872_);
  and _56046_ (_23399_, _22743_, _22518_);
  and _56047_ (_23400_, _22755_, _21873_);
  or _56048_ (_23401_, _23400_, _23399_);
  or _56049_ (_23402_, _23401_, _23398_);
  or _56050_ (_23403_, _23402_, _23397_);
  and _56051_ (_23404_, _23403_, _23395_);
  and _56052_ (_23405_, _23404_, _23024_);
  or _56053_ (_23406_, _23405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _56054_ (_23407_, _23405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _56055_ (_23408_, _23407_, _23406_);
  and _56056_ (_23409_, _22789_, _21872_);
  or _56057_ (_23410_, _23409_, _21868_);
  and _56058_ (_23411_, _22785_, _22518_);
  and _56059_ (_23412_, _22793_, _21846_);
  or _56060_ (_23413_, _23412_, _23411_);
  and _56061_ (_23414_, _22797_, _21873_);
  or _56062_ (_23415_, _23414_, _23413_);
  or _56063_ (_23416_, _23415_, _23410_);
  and _56064_ (_23417_, _22773_, _21846_);
  or _56065_ (_23418_, _23417_, _22142_);
  and _56066_ (_23419_, _22769_, _21872_);
  and _56067_ (_23420_, _22765_, _22518_);
  and _56068_ (_23421_, _22777_, _21873_);
  or _56069_ (_23422_, _23421_, _23420_);
  or _56070_ (_23423_, _23422_, _23419_);
  or _56071_ (_23424_, _23423_, _23418_);
  and _56072_ (_23425_, _23424_, _23416_);
  and _56073_ (_23426_, _23425_, _23024_);
  nor _56074_ (_23427_, _23426_, _16475_);
  and _56075_ (_23428_, _23426_, _16475_);
  or _56076_ (_23429_, _23428_, _23427_);
  or _56077_ (_23430_, _23429_, _23408_);
  and _56078_ (_23431_, _23080_, _21872_);
  or _56079_ (_23432_, _23431_, _22142_);
  and _56080_ (_23433_, _23075_, _21846_);
  and _56081_ (_23434_, _23085_, _22518_);
  or _56082_ (_23435_, _23434_, _23433_);
  and _56083_ (_23436_, _23089_, _21873_);
  or _56084_ (_23437_, _23436_, _23435_);
  or _56085_ (_23438_, _23437_, _23432_);
  and _56086_ (_23439_, _23101_, _21872_);
  or _56087_ (_23440_, _23439_, _21868_);
  and _56088_ (_23441_, _23096_, _21846_);
  and _56089_ (_23442_, _23106_, _22518_);
  and _56090_ (_23443_, _23110_, _21873_);
  or _56091_ (_23444_, _23443_, _23442_);
  or _56092_ (_23445_, _23444_, _23441_);
  or _56093_ (_23446_, _23445_, _23440_);
  and _56094_ (_23447_, _23446_, _23438_);
  and _56095_ (_23448_, _23447_, _23024_);
  nand _56096_ (_23449_, _23448_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _56097_ (_23450_, _23448_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _56098_ (_23451_, _23450_, _23449_);
  and _56099_ (_23452_, _23045_, _21873_);
  or _56100_ (_23453_, _23452_, _22142_);
  and _56101_ (_23454_, _23041_, _21846_);
  and _56102_ (_23455_, _23033_, _22518_);
  and _56103_ (_23456_, _23037_, _21872_);
  or _56104_ (_23457_, _23456_, _23455_);
  or _56105_ (_23458_, _23457_, _23454_);
  or _56106_ (_23459_, _23458_, _23453_);
  and _56107_ (_23460_, _23061_, _21846_);
  or _56108_ (_23461_, _23460_, _21868_);
  and _56109_ (_23462_, _23057_, _21872_);
  and _56110_ (_23463_, _23053_, _22518_);
  and _56111_ (_23464_, _23065_, _21873_);
  or _56112_ (_23465_, _23464_, _23463_);
  or _56113_ (_23466_, _23465_, _23462_);
  or _56114_ (_23467_, _23466_, _23461_);
  and _56115_ (_23468_, _23467_, _23459_);
  and _56116_ (_23469_, _23468_, _23024_);
  nor _56117_ (_23470_, _23469_, _16479_);
  and _56118_ (_23471_, _23469_, _16479_);
  or _56119_ (_23472_, _23471_, _23470_);
  or _56120_ (_23473_, _23472_, _23451_);
  or _56121_ (_23474_, _23473_, _23430_);
  or _56122_ (_23475_, _23474_, _23387_);
  or _56123_ (_23476_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _56124_ (_23477_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _56125_ (_23478_, _23477_, _23476_);
  and _56126_ (_23479_, _22301_, _16487_);
  nor _56127_ (_23480_, _22301_, _16487_);
  or _56128_ (_23481_, _23480_, _23479_);
  or _56129_ (_23482_, _23481_, _23478_);
  or _56130_ (_23483_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _56131_ (_23484_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _56132_ (_23485_, _23484_, _23483_);
  nor _56133_ (_23486_, _22223_, _16495_);
  and _56134_ (_23487_, _22223_, _16495_);
  or _56135_ (_23488_, _23487_, _23486_);
  or _56136_ (_23489_, _23488_, _23485_);
  or _56137_ (_23490_, _23489_, _23482_);
  or _56138_ (_23491_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _56139_ (_23492_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _56140_ (_23493_, _23492_, _23491_);
  nor _56141_ (_23494_, _22138_, _16503_);
  and _56142_ (_23495_, _22138_, _16503_);
  or _56143_ (_23496_, _23495_, _23494_);
  or _56144_ (_23497_, _23496_, _23493_);
  nor _56145_ (_23498_, _21967_, _15859_);
  and _56146_ (_23499_, _21967_, _15859_);
  or _56147_ (_23500_, _23499_, _23498_);
  and _56148_ (_23501_, _22048_, _16511_);
  nor _56149_ (_23502_, _22048_, _16511_);
  or _56150_ (_23503_, _23502_, _23501_);
  or _56151_ (_23504_, _23503_, _23500_);
  or _56152_ (_23505_, _23504_, _23497_);
  or _56153_ (_23506_, _23505_, _23490_);
  or _56154_ (_23507_, _23506_, _23475_);
  nor _56155_ (_23508_, _23274_, _23072_);
  not _56156_ (_23509_, _22718_);
  and _56157_ (_23510_, _23509_, _22632_);
  and _56158_ (_23511_, _22805_, _23510_);
  and _56159_ (_23512_, _23511_, _22674_);
  and _56160_ (_23513_, _23512_, _23508_);
  and _56161_ (_23514_, _23513_, _23030_);
  and _56162_ (property_invalid_ljmp, _23514_, _23507_);
  and _56163_ (_23515_, _22348_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _56164_ (_23516_, _22348_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or _56165_ (_23517_, _22356_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _56166_ (_23518_, _22356_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _56167_ (_23519_, _23518_, _23517_);
  or _56168_ (_23520_, _22364_, _16507_);
  nand _56169_ (_23521_, _22364_, _16507_);
  and _56170_ (_23522_, _23521_, _23520_);
  or _56171_ (_23523_, _22371_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _56172_ (_23524_, _22371_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _56173_ (_23525_, _23524_, _23523_);
  and _56174_ (_23526_, _22381_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _56175_ (_23527_, _22381_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _56176_ (_23528_, _22389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _56177_ (_23529_, _22389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _56178_ (_23531_, _22421_, _16479_);
  nor _56179_ (_23532_, _22421_, _16479_);
  nor _56180_ (_23533_, _22427_, _16475_);
  and _56181_ (_23534_, _22427_, _16475_);
  and _56182_ (_23535_, _22435_, _16471_);
  nor _56183_ (_23536_, _22435_, _16471_);
  and _56184_ (_23537_, _22441_, _16467_);
  nor _56185_ (_23538_, _22441_, _16467_);
  and _56186_ (_23539_, _22465_, _16463_);
  or _56187_ (_23540_, _22449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56188_ (_23541_, _22449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _56189_ (_23542_, _23541_, _23540_);
  or _56190_ (_23543_, _23542_, _23189_);
  nor _56191_ (_23544_, _22465_, _16463_);
  or _56192_ (_23545_, _23544_, _23543_);
  or _56193_ (_23546_, _23545_, _23539_);
  or _56194_ (_23547_, _23546_, _23538_);
  or _56195_ (_23548_, _23547_, _23537_);
  or _56196_ (_23549_, _23548_, _23536_);
  or _56197_ (_23550_, _23549_, _23535_);
  or _56198_ (_23551_, _23550_, _23534_);
  or _56199_ (_23552_, _23551_, _23533_);
  or _56200_ (_23553_, _23552_, _23532_);
  or _56201_ (_23554_, _23553_, _23531_);
  or _56202_ (_23555_, _23554_, _22415_);
  or _56203_ (_23556_, _23555_, _22408_);
  or _56204_ (_23557_, _23556_, _23529_);
  or _56205_ (_23558_, _23557_, _23528_);
  nor _56206_ (_23559_, _22485_, _16495_);
  and _56207_ (_23560_, _22485_, _16495_);
  or _56208_ (_23561_, _23560_, _23559_);
  or _56209_ (_23562_, _23561_, _23558_);
  or _56210_ (_23563_, _23562_, _23527_);
  or _56211_ (_23564_, _23563_, _23526_);
  or _56212_ (_23565_, _23564_, _23525_);
  or _56213_ (_23566_, _23565_, _23522_);
  or _56214_ (_23567_, _23566_, _23519_);
  or _56215_ (_23568_, _23567_, _23516_);
  or _56216_ (_23569_, _23568_, _23515_);
  not _56217_ (_23570_, _23072_);
  and _56218_ (_23571_, _23274_, _23570_);
  and _56219_ (_23572_, _23571_, _23230_);
  and _56220_ (_23573_, _23572_, _22720_);
  and _56221_ (_23574_, _23573_, _23030_);
  and _56222_ (property_invalid_sjmp, _23574_, _23569_);
  and _56223_ (_23575_, _22961_, _21850_);
  and _56224_ (_23576_, _23575_, _21854_);
  and _56225_ (_23577_, _23576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _56226_ (_23578_, _23577_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _56227_ (_23579_, _23578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _56228_ (_23580_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _56229_ (_23581_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _56230_ (_23582_, _23581_, _23580_);
  not _56231_ (_23583_, _23582_);
  nor _56232_ (_23584_, _23583_, _23579_);
  and _56233_ (_23585_, _23583_, _23579_);
  not _56234_ (_23586_, _23577_);
  nor _56235_ (_23587_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _56236_ (_23588_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _56237_ (_23589_, _23588_, _23587_);
  nor _56238_ (_23590_, _23589_, _23586_);
  and _56239_ (_23591_, _23575_, _21852_);
  and _56240_ (_23592_, _23575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _56241_ (_23593_, _23592_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _56242_ (_23594_, _23593_, _23591_);
  and _56243_ (_23595_, _23594_, _16491_);
  and _56244_ (_23596_, _22961_, _21849_);
  and _56245_ (_23597_, _22961_, _21848_);
  nor _56246_ (_23598_, _23597_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _56247_ (_23599_, _23598_, _23596_);
  nor _56248_ (_23600_, _23599_, _16479_);
  or _56249_ (_23601_, _23600_, _23595_);
  nor _56250_ (_23602_, _23594_, _16491_);
  and _56251_ (_23603_, _23599_, _16479_);
  or _56252_ (_23604_, _23603_, _23602_);
  or _56253_ (_23605_, _23604_, _23601_);
  or _56254_ (_23606_, _23605_, _23590_);
  nor _56255_ (_23607_, _23596_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _56256_ (_23608_, _23607_, _23575_);
  nand _56257_ (_23609_, _23608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _56258_ (_23610_, _23608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _56259_ (_23611_, _23610_, _23609_);
  and _56260_ (_23612_, _23589_, _23586_);
  or _56261_ (_23613_, _23612_, _23611_);
  or _56262_ (_23614_, _23613_, _23606_);
  or _56263_ (_23615_, _23614_, _23585_);
  or _56264_ (_23616_, _23615_, _23584_);
  nor _56265_ (_23617_, _23578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _56266_ (_23618_, _23617_, _23579_);
  and _56267_ (_23619_, _23618_, _16511_);
  nor _56268_ (_23620_, _23618_, _16511_);
  nor _56269_ (_23621_, _23576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _56270_ (_23622_, _23621_, _23577_);
  and _56271_ (_23623_, _23622_, _16503_);
  nor _56272_ (_23624_, _23622_, _16503_);
  and _56273_ (_23625_, _23575_, _21853_);
  nor _56274_ (_23626_, _23591_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _56275_ (_23627_, _23626_, _23625_);
  and _56276_ (_23628_, _23627_, _16495_);
  and _56277_ (_23629_, _22961_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _56278_ (_23630_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _56279_ (_23631_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _56280_ (_23632_, _23631_, _23630_);
  not _56281_ (_23633_, _23632_);
  nor _56282_ (_23634_, _23633_, _23629_);
  and _56283_ (_23635_, _22963_, _16467_);
  and _56284_ (_23636_, _23633_, _23629_);
  or _56285_ (_23637_, _23636_, _23635_);
  or _56286_ (_23638_, _23637_, _23634_);
  and _56287_ (_23639_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _56288_ (_23640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _56289_ (_23641_, _23640_, _23639_);
  nand _56290_ (_23642_, _23641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _56291_ (_23643_, _23641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _56292_ (_23644_, _23643_, _23642_);
  nand _56293_ (_23645_, _22966_, _16463_);
  nand _56294_ (_23646_, _23645_, _23644_);
  nor _56295_ (_23647_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _56296_ (_23648_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _56297_ (_23649_, _23648_, _23647_);
  not _56298_ (_23650_, _23649_);
  nor _56299_ (_23651_, _23650_, _22961_);
  nor _56300_ (_23652_, _22966_, _16463_);
  or _56301_ (_23653_, _23652_, _23651_);
  or _56302_ (_23654_, _23653_, _23646_);
  nor _56303_ (_23655_, _22963_, _16467_);
  and _56304_ (_23656_, _23650_, _22961_);
  or _56305_ (_23657_, _23656_, _22456_);
  or _56306_ (_23658_, _23657_, _23655_);
  or _56307_ (_23659_, _23658_, _23654_);
  or _56308_ (_23660_, _23659_, _23638_);
  nor _56309_ (_23661_, _23575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _56310_ (_23662_, _23661_, _23592_);
  nor _56311_ (_23663_, _23662_, _16487_);
  and _56312_ (_23664_, _23662_, _16487_);
  or _56313_ (_23665_, _23664_, _23663_);
  or _56314_ (_23666_, _23665_, _23660_);
  or _56315_ (_23667_, _23666_, _23628_);
  nor _56316_ (_23668_, _23627_, _16495_);
  nor _56317_ (_23669_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _56318_ (_23670_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _56319_ (_23671_, _23670_, _23669_);
  or _56320_ (_23672_, _23671_, _23625_);
  nand _56321_ (_23673_, _23671_, _23625_);
  and _56322_ (_23674_, _23673_, _23672_);
  or _56323_ (_23675_, _23674_, _23668_);
  or _56324_ (_23676_, _23675_, _23667_);
  or _56325_ (_23677_, _23676_, _23624_);
  or _56326_ (_23678_, _23677_, _23623_);
  or _56327_ (_23679_, _23678_, _23620_);
  or _56328_ (_23680_, _23679_, _23619_);
  or _56329_ (_23681_, _23680_, _23616_);
  not _56330_ (_23682_, _22762_);
  nor _56331_ (_23683_, _22673_, _22588_);
  and _56332_ (_23684_, _23683_, _22631_);
  and _56333_ (_23685_, _23684_, _22718_);
  and _56334_ (_23686_, _23685_, _23682_);
  and _56335_ (_23687_, _23686_, _22805_);
  or _56336_ (_23688_, _23687_, _22807_);
  and _56337_ (_23689_, _23688_, _23571_);
  and _56338_ (_23690_, _23685_, _22804_);
  and _56339_ (_23691_, _23690_, _22762_);
  and _56340_ (_23692_, _23298_, _22673_);
  nand _56341_ (_23693_, _22804_, _22761_);
  and _56342_ (_23694_, _23693_, _23692_);
  or _56343_ (_23695_, _23694_, _23691_);
  and _56344_ (_23696_, _23695_, _23117_);
  or _56345_ (_23697_, _23696_, _23689_);
  and _56346_ (_23698_, _23697_, _23030_);
  and _56347_ (property_invalid_pcp3, _23698_, _23681_);
  not _56348_ (_23699_, _22717_);
  and _56349_ (_23700_, _23684_, _23699_);
  and _56350_ (_23701_, _22674_, _22631_);
  and _56351_ (_23702_, _23701_, _22762_);
  and _56352_ (_23703_, _23702_, _22804_);
  or _56353_ (_23704_, _23703_, _23700_);
  and _56354_ (_23705_, _23704_, _23116_);
  or _56355_ (_23706_, _23705_, _23686_);
  and _56356_ (_23707_, _23706_, _23072_);
  or _56357_ (_23708_, _23512_, _23072_);
  or _56358_ (_23709_, _23690_, _23511_);
  and _56359_ (_23710_, _23709_, _23274_);
  and _56360_ (_23711_, _23710_, _23708_);
  and _56361_ (_23712_, _23684_, _22806_);
  not _56362_ (_23713_, _22761_);
  or _56363_ (_23714_, _23701_, _22589_);
  and _56364_ (_23715_, _23714_, _23713_);
  or _56365_ (_23716_, _23715_, _23712_);
  and _56366_ (_23717_, _23716_, _23571_);
  not _56367_ (_23718_, _23274_);
  and _56368_ (_23719_, _23685_, _22805_);
  and _56369_ (_23720_, _23071_, _22588_);
  and _56370_ (_23721_, _23720_, _22804_);
  and _56371_ (_23722_, _23721_, _22761_);
  or _56372_ (_23723_, _23722_, _23719_);
  and _56373_ (_23724_, _23723_, _23718_);
  and _56374_ (_23725_, _23571_, _22803_);
  and _56375_ (_23726_, _23117_, _22674_);
  or _56376_ (_23727_, _23726_, _23725_);
  and _56377_ (_23728_, _23727_, _23510_);
  and _56378_ (_23729_, _23508_, _22804_);
  and _56379_ (_23730_, _23729_, _23684_);
  or _56380_ (_23731_, _23730_, _23728_);
  or _56381_ (_23732_, _23731_, _23724_);
  or _56382_ (_23733_, _23732_, _23717_);
  or _56383_ (_23734_, _23733_, _23711_);
  or _56384_ (_23735_, _23734_, _23707_);
  and _56385_ (_23736_, _21997_, _16491_);
  or _56386_ (_23737_, _22051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _56387_ (_23738_, _22051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _56388_ (_23739_, _23738_, _23737_);
  nor _56389_ (_23740_, _21997_, _16491_);
  or _56390_ (_23741_, _23740_, _23739_);
  or _56391_ (_23742_, _23741_, _23736_);
  and _56392_ (_23743_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _56393_ (_23744_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _56394_ (_23745_, _23744_, _23743_);
  or _56395_ (_23746_, _23649_, _21847_);
  nand _56396_ (_23747_, _23649_, _21847_);
  and _56397_ (_23748_, _23747_, _23746_);
  nand _56398_ (_23749_, _23641_, _22456_);
  or _56399_ (_23750_, _23749_, _23748_);
  or _56400_ (_23751_, _23750_, _23745_);
  or _56401_ (_23752_, _23632_, _22094_);
  nand _56402_ (_23753_, _23632_, _22094_);
  and _56403_ (_23754_, _23753_, _23752_);
  or _56404_ (_23755_, _21868_, _16467_);
  nand _56405_ (_23756_, _21868_, _16467_);
  and _56406_ (_23757_, _23756_, _23755_);
  or _56407_ (_23758_, _23757_, _23754_);
  or _56408_ (_23759_, _23758_, _23751_);
  or _56409_ (_23760_, _23759_, _22401_);
  or _56410_ (_23761_, _23760_, _22398_);
  or _56411_ (_23762_, _23761_, _23273_);
  nor _56412_ (_23763_, _21991_, _16495_);
  and _56413_ (_23764_, _21991_, _16495_);
  or _56414_ (_23765_, _23764_, _23763_);
  or _56415_ (_23766_, _23765_, _23762_);
  or _56416_ (_23767_, _23766_, _23742_);
  or _56417_ (_23768_, _23767_, _23255_);
  and _56418_ (_23769_, _23768_, _23030_);
  and _56419_ (property_invalid_pcp2, _23769_, _23735_);
  and _56420_ (_23770_, _22806_, _22588_);
  and _56421_ (_23771_, _23230_, _22719_);
  and _56422_ (_23772_, _23699_, _22631_);
  and _56423_ (_23773_, _23772_, _22805_);
  or _56424_ (_23774_, _23773_, _23771_);
  and _56425_ (_23775_, _23774_, _23718_);
  and _56426_ (_23776_, _23700_, _23230_);
  or _56427_ (_23777_, _23776_, _23692_);
  or _56428_ (_23778_, _23777_, _23775_);
  or _56429_ (_23779_, _23778_, _23770_);
  and _56430_ (_23780_, _23779_, _23570_);
  and _56431_ (_23781_, _23115_, _23699_);
  and _56432_ (_23782_, _23781_, _22804_);
  or _56433_ (_23783_, _23782_, _23715_);
  and _56434_ (_23784_, _22718_, _22674_);
  or _56435_ (_23785_, _23772_, _23784_);
  nor _56436_ (_23786_, _23116_, _22589_);
  and _56437_ (_23787_, _23786_, _23785_);
  or _56438_ (_23788_, _23787_, _23783_);
  and _56439_ (_23789_, _23788_, _23072_);
  and _56440_ (_23790_, _23684_, _23682_);
  and _56441_ (_23791_, _23725_, _23790_);
  nor _56442_ (_23792_, _23115_, _22803_);
  and _56443_ (_23793_, _23792_, _22589_);
  and _56444_ (_23794_, _23721_, _23274_);
  or _56445_ (_23795_, _23794_, _23793_);
  or _56446_ (_23796_, _23795_, _23791_);
  nor _56447_ (_23797_, _22804_, _22589_);
  and _56448_ (_23798_, _23797_, _23702_);
  and _56449_ (_23799_, _23714_, _23508_);
  or _56450_ (_23800_, _23799_, _23798_);
  or _56451_ (_23801_, _23800_, _23796_);
  or _56452_ (_23802_, _23801_, _23789_);
  or _56453_ (_23803_, _23802_, _23780_);
  and _56454_ (_23804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _16515_);
  and _56455_ (_23805_, _21975_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _56456_ (_23806_, _23805_, _23804_);
  nor _56457_ (_23807_, _23806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _56458_ (_23808_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _56459_ (_23809_, _23808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _56460_ (_23810_, _23808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _56461_ (_23811_, _23810_, _23809_);
  and _56462_ (_23812_, _23811_, _16511_);
  and _56463_ (_23813_, _23806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or _56464_ (_23814_, _23813_, _23812_);
  or _56465_ (_23815_, _23814_, _23807_);
  or _56466_ (_23816_, _16547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _56467_ (_23817_, _21997_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _56468_ (_23818_, _23817_, _23816_);
  and _56469_ (_23819_, _23818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _56470_ (_23820_, _23818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _56471_ (_23821_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _56472_ (_23822_, _23821_, _21850_);
  and _56473_ (_23823_, _23822_, _21853_);
  or _56474_ (_23824_, _23823_, _23671_);
  nand _56475_ (_23825_, _23823_, _23671_);
  and _56476_ (_23826_, _23825_, _23824_);
  nor _56477_ (_23827_, _21877_, _16463_);
  and _56478_ (_23828_, _21877_, _16463_);
  or _56479_ (_23829_, _23828_, _23827_);
  not _56480_ (_23830_, _23822_);
  nor _56481_ (_23831_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _56482_ (_23832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _56483_ (_23833_, _23832_, _23831_);
  nor _56484_ (_23834_, _23833_, _23830_);
  and _56485_ (_23835_, _23833_, _23830_);
  or _56486_ (_23836_, _23835_, _23834_);
  or _56487_ (_23837_, _23836_, _23829_);
  and _56488_ (_23838_, _22004_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _56489_ (_23839_, _23838_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _56490_ (_23840_, _23839_, _23822_);
  and _56491_ (_23841_, _23840_, _16483_);
  nor _56492_ (_23842_, _23821_, _23650_);
  and _56493_ (_23843_, _23821_, _23650_);
  or _56494_ (_23844_, _23843_, _22456_);
  or _56495_ (_23845_, _23844_, _23842_);
  or _56496_ (_23846_, _23845_, _23644_);
  or _56497_ (_23847_, _23846_, _23841_);
  or _56498_ (_23848_, _23847_, _23837_);
  or _56499_ (_23849_, _23848_, _23826_);
  not _56500_ (_23850_, _22050_);
  nor _56501_ (_23851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _56502_ (_23852_, _23851_, _23838_);
  and _56503_ (_23853_, _23852_, _23850_);
  or _56504_ (_23854_, _23853_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _56505_ (_23855_, _23853_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _56506_ (_23856_, _23855_, _23854_);
  nor _56507_ (_23857_, _23840_, _16483_);
  nor _56508_ (_23858_, _21870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _56509_ (_23859_, _21870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _56510_ (_23860_, _23859_, _23858_);
  or _56511_ (_23861_, _23860_, _23857_);
  or _56512_ (_23862_, _23861_, _23856_);
  or _56513_ (_23863_, _23862_, _23849_);
  or _56514_ (_23864_, _23863_, _23820_);
  or _56515_ (_23865_, _23864_, _23819_);
  nor _56516_ (_23866_, _23811_, _16511_);
  and _56517_ (_23867_, _23822_, _21854_);
  and _56518_ (_23868_, _23867_, _16558_);
  nor _56519_ (_23869_, _23867_, _16558_);
  or _56520_ (_23870_, _23869_, _23868_);
  nand _56521_ (_23871_, _23870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or _56522_ (_23872_, _23870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _56523_ (_23873_, _23872_, _23871_);
  and _56524_ (_23874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _16515_);
  and _56525_ (_23875_, _22096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _56526_ (_23876_, _23875_, _23874_);
  or _56527_ (_23877_, _23876_, _16475_);
  nand _56528_ (_23878_, _23876_, _16475_);
  and _56529_ (_23879_, _23878_, _23877_);
  or _56530_ (_23880_, _23879_, _23873_);
  nor _56531_ (_23881_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _56532_ (_23882_, _23881_, _23823_);
  nor _56533_ (_23883_, _23882_, _21990_);
  nor _56534_ (_23884_, _23883_, _16495_);
  and _56535_ (_23885_, _23883_, _16495_);
  or _56536_ (_23886_, _23885_, _23884_);
  or _56537_ (_23887_, _23886_, _23880_);
  or _56538_ (_23888_, _23887_, _23866_);
  or _56539_ (_23889_, _23888_, _23865_);
  nor _56540_ (_23890_, _23809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _56541_ (_23891_, _23809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _56542_ (_23892_, _23891_, _23890_);
  and _56543_ (_23893_, _23892_, _15859_);
  nor _56544_ (_23894_, _23892_, _15859_);
  or _56545_ (_23895_, _23894_, _23893_);
  or _56546_ (_23896_, _23895_, _23889_);
  or _56547_ (_23897_, _23896_, _23815_);
  and _56548_ (_23898_, _23897_, _23030_);
  and _56549_ (property_invalid_pcp1, _23898_, _23803_);
  buf _56550_ (_00587_, _27357_);
  buf _56551_ (_02706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7]);
  buf _56552_ (_10034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0]);
  buf _56553_ (_10038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1]);
  buf _56554_ (_10042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2]);
  buf _56555_ (_10046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3]);
  buf _56556_ (_10050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4]);
  buf _56557_ (_10054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5]);
  buf _56558_ (_10058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6]);
  buf _56559_ (_24407_, _24307_);
  buf _56560_ (_24409_, _24308_);
  buf _56561_ (_24421_, _24307_);
  buf _56562_ (_24422_, _24308_);
  buf _56563_ (_24739_, _24328_);
  buf _56564_ (_24740_, _24329_);
  buf _56565_ (_24741_, _24330_);
  buf _56566_ (_24743_, _24331_);
  buf _56567_ (_24744_, _24333_);
  buf _56568_ (_24745_, _24334_);
  buf _56569_ (_24746_, _24335_);
  buf _56570_ (_24747_, _24336_);
  buf _56571_ (_24748_, _24337_);
  buf _56572_ (_24749_, _24339_);
  buf _56573_ (_24750_, _24340_);
  buf _56574_ (_24751_, _24341_);
  buf _56575_ (_24752_, _24342_);
  buf _56576_ (_24754_, _24343_);
  buf _56577_ (_24805_, _24328_);
  buf _56578_ (_24806_, _24329_);
  buf _56579_ (_24807_, _24330_);
  buf _56580_ (_24809_, _24331_);
  buf _56581_ (_24810_, _24333_);
  buf _56582_ (_24811_, _24334_);
  buf _56583_ (_24812_, _24335_);
  buf _56584_ (_24813_, _24336_);
  buf _56585_ (_24814_, _24337_);
  buf _56586_ (_24815_, _24339_);
  buf _56587_ (_24816_, _24340_);
  buf _56588_ (_24817_, _24341_);
  buf _56589_ (_24818_, _24342_);
  buf _56590_ (_24820_, _24343_);
  buf _56591_ (_25393_, _25154_);
  buf _56592_ (_25569_, _25154_);
  dff _56593_ (cy_reg, _00000_, clk);
  dff _56594_ (pc_log_change_r, pc_log_change, clk);
  dff _56595_ (first_instr, _00001_, clk);
  dff _56596_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _28202_[0], clk);
  dff _56597_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _28202_[1], clk);
  dff _56598_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _28202_[2], clk);
  dff _56599_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _28202_[3], clk);
  dff _56600_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _28202_[4], clk);
  dff _56601_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _28202_[5], clk);
  dff _56602_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _28202_[6], clk);
  dff _56603_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _28202_[7], clk);
  dff _56604_ (\oc8051_symbolic_cxrom1.regvalid [0], _25625_, clk);
  dff _56605_ (\oc8051_symbolic_cxrom1.regvalid [1], _25629_, clk);
  dff _56606_ (\oc8051_symbolic_cxrom1.regvalid [2], _25634_, clk);
  dff _56607_ (\oc8051_symbolic_cxrom1.regvalid [3], _25640_, clk);
  dff _56608_ (\oc8051_symbolic_cxrom1.regvalid [4], _25647_, clk);
  dff _56609_ (\oc8051_symbolic_cxrom1.regvalid [5], _25655_, clk);
  dff _56610_ (\oc8051_symbolic_cxrom1.regvalid [6], _25663_, clk);
  dff _56611_ (\oc8051_symbolic_cxrom1.regvalid [7], _25673_, clk);
  dff _56612_ (\oc8051_symbolic_cxrom1.regvalid [8], _25683_, clk);
  dff _56613_ (\oc8051_symbolic_cxrom1.regvalid [9], _28201_[9], clk);
  dff _56614_ (\oc8051_symbolic_cxrom1.regvalid [10], _28201_[10], clk);
  dff _56615_ (\oc8051_symbolic_cxrom1.regvalid [11], _28201_[11], clk);
  dff _56616_ (\oc8051_symbolic_cxrom1.regvalid [12], _28201_[12], clk);
  dff _56617_ (\oc8051_symbolic_cxrom1.regvalid [13], _28201_[13], clk);
  dff _56618_ (\oc8051_symbolic_cxrom1.regvalid [14], _28201_[14], clk);
  dff _56619_ (\oc8051_symbolic_cxrom1.regvalid [15], _25618_, clk);
  dff _56620_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _28209_[0], clk);
  dff _56621_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _28209_[1], clk);
  dff _56622_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _28209_[2], clk);
  dff _56623_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _28209_[3], clk);
  dff _56624_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _28209_[4], clk);
  dff _56625_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _28209_[5], clk);
  dff _56626_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _28209_[6], clk);
  dff _56627_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _28209_[7], clk);
  dff _56628_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _28210_[0], clk);
  dff _56629_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _28210_[1], clk);
  dff _56630_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _28210_[2], clk);
  dff _56631_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _28210_[3], clk);
  dff _56632_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _28210_[4], clk);
  dff _56633_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _28210_[5], clk);
  dff _56634_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _28210_[6], clk);
  dff _56635_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _28210_[7], clk);
  dff _56636_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _28211_[0], clk);
  dff _56637_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _28211_[1], clk);
  dff _56638_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _28211_[2], clk);
  dff _56639_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _28211_[3], clk);
  dff _56640_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _28211_[4], clk);
  dff _56641_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _28211_[5], clk);
  dff _56642_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _28211_[6], clk);
  dff _56643_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _28211_[7], clk);
  dff _56644_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _28212_[0], clk);
  dff _56645_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _28212_[1], clk);
  dff _56646_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _28212_[2], clk);
  dff _56647_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _28212_[3], clk);
  dff _56648_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _28212_[4], clk);
  dff _56649_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _28212_[5], clk);
  dff _56650_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _28212_[6], clk);
  dff _56651_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _28212_[7], clk);
  dff _56652_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _28213_[0], clk);
  dff _56653_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _28213_[1], clk);
  dff _56654_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _28213_[2], clk);
  dff _56655_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _28213_[3], clk);
  dff _56656_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _28213_[4], clk);
  dff _56657_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _28213_[5], clk);
  dff _56658_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _28213_[6], clk);
  dff _56659_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _28213_[7], clk);
  dff _56660_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _28214_[0], clk);
  dff _56661_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _28214_[1], clk);
  dff _56662_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _28214_[2], clk);
  dff _56663_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _28214_[3], clk);
  dff _56664_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _28214_[4], clk);
  dff _56665_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _28214_[5], clk);
  dff _56666_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _28214_[6], clk);
  dff _56667_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _28214_[7], clk);
  dff _56668_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _28215_[0], clk);
  dff _56669_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _28215_[1], clk);
  dff _56670_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _28215_[2], clk);
  dff _56671_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _28215_[3], clk);
  dff _56672_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _28215_[4], clk);
  dff _56673_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _28215_[5], clk);
  dff _56674_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _28215_[6], clk);
  dff _56675_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _28215_[7], clk);
  dff _56676_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _28216_[0], clk);
  dff _56677_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _28216_[1], clk);
  dff _56678_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _28216_[2], clk);
  dff _56679_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _28216_[3], clk);
  dff _56680_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _28216_[4], clk);
  dff _56681_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _28216_[5], clk);
  dff _56682_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _28216_[6], clk);
  dff _56683_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _28216_[7], clk);
  dff _56684_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _28217_[0], clk);
  dff _56685_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _28217_[1], clk);
  dff _56686_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _28217_[2], clk);
  dff _56687_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _28217_[3], clk);
  dff _56688_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _28217_[4], clk);
  dff _56689_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _28217_[5], clk);
  dff _56690_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _28217_[6], clk);
  dff _56691_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _28217_[7], clk);
  dff _56692_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _28203_[0], clk);
  dff _56693_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _28203_[1], clk);
  dff _56694_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _28203_[2], clk);
  dff _56695_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _28203_[3], clk);
  dff _56696_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _28203_[4], clk);
  dff _56697_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _28203_[5], clk);
  dff _56698_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _28203_[6], clk);
  dff _56699_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _28203_[7], clk);
  dff _56700_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _28204_[0], clk);
  dff _56701_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _28204_[1], clk);
  dff _56702_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _28204_[2], clk);
  dff _56703_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _28204_[3], clk);
  dff _56704_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _28204_[4], clk);
  dff _56705_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _28204_[5], clk);
  dff _56706_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _28204_[6], clk);
  dff _56707_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _28204_[7], clk);
  dff _56708_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _28205_[0], clk);
  dff _56709_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _28205_[1], clk);
  dff _56710_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _28205_[2], clk);
  dff _56711_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _28205_[3], clk);
  dff _56712_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _28205_[4], clk);
  dff _56713_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _28205_[5], clk);
  dff _56714_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _28205_[6], clk);
  dff _56715_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _28205_[7], clk);
  dff _56716_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _28206_[0], clk);
  dff _56717_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _28206_[1], clk);
  dff _56718_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _28206_[2], clk);
  dff _56719_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _28206_[3], clk);
  dff _56720_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _28206_[4], clk);
  dff _56721_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _28206_[5], clk);
  dff _56722_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _28206_[6], clk);
  dff _56723_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _28206_[7], clk);
  dff _56724_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _28207_[0], clk);
  dff _56725_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _28207_[1], clk);
  dff _56726_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _28207_[2], clk);
  dff _56727_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _28207_[3], clk);
  dff _56728_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _28207_[4], clk);
  dff _56729_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _28207_[5], clk);
  dff _56730_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _28207_[6], clk);
  dff _56731_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _28207_[7], clk);
  dff _56732_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _28208_[0], clk);
  dff _56733_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _28208_[1], clk);
  dff _56734_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _28208_[2], clk);
  dff _56735_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _28208_[3], clk);
  dff _56736_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _28208_[4], clk);
  dff _56737_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _28208_[5], clk);
  dff _56738_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _28208_[6], clk);
  dff _56739_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _25622_, clk);
  dff _56740_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03039_, clk);
  dff _56741_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03049_, clk);
  dff _56742_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03068_, clk);
  dff _56743_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03084_, clk);
  dff _56744_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03100_, clk);
  dff _56745_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00985_, clk);
  dff _56746_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03108_, clk);
  dff _56747_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00958_, clk);
  dff _56748_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03117_, clk);
  dff _56749_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03125_, clk);
  dff _56750_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03132_, clk);
  dff _56751_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03141_, clk);
  dff _56752_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03149_, clk);
  dff _56753_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03158_, clk);
  dff _56754_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03166_, clk);
  dff _56755_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01001_, clk);
  dff _56756_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02784_, clk);
  dff _56757_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _23530_, clk);
  dff _56758_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02984_, clk);
  dff _56759_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03157_, clk);
  dff _56760_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03302_, clk);
  dff _56761_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03443_, clk);
  dff _56762_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03584_, clk);
  dff _56763_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03782_, clk);
  dff _56764_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03985_, clk);
  dff _56765_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04190_, clk);
  dff _56766_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04293_, clk);
  dff _56767_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04397_, clk);
  dff _56768_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04499_, clk);
  dff _56769_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04604_, clk);
  dff _56770_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04707_, clk);
  dff _56771_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04810_, clk);
  dff _56772_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04914_, clk);
  dff _56773_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _23899_, clk);
  dff _56774_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _24320_, clk);
  dff _56775_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _24321_, clk);
  dff _56776_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _24322_, clk);
  dff _56777_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _24323_, clk);
  dff _56778_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _24324_, clk);
  dff _56779_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _24325_, clk);
  dff _56780_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _24327_, clk);
  dff _56781_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _24306_, clk);
  dff _56782_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _24328_, clk);
  dff _56783_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _24329_, clk);
  dff _56784_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _24330_, clk);
  dff _56785_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _24331_, clk);
  dff _56786_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _24333_, clk);
  dff _56787_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _24334_, clk);
  dff _56788_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _24335_, clk);
  dff _56789_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _24307_, clk);
  dff _56790_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _24336_, clk);
  dff _56791_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _24337_, clk);
  dff _56792_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _24339_, clk);
  dff _56793_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _24340_, clk);
  dff _56794_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _24341_, clk);
  dff _56795_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _24342_, clk);
  dff _56796_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _24343_, clk);
  dff _56797_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _24308_, clk);
  dff _56798_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _23904_, clk);
  dff _56799_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _18908_, clk);
  dff _56800_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _23905_, clk);
  dff _56801_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _23906_, clk);
  dff _56802_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _18911_, clk);
  dff _56803_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _23907_, clk);
  dff _56804_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _23908_, clk);
  dff _56805_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18914_, clk);
  dff _56806_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _23909_, clk);
  dff _56807_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _18917_, clk);
  dff _56808_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _23910_, clk);
  dff _56809_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _23911_, clk);
  dff _56810_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _23912_, clk);
  dff _56811_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _18920_, clk);
  dff _56812_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _23913_, clk);
  dff _56813_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _18923_, clk);
  dff _56814_ (\oc8051_top_1.oc8051_decoder1.wr , _18926_, clk);
  dff _56815_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _18984_, clk);
  dff _56816_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _18986_, clk);
  dff _56817_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _18890_, clk);
  dff _56818_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _18989_, clk);
  dff _56819_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _18992_, clk);
  dff _56820_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _18893_, clk);
  dff _56821_ (\oc8051_top_1.oc8051_decoder1.state [0], _18995_, clk);
  dff _56822_ (\oc8051_top_1.oc8051_decoder1.state [1], _18896_, clk);
  dff _56823_ (\oc8051_top_1.oc8051_decoder1.op [0], _18998_, clk);
  dff _56824_ (\oc8051_top_1.oc8051_decoder1.op [1], _19001_, clk);
  dff _56825_ (\oc8051_top_1.oc8051_decoder1.op [2], _19004_, clk);
  dff _56826_ (\oc8051_top_1.oc8051_decoder1.op [3], _19007_, clk);
  dff _56827_ (\oc8051_top_1.oc8051_decoder1.op [4], _19010_, clk);
  dff _56828_ (\oc8051_top_1.oc8051_decoder1.op [5], _19013_, clk);
  dff _56829_ (\oc8051_top_1.oc8051_decoder1.op [6], _19016_, clk);
  dff _56830_ (\oc8051_top_1.oc8051_decoder1.op [7], _18899_, clk);
  dff _56831_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _18902_, clk);
  dff _56832_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _19019_, clk);
  dff _56833_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18905_, clk);
  dff _56834_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _25154_, clk);
  dff _56835_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _25261_, clk);
  dff _56836_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _25262_, clk);
  dff _56837_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _25263_, clk);
  dff _56838_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _25264_, clk);
  dff _56839_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _25265_, clk);
  dff _56840_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _25267_, clk);
  dff _56841_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _25268_, clk);
  dff _56842_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _25156_, clk);
  dff _56843_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _25269_, clk);
  dff _56844_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _25270_, clk);
  dff _56845_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _25271_, clk);
  dff _56846_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _25272_, clk);
  dff _56847_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _25273_, clk);
  dff _56848_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _25274_, clk);
  dff _56849_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _25275_, clk);
  dff _56850_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _25157_, clk);
  dff _56851_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _25276_, clk);
  dff _56852_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _25278_, clk);
  dff _56853_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _25279_, clk);
  dff _56854_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _25280_, clk);
  dff _56855_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _25281_, clk);
  dff _56856_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _25282_, clk);
  dff _56857_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _25283_, clk);
  dff _56858_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _25158_, clk);
  dff _56859_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _25284_, clk);
  dff _56860_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _25285_, clk);
  dff _56861_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _25286_, clk);
  dff _56862_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _25287_, clk);
  dff _56863_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _25289_, clk);
  dff _56864_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _25290_, clk);
  dff _56865_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _25291_, clk);
  dff _56866_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _25159_, clk);
  dff _56867_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _25292_, clk);
  dff _56868_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _25293_, clk);
  dff _56869_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _25294_, clk);
  dff _56870_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _25295_, clk);
  dff _56871_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _25296_, clk);
  dff _56872_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _25297_, clk);
  dff _56873_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _25298_, clk);
  dff _56874_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _25160_, clk);
  dff _56875_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _25300_, clk);
  dff _56876_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _25301_, clk);
  dff _56877_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _25302_, clk);
  dff _56878_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _25303_, clk);
  dff _56879_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _25304_, clk);
  dff _56880_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _25305_, clk);
  dff _56881_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _25306_, clk);
  dff _56882_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _25161_, clk);
  dff _56883_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _25307_, clk);
  dff _56884_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _25308_, clk);
  dff _56885_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _25309_, clk);
  dff _56886_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _25311_, clk);
  dff _56887_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _25312_, clk);
  dff _56888_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _25313_, clk);
  dff _56889_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _25314_, clk);
  dff _56890_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _25162_, clk);
  dff _56891_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _25315_, clk);
  dff _56892_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _25316_, clk);
  dff _56893_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _25317_, clk);
  dff _56894_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _25318_, clk);
  dff _56895_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _25319_, clk);
  dff _56896_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _25320_, clk);
  dff _56897_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _25322_, clk);
  dff _56898_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _25163_, clk);
  dff _56899_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _24692_, clk);
  dff _56900_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _24693_, clk);
  dff _56901_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _24695_, clk);
  dff _56902_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _24696_, clk);
  dff _56903_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _24405_, clk);
  dff _56904_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _24470_, clk);
  dff _56905_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _24472_, clk);
  dff _56906_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _24473_, clk);
  dff _56907_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _24474_, clk);
  dff _56908_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _24475_, clk);
  dff _56909_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _24476_, clk);
  dff _56910_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _24477_, clk);
  dff _56911_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _24478_, clk);
  dff _56912_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _24479_, clk);
  dff _56913_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _24480_, clk);
  dff _56914_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _24481_, clk);
  dff _56915_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _24483_, clk);
  dff _56916_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _24484_, clk);
  dff _56917_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _24485_, clk);
  dff _56918_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _24486_, clk);
  dff _56919_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _24370_, clk);
  dff _56920_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _24490_, clk);
  dff _56921_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _24491_, clk);
  dff _56922_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _24492_, clk);
  dff _56923_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _24493_, clk);
  dff _56924_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _24494_, clk);
  dff _56925_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _24495_, clk);
  dff _56926_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _24497_, clk);
  dff _56927_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _24498_, clk);
  dff _56928_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _24499_, clk);
  dff _56929_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _24500_, clk);
  dff _56930_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _24501_, clk);
  dff _56931_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _24502_, clk);
  dff _56932_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _24503_, clk);
  dff _56933_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _24504_, clk);
  dff _56934_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _24505_, clk);
  dff _56935_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _24372_, clk);
  dff _56936_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _24697_, clk);
  dff _56937_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _24698_, clk);
  dff _56938_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _24699_, clk);
  dff _56939_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _24700_, clk);
  dff _56940_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _24701_, clk);
  dff _56941_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _24702_, clk);
  dff _56942_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _24703_, clk);
  dff _56943_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _24704_, clk);
  dff _56944_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _24706_, clk);
  dff _56945_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _24707_, clk);
  dff _56946_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _24708_, clk);
  dff _56947_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _24709_, clk);
  dff _56948_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _24710_, clk);
  dff _56949_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _24711_, clk);
  dff _56950_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _24712_, clk);
  dff _56951_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _24713_, clk);
  dff _56952_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _24714_, clk);
  dff _56953_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _24715_, clk);
  dff _56954_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _24717_, clk);
  dff _56955_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _24718_, clk);
  dff _56956_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _24719_, clk);
  dff _56957_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _24720_, clk);
  dff _56958_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _24721_, clk);
  dff _56959_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _24722_, clk);
  dff _56960_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _24723_, clk);
  dff _56961_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _24724_, clk);
  dff _56962_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _24725_, clk);
  dff _56963_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _24726_, clk);
  dff _56964_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _24728_, clk);
  dff _56965_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _24729_, clk);
  dff _56966_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _24730_, clk);
  dff _56967_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _24429_, clk);
  dff _56968_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _24404_, clk);
  dff _56969_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _56970_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _24731_, clk);
  dff _56971_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _24732_, clk);
  dff _56972_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _24733_, clk);
  dff _56973_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _24735_, clk);
  dff _56974_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _24736_, clk);
  dff _56975_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _24737_, clk);
  dff _56976_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _24738_, clk);
  dff _56977_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _24406_, clk);
  dff _56978_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _24739_, clk);
  dff _56979_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _24740_, clk);
  dff _56980_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _24741_, clk);
  dff _56981_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _24743_, clk);
  dff _56982_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _24744_, clk);
  dff _56983_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _24745_, clk);
  dff _56984_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _24746_, clk);
  dff _56985_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _24407_, clk);
  dff _56986_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _24747_, clk);
  dff _56987_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _24748_, clk);
  dff _56988_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _24749_, clk);
  dff _56989_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _24750_, clk);
  dff _56990_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _24751_, clk);
  dff _56991_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _24752_, clk);
  dff _56992_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _24754_, clk);
  dff _56993_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _24409_, clk);
  dff _56994_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _24410_, clk);
  dff _56995_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _24411_, clk);
  dff _56996_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _24755_, clk);
  dff _56997_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _24756_, clk);
  dff _56998_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _24757_, clk);
  dff _56999_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _24758_, clk);
  dff _57000_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _24759_, clk);
  dff _57001_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _24760_, clk);
  dff _57002_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _24761_, clk);
  dff _57003_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _24412_, clk);
  dff _57004_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _24762_, clk);
  dff _57005_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _24763_, clk);
  dff _57006_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _24765_, clk);
  dff _57007_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _24766_, clk);
  dff _57008_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _24767_, clk);
  dff _57009_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _24768_, clk);
  dff _57010_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _24769_, clk);
  dff _57011_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _24770_, clk);
  dff _57012_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _24771_, clk);
  dff _57013_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _24772_, clk);
  dff _57014_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _24773_, clk);
  dff _57015_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _24774_, clk);
  dff _57016_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _24776_, clk);
  dff _57017_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _24777_, clk);
  dff _57018_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _24778_, clk);
  dff _57019_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _24414_, clk);
  dff _57020_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _24779_, clk);
  dff _57021_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _24780_, clk);
  dff _57022_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _24781_, clk);
  dff _57023_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _24782_, clk);
  dff _57024_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _24783_, clk);
  dff _57025_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _24784_, clk);
  dff _57026_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _24785_, clk);
  dff _57027_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _24787_, clk);
  dff _57028_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _24788_, clk);
  dff _57029_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _24789_, clk);
  dff _57030_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _24790_, clk);
  dff _57031_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _24791_, clk);
  dff _57032_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _24792_, clk);
  dff _57033_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _24793_, clk);
  dff _57034_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _24794_, clk);
  dff _57035_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _24415_, clk);
  dff _57036_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _24416_, clk);
  dff _57037_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _24418_, clk);
  dff _57038_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _24417_, clk);
  dff _57039_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _24795_, clk);
  dff _57040_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _24796_, clk);
  dff _57041_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _24798_, clk);
  dff _57042_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _24799_, clk);
  dff _57043_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _24800_, clk);
  dff _57044_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _24801_, clk);
  dff _57045_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _24802_, clk);
  dff _57046_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _24419_, clk);
  dff _57047_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _24803_, clk);
  dff _57048_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _24804_, clk);
  dff _57049_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _24420_, clk);
  dff _57050_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _24805_, clk);
  dff _57051_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _24806_, clk);
  dff _57052_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _24807_, clk);
  dff _57053_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _24809_, clk);
  dff _57054_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _24810_, clk);
  dff _57055_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _24811_, clk);
  dff _57056_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _24812_, clk);
  dff _57057_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _24421_, clk);
  dff _57058_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _24813_, clk);
  dff _57059_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _24814_, clk);
  dff _57060_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _24815_, clk);
  dff _57061_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _24816_, clk);
  dff _57062_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _24817_, clk);
  dff _57063_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _24818_, clk);
  dff _57064_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _24820_, clk);
  dff _57065_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _24422_, clk);
  dff _57066_ (\oc8051_top_1.oc8051_memory_interface1.reti , _24423_, clk);
  dff _57067_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _24821_, clk);
  dff _57068_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _24822_, clk);
  dff _57069_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _24823_, clk);
  dff _57070_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _24824_, clk);
  dff _57071_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _24825_, clk);
  dff _57072_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _24826_, clk);
  dff _57073_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _24827_, clk);
  dff _57074_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _24424_, clk);
  dff _57075_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _24426_, clk);
  dff _57076_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _24427_, clk);
  dff _57077_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _24828_, clk);
  dff _57078_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _24829_, clk);
  dff _57079_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _24831_, clk);
  dff _57080_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _24428_, clk);
  dff _57081_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _24832_, clk);
  dff _57082_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _24833_, clk);
  dff _57083_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _24834_, clk);
  dff _57084_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _24835_, clk);
  dff _57085_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _24836_, clk);
  dff _57086_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _24837_, clk);
  dff _57087_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _24838_, clk);
  dff _57088_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _24839_, clk);
  dff _57089_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _24840_, clk);
  dff _57090_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _24842_, clk);
  dff _57091_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _24843_, clk);
  dff _57092_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _24844_, clk);
  dff _57093_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _24845_, clk);
  dff _57094_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _24846_, clk);
  dff _57095_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _24847_, clk);
  dff _57096_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _24848_, clk);
  dff _57097_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _24849_, clk);
  dff _57098_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _24850_, clk);
  dff _57099_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _24851_, clk);
  dff _57100_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _24853_, clk);
  dff _57101_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _24854_, clk);
  dff _57102_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _24855_, clk);
  dff _57103_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _24856_, clk);
  dff _57104_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _24857_, clk);
  dff _57105_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _24858_, clk);
  dff _57106_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _24859_, clk);
  dff _57107_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _24860_, clk);
  dff _57108_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _24861_, clk);
  dff _57109_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _24862_, clk);
  dff _57110_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _24864_, clk);
  dff _57111_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _24865_, clk);
  dff _57112_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _24430_, clk);
  dff _57113_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _24866_, clk);
  dff _57114_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _24867_, clk);
  dff _57115_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _24868_, clk);
  dff _57116_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _24869_, clk);
  dff _57117_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _24870_, clk);
  dff _57118_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _24871_, clk);
  dff _57119_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _24872_, clk);
  dff _57120_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _24431_, clk);
  dff _57121_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _24433_, clk);
  dff _57122_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _24434_, clk);
  dff _57123_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _24873_, clk);
  dff _57124_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _24875_, clk);
  dff _57125_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _24876_, clk);
  dff _57126_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _24877_, clk);
  dff _57127_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _24878_, clk);
  dff _57128_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _24879_, clk);
  dff _57129_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _24880_, clk);
  dff _57130_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _24881_, clk);
  dff _57131_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _24882_, clk);
  dff _57132_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _24883_, clk);
  dff _57133_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _24884_, clk);
  dff _57134_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _24886_, clk);
  dff _57135_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _24887_, clk);
  dff _57136_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _24888_, clk);
  dff _57137_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _24889_, clk);
  dff _57138_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _24435_, clk);
  dff _57139_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _24436_, clk);
  dff _57140_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _24437_, clk);
  dff _57141_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _24438_, clk);
  dff _57142_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _24890_, clk);
  dff _57143_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _24891_, clk);
  dff _57144_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _24892_, clk);
  dff _57145_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _24893_, clk);
  dff _57146_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _24894_, clk);
  dff _57147_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _24895_, clk);
  dff _57148_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _24897_, clk);
  dff _57149_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _24898_, clk);
  dff _57150_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _24899_, clk);
  dff _57151_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _24900_, clk);
  dff _57152_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _24901_, clk);
  dff _57153_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _24902_, clk);
  dff _57154_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _24903_, clk);
  dff _57155_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _24904_, clk);
  dff _57156_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _24905_, clk);
  dff _57157_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _24439_, clk);
  dff _57158_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _24440_, clk);
  dff _57159_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _25567_, clk);
  dff _57160_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _25586_, clk);
  dff _57161_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _25587_, clk);
  dff _57162_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _25588_, clk);
  dff _57163_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _25589_, clk);
  dff _57164_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _25590_, clk);
  dff _57165_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _25591_, clk);
  dff _57166_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _25592_, clk);
  dff _57167_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _25568_, clk);
  dff _57168_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25569_, clk);
  dff _57169_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _25593_, clk);
  dff _57170_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _25594_, clk);
  dff _57171_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _25571_, clk);
  dff _57172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _04005_, clk);
  dff _57173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _04008_, clk);
  dff _57174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _04011_, clk);
  dff _57175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _04014_, clk);
  dff _57176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _04017_, clk);
  dff _57177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _04021_, clk);
  dff _57178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _04024_, clk);
  dff _57179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _04026_, clk);
  dff _57180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03977_, clk);
  dff _57181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03980_, clk);
  dff _57182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03983_, clk);
  dff _57183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03987_, clk);
  dff _57184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03990_, clk);
  dff _57185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03993_, clk);
  dff _57186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03997_, clk);
  dff _57187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _03999_, clk);
  dff _57188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03952_, clk);
  dff _57189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03955_, clk);
  dff _57190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03958_, clk);
  dff _57191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03961_, clk);
  dff _57192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03964_, clk);
  dff _57193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03967_, clk);
  dff _57194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03970_, clk);
  dff _57195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03973_, clk);
  dff _57196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03926_, clk);
  dff _57197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03929_, clk);
  dff _57198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03932_, clk);
  dff _57199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03935_, clk);
  dff _57200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03938_, clk);
  dff _57201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03942_, clk);
  dff _57202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03945_, clk);
  dff _57203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03947_, clk);
  dff _57204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _04030_, clk);
  dff _57205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _04033_, clk);
  dff _57206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _04036_, clk);
  dff _57207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _04039_, clk);
  dff _57208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _04042_, clk);
  dff _57209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _04045_, clk);
  dff _57210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _04049_, clk);
  dff _57211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _04051_, clk);
  dff _57212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03901_, clk);
  dff _57213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03904_, clk);
  dff _57214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03907_, clk);
  dff _57215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03910_, clk);
  dff _57216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03913_, clk);
  dff _57217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03917_, clk);
  dff _57218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03920_, clk);
  dff _57219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03922_, clk);
  dff _57220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03875_, clk);
  dff _57221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03878_, clk);
  dff _57222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03881_, clk);
  dff _57223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03884_, clk);
  dff _57224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03887_, clk);
  dff _57225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03891_, clk);
  dff _57226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03894_, clk);
  dff _57227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03896_, clk);
  dff _57228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03850_, clk);
  dff _57229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03853_, clk);
  dff _57230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03856_, clk);
  dff _57231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03859_, clk);
  dff _57232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03862_, clk);
  dff _57233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03865_, clk);
  dff _57234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03868_, clk);
  dff _57235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03871_, clk);
  dff _57236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03824_, clk);
  dff _57237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03827_, clk);
  dff _57238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03830_, clk);
  dff _57239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03833_, clk);
  dff _57240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03837_, clk);
  dff _57241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03840_, clk);
  dff _57242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03843_, clk);
  dff _57243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03845_, clk);
  dff _57244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _04055_, clk);
  dff _57245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _04058_, clk);
  dff _57246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _04061_, clk);
  dff _57247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _04064_, clk);
  dff _57248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _04067_, clk);
  dff _57249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _04070_, clk);
  dff _57250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _04073_, clk);
  dff _57251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _04076_, clk);
  dff _57252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _04278_, clk);
  dff _57253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _04281_, clk);
  dff _57254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _04284_, clk);
  dff _57255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _04287_, clk);
  dff _57256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _04290_, clk);
  dff _57257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _04294_, clk);
  dff _57258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04297_, clk);
  dff _57259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _04300_, clk);
  dff _57260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _04253_, clk);
  dff _57261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _04256_, clk);
  dff _57262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _04259_, clk);
  dff _57263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _04262_, clk);
  dff _57264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _04266_, clk);
  dff _57265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _04269_, clk);
  dff _57266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _04272_, clk);
  dff _57267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _04274_, clk);
  dff _57268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _04228_, clk);
  dff _57269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _04231_, clk);
  dff _57270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _04234_, clk);
  dff _57271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _04238_, clk);
  dff _57272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04241_, clk);
  dff _57273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _04244_, clk);
  dff _57274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _04247_, clk);
  dff _57275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _04249_, clk);
  dff _57276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _04855_, clk);
  dff _57277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _04858_, clk);
  dff _57278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _04861_, clk);
  dff _57279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _04864_, clk);
  dff _57280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _04867_, clk);
  dff _57281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _04870_, clk);
  dff _57282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _04873_, clk);
  dff _57283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _04876_, clk);
  dff _57284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _04830_, clk);
  dff _57285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _04834_, clk);
  dff _57286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _04837_, clk);
  dff _57287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _04840_, clk);
  dff _57288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _04843_, clk);
  dff _57289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _04846_, clk);
  dff _57290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _04849_, clk);
  dff _57291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _04851_, clk);
  dff _57292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _04805_, clk);
  dff _57293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _04808_, clk);
  dff _57294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _04812_, clk);
  dff _57295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _04815_, clk);
  dff _57296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _04818_, clk);
  dff _57297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _04821_, clk);
  dff _57298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _04824_, clk);
  dff _57299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _04826_, clk);
  dff _57300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _04779_, clk);
  dff _57301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _04782_, clk);
  dff _57302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _04785_, clk);
  dff _57303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _04788_, clk);
  dff _57304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _04791_, clk);
  dff _57305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _04794_, clk);
  dff _57306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _04797_, clk);
  dff _57307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _04799_, clk);
  dff _57308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _04754_, clk);
  dff _57309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _04757_, clk);
  dff _57310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _04760_, clk);
  dff _57311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _04763_, clk);
  dff _57312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _04766_, clk);
  dff _57313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _04769_, clk);
  dff _57314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _04772_, clk);
  dff _57315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _04775_, clk);
  dff _57316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _04730_, clk);
  dff _57317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _04733_, clk);
  dff _57318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _04736_, clk);
  dff _57319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _04739_, clk);
  dff _57320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _04742_, clk);
  dff _57321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _04745_, clk);
  dff _57322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _04748_, clk);
  dff _57323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _04750_, clk);
  dff _57324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _04704_, clk);
  dff _57325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _04708_, clk);
  dff _57326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _04711_, clk);
  dff _57327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _04714_, clk);
  dff _57328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _04717_, clk);
  dff _57329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _04720_, clk);
  dff _57330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _04723_, clk);
  dff _57331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _04726_, clk);
  dff _57332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _04679_, clk);
  dff _57333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _04682_, clk);
  dff _57334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _04685_, clk);
  dff _57335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _04688_, clk);
  dff _57336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _04691_, clk);
  dff _57337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _04694_, clk);
  dff _57338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _04698_, clk);
  dff _57339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _04700_, clk);
  dff _57340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _04655_, clk);
  dff _57341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _04658_, clk);
  dff _57342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _04661_, clk);
  dff _57343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _04664_, clk);
  dff _57344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _04667_, clk);
  dff _57345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _04670_, clk);
  dff _57346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _04673_, clk);
  dff _57347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _04676_, clk);
  dff _57348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _04630_, clk);
  dff _57349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _04633_, clk);
  dff _57350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _04636_, clk);
  dff _57351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _04639_, clk);
  dff _57352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _04642_, clk);
  dff _57353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _04646_, clk);
  dff _57354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _04649_, clk);
  dff _57355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _04651_, clk);
  dff _57356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _04605_, clk);
  dff _57357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _04608_, clk);
  dff _57358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _04611_, clk);
  dff _57359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _04614_, clk);
  dff _57360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _04618_, clk);
  dff _57361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _04621_, clk);
  dff _57362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _04624_, clk);
  dff _57363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _04626_, clk);
  dff _57364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _06067_, clk);
  dff _57365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _06070_, clk);
  dff _57366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _06073_, clk);
  dff _57367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _06076_, clk);
  dff _57368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _06079_, clk);
  dff _57369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _06082_, clk);
  dff _57370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _06085_, clk);
  dff _57371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _06088_, clk);
  dff _57372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _06043_, clk);
  dff _57373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _06046_, clk);
  dff _57374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _06049_, clk);
  dff _57375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _06052_, clk);
  dff _57376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _06055_, clk);
  dff _57377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _06058_, clk);
  dff _57378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _06061_, clk);
  dff _57379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _06064_, clk);
  dff _57380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _06018_, clk);
  dff _57381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _06021_, clk);
  dff _57382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _06024_, clk);
  dff _57383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _06027_, clk);
  dff _57384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _06030_, clk);
  dff _57385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _06033_, clk);
  dff _57386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _06037_, clk);
  dff _57387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _06039_, clk);
  dff _57388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _05993_, clk);
  dff _57389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _05996_, clk);
  dff _57390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _05999_, clk);
  dff _57391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _06002_, clk);
  dff _57392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _06005_, clk);
  dff _57393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _06009_, clk);
  dff _57394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _06012_, clk);
  dff _57395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _06014_, clk);
  dff _57396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _05968_, clk);
  dff _57397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _05971_, clk);
  dff _57398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _05974_, clk);
  dff _57399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _05977_, clk);
  dff _57400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _05980_, clk);
  dff _57401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _05984_, clk);
  dff _57402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _05987_, clk);
  dff _57403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _05989_, clk);
  dff _57404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _05943_, clk);
  dff _57405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _05946_, clk);
  dff _57406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _05949_, clk);
  dff _57407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _05952_, clk);
  dff _57408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _05956_, clk);
  dff _57409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _05959_, clk);
  dff _57410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _05962_, clk);
  dff _57411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _05964_, clk);
  dff _57412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _05919_, clk);
  dff _57413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _05922_, clk);
  dff _57414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _05925_, clk);
  dff _57415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _05928_, clk);
  dff _57416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _05931_, clk);
  dff _57417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _05934_, clk);
  dff _57418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _05937_, clk);
  dff _57419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _05940_, clk);
  dff _57420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _05894_, clk);
  dff _57421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _05897_, clk);
  dff _57422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _05900_, clk);
  dff _57423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _05904_, clk);
  dff _57424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _05907_, clk);
  dff _57425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _05910_, clk);
  dff _57426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _05913_, clk);
  dff _57427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _05915_, clk);
  dff _57428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _06314_, clk);
  dff _57429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _06317_, clk);
  dff _57430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _06320_, clk);
  dff _57431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _06323_, clk);
  dff _57432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _06326_, clk);
  dff _57433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _06329_, clk);
  dff _57434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _06333_, clk);
  dff _57435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _06335_, clk);
  dff _57436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _06289_, clk);
  dff _57437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _06292_, clk);
  dff _57438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _06295_, clk);
  dff _57439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _06298_, clk);
  dff _57440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _06301_, clk);
  dff _57441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _06305_, clk);
  dff _57442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _06308_, clk);
  dff _57443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _06310_, clk);
  dff _57444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _06264_, clk);
  dff _57445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _06267_, clk);
  dff _57446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _06270_, clk);
  dff _57447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _06273_, clk);
  dff _57448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _06277_, clk);
  dff _57449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _06280_, clk);
  dff _57450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _06283_, clk);
  dff _57451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _06286_, clk);
  dff _57452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _06239_, clk);
  dff _57453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _06242_, clk);
  dff _57454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _06245_, clk);
  dff _57455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _06249_, clk);
  dff _57456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _06252_, clk);
  dff _57457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _06255_, clk);
  dff _57458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _06258_, clk);
  dff _57459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _06260_, clk);
  dff _57460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _06339_, clk);
  dff _57461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _06342_, clk);
  dff _57462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _06345_, clk);
  dff _57463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _06348_, clk);
  dff _57464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _06351_, clk);
  dff _57465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _06354_, clk);
  dff _57466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _06357_, clk);
  dff _57467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _06360_, clk);
  dff _57468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _06487_, clk);
  dff _57469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _06490_, clk);
  dff _57470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _06493_, clk);
  dff _57471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _06496_, clk);
  dff _57472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _06499_, clk);
  dff _57473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _06502_, clk);
  dff _57474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _06505_, clk);
  dff _57475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _06508_, clk);
  dff _57476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _06462_, clk);
  dff _57477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _06466_, clk);
  dff _57478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _06469_, clk);
  dff _57479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _06472_, clk);
  dff _57480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _06475_, clk);
  dff _57481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _06478_, clk);
  dff _57482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _06481_, clk);
  dff _57483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _06483_, clk);
  dff _57484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _06438_, clk);
  dff _57485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _06441_, clk);
  dff _57486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06444_, clk);
  dff _57487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _06447_, clk);
  dff _57488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06450_, clk);
  dff _57489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _06453_, clk);
  dff _57490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _06456_, clk);
  dff _57491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06458_, clk);
  dff _57492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0], _10034_, clk);
  dff _57493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1], _10038_, clk);
  dff _57494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2], _10042_, clk);
  dff _57495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3], _10046_, clk);
  dff _57496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4], _10050_, clk);
  dff _57497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5], _10054_, clk);
  dff _57498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6], _10058_, clk);
  dff _57499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7], _02706_, clk);
  dff _57500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _09997_, clk);
  dff _57501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _10001_, clk);
  dff _57502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _10005_, clk);
  dff _57503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _10009_, clk);
  dff _57504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _10013_, clk);
  dff _57505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _10017_, clk);
  dff _57506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _10021_, clk);
  dff _57507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _10024_, clk);
  dff _57508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _09965_, clk);
  dff _57509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _09969_, clk);
  dff _57510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _09973_, clk);
  dff _57511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _09977_, clk);
  dff _57512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _09981_, clk);
  dff _57513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _09985_, clk);
  dff _57514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _09989_, clk);
  dff _57515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _09992_, clk);
  dff _57516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _09933_, clk);
  dff _57517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _09937_, clk);
  dff _57518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _09941_, clk);
  dff _57519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _09945_, clk);
  dff _57520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _09949_, clk);
  dff _57521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _09953_, clk);
  dff _57522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _09957_, clk);
  dff _57523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _09960_, clk);
  dff _57524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _09901_, clk);
  dff _57525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _09905_, clk);
  dff _57526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _09909_, clk);
  dff _57527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _09913_, clk);
  dff _57528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _09917_, clk);
  dff _57529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _09921_, clk);
  dff _57530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _09925_, clk);
  dff _57531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _09928_, clk);
  dff _57532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _09869_, clk);
  dff _57533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _09873_, clk);
  dff _57534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _09877_, clk);
  dff _57535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _09881_, clk);
  dff _57536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _09885_, clk);
  dff _57537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _09889_, clk);
  dff _57538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _09893_, clk);
  dff _57539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _09896_, clk);
  dff _57540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _05475_, clk);
  dff _57541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _05478_, clk);
  dff _57542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _05481_, clk);
  dff _57543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _05484_, clk);
  dff _57544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _05487_, clk);
  dff _57545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _05490_, clk);
  dff _57546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _05493_, clk);
  dff _57547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _05495_, clk);
  dff _57548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _09837_, clk);
  dff _57549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _09841_, clk);
  dff _57550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _09845_, clk);
  dff _57551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _09849_, clk);
  dff _57552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _09853_, clk);
  dff _57553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _09857_, clk);
  dff _57554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _09861_, clk);
  dff _57555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _09864_, clk);
  dff _57556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _09805_, clk);
  dff _57557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _09809_, clk);
  dff _57558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _09813_, clk);
  dff _57559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _09817_, clk);
  dff _57560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _09821_, clk);
  dff _57561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _09825_, clk);
  dff _57562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _09829_, clk);
  dff _57563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _09832_, clk);
  dff _57564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _09773_, clk);
  dff _57565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _09777_, clk);
  dff _57566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _09781_, clk);
  dff _57567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _09785_, clk);
  dff _57568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _09789_, clk);
  dff _57569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _09793_, clk);
  dff _57570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _09797_, clk);
  dff _57571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _09800_, clk);
  dff _57572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _09741_, clk);
  dff _57573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _09745_, clk);
  dff _57574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _09749_, clk);
  dff _57575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _09753_, clk);
  dff _57576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _09757_, clk);
  dff _57577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _09761_, clk);
  dff _57578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _09765_, clk);
  dff _57579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _09768_, clk);
  dff _57580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _09709_, clk);
  dff _57581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _09713_, clk);
  dff _57582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _09717_, clk);
  dff _57583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _09721_, clk);
  dff _57584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _09725_, clk);
  dff _57585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _09729_, clk);
  dff _57586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _09733_, clk);
  dff _57587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _09736_, clk);
  dff _57588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _09684_, clk);
  dff _57589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _09687_, clk);
  dff _57590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _09690_, clk);
  dff _57591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _09693_, clk);
  dff _57592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _09696_, clk);
  dff _57593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _09699_, clk);
  dff _57594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _09702_, clk);
  dff _57595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _09704_, clk);
  dff _57596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _09659_, clk);
  dff _57597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _09662_, clk);
  dff _57598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _09665_, clk);
  dff _57599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _09668_, clk);
  dff _57600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _09671_, clk);
  dff _57601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _09674_, clk);
  dff _57602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _09677_, clk);
  dff _57603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _09680_, clk);
  dff _57604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _09635_, clk);
  dff _57605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _09638_, clk);
  dff _57606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _09641_, clk);
  dff _57607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _09644_, clk);
  dff _57608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _09647_, clk);
  dff _57609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _09650_, clk);
  dff _57610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _09653_, clk);
  dff _57611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _09656_, clk);
  dff _57612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _09610_, clk);
  dff _57613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _09613_, clk);
  dff _57614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _09616_, clk);
  dff _57615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _09619_, clk);
  dff _57616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _09622_, clk);
  dff _57617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _09625_, clk);
  dff _57618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _09629_, clk);
  dff _57619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _09631_, clk);
  dff _57620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _09585_, clk);
  dff _57621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _09588_, clk);
  dff _57622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _09591_, clk);
  dff _57623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _09594_, clk);
  dff _57624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _09597_, clk);
  dff _57625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _09601_, clk);
  dff _57626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _09604_, clk);
  dff _57627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _09606_, clk);
  dff _57628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _09561_, clk);
  dff _57629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _09564_, clk);
  dff _57630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _09567_, clk);
  dff _57631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _09570_, clk);
  dff _57632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _09573_, clk);
  dff _57633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _09576_, clk);
  dff _57634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _09579_, clk);
  dff _57635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _09582_, clk);
  dff _57636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _09535_, clk);
  dff _57637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _09538_, clk);
  dff _57638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _09541_, clk);
  dff _57639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _09544_, clk);
  dff _57640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _09548_, clk);
  dff _57641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _09551_, clk);
  dff _57642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _09554_, clk);
  dff _57643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _09556_, clk);
  dff _57644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _09511_, clk);
  dff _57645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _09514_, clk);
  dff _57646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _09517_, clk);
  dff _57647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _09520_, clk);
  dff _57648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _09523_, clk);
  dff _57649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _09526_, clk);
  dff _57650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _09529_, clk);
  dff _57651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _09532_, clk);
  dff _57652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _09485_, clk);
  dff _57653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _09488_, clk);
  dff _57654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _09491_, clk);
  dff _57655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _09495_, clk);
  dff _57656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _09499_, clk);
  dff _57657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _09502_, clk);
  dff _57658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _09505_, clk);
  dff _57659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _09507_, clk);
  dff _57660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _05426_, clk);
  dff _57661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _05429_, clk);
  dff _57662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _05432_, clk);
  dff _57663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _05435_, clk);
  dff _57664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _05438_, clk);
  dff _57665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _05441_, clk);
  dff _57666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _05444_, clk);
  dff _57667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _05446_, clk);
  dff _57668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _09459_, clk);
  dff _57669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _09462_, clk);
  dff _57670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _09466_, clk);
  dff _57671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _09469_, clk);
  dff _57672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _09472_, clk);
  dff _57673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _09476_, clk);
  dff _57674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _09479_, clk);
  dff _57675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _09481_, clk);
  dff _57676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _05450_, clk);
  dff _57677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _05453_, clk);
  dff _57678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _05456_, clk);
  dff _57679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _05459_, clk);
  dff _57680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _05462_, clk);
  dff _57681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _05465_, clk);
  dff _57682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _05468_, clk);
  dff _57683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _05471_, clk);
  dff _57684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _09435_, clk);
  dff _57685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _09438_, clk);
  dff _57686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _09441_, clk);
  dff _57687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _09444_, clk);
  dff _57688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _09447_, clk);
  dff _57689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _09450_, clk);
  dff _57690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _09453_, clk);
  dff _57691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _09456_, clk);
  dff _57692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _09410_, clk);
  dff _57693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _09414_, clk);
  dff _57694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _09417_, clk);
  dff _57695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _09420_, clk);
  dff _57696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _09423_, clk);
  dff _57697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _09426_, clk);
  dff _57698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _09429_, clk);
  dff _57699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _09431_, clk);
  dff _57700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _09386_, clk);
  dff _57701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _09389_, clk);
  dff _57702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _09392_, clk);
  dff _57703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _09395_, clk);
  dff _57704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _09398_, clk);
  dff _57705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _09401_, clk);
  dff _57706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _09404_, clk);
  dff _57707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _09406_, clk);
  dff _57708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _09361_, clk);
  dff _57709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _09364_, clk);
  dff _57710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _09367_, clk);
  dff _57711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _09370_, clk);
  dff _57712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _09373_, clk);
  dff _57713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _09376_, clk);
  dff _57714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _09379_, clk);
  dff _57715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _09382_, clk);
  dff _57716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _09337_, clk);
  dff _57717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _09340_, clk);
  dff _57718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _09343_, clk);
  dff _57719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _09346_, clk);
  dff _57720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _09349_, clk);
  dff _57721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _09352_, clk);
  dff _57722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _09355_, clk);
  dff _57723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _09357_, clk);
  dff _57724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _09312_, clk);
  dff _57725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _09315_, clk);
  dff _57726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _09318_, clk);
  dff _57727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _09321_, clk);
  dff _57728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _09324_, clk);
  dff _57729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _09327_, clk);
  dff _57730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _09330_, clk);
  dff _57731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _09333_, clk);
  dff _57732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _05401_, clk);
  dff _57733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _05404_, clk);
  dff _57734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _05407_, clk);
  dff _57735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _05410_, clk);
  dff _57736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _05413_, clk);
  dff _57737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _05416_, clk);
  dff _57738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _05419_, clk);
  dff _57739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _05422_, clk);
  dff _57740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _05376_, clk);
  dff _57741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _05379_, clk);
  dff _57742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _05382_, clk);
  dff _57743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _05385_, clk);
  dff _57744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _05388_, clk);
  dff _57745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _05391_, clk);
  dff _57746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _05395_, clk);
  dff _57747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _05397_, clk);
  dff _57748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _05327_, clk);
  dff _57749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _05330_, clk);
  dff _57750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _05333_, clk);
  dff _57751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _05336_, clk);
  dff _57752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _05339_, clk);
  dff _57753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _05342_, clk);
  dff _57754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _05345_, clk);
  dff _57755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _05348_, clk);
  dff _57756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _05302_, clk);
  dff _57757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _05305_, clk);
  dff _57758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _05308_, clk);
  dff _57759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _05311_, clk);
  dff _57760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _05315_, clk);
  dff _57761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _05318_, clk);
  dff _57762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _05321_, clk);
  dff _57763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _05323_, clk);
  dff _57764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _05277_, clk);
  dff _57765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _05280_, clk);
  dff _57766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _05283_, clk);
  dff _57767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _05287_, clk);
  dff _57768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _05290_, clk);
  dff _57769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _05293_, clk);
  dff _57770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _05296_, clk);
  dff _57771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _05298_, clk);
  dff _57772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _03613_, clk);
  dff _57773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _03616_, clk);
  dff _57774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _03619_, clk);
  dff _57775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _03622_, clk);
  dff _57776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _03626_, clk);
  dff _57777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _03629_, clk);
  dff _57778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _03632_, clk);
  dff _57779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _03634_, clk);
  dff _57780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _05228_, clk);
  dff _57781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _05231_, clk);
  dff _57782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _05235_, clk);
  dff _57783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _05238_, clk);
  dff _57784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _05241_, clk);
  dff _57785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _05244_, clk);
  dff _57786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _05247_, clk);
  dff _57787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _05249_, clk);
  dff _57788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _03577_, clk);
  dff _57789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _03581_, clk);
  dff _57790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _03587_, clk);
  dff _57791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _03591_, clk);
  dff _57792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _03595_, clk);
  dff _57793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _03600_, clk);
  dff _57794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _03605_, clk);
  dff _57795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _03607_, clk);
  dff _57796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _03694_, clk);
  dff _57797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _03697_, clk);
  dff _57798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _03700_, clk);
  dff _57799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _03704_, clk);
  dff _57800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _03707_, clk);
  dff _57801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _03710_, clk);
  dff _57802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _03713_, clk);
  dff _57803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _03716_, clk);
  dff _57804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _03667_, clk);
  dff _57805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _03670_, clk);
  dff _57806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _03673_, clk);
  dff _57807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _03676_, clk);
  dff _57808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _03679_, clk);
  dff _57809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _03682_, clk);
  dff _57810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _03685_, clk);
  dff _57811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _03688_, clk);
  dff _57812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _03641_, clk);
  dff _57813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _03644_, clk);
  dff _57814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _03647_, clk);
  dff _57815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _03650_, clk);
  dff _57816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _03653_, clk);
  dff _57817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _03656_, clk);
  dff _57818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _03659_, clk);
  dff _57819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _03662_, clk);
  dff _57820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03771_, clk);
  dff _57821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03774_, clk);
  dff _57822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03777_, clk);
  dff _57823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03780_, clk);
  dff _57824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03784_, clk);
  dff _57825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03787_, clk);
  dff _57826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03790_, clk);
  dff _57827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03793_, clk);
  dff _57828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _03745_, clk);
  dff _57829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _03748_, clk);
  dff _57830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03751_, clk);
  dff _57831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03754_, clk);
  dff _57832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03758_, clk);
  dff _57833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03761_, clk);
  dff _57834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03764_, clk);
  dff _57835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03766_, clk);
  dff _57836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _03720_, clk);
  dff _57837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _03723_, clk);
  dff _57838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _03726_, clk);
  dff _57839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _03729_, clk);
  dff _57840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _03733_, clk);
  dff _57841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _03736_, clk);
  dff _57842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _03739_, clk);
  dff _57843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _03741_, clk);
  dff _57844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _05253_, clk);
  dff _57845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _05256_, clk);
  dff _57846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _05259_, clk);
  dff _57847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _05262_, clk);
  dff _57848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _05265_, clk);
  dff _57849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _05268_, clk);
  dff _57850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _05271_, clk);
  dff _57851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _05274_, clk);
  dff _57852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03799_, clk);
  dff _57853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03802_, clk);
  dff _57854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03805_, clk);
  dff _57855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03808_, clk);
  dff _57856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03812_, clk);
  dff _57857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03815_, clk);
  dff _57858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03818_, clk);
  dff _57859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03820_, clk);
  dff _57860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _09287_, clk);
  dff _57861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _09290_, clk);
  dff _57862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _09293_, clk);
  dff _57863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _09296_, clk);
  dff _57864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _09299_, clk);
  dff _57865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _09302_, clk);
  dff _57866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _09306_, clk);
  dff _57867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _09308_, clk);
  dff _57868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _09262_, clk);
  dff _57869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _09265_, clk);
  dff _57870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _09268_, clk);
  dff _57871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _09271_, clk);
  dff _57872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _09274_, clk);
  dff _57873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _09278_, clk);
  dff _57874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _09281_, clk);
  dff _57875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _09284_, clk);
  dff _57876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _09238_, clk);
  dff _57877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _09241_, clk);
  dff _57878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _09244_, clk);
  dff _57879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _09247_, clk);
  dff _57880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _09250_, clk);
  dff _57881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _09253_, clk);
  dff _57882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _09256_, clk);
  dff _57883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _09259_, clk);
  dff _57884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _09213_, clk);
  dff _57885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _09216_, clk);
  dff _57886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _09219_, clk);
  dff _57887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _09222_, clk);
  dff _57888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _09226_, clk);
  dff _57889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _09229_, clk);
  dff _57890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _09232_, clk);
  dff _57891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _09234_, clk);
  dff _57892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _09188_, clk);
  dff _57893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _09191_, clk);
  dff _57894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _09194_, clk);
  dff _57895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _09198_, clk);
  dff _57896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _09201_, clk);
  dff _57897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _09204_, clk);
  dff _57898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _09207_, clk);
  dff _57899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _09209_, clk);
  dff _57900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _09164_, clk);
  dff _57901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _09167_, clk);
  dff _57902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _09170_, clk);
  dff _57903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _09173_, clk);
  dff _57904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _09176_, clk);
  dff _57905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _09179_, clk);
  dff _57906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _09182_, clk);
  dff _57907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _09185_, clk);
  dff _57908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _09138_, clk);
  dff _57909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _09141_, clk);
  dff _57910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _09145_, clk);
  dff _57911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _09148_, clk);
  dff _57912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _09151_, clk);
  dff _57913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _09154_, clk);
  dff _57914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _09157_, clk);
  dff _57915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _09159_, clk);
  dff _57916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _09114_, clk);
  dff _57917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _09117_, clk);
  dff _57918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _09120_, clk);
  dff _57919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _09123_, clk);
  dff _57920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _09126_, clk);
  dff _57921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _09129_, clk);
  dff _57922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _09132_, clk);
  dff _57923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _09135_, clk);
  dff _57924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _09089_, clk);
  dff _57925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _09093_, clk);
  dff _57926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _09096_, clk);
  dff _57927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _09099_, clk);
  dff _57928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _09102_, clk);
  dff _57929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _09105_, clk);
  dff _57930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _09108_, clk);
  dff _57931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _09110_, clk);
  dff _57932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _09065_, clk);
  dff _57933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _09068_, clk);
  dff _57934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _09071_, clk);
  dff _57935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _09074_, clk);
  dff _57936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _09077_, clk);
  dff _57937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _09080_, clk);
  dff _57938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _09083_, clk);
  dff _57939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _09085_, clk);
  dff _57940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _09040_, clk);
  dff _57941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _09043_, clk);
  dff _57942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _09046_, clk);
  dff _57943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _09049_, clk);
  dff _57944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _09052_, clk);
  dff _57945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _09055_, clk);
  dff _57946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _09058_, clk);
  dff _57947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _09061_, clk);
  dff _57948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _09016_, clk);
  dff _57949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _09019_, clk);
  dff _57950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _09022_, clk);
  dff _57951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _09025_, clk);
  dff _57952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _09028_, clk);
  dff _57953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _09031_, clk);
  dff _57954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _09034_, clk);
  dff _57955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _09036_, clk);
  dff _57956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _08991_, clk);
  dff _57957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _08994_, clk);
  dff _57958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _08997_, clk);
  dff _57959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _09000_, clk);
  dff _57960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _09003_, clk);
  dff _57961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _09006_, clk);
  dff _57962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _09009_, clk);
  dff _57963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _09012_, clk);
  dff _57964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _08966_, clk);
  dff _57965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _08969_, clk);
  dff _57966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _08972_, clk);
  dff _57967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _08975_, clk);
  dff _57968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _08978_, clk);
  dff _57969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _08981_, clk);
  dff _57970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _08985_, clk);
  dff _57971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _08987_, clk);
  dff _57972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _08942_, clk);
  dff _57973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _08945_, clk);
  dff _57974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _08948_, clk);
  dff _57975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _08951_, clk);
  dff _57976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _08954_, clk);
  dff _57977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _08957_, clk);
  dff _57978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _08960_, clk);
  dff _57979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _08963_, clk);
  dff _57980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _08917_, clk);
  dff _57981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _08920_, clk);
  dff _57982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _08923_, clk);
  dff _57983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _08926_, clk);
  dff _57984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _08929_, clk);
  dff _57985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _08933_, clk);
  dff _57986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _08936_, clk);
  dff _57987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _08938_, clk);
  dff _57988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _08890_, clk);
  dff _57989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _08893_, clk);
  dff _57990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _08896_, clk);
  dff _57991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _08900_, clk);
  dff _57992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _08904_, clk);
  dff _57993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _08907_, clk);
  dff _57994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _08911_, clk);
  dff _57995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _08913_, clk);
  dff _57996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _08863_, clk);
  dff _57997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _08867_, clk);
  dff _57998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _08870_, clk);
  dff _57999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _08873_, clk);
  dff _58000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _08877_, clk);
  dff _58001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _08880_, clk);
  dff _58002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _08883_, clk);
  dff _58003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _08886_, clk);
  dff _58004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _08836_, clk);
  dff _58005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _08839_, clk);
  dff _58006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _08843_, clk);
  dff _58007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _08847_, clk);
  dff _58008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _08850_, clk);
  dff _58009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _08854_, clk);
  dff _58010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _08857_, clk);
  dff _58011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _08859_, clk);
  dff _58012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _08811_, clk);
  dff _58013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _08814_, clk);
  dff _58014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _08818_, clk);
  dff _58015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _08821_, clk);
  dff _58016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _08824_, clk);
  dff _58017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _08827_, clk);
  dff _58018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _08830_, clk);
  dff _58019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _08832_, clk);
  dff _58020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _08786_, clk);
  dff _58021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _08790_, clk);
  dff _58022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _08793_, clk);
  dff _58023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _08796_, clk);
  dff _58024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _08799_, clk);
  dff _58025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _08802_, clk);
  dff _58026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _08805_, clk);
  dff _58027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _08807_, clk);
  dff _58028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _08762_, clk);
  dff _58029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _08765_, clk);
  dff _58030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _08768_, clk);
  dff _58031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _08771_, clk);
  dff _58032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _08774_, clk);
  dff _58033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _08777_, clk);
  dff _58034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _08780_, clk);
  dff _58035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _08783_, clk);
  dff _58036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _08737_, clk);
  dff _58037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _08740_, clk);
  dff _58038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _08743_, clk);
  dff _58039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _08746_, clk);
  dff _58040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _08749_, clk);
  dff _58041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _08752_, clk);
  dff _58042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _08755_, clk);
  dff _58043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _08757_, clk);
  dff _58044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _08712_, clk);
  dff _58045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _08715_, clk);
  dff _58046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _08718_, clk);
  dff _58047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _08721_, clk);
  dff _58048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _08724_, clk);
  dff _58049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _08727_, clk);
  dff _58050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _08730_, clk);
  dff _58051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _08733_, clk);
  dff _58052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _08688_, clk);
  dff _58053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _08691_, clk);
  dff _58054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _08694_, clk);
  dff _58055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _08697_, clk);
  dff _58056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _08700_, clk);
  dff _58057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _08703_, clk);
  dff _58058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _08706_, clk);
  dff _58059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _08708_, clk);
  dff _58060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _08663_, clk);
  dff _58061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _08666_, clk);
  dff _58062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _08669_, clk);
  dff _58063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _08672_, clk);
  dff _58064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _08675_, clk);
  dff _58065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _08678_, clk);
  dff _58066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _08681_, clk);
  dff _58067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _08684_, clk);
  dff _58068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _08638_, clk);
  dff _58069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _08641_, clk);
  dff _58070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _08644_, clk);
  dff _58071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _08647_, clk);
  dff _58072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _08650_, clk);
  dff _58073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _08653_, clk);
  dff _58074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _08657_, clk);
  dff _58075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _08659_, clk);
  dff _58076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _08614_, clk);
  dff _58077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _08617_, clk);
  dff _58078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _08620_, clk);
  dff _58079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _08623_, clk);
  dff _58080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _08626_, clk);
  dff _58081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _08629_, clk);
  dff _58082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _08632_, clk);
  dff _58083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _08635_, clk);
  dff _58084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _08589_, clk);
  dff _58085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _08592_, clk);
  dff _58086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _08595_, clk);
  dff _58087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _08598_, clk);
  dff _58088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _08601_, clk);
  dff _58089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _08605_, clk);
  dff _58090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _08608_, clk);
  dff _58091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _08610_, clk);
  dff _58092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _08564_, clk);
  dff _58093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _08567_, clk);
  dff _58094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _08570_, clk);
  dff _58095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _08573_, clk);
  dff _58096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _08577_, clk);
  dff _58097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _08580_, clk);
  dff _58098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _08583_, clk);
  dff _58099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _08585_, clk);
  dff _58100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _08540_, clk);
  dff _58101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _08543_, clk);
  dff _58102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _08546_, clk);
  dff _58103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _08549_, clk);
  dff _58104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _08552_, clk);
  dff _58105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _08555_, clk);
  dff _58106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _08558_, clk);
  dff _58107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _08561_, clk);
  dff _58108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _08515_, clk);
  dff _58109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _08518_, clk);
  dff _58110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _08521_, clk);
  dff _58111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _08525_, clk);
  dff _58112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _08528_, clk);
  dff _58113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _08531_, clk);
  dff _58114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _08534_, clk);
  dff _58115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _08536_, clk);
  dff _58116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _08490_, clk);
  dff _58117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _08493_, clk);
  dff _58118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _08497_, clk);
  dff _58119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _08500_, clk);
  dff _58120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _08503_, clk);
  dff _58121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _08506_, clk);
  dff _58122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _08509_, clk);
  dff _58123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _08511_, clk);
  dff _58124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _08466_, clk);
  dff _58125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _08469_, clk);
  dff _58126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _08472_, clk);
  dff _58127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _08475_, clk);
  dff _58128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _08478_, clk);
  dff _58129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _08481_, clk);
  dff _58130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _08484_, clk);
  dff _58131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _08487_, clk);
  dff _58132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _08441_, clk);
  dff _58133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _08445_, clk);
  dff _58134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _08448_, clk);
  dff _58135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _08451_, clk);
  dff _58136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _08454_, clk);
  dff _58137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _08457_, clk);
  dff _58138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _08460_, clk);
  dff _58139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _08462_, clk);
  dff _58140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _08417_, clk);
  dff _58141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _08420_, clk);
  dff _58142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _08423_, clk);
  dff _58143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _08426_, clk);
  dff _58144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _08429_, clk);
  dff _58145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _08432_, clk);
  dff _58146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _08435_, clk);
  dff _58147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _08437_, clk);
  dff _58148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _08392_, clk);
  dff _58149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _08395_, clk);
  dff _58150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _08398_, clk);
  dff _58151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _08401_, clk);
  dff _58152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _08404_, clk);
  dff _58153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _08407_, clk);
  dff _58154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _08410_, clk);
  dff _58155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _08412_, clk);
  dff _58156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _08367_, clk);
  dff _58157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _08370_, clk);
  dff _58158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _08373_, clk);
  dff _58159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _08376_, clk);
  dff _58160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _08379_, clk);
  dff _58161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _08382_, clk);
  dff _58162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _08385_, clk);
  dff _58163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _08388_, clk);
  dff _58164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _08341_, clk);
  dff _58165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _08344_, clk);
  dff _58166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _08347_, clk);
  dff _58167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _08350_, clk);
  dff _58168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _08353_, clk);
  dff _58169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _08356_, clk);
  dff _58170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _08359_, clk);
  dff _58171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _08362_, clk);
  dff _58172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _08317_, clk);
  dff _58173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _08320_, clk);
  dff _58174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _08323_, clk);
  dff _58175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _08326_, clk);
  dff _58176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _08329_, clk);
  dff _58177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _08332_, clk);
  dff _58178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _08335_, clk);
  dff _58179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _08338_, clk);
  dff _58180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _08292_, clk);
  dff _58181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _08295_, clk);
  dff _58182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _08298_, clk);
  dff _58183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _08301_, clk);
  dff _58184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _08304_, clk);
  dff _58185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _08307_, clk);
  dff _58186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _08311_, clk);
  dff _58187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _08313_, clk);
  dff _58188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _08267_, clk);
  dff _58189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _08270_, clk);
  dff _58190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _08273_, clk);
  dff _58191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _08276_, clk);
  dff _58192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _08279_, clk);
  dff _58193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _08283_, clk);
  dff _58194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _08286_, clk);
  dff _58195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _08288_, clk);
  dff _58196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _06413_, clk);
  dff _58197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _06416_, clk);
  dff _58198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _06419_, clk);
  dff _58199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _06422_, clk);
  dff _58200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _06425_, clk);
  dff _58201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _06428_, clk);
  dff _58202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _06431_, clk);
  dff _58203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _06434_, clk);
  dff _58204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _06215_, clk);
  dff _58205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _06218_, clk);
  dff _58206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _06221_, clk);
  dff _58207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _06224_, clk);
  dff _58208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _06227_, clk);
  dff _58209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _06230_, clk);
  dff _58210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _06233_, clk);
  dff _58211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _06236_, clk);
  dff _58212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _05869_, clk);
  dff _58213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _05872_, clk);
  dff _58214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _05876_, clk);
  dff _58215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _05879_, clk);
  dff _58216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _05882_, clk);
  dff _58217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _05885_, clk);
  dff _58218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _05888_, clk);
  dff _58219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _05890_, clk);
  dff _58220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _05844_, clk);
  dff _58221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _05848_, clk);
  dff _58222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _05851_, clk);
  dff _58223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _05854_, clk);
  dff _58224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _05857_, clk);
  dff _58225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _05860_, clk);
  dff _58226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _05863_, clk);
  dff _58227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _05866_, clk);
  dff _58228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _05820_, clk);
  dff _58229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _05823_, clk);
  dff _58230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _05826_, clk);
  dff _58231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _05829_, clk);
  dff _58232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _05832_, clk);
  dff _58233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _05835_, clk);
  dff _58234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _05838_, clk);
  dff _58235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _05841_, clk);
  dff _58236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _05796_, clk);
  dff _58237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _05799_, clk);
  dff _58238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _05802_, clk);
  dff _58239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _05805_, clk);
  dff _58240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _05808_, clk);
  dff _58241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _05811_, clk);
  dff _58242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _05814_, clk);
  dff _58243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _05816_, clk);
  dff _58244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _05771_, clk);
  dff _58245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _05774_, clk);
  dff _58246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _05777_, clk);
  dff _58247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _05780_, clk);
  dff _58248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _05783_, clk);
  dff _58249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _05786_, clk);
  dff _58250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _05789_, clk);
  dff _58251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _05791_, clk);
  dff _58252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _05746_, clk);
  dff _58253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _05749_, clk);
  dff _58254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _05752_, clk);
  dff _58255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _05755_, clk);
  dff _58256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _05758_, clk);
  dff _58257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _05761_, clk);
  dff _58258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _05764_, clk);
  dff _58259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _05767_, clk);
  dff _58260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _05722_, clk);
  dff _58261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _05725_, clk);
  dff _58262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _05728_, clk);
  dff _58263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _05731_, clk);
  dff _58264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _05734_, clk);
  dff _58265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _05737_, clk);
  dff _58266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _05740_, clk);
  dff _58267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _05743_, clk);
  dff _58268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _05697_, clk);
  dff _58269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _05700_, clk);
  dff _58270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _05703_, clk);
  dff _58271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _05706_, clk);
  dff _58272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _05709_, clk);
  dff _58273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _05712_, clk);
  dff _58274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _05716_, clk);
  dff _58275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _05718_, clk);
  dff _58276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _05672_, clk);
  dff _58277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _05675_, clk);
  dff _58278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _05678_, clk);
  dff _58279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _05681_, clk);
  dff _58280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _05684_, clk);
  dff _58281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _05688_, clk);
  dff _58282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _05691_, clk);
  dff _58283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _05693_, clk);
  dff _58284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _05648_, clk);
  dff _58285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _05651_, clk);
  dff _58286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _05654_, clk);
  dff _58287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _05657_, clk);
  dff _58288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _05660_, clk);
  dff _58289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _05663_, clk);
  dff _58290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _05666_, clk);
  dff _58291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _05669_, clk);
  dff _58292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _05623_, clk);
  dff _58293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _05626_, clk);
  dff _58294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _05629_, clk);
  dff _58295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _05632_, clk);
  dff _58296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _05636_, clk);
  dff _58297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _05639_, clk);
  dff _58298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _05642_, clk);
  dff _58299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _05644_, clk);
  dff _58300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _05598_, clk);
  dff _58301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _05601_, clk);
  dff _58302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _05604_, clk);
  dff _58303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _05608_, clk);
  dff _58304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _05611_, clk);
  dff _58305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _05614_, clk);
  dff _58306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _05617_, clk);
  dff _58307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _05619_, clk);
  dff _58308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _05573_, clk);
  dff _58309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _05576_, clk);
  dff _58310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _05579_, clk);
  dff _58311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _05583_, clk);
  dff _58312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _05586_, clk);
  dff _58313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _05589_, clk);
  dff _58314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _05592_, clk);
  dff _58315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _05594_, clk);
  dff _58316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _05548_, clk);
  dff _58317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _05551_, clk);
  dff _58318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _05555_, clk);
  dff _58319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _05558_, clk);
  dff _58320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _05561_, clk);
  dff _58321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _05564_, clk);
  dff _58322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _05567_, clk);
  dff _58323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _05569_, clk);
  dff _58324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _05524_, clk);
  dff _58325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _05527_, clk);
  dff _58326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _05530_, clk);
  dff _58327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _05533_, clk);
  dff _58328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _05536_, clk);
  dff _58329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _05539_, clk);
  dff _58330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _05542_, clk);
  dff _58331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _05545_, clk);
  dff _58332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _05499_, clk);
  dff _58333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _05503_, clk);
  dff _58334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _05506_, clk);
  dff _58335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _05509_, clk);
  dff _58336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _05512_, clk);
  dff _58337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _05515_, clk);
  dff _58338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _05518_, clk);
  dff _58339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _05520_, clk);
  dff _58340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _04580_, clk);
  dff _58341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _04583_, clk);
  dff _58342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _04586_, clk);
  dff _58343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _04589_, clk);
  dff _58344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _04592_, clk);
  dff _58345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _04595_, clk);
  dff _58346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _04598_, clk);
  dff _58347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _04601_, clk);
  dff _58348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _04930_, clk);
  dff _58349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _04933_, clk);
  dff _58350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _04936_, clk);
  dff _58351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _04939_, clk);
  dff _58352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _04942_, clk);
  dff _58353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _04945_, clk);
  dff _58354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _04948_, clk);
  dff _58355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _04951_, clk);
  dff _58356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _04554_, clk);
  dff _58357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _04557_, clk);
  dff _58358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _04561_, clk);
  dff _58359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _04565_, clk);
  dff _58360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _04568_, clk);
  dff _58361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _04571_, clk);
  dff _58362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _04574_, clk);
  dff _58363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _04576_, clk);
  dff _58364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _04904_, clk);
  dff _58365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _04907_, clk);
  dff _58366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _04910_, clk);
  dff _58367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _04915_, clk);
  dff _58368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _04918_, clk);
  dff _58369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _04921_, clk);
  dff _58370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _04924_, clk);
  dff _58371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _04926_, clk);
  dff _58372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _04529_, clk);
  dff _58373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _04533_, clk);
  dff _58374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _04536_, clk);
  dff _58375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _04539_, clk);
  dff _58376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _04542_, clk);
  dff _58377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _04545_, clk);
  dff _58378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _04548_, clk);
  dff _58379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _04550_, clk);
  dff _58380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _04879_, clk);
  dff _58381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _04882_, clk);
  dff _58382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _04886_, clk);
  dff _58383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _04889_, clk);
  dff _58384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _04892_, clk);
  dff _58385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _04895_, clk);
  dff _58386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _04898_, clk);
  dff _58387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _04900_, clk);
  dff _58388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _04505_, clk);
  dff _58389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _04508_, clk);
  dff _58390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _04511_, clk);
  dff _58391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _04514_, clk);
  dff _58392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _04517_, clk);
  dff _58393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _04520_, clk);
  dff _58394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _04523_, clk);
  dff _58395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _04526_, clk);
  dff _58396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _04480_, clk);
  dff _58397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _04483_, clk);
  dff _58398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _04486_, clk);
  dff _58399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _04489_, clk);
  dff _58400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _04492_, clk);
  dff _58401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _04495_, clk);
  dff _58402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _04498_, clk);
  dff _58403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _04501_, clk);
  dff _58404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _04455_, clk);
  dff _58405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _04458_, clk);
  dff _58406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _04461_, clk);
  dff _58407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _04464_, clk);
  dff _58408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _04467_, clk);
  dff _58409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _04470_, clk);
  dff _58410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _04473_, clk);
  dff _58411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _04475_, clk);
  dff _58412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _04430_, clk);
  dff _58413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _04433_, clk);
  dff _58414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _04436_, clk);
  dff _58415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _04439_, clk);
  dff _58416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _04442_, clk);
  dff _58417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _04445_, clk);
  dff _58418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _04448_, clk);
  dff _58419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _04451_, clk);
  dff _58420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _04406_, clk);
  dff _58421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _04409_, clk);
  dff _58422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _04412_, clk);
  dff _58423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _04415_, clk);
  dff _58424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _04418_, clk);
  dff _58425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _04421_, clk);
  dff _58426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _04424_, clk);
  dff _58427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _04427_, clk);
  dff _58428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _04377_, clk);
  dff _58429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _04380_, clk);
  dff _58430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _04383_, clk);
  dff _58431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _04386_, clk);
  dff _58432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _04389_, clk);
  dff _58433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _04392_, clk);
  dff _58434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _04395_, clk);
  dff _58435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _04399_, clk);
  dff _58436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _04353_, clk);
  dff _58437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _04356_, clk);
  dff _58438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _04359_, clk);
  dff _58439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _04362_, clk);
  dff _58440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _04365_, clk);
  dff _58441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _04368_, clk);
  dff _58442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _04371_, clk);
  dff _58443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _04374_, clk);
  dff _58444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _04328_, clk);
  dff _58445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _04331_, clk);
  dff _58446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _04334_, clk);
  dff _58447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _04337_, clk);
  dff _58448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _04340_, clk);
  dff _58449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _04343_, clk);
  dff _58450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _04347_, clk);
  dff _58451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _04349_, clk);
  dff _58452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _04303_, clk);
  dff _58453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04306_, clk);
  dff _58454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04309_, clk);
  dff _58455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04312_, clk);
  dff _58456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _04315_, clk);
  dff _58457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _04319_, clk);
  dff _58458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _04322_, clk);
  dff _58459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _04324_, clk);
  dff _58460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04204_, clk);
  dff _58461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _04207_, clk);
  dff _58462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _04210_, clk);
  dff _58463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _04213_, clk);
  dff _58464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _04216_, clk);
  dff _58465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _04219_, clk);
  dff _58466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _04222_, clk);
  dff _58467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _04225_, clk);
  dff _58468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _06117_, clk);
  dff _58469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _06120_, clk);
  dff _58470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _06123_, clk);
  dff _58471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _06126_, clk);
  dff _58472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _06129_, clk);
  dff _58473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _06132_, clk);
  dff _58474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _06135_, clk);
  dff _58475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _06137_, clk);
  dff _58476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _07946_, clk);
  dff _58477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _07949_, clk);
  dff _58478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _07952_, clk);
  dff _58479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _07955_, clk);
  dff _58480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _07958_, clk);
  dff _58481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _07962_, clk);
  dff _58482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _07965_, clk);
  dff _58483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _07967_, clk);
  dff _58484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _07675_, clk);
  dff _58485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _07678_, clk);
  dff _58486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _07681_, clk);
  dff _58487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _07684_, clk);
  dff _58488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _07687_, clk);
  dff _58489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _07690_, clk);
  dff _58490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _07694_, clk);
  dff _58491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _07696_, clk);
  dff _58492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _07651_, clk);
  dff _58493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _07654_, clk);
  dff _58494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _07657_, clk);
  dff _58495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _07660_, clk);
  dff _58496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _07663_, clk);
  dff _58497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _07666_, clk);
  dff _58498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _07669_, clk);
  dff _58499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _07672_, clk);
  dff _58500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _06935_, clk);
  dff _58501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _06938_, clk);
  dff _58502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _06941_, clk);
  dff _58503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _06944_, clk);
  dff _58504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06947_, clk);
  dff _58505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06950_, clk);
  dff _58506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _06953_, clk);
  dff _58507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _06956_, clk);
  dff _58508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _06984_, clk);
  dff _58509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06987_, clk);
  dff _58510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _06990_, clk);
  dff _58511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06993_, clk);
  dff _58512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _06996_, clk);
  dff _58513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _07000_, clk);
  dff _58514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07003_, clk);
  dff _58515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _07005_, clk);
  dff _58516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _06959_, clk);
  dff _58517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06962_, clk);
  dff _58518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _06965_, clk);
  dff _58519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _06968_, clk);
  dff _58520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06972_, clk);
  dff _58521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _06975_, clk);
  dff _58522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _06978_, clk);
  dff _58523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _06980_, clk);
  dff _58524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _06685_, clk);
  dff _58525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _06688_, clk);
  dff _58526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06691_, clk);
  dff _58527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _06694_, clk);
  dff _58528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _06697_, clk);
  dff _58529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _06700_, clk);
  dff _58530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _06703_, clk);
  dff _58531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _06706_, clk);
  dff _58532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _06660_, clk);
  dff _58533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _06663_, clk);
  dff _58534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _06666_, clk);
  dff _58535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _06669_, clk);
  dff _58536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _06672_, clk);
  dff _58537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _06675_, clk);
  dff _58538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _06679_, clk);
  dff _58539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _06681_, clk);
  dff _58540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _06092_, clk);
  dff _58541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _06095_, clk);
  dff _58542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _06098_, clk);
  dff _58543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _06101_, clk);
  dff _58544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _06104_, clk);
  dff _58545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _06107_, clk);
  dff _58546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _06110_, clk);
  dff _58547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _06112_, clk);
  dff _58548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _06141_, clk);
  dff _58549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _06144_, clk);
  dff _58550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _06147_, clk);
  dff _58551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _06150_, clk);
  dff _58552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _06153_, clk);
  dff _58553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _06156_, clk);
  dff _58554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _06159_, clk);
  dff _58555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _06162_, clk);
  dff _58556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _05351_, clk);
  dff _58557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _05354_, clk);
  dff _58558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _05357_, clk);
  dff _58559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _05360_, clk);
  dff _58560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _05363_, clk);
  dff _58561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _05367_, clk);
  dff _58562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _05370_, clk);
  dff _58563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _05372_, clk);
  dff _58564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _05203_, clk);
  dff _58565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _05207_, clk);
  dff _58566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _05210_, clk);
  dff _58567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _05213_, clk);
  dff _58568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _05216_, clk);
  dff _58569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _05219_, clk);
  dff _58570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _05222_, clk);
  dff _58571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _05224_, clk);
  dff _58572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _05053_, clk);
  dff _58573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _05056_, clk);
  dff _58574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _05059_, clk);
  dff _58575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _05062_, clk);
  dff _58576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _05065_, clk);
  dff _58577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _05068_, clk);
  dff _58578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _05071_, clk);
  dff _58579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _05074_, clk);
  dff _58580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _05176_, clk);
  dff _58581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _05179_, clk);
  dff _58582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _05183_, clk);
  dff _58583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _05186_, clk);
  dff _58584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _05189_, clk);
  dff _58585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _05192_, clk);
  dff _58586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _05195_, clk);
  dff _58587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _05197_, clk);
  dff _58588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _05151_, clk);
  dff _58589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _05155_, clk);
  dff _58590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _05158_, clk);
  dff _58591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _05161_, clk);
  dff _58592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _05164_, clk);
  dff _58593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _05167_, clk);
  dff _58594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _05170_, clk);
  dff _58595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _05172_, clk);
  dff _58596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _05127_, clk);
  dff _58597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _05130_, clk);
  dff _58598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _05133_, clk);
  dff _58599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _05136_, clk);
  dff _58600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _05139_, clk);
  dff _58601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _05142_, clk);
  dff _58602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _05145_, clk);
  dff _58603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _05148_, clk);
  dff _58604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _05103_, clk);
  dff _58605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _05106_, clk);
  dff _58606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _05109_, clk);
  dff _58607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _05112_, clk);
  dff _58608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _05115_, clk);
  dff _58609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _05118_, clk);
  dff _58610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _05121_, clk);
  dff _58611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _05123_, clk);
  dff _58612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _05078_, clk);
  dff _58613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _05081_, clk);
  dff _58614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _05084_, clk);
  dff _58615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _05087_, clk);
  dff _58616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _05090_, clk);
  dff _58617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _05093_, clk);
  dff _58618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _05096_, clk);
  dff _58619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _05098_, clk);
  dff _58620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _05029_, clk);
  dff _58621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _05032_, clk);
  dff _58622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _05035_, clk);
  dff _58623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _05038_, clk);
  dff _58624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _05041_, clk);
  dff _58625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _05044_, clk);
  dff _58626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _05047_, clk);
  dff _58627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _05050_, clk);
  dff _58628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _05004_, clk);
  dff _58629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _05007_, clk);
  dff _58630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _05010_, clk);
  dff _58631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _05013_, clk);
  dff _58632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _05016_, clk);
  dff _58633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _05019_, clk);
  dff _58634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _05023_, clk);
  dff _58635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _05025_, clk);
  dff _58636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _04979_, clk);
  dff _58637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _04982_, clk);
  dff _58638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _04985_, clk);
  dff _58639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _04988_, clk);
  dff _58640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _04991_, clk);
  dff _58641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _04995_, clk);
  dff _58642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _04998_, clk);
  dff _58643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _05000_, clk);
  dff _58644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _04954_, clk);
  dff _58645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _04957_, clk);
  dff _58646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _04960_, clk);
  dff _58647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _04963_, clk);
  dff _58648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _04967_, clk);
  dff _58649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _04970_, clk);
  dff _58650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _04973_, clk);
  dff _58651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _04975_, clk);
  dff _58652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _04178_, clk);
  dff _58653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _04181_, clk);
  dff _58654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _04185_, clk);
  dff _58655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _04188_, clk);
  dff _58656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _04192_, clk);
  dff _58657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _04195_, clk);
  dff _58658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _04198_, clk);
  dff _58659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _04200_, clk);
  dff _58660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _04153_, clk);
  dff _58661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _04157_, clk);
  dff _58662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _04160_, clk);
  dff _58663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _04163_, clk);
  dff _58664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _04166_, clk);
  dff _58665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _04169_, clk);
  dff _58666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _04172_, clk);
  dff _58667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _04174_, clk);
  dff _58668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _04129_, clk);
  dff _58669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _04132_, clk);
  dff _58670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _04135_, clk);
  dff _58671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _04138_, clk);
  dff _58672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _04141_, clk);
  dff _58673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _04144_, clk);
  dff _58674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _04147_, clk);
  dff _58675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _04150_, clk);
  dff _58676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _04104_, clk);
  dff _58677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _04107_, clk);
  dff _58678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _04110_, clk);
  dff _58679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _04113_, clk);
  dff _58680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _04116_, clk);
  dff _58681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _04119_, clk);
  dff _58682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _04122_, clk);
  dff _58683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _04124_, clk);
  dff _58684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _04079_, clk);
  dff _58685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _04082_, clk);
  dff _58686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _04085_, clk);
  dff _58687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _04088_, clk);
  dff _58688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _04091_, clk);
  dff _58689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _04094_, clk);
  dff _58690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _04097_, clk);
  dff _58691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _04100_, clk);
  dff _58692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _08243_, clk);
  dff _58693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _08246_, clk);
  dff _58694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _08249_, clk);
  dff _58695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _08252_, clk);
  dff _58696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _08255_, clk);
  dff _58697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _08258_, clk);
  dff _58698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _08261_, clk);
  dff _58699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _08264_, clk);
  dff _58700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _08218_, clk);
  dff _58701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _08221_, clk);
  dff _58702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _08224_, clk);
  dff _58703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _08227_, clk);
  dff _58704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _08231_, clk);
  dff _58705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _08234_, clk);
  dff _58706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _08237_, clk);
  dff _58707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _08239_, clk);
  dff _58708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _08193_, clk);
  dff _58709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _08196_, clk);
  dff _58710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _08199_, clk);
  dff _58711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _08203_, clk);
  dff _58712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _08206_, clk);
  dff _58713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _08209_, clk);
  dff _58714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _08212_, clk);
  dff _58715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _08214_, clk);
  dff _58716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _08169_, clk);
  dff _58717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _08172_, clk);
  dff _58718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _08175_, clk);
  dff _58719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _08178_, clk);
  dff _58720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _08181_, clk);
  dff _58721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _08184_, clk);
  dff _58722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _08187_, clk);
  dff _58723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _08190_, clk);
  dff _58724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _08144_, clk);
  dff _58725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _08147_, clk);
  dff _58726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _08151_, clk);
  dff _58727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _08154_, clk);
  dff _58728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _08157_, clk);
  dff _58729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _08160_, clk);
  dff _58730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _08163_, clk);
  dff _58731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _08165_, clk);
  dff _58732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _08119_, clk);
  dff _58733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _08123_, clk);
  dff _58734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _08126_, clk);
  dff _58735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _08129_, clk);
  dff _58736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _08132_, clk);
  dff _58737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _08135_, clk);
  dff _58738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _08138_, clk);
  dff _58739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _08140_, clk);
  dff _58740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _08095_, clk);
  dff _58741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _08098_, clk);
  dff _58742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _08101_, clk);
  dff _58743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _08104_, clk);
  dff _58744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _08107_, clk);
  dff _58745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _08110_, clk);
  dff _58746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _08113_, clk);
  dff _58747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _08116_, clk);
  dff _58748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _08071_, clk);
  dff _58749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _08074_, clk);
  dff _58750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _08077_, clk);
  dff _58751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _08080_, clk);
  dff _58752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _08083_, clk);
  dff _58753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _08086_, clk);
  dff _58754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _08089_, clk);
  dff _58755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _08091_, clk);
  dff _58756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _07921_, clk);
  dff _58757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _07924_, clk);
  dff _58758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _07927_, clk);
  dff _58759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _07930_, clk);
  dff _58760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _07934_, clk);
  dff _58761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _07937_, clk);
  dff _58762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _07940_, clk);
  dff _58763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _07942_, clk);
  dff _58764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _08046_, clk);
  dff _58765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _08049_, clk);
  dff _58766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _08052_, clk);
  dff _58767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _08055_, clk);
  dff _58768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _08058_, clk);
  dff _58769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _08061_, clk);
  dff _58770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _08064_, clk);
  dff _58771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _08066_, clk);
  dff _58772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _08021_, clk);
  dff _58773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _08024_, clk);
  dff _58774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _08027_, clk);
  dff _58775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _08030_, clk);
  dff _58776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _08033_, clk);
  dff _58777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _08036_, clk);
  dff _58778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _08039_, clk);
  dff _58779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _08042_, clk);
  dff _58780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _07971_, clk);
  dff _58781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _07974_, clk);
  dff _58782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _07977_, clk);
  dff _58783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _07980_, clk);
  dff _58784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _07983_, clk);
  dff _58785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _07987_, clk);
  dff _58786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _07991_, clk);
  dff _58787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _07993_, clk);
  dff _58788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _07997_, clk);
  dff _58789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _08000_, clk);
  dff _58790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _08003_, clk);
  dff _58791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _08006_, clk);
  dff _58792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _08009_, clk);
  dff _58793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _08012_, clk);
  dff _58794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _08015_, clk);
  dff _58795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _08018_, clk);
  dff _58796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _07897_, clk);
  dff _58797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _07900_, clk);
  dff _58798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _07903_, clk);
  dff _58799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _07906_, clk);
  dff _58800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _07909_, clk);
  dff _58801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _07912_, clk);
  dff _58802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _07915_, clk);
  dff _58803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _07918_, clk);
  dff _58804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _07872_, clk);
  dff _58805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _07875_, clk);
  dff _58806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _07878_, clk);
  dff _58807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _07882_, clk);
  dff _58808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _07885_, clk);
  dff _58809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _07888_, clk);
  dff _58810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _07891_, clk);
  dff _58811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _07893_, clk);
  dff _58812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _07823_, clk);
  dff _58813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _07826_, clk);
  dff _58814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _07829_, clk);
  dff _58815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _07832_, clk);
  dff _58816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _07835_, clk);
  dff _58817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _07838_, clk);
  dff _58818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _07841_, clk);
  dff _58819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _07844_, clk);
  dff _58820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _07847_, clk);
  dff _58821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _07850_, clk);
  dff _58822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _07854_, clk);
  dff _58823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _07857_, clk);
  dff _58824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _07860_, clk);
  dff _58825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _07863_, clk);
  dff _58826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _07866_, clk);
  dff _58827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _07868_, clk);
  dff _58828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _07798_, clk);
  dff _58829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _07802_, clk);
  dff _58830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _07805_, clk);
  dff _58831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _07808_, clk);
  dff _58832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _07811_, clk);
  dff _58833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _07814_, clk);
  dff _58834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _07817_, clk);
  dff _58835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _07819_, clk);
  dff _58836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _07774_, clk);
  dff _58837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _07777_, clk);
  dff _58838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _07780_, clk);
  dff _58839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _07783_, clk);
  dff _58840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _07786_, clk);
  dff _58841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _07789_, clk);
  dff _58842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _07792_, clk);
  dff _58843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _07794_, clk);
  dff _58844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _07749_, clk);
  dff _58845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _07752_, clk);
  dff _58846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _07755_, clk);
  dff _58847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _07758_, clk);
  dff _58848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _07761_, clk);
  dff _58849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _07764_, clk);
  dff _58850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _07767_, clk);
  dff _58851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _07770_, clk);
  dff _58852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _07725_, clk);
  dff _58853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _07728_, clk);
  dff _58854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _07731_, clk);
  dff _58855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _07734_, clk);
  dff _58856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _07737_, clk);
  dff _58857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _07740_, clk);
  dff _58858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _07743_, clk);
  dff _58859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _07745_, clk);
  dff _58860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _07700_, clk);
  dff _58861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _07703_, clk);
  dff _58862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _07706_, clk);
  dff _58863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _07709_, clk);
  dff _58864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _07712_, clk);
  dff _58865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _07715_, clk);
  dff _58866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _07718_, clk);
  dff _58867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _07721_, clk);
  dff _58868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _07626_, clk);
  dff _58869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _07629_, clk);
  dff _58870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _07632_, clk);
  dff _58871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _07635_, clk);
  dff _58872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _07638_, clk);
  dff _58873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _07642_, clk);
  dff _58874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _07645_, clk);
  dff _58875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _07647_, clk);
  dff _58876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _07601_, clk);
  dff _58877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _07604_, clk);
  dff _58878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _07607_, clk);
  dff _58879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _07610_, clk);
  dff _58880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _07614_, clk);
  dff _58881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _07617_, clk);
  dff _58882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _07620_, clk);
  dff _58883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _07622_, clk);
  dff _58884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _07551_, clk);
  dff _58885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _07554_, clk);
  dff _58886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _07557_, clk);
  dff _58887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _07561_, clk);
  dff _58888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _07564_, clk);
  dff _58889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _07567_, clk);
  dff _58890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _07570_, clk);
  dff _58891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _07572_, clk);
  dff _58892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _07577_, clk);
  dff _58893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _07580_, clk);
  dff _58894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _07583_, clk);
  dff _58895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _07586_, clk);
  dff _58896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _07589_, clk);
  dff _58897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _07592_, clk);
  dff _58898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _07595_, clk);
  dff _58899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _07598_, clk);
  dff _58900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _07502_, clk);
  dff _58901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _07505_, clk);
  dff _58902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _07508_, clk);
  dff _58903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _07511_, clk);
  dff _58904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _07514_, clk);
  dff _58905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _07517_, clk);
  dff _58906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _07520_, clk);
  dff _58907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _07523_, clk);
  dff _58908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _07526_, clk);
  dff _58909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _07529_, clk);
  dff _58910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _07533_, clk);
  dff _58911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _07536_, clk);
  dff _58912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _07539_, clk);
  dff _58913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _07542_, clk);
  dff _58914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _07545_, clk);
  dff _58915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _07547_, clk);
  dff _58916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _07477_, clk);
  dff _58917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _07481_, clk);
  dff _58918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _07484_, clk);
  dff _58919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _07487_, clk);
  dff _58920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _07490_, clk);
  dff _58921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _07493_, clk);
  dff _58922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _07496_, clk);
  dff _58923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _07498_, clk);
  dff _58924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _07453_, clk);
  dff _58925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _07456_, clk);
  dff _58926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _07459_, clk);
  dff _58927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _07462_, clk);
  dff _58928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _07465_, clk);
  dff _58929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _07468_, clk);
  dff _58930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _07471_, clk);
  dff _58931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _07473_, clk);
  dff _58932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _07428_, clk);
  dff _58933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _07431_, clk);
  dff _58934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _07434_, clk);
  dff _58935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _07437_, clk);
  dff _58936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _07440_, clk);
  dff _58937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _07443_, clk);
  dff _58938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _07446_, clk);
  dff _58939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _07449_, clk);
  dff _58940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _07379_, clk);
  dff _58941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _07382_, clk);
  dff _58942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _07385_, clk);
  dff _58943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _07388_, clk);
  dff _58944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _07391_, clk);
  dff _58945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _07394_, clk);
  dff _58946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _07397_, clk);
  dff _58947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _07400_, clk);
  dff _58948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _07404_, clk);
  dff _58949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _07407_, clk);
  dff _58950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _07410_, clk);
  dff _58951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _07413_, clk);
  dff _58952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _07416_, clk);
  dff _58953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _07419_, clk);
  dff _58954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _07422_, clk);
  dff _58955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _07424_, clk);
  dff _58956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _07354_, clk);
  dff _58957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _07357_, clk);
  dff _58958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _07360_, clk);
  dff _58959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _07363_, clk);
  dff _58960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _07366_, clk);
  dff _58961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _07369_, clk);
  dff _58962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _07373_, clk);
  dff _58963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _07375_, clk);
  dff _58964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _07330_, clk);
  dff _58965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _07333_, clk);
  dff _58966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _07336_, clk);
  dff _58967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _07339_, clk);
  dff _58968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _07342_, clk);
  dff _58969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _07345_, clk);
  dff _58970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _07348_, clk);
  dff _58971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _07351_, clk);
  dff _58972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _07305_, clk);
  dff _58973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _07308_, clk);
  dff _58974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _07311_, clk);
  dff _58975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _07314_, clk);
  dff _58976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _07317_, clk);
  dff _58977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _07321_, clk);
  dff _58978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _07324_, clk);
  dff _58979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _07326_, clk);
  dff _58980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _07256_, clk);
  dff _58981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _07259_, clk);
  dff _58982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _07262_, clk);
  dff _58983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _07265_, clk);
  dff _58984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _07268_, clk);
  dff _58985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _07271_, clk);
  dff _58986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _07274_, clk);
  dff _58987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _07277_, clk);
  dff _58988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _07280_, clk);
  dff _58989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _07283_, clk);
  dff _58990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _07286_, clk);
  dff _58991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _07289_, clk);
  dff _58992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _07293_, clk);
  dff _58993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _07296_, clk);
  dff _58994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _07299_, clk);
  dff _58995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _07301_, clk);
  dff _58996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _07231_, clk);
  dff _58997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _07234_, clk);
  dff _58998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _07237_, clk);
  dff _58999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _07241_, clk);
  dff _59000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _07244_, clk);
  dff _59001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _07247_, clk);
  dff _59002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _07250_, clk);
  dff _59003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _07252_, clk);
  dff _59004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _07206_, clk);
  dff _59005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _07209_, clk);
  dff _59006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _07213_, clk);
  dff _59007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _07216_, clk);
  dff _59008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _07219_, clk);
  dff _59009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _07222_, clk);
  dff _59010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _07225_, clk);
  dff _59011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _07227_, clk);
  dff _59012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _07182_, clk);
  dff _59013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _07185_, clk);
  dff _59014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _07188_, clk);
  dff _59015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _07191_, clk);
  dff _59016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _07194_, clk);
  dff _59017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _07197_, clk);
  dff _59018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _07200_, clk);
  dff _59019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _07203_, clk);
  dff _59020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _07132_, clk);
  dff _59021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _07135_, clk);
  dff _59022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _07138_, clk);
  dff _59023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _07141_, clk);
  dff _59024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _07144_, clk);
  dff _59025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _07147_, clk);
  dff _59026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _07150_, clk);
  dff _59027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _07153_, clk);
  dff _59028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _07156_, clk);
  dff _59029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _07160_, clk);
  dff _59030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _07163_, clk);
  dff _59031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _07166_, clk);
  dff _59032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _07169_, clk);
  dff _59033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _07172_, clk);
  dff _59034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _07175_, clk);
  dff _59035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _07177_, clk);
  dff _59036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _07107_, clk);
  dff _59037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _07110_, clk);
  dff _59038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _07113_, clk);
  dff _59039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _07116_, clk);
  dff _59040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _07119_, clk);
  dff _59041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _07122_, clk);
  dff _59042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _07125_, clk);
  dff _59043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _07128_, clk);
  dff _59044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07083_, clk);
  dff _59045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _07086_, clk);
  dff _59046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _07089_, clk);
  dff _59047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _07092_, clk);
  dff _59048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _07095_, clk);
  dff _59049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07098_, clk);
  dff _59050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _07101_, clk);
  dff _59051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07103_, clk);
  dff _59052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _07058_, clk);
  dff _59053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07061_, clk);
  dff _59054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _07064_, clk);
  dff _59055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07067_, clk);
  dff _59056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _07070_, clk);
  dff _59057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _07073_, clk);
  dff _59058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07076_, clk);
  dff _59059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07079_, clk);
  dff _59060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _07033_, clk);
  dff _59061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _07036_, clk);
  dff _59062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _07039_, clk);
  dff _59063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _07042_, clk);
  dff _59064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _07045_, clk);
  dff _59065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _07048_, clk);
  dff _59066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _07052_, clk);
  dff _59067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _07054_, clk);
  dff _59068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _07009_, clk);
  dff _59069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _07012_, clk);
  dff _59070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _07015_, clk);
  dff _59071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _07018_, clk);
  dff _59072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _07021_, clk);
  dff _59073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _07024_, clk);
  dff _59074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _07027_, clk);
  dff _59075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _07030_, clk);
  dff _59076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _06885_, clk);
  dff _59077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06888_, clk);
  dff _59078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06892_, clk);
  dff _59079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _06895_, clk);
  dff _59080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _06898_, clk);
  dff _59081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _06901_, clk);
  dff _59082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _06904_, clk);
  dff _59083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _06906_, clk);
  dff _59084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _06910_, clk);
  dff _59085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _06913_, clk);
  dff _59086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06916_, clk);
  dff _59087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _06920_, clk);
  dff _59088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _06923_, clk);
  dff _59089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _06926_, clk);
  dff _59090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06929_, clk);
  dff _59091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _06931_, clk);
  dff _59092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _06861_, clk);
  dff _59093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _06864_, clk);
  dff _59094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _06867_, clk);
  dff _59095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _06870_, clk);
  dff _59096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _06873_, clk);
  dff _59097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _06876_, clk);
  dff _59098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _06879_, clk);
  dff _59099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _06882_, clk);
  dff _59100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _06836_, clk);
  dff _59101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _06840_, clk);
  dff _59102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _06843_, clk);
  dff _59103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _06846_, clk);
  dff _59104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _06849_, clk);
  dff _59105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _06852_, clk);
  dff _59106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _06855_, clk);
  dff _59107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _06857_, clk);
  dff _59108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _06812_, clk);
  dff _59109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _06815_, clk);
  dff _59110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _06818_, clk);
  dff _59111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _06821_, clk);
  dff _59112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _06824_, clk);
  dff _59113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _06827_, clk);
  dff _59114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _06830_, clk);
  dff _59115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _06832_, clk);
  dff _59116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _06759_, clk);
  dff _59117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _06762_, clk);
  dff _59118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _06765_, clk);
  dff _59119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _06768_, clk);
  dff _59120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _06771_, clk);
  dff _59121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _06774_, clk);
  dff _59122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _06777_, clk);
  dff _59123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _06780_, clk);
  dff _59124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _06787_, clk);
  dff _59125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _06790_, clk);
  dff _59126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _06793_, clk);
  dff _59127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _06796_, clk);
  dff _59128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _06799_, clk);
  dff _59129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _06802_, clk);
  dff _59130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06805_, clk);
  dff _59131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _06808_, clk);
  dff _59132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _06735_, clk);
  dff _59133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06738_, clk);
  dff _59134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _06741_, clk);
  dff _59135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06744_, clk);
  dff _59136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _06747_, clk);
  dff _59137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _06750_, clk);
  dff _59138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _06753_, clk);
  dff _59139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _06755_, clk);
  dff _59140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _06710_, clk);
  dff _59141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06713_, clk);
  dff _59142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _06716_, clk);
  dff _59143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _06719_, clk);
  dff _59144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _06722_, clk);
  dff _59145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _06725_, clk);
  dff _59146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _06728_, clk);
  dff _59147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _06730_, clk);
  dff _59148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _06511_, clk);
  dff _59149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _06514_, clk);
  dff _59150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _06518_, clk);
  dff _59151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _06521_, clk);
  dff _59152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _06525_, clk);
  dff _59153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _06528_, clk);
  dff _59154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _06531_, clk);
  dff _59155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _06533_, clk);
  dff _59156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06636_, clk);
  dff _59157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _06639_, clk);
  dff _59158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _06642_, clk);
  dff _59159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _06645_, clk);
  dff _59160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _06648_, clk);
  dff _59161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _06651_, clk);
  dff _59162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _06654_, clk);
  dff _59163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _06657_, clk);
  dff _59164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _06611_, clk);
  dff _59165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _06614_, clk);
  dff _59166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06617_, clk);
  dff _59167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06620_, clk);
  dff _59168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _06623_, clk);
  dff _59169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06627_, clk);
  dff _59170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _06630_, clk);
  dff _59171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _06632_, clk);
  dff _59172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _06586_, clk);
  dff _59173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _06589_, clk);
  dff _59174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _06592_, clk);
  dff _59175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _06595_, clk);
  dff _59176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _06599_, clk);
  dff _59177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _06602_, clk);
  dff _59178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _06605_, clk);
  dff _59179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _06607_, clk);
  dff _59180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _06537_, clk);
  dff _59181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _06540_, clk);
  dff _59182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _06543_, clk);
  dff _59183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _06547_, clk);
  dff _59184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _06550_, clk);
  dff _59185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _06553_, clk);
  dff _59186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _06556_, clk);
  dff _59187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _06558_, clk);
  dff _59188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _06562_, clk);
  dff _59189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _06565_, clk);
  dff _59190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _06568_, clk);
  dff _59191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _06571_, clk);
  dff _59192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _06574_, clk);
  dff _59193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _06577_, clk);
  dff _59194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _06580_, clk);
  dff _59195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _06583_, clk);
  dff _59196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _06363_, clk);
  dff _59197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _06366_, clk);
  dff _59198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _06369_, clk);
  dff _59199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _06372_, clk);
  dff _59200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _06375_, clk);
  dff _59201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _06378_, clk);
  dff _59202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _06381_, clk);
  dff _59203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _06384_, clk);
  dff _59204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _06389_, clk);
  dff _59205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _06392_, clk);
  dff _59206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _06395_, clk);
  dff _59207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _06398_, clk);
  dff _59208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _06401_, clk);
  dff _59209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _06404_, clk);
  dff _59210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _06407_, clk);
  dff _59211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _06409_, clk);
  dff _59212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _06190_, clk);
  dff _59213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _06193_, clk);
  dff _59214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _06197_, clk);
  dff _59215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _06200_, clk);
  dff _59216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _06203_, clk);
  dff _59217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _06206_, clk);
  dff _59218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _06209_, clk);
  dff _59219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _06211_, clk);
  dff _59220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _06165_, clk);
  dff _59221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _06169_, clk);
  dff _59222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _06172_, clk);
  dff _59223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _06175_, clk);
  dff _59224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _06178_, clk);
  dff _59225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _06181_, clk);
  dff _59226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _06184_, clk);
  dff _59227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _06186_, clk);
  dff _59228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _15236_, clk);
  dff _59229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _15238_, clk);
  dff _59230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _15240_, clk);
  dff _59231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _15242_, clk);
  dff _59232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _15244_, clk);
  dff _59233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _15246_, clk);
  dff _59234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _15248_, clk);
  dff _59235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02715_, clk);
  dff _59236_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _59237_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _59238_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _59239_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _59240_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _59241_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _59242_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _59243_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _59244_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _59245_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _59246_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _59247_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _59248_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _59249_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _59250_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _59251_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _59252_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _59253_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _59254_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _59255_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _59256_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _59257_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _59258_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _59259_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _59260_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _59261_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _59262_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _59263_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _59264_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _59265_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _59266_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _59267_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _59268_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _59269_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _25387_, clk);
  dff _59270_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _25485_, clk);
  dff _59271_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _25486_, clk);
  dff _59272_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _25487_, clk);
  dff _59273_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _25388_, clk);
  dff _59274_ (\oc8051_top_1.oc8051_sfr1.bit_out , _25389_, clk);
  dff _59275_ (\oc8051_top_1.oc8051_sfr1.wait_data , _25391_, clk);
  dff _59276_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _25488_, clk);
  dff _59277_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _25489_, clk);
  dff _59278_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _25490_, clk);
  dff _59279_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _25492_, clk);
  dff _59280_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _25493_, clk);
  dff _59281_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _25494_, clk);
  dff _59282_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _25495_, clk);
  dff _59283_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _25392_, clk);
  dff _59284_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _25393_, clk);
  dff _59285_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19498_, clk);
  dff _59286_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19508_, clk);
  dff _59287_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19518_, clk);
  dff _59288_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19528_, clk);
  dff _59289_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19539_, clk);
  dff _59290_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19549_, clk);
  dff _59291_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19559_, clk);
  dff _59292_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17824_, clk);
  dff _59293_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08841_, clk);
  dff _59294_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08853_, clk);
  dff _59295_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08864_, clk);
  dff _59296_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08876_, clk);
  dff _59297_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08887_, clk);
  dff _59298_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08898_, clk);
  dff _59299_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08909_, clk);
  dff _59300_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06524_, clk);
  dff _59301_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13683_, clk);
  dff _59302_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13694_, clk);
  dff _59303_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13705_, clk);
  dff _59304_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13716_, clk);
  dff _59305_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13727_, clk);
  dff _59306_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13738_, clk);
  dff _59307_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13749_, clk);
  dff _59308_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12743_, clk);
  dff _59309_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13760_, clk);
  dff _59310_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13771_, clk);
  dff _59311_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13782_, clk);
  dff _59312_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13793_, clk);
  dff _59313_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13804_, clk);
  dff _59314_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13815_, clk);
  dff _59315_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13826_, clk);
  dff _59316_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12764_, clk);
  dff _59317_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _27359_, clk);
  dff _59318_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _27357_, clk);
  dff _59319_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _59320_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _27355_, clk);
  dff _59321_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00142_, clk);
  dff _59322_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00144_, clk);
  dff _59323_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00146_, clk);
  dff _59324_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00148_, clk);
  dff _59325_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00150_, clk);
  dff _59326_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00152_, clk);
  dff _59327_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00154_, clk);
  dff _59328_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27353_, clk);
  dff _59329_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00156_, clk);
  dff _59330_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _27351_, clk);
  dff _59331_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _27349_, clk);
  dff _59332_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00158_, clk);
  dff _59333_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00160_, clk);
  dff _59334_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _27347_, clk);
  dff _59335_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00162_, clk);
  dff _59336_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00164_, clk);
  dff _59337_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _27345_, clk);
  dff _59338_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00166_, clk);
  dff _59339_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27343_, clk);
  dff _59340_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00168_, clk);
  dff _59341_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27341_, clk);
  dff _59342_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _27307_, clk);
  dff _59343_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _27305_, clk);
  dff _59344_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _27303_, clk);
  dff _59345_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _27301_, clk);
  dff _59346_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00170_, clk);
  dff _59347_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00172_, clk);
  dff _59348_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00174_, clk);
  dff _59349_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _27298_, clk);
  dff _59350_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00176_, clk);
  dff _59351_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00178_, clk);
  dff _59352_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00180_, clk);
  dff _59353_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00182_, clk);
  dff _59354_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00184_, clk);
  dff _59355_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00186_, clk);
  dff _59356_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00188_, clk);
  dff _59357_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _27296_, clk);
  dff _59358_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00190_, clk);
  dff _59359_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00192_, clk);
  dff _59360_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00194_, clk);
  dff _59361_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00196_, clk);
  dff _59362_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00198_, clk);
  dff _59363_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00200_, clk);
  dff _59364_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00202_, clk);
  dff _59365_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _27294_, clk);
  dff _59366_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _24987_, clk);
  dff _59367_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _24989_, clk);
  dff _59368_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _24991_, clk);
  dff _59369_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _24993_, clk);
  dff _59370_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _24995_, clk);
  dff _59371_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _24997_, clk);
  dff _59372_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _24999_, clk);
  dff _59373_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _23900_, clk);
  dff _59374_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _25001_, clk);
  dff _59375_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _25003_, clk);
  dff _59376_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _25005_, clk);
  dff _59377_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _25007_, clk);
  dff _59378_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _25009_, clk);
  dff _59379_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _25011_, clk);
  dff _59380_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _25013_, clk);
  dff _59381_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _23901_, clk);
  dff _59382_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _25015_, clk);
  dff _59383_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _25017_, clk);
  dff _59384_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _25019_, clk);
  dff _59385_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _25021_, clk);
  dff _59386_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _25023_, clk);
  dff _59387_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _25025_, clk);
  dff _59388_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _25027_, clk);
  dff _59389_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _23902_, clk);
  dff _59390_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _25029_, clk);
  dff _59391_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _25031_, clk);
  dff _59392_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _25033_, clk);
  dff _59393_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _25035_, clk);
  dff _59394_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _25037_, clk);
  dff _59395_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _25039_, clk);
  dff _59396_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _25041_, clk);
  dff _59397_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _23903_, clk);
  dff _59398_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17288_, clk);
  dff _59399_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17297_, clk);
  dff _59400_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17306_, clk);
  dff _59401_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17315_, clk);
  dff _59402_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17324_, clk);
  dff _59403_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17332_, clk);
  dff _59404_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15222_, clk);
  dff _59405_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09474_, clk);
  dff _59406_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10718_, clk);
  dff _59407_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10729_, clk);
  dff _59408_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10740_, clk);
  dff _59409_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10751_, clk);
  dff _59410_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10762_, clk);
  dff _59411_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10773_, clk);
  dff _59412_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10784_, clk);
  dff _59413_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09496_, clk);
  dff _59414_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _25436_, clk);
  dff _59415_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _25439_, clk);
  dff _59416_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _26040_, clk);
  dff _59417_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _26042_, clk);
  dff _59418_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _26044_, clk);
  dff _59419_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _26046_, clk);
  dff _59420_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _26048_, clk);
  dff _59421_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _26050_, clk);
  dff _59422_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _26052_, clk);
  dff _59423_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _25442_, clk);
  dff _59424_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _26054_, clk);
  dff _59425_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _26056_, clk);
  dff _59426_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _26058_, clk);
  dff _59427_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _26060_, clk);
  dff _59428_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _26062_, clk);
  dff _59429_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _26064_, clk);
  dff _59430_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _26066_, clk);
  dff _59431_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _25445_, clk);
  dff _59432_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _25448_, clk);
  dff _59433_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _25451_, clk);
  dff _59434_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _26068_, clk);
  dff _59435_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _26070_, clk);
  dff _59436_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _26072_, clk);
  dff _59437_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _26074_, clk);
  dff _59438_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _26076_, clk);
  dff _59439_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _26078_, clk);
  dff _59440_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _26080_, clk);
  dff _59441_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _25454_, clk);
  dff _59442_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _26082_, clk);
  dff _59443_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _26084_, clk);
  dff _59444_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _26086_, clk);
  dff _59445_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _26088_, clk);
  dff _59446_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _26090_, clk);
  dff _59447_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _26092_, clk);
  dff _59448_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _26094_, clk);
  dff _59449_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _25457_, clk);
  dff _59450_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _25460_, clk);
  dff _59451_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _26096_, clk);
  dff _59452_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _26098_, clk);
  dff _59453_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _26100_, clk);
  dff _59454_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _26102_, clk);
  dff _59455_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _26104_, clk);
  dff _59456_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _26106_, clk);
  dff _59457_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _26108_, clk);
  dff _59458_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _25463_, clk);
  dff _59459_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01640_, clk);
  dff _59460_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01643_, clk);
  dff _59461_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01646_, clk);
  dff _59462_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01649_, clk);
  dff _59463_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02203_, clk);
  dff _59464_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02205_, clk);
  dff _59465_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02207_, clk);
  dff _59466_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02209_, clk);
  dff _59467_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02211_, clk);
  dff _59468_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02213_, clk);
  dff _59469_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02215_, clk);
  dff _59470_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01652_, clk);
  dff _59471_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02217_, clk);
  dff _59472_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02219_, clk);
  dff _59473_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02221_, clk);
  dff _59474_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02223_, clk);
  dff _59475_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02225_, clk);
  dff _59476_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02227_, clk);
  dff _59477_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02229_, clk);
  dff _59478_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01655_, clk);
  dff _59479_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01658_, clk);
  dff _59480_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02231_, clk);
  dff _59481_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02233_, clk);
  dff _59482_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02235_, clk);
  dff _59483_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02237_, clk);
  dff _59484_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02239_, clk);
  dff _59485_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02241_, clk);
  dff _59486_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02243_, clk);
  dff _59487_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01661_, clk);
  dff _59488_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02245_, clk);
  dff _59489_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02247_, clk);
  dff _59490_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02249_, clk);
  dff _59491_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02251_, clk);
  dff _59492_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02253_, clk);
  dff _59493_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02255_, clk);
  dff _59494_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02257_, clk);
  dff _59495_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01664_, clk);
  dff _59496_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01667_, clk);
  dff _59497_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02259_, clk);
  dff _59498_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02261_, clk);
  dff _59499_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02263_, clk);
  dff _59500_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02265_, clk);
  dff _59501_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02267_, clk);
  dff _59502_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02269_, clk);
  dff _59503_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02271_, clk);
  dff _59504_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01670_, clk);
  dff _59505_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01239_, clk);
  dff _59506_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01241_, clk);
  dff _59507_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01243_, clk);
  dff _59508_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01245_, clk);
  dff _59509_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01247_, clk);
  dff _59510_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01248_, clk);
  dff _59511_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01250_, clk);
  dff _59512_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01252_, clk);
  dff _59513_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01254_, clk);
  dff _59514_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01256_, clk);
  dff _59515_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01258_, clk);
  dff _59516_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00612_, clk);
  dff _59517_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00587_, clk);
  dff _59518_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00590_, clk);
  dff _59519_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00593_, clk);
  dff _59520_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00595_, clk);
  dff _59521_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00598_, clk);
  dff _59522_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00601_, clk);
  dff _59523_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01260_, clk);
  dff _59524_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00604_, clk);
  dff _59525_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01262_, clk);
  dff _59526_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01264_, clk);
  dff _59527_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01266_, clk);
  dff _59528_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00607_, clk);
  dff _59529_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01267_, clk);
  dff _59530_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01269_, clk);
  dff _59531_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01271_, clk);
  dff _59532_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01273_, clk);
  dff _59533_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01275_, clk);
  dff _59534_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01277_, clk);
  dff _59535_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01279_, clk);
  dff _59536_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00610_, clk);
  dff _59537_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00615_, clk);
  dff _59538_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00617_, clk);
  dff _59539_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00620_, clk);
  dff _59540_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00623_, clk);
  dff _59541_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00626_, clk);
  dff _59542_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01281_, clk);
  dff _59543_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01282_, clk);
  dff _59544_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01284_, clk);
  dff _59545_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00629_, clk);
  dff _59546_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01286_, clk);
  dff _59547_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01288_, clk);
  dff _59548_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01290_, clk);
  dff _59549_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01292_, clk);
  dff _59550_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01294_, clk);
  dff _59551_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01296_, clk);
  dff _59552_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01297_, clk);
  dff _59553_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01299_, clk);
  dff _59554_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01301_, clk);
  dff _59555_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01303_, clk);
  dff _59556_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00632_, clk);
  dff _59557_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01305_, clk);
  dff _59558_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01307_, clk);
  dff _59559_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01309_, clk);
  dff _59560_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01310_, clk);
  dff _59561_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01312_, clk);
  dff _59562_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01314_, clk);
  dff _59563_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01316_, clk);
  dff _59564_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00635_, clk);
  dff _59565_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01318_, clk);
  dff _59566_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01320_, clk);
  dff _59567_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01322_, clk);
  dff _59568_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01323_, clk);
  dff _59569_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01325_, clk);
  dff _59570_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01327_, clk);
  dff _59571_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01329_, clk);
  dff _59572_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00637_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
