module oc8051_golden_model(
  clk,
  rst,
  step,
  RD_ROM_0_ADDR,
  RD_ROM_1_ADDR,
  RD_ROM_2_ADDR,
  ACC,
  ACC_next,
  P2,
  P2_next,
  P0,
  P0_next,
  P1,
  P1_next,
  P3,
  P3_next,
  SP,
  SP_next,
  PC,
  PC_next,
  B,
  B_next,
  DPL,
  DPL_next,
  PSW,
  PSW_next,
  DPH,
  DPH_next,
  IRAM_full,
  SBUF,
  SBUF_next,
  SCON,
  SCON_next,
  PCON,
  PCON_next,
  TCON,
  TCON_next,
  TL0,
  TL0_next,
  TL1,
  TL1_next,
  TH0,
  TH0_next,
  TH1,
  TH1_next,
  TMOD,
  TMOD_next,
  IE,
  IE_next,
  IP,
  IP_next,
  P0IN,
  P1IN,
  P2IN,
  P3IN,
  RD_ROM_0,
  RD_ROM_1,
  RD_ROM_2,
  RD_IRAM_0_ABSTR_ADDR,
  RD_IRAM_1_ABSTR_ADDR,
  RD_ROM_1_ABSTR_ADDR,
  RD_ROM_2_ABSTR_ADDR,
  RD_XRAM_0_ABSTR_ADDR,
  ACC_abstr,
  P2_abstr,
  P0_abstr,
  P1_abstr,
  P3_abstr,
  SP_abstr,
  PC_abstr,
  B_abstr,
  DPL_abstr,
  PSW_abstr,
  DPH_abstr,
  WR_COND_ABSTR_IRAM_0,
  WR_ADDR_ABSTR_IRAM_0,
  WR_DATA_ABSTR_IRAM_0,
  WR_COND_ABSTR_IRAM_1,
  WR_ADDR_ABSTR_IRAM_1,
  WR_DATA_ABSTR_IRAM_1
);
output [15:0] RD_ROM_0_ADDR;
output [15:0] RD_ROM_1_ADDR;
output [15:0] RD_ROM_2_ADDR;
output [7:0] ACC;
output [7:0] ACC_next;
output [7:0] P2;
output [7:0] P2_next;
output [7:0] P0;
output [7:0] P0_next;
output [7:0] P1;
output [7:0] P1_next;
output [7:0] P3;
output [7:0] P3_next;
output [7:0] SP;
output [7:0] SP_next;
output [15:0] PC;
output [15:0] PC_next;
output [7:0] B;
output [7:0] B_next;
output [7:0] DPL;
output [7:0] DPL_next;
output [7:0] PSW;
output [7:0] PSW_next;
output [7:0] DPH;
output [7:0] DPH_next;
output [127:0] IRAM_full;
output [7:0] SBUF;
output [7:0] SBUF_next;
output [7:0] SCON;
output [7:0] SCON_next;
output [7:0] PCON;
output [7:0] PCON_next;
output [7:0] TCON;
output [7:0] TCON_next;
output [7:0] TL0;
output [7:0] TL0_next;
output [7:0] TL1;
output [7:0] TL1_next;
output [7:0] TH0;
output [7:0] TH0_next;
output [7:0] TH1;
output [7:0] TH1_next;
output [7:0] TMOD;
output [7:0] TMOD_next;
output [7:0] IE;
output [7:0] IE_next;
output [7:0] IP;
output [7:0] IP_next;

input clk, rst, step;
input [7:0] P0IN;
input [7:0] P1IN;
input [7:0] P2IN;
input [7:0] P3IN;
input [7:0] RD_ROM_0;
input [7:0] RD_ROM_1;
input [7:0] RD_ROM_2;
input [7:0] RD_IRAM_0_ABSTR_ADDR;
input [7:0] RD_IRAM_1_ABSTR_ADDR;
input [15:0] RD_ROM_1_ABSTR_ADDR;
input [15:0] RD_ROM_2_ABSTR_ADDR;
input [15:0] RD_XRAM_0_ABSTR_ADDR;
input [7:0] ACC_abstr;
input [7:0] P2_abstr;
input [7:0] P0_abstr;
input [7:0] P1_abstr;
input [7:0] P3_abstr;
input [7:0] SP_abstr;
input [15:0] PC_abstr;
input [7:0] B_abstr;
input [7:0] DPL_abstr;
input [7:0] PSW_abstr;
input [7:0] DPH_abstr;
input WR_COND_ABSTR_IRAM_0;
input [3:0] WR_ADDR_ABSTR_IRAM_0;
input [7:0] WR_DATA_ABSTR_IRAM_0;
input WR_COND_ABSTR_IRAM_1;
input [3:0] WR_ADDR_ABSTR_IRAM_1;
input [7:0] WR_DATA_ABSTR_IRAM_1;

reg [7:0] ACC;
reg [7:0] B;
reg [7:0] DPH;
reg [7:0] DPL;
reg [7:0] IE;
reg [7:0] IP;
reg [7:0] P0;
reg [7:0] P0INREG;
reg [7:0] P1;
reg [7:0] P1INREG;
reg [7:0] P2;
reg [7:0] P2INREG;
reg [7:0] P3;
reg [7:0] P3INREG;
reg [15:0] PC;
reg [7:0] PCON;
reg [7:0] PSW;
reg [7:0] SBUF;
reg [7:0] SCON;
reg [7:0] SP;
reg [7:0] TCON;
reg [7:0] TH0;
reg [7:0] TH1;
reg [7:0] TL0;
reg [7:0] TL1;
reg [7:0] TMOD;

wire [7:0] ACC_4b;
wire [7:0] ACC_next;
wire [7:0] B_4b;
wire [7:0] B_next;
wire [7:0] DPH_4b;
wire [7:0] DPH_next;
wire [7:0] DPL_4b;
wire [7:0] DPL_next;
wire [7:0] IE_next;
wire [7:0] IP_next;
wire [7:0] P0_4b;
wire [7:0] P0_next;
wire [7:0] P1_4b;
wire [7:0] P1_next;
wire [7:0] P2_4b;
wire [7:0] P2_next;
wire [7:0] P3_4b;
wire [7:0] P3_next;
wire [7:0] PCON_next;
wire [15:0] PC_4b;
wire [15:0] PC_next;
wire [7:0] PSW_4b;
wire [7:0] PSW_next;
wire [7:0] RD_IRAM_0;
wire [7:0] RD_IRAM_0_ADDR;
wire [7:0] RD_IRAM_1;
wire [7:0] RD_IRAM_1_ADDR;
wire [7:0] RD_ROM_0;
wire [15:0] RD_ROM_0_ADDR;
wire [7:0] RD_ROM_1;
wire [15:0] RD_ROM_1_ADDR;
wire [7:0] RD_ROM_2;
wire [15:0] RD_ROM_2_ADDR;
wire [7:0] RD_XRAM_0;
wire [15:0] RD_XRAM_0_ADDR;
wire [7:0] SBUF_next;
wire [7:0] SCON_next;
wire [7:0] SP_4b;
wire [7:0] SP_next;
wire [7:0] TCON_next;
wire [7:0] TH0_next;
wire [7:0] TH1_next;
wire [7:0] TL0_next;
wire [7:0] TL1_next;
wire [7:0] TMOD_next;
wire [3:0] WR_ADDR_0_IRAM;
wire [3:0] WR_ADDR_1_IRAM;
wire WR_COND_0_IRAM;
wire WR_COND_1_IRAM;
wire [7:0] WR_DATA_0_IRAM;
wire [7:0] WR_DATA_1_IRAM;
wire [7:0] n0001;
wire n0002;
wire [2:0] n0003;
wire [1:0] n0004;
wire [2:0] n0005;
wire [7:0] n0006;
wire [7:0] n0007;
wire [3:0] n0008;
wire [7:0] n0009;
wire [3:0] n0010;
wire [7:0] n0011;
wire [7:0] n0012;
wire [0:0] n0013;
wire [0:0] n0014;
wire n0015;
wire [3:0] n0016;
wire [7:0] n0017;
wire n0018;
wire [7:0] n0019;
wire n0020;
wire [7:0] n0021;
wire n0022;
wire [7:0] n0023;
wire n0024;
wire [7:0] n0025;
wire n0026;
wire [7:0] n0027;
wire n0028;
wire [7:0] n0029;
wire n0030;
wire [7:0] n0031;
wire n0032;
wire [7:0] n0033;
wire n0034;
wire [7:0] n0035;
wire n0036;
wire [7:0] n0037;
wire n0038;
wire [7:0] n0039;
wire n0040;
wire [7:0] n0041;
wire n0042;
wire [7:0] n0043;
wire n0044;
wire [7:0] n0045;
wire n0046;
wire [7:0] n0047;
wire n0048;
wire [7:0] n0049;
wire n0050;
wire [7:0] n0051;
wire n0052;
wire [7:0] n0053;
wire n0054;
wire [7:0] n0055;
wire n0056;
wire [7:0] n0057;
wire n0058;
wire [7:0] n0059;
wire [7:0] n0060;
wire [7:0] n0061;
wire [7:0] n0062;
wire [7:0] n0063;
wire [7:0] n0064;
wire [7:0] n0065;
wire [7:0] n0066;
wire [7:0] n0067;
wire [7:0] n0068;
wire [7:0] n0069;
wire [7:0] n0070;
wire [7:0] n0071;
wire [7:0] n0072;
wire [7:0] n0073;
wire [7:0] n0074;
wire [7:0] n0075;
wire [7:0] n0076;
wire [7:0] n0077;
wire [7:0] n0078;
wire [7:0] n0079;
wire [7:0] n0080;
wire [7:0] n0081;
wire [7:0] n0082;
wire [7:0] n0083;
wire [3:0] n0084;
wire [7:0] n0085;
wire [7:0] n0086;
wire [3:0] n0087;
wire [7:0] n0088;
wire [2:0] n0089;
wire [7:0] n0090;
wire [3:0] n0091;
wire [2:0] n0092;
wire [7:0] n0093;
wire [3:0] n0094;
wire [3:0] n0095;
wire [2:0] n0096;
wire [7:0] n0097;
wire [3:0] n0098;
wire [2:0] n0099;
wire [7:0] n0100;
wire [3:0] n0101;
wire [2:0] n0102;
wire [7:0] n0103;
wire [3:0] n0104;
wire [2:0] n0105;
wire [7:0] n0106;
wire [3:0] n0107;
wire [0:0] n0108;
wire n0109;
wire [4:0] n0110;
wire [7:0] n0111;
wire [7:0] n0112;
wire [7:0] n0113;
wire [7:0] n0114;
wire [7:0] n0115;
wire [0:0] n0116;
wire n0117;
wire [3:0] n0118;
wire [2:0] n0119;
wire [7:0] n0120;
wire [7:0] n0121;
wire [7:0] n0122;
wire n0123;
wire n0124;
wire n0125;
wire n0126;
wire n0127;
wire n0128;
wire n0129;
wire n0130;
wire n0131;
wire n0132;
wire n0133;
wire [7:0] n0134;
wire [7:0] n0135;
wire [7:0] n0136;
wire [7:0] n0137;
wire [7:0] n0138;
wire [7:0] n0139;
wire [7:0] n0140;
wire [7:0] n0141;
wire [7:0] n0142;
wire [7:0] n0143;
wire [7:0] n0144;
wire [7:0] n0145;
wire [7:0] n0146;
wire [7:0] n0147;
wire [7:0] n0148;
wire [7:0] n0149;
wire [7:0] n0150;
wire [3:0] n0151;
wire [15:0] n0152;
wire [15:0] n0153;
wire [7:0] n0154;
wire [7:0] n0155;
wire [3:0] n0156;
wire [7:0] n0157;
wire [15:0] n0158;
wire [15:0] n0159;
wire [7:0] n0160;
wire [7:0] n0161;
wire [7:0] n0162;
wire [7:0] n0163;
wire [7:0] n0164;
wire [7:0] n0165;
wire [7:0] n0166;
wire [7:0] n0167;
wire [15:0] n0168;
wire [15:0] n0169;
wire [6:0] n0170;
wire [0:0] n0171;
wire [0:0] n0172;
wire [0:0] n0173;
wire [0:0] n0174;
wire [0:0] n0175;
wire [0:0] n0176;
wire [0:0] n0177;
wire [0:0] n0178;
wire [0:0] n0179;
wire [0:0] n0180;
wire [0:0] n0181;
wire [0:0] n0182;
wire [0:0] n0183;
wire [0:0] n0184;
wire [0:0] n0185;
wire [7:0] n0186;
wire [7:0] n0187;
wire [7:0] n0188;
wire [7:0] n0189;
wire [7:0] n0190;
wire [0:0] n0191;
wire n0192;
wire n0193;
wire n0194;
wire n0195;
wire n0196;
wire n0197;
wire n0198;
wire n0199;
wire n0200;
wire n0201;
wire n0202;
wire n0203;
wire n0204;
wire n0205;
wire n0206;
wire n0207;
wire n0208;
wire n0209;
wire n0210;
wire n0211;
wire n0212;
wire n0213;
wire [7:0] n0214;
wire [7:0] n0215;
wire [7:0] n0216;
wire [7:0] n0217;
wire [7:0] n0218;
wire [7:0] n0219;
wire [7:0] n0220;
wire [7:0] n0221;
wire [7:0] n0222;
wire [7:0] n0223;
wire [7:0] n0224;
wire [7:0] n0225;
wire [7:0] n0226;
wire [7:0] n0227;
wire [7:0] n0228;
wire [7:0] n0229;
wire [7:0] n0230;
wire [7:0] n0231;
wire [7:0] n0232;
wire [7:0] n0233;
wire [7:0] n0234;
wire [7:0] n0235;
wire [0:0] n0236;
wire [7:0] n0237;
wire [7:0] n0238;
wire [7:0] n0239;
wire [7:0] n0240;
wire [7:0] n0241;
wire [7:0] n0242;
wire [7:0] n0243;
wire [7:0] n0244;
wire [7:0] n0245;
wire [7:0] n0246;
wire [7:0] n0247;
wire [7:0] n0248;
wire [7:0] n0249;
wire [7:0] n0250;
wire [7:0] n0251;
wire [7:0] n0252;
wire [7:0] n0253;
wire [7:0] n0254;
wire [7:0] n0255;
wire [7:0] n0256;
wire [7:0] n0257;
wire [7:0] n0258;
wire [7:0] n0259;
wire [7:0] n0260;
wire [7:0] n0261;
wire [7:0] n0262;
wire [7:0] n0263;
wire [7:0] n0264;
wire [7:0] n0265;
wire [7:0] n0266;
wire [7:0] n0267;
wire [0:0] n0268;
wire [0:0] n0269;
wire [7:0] n0270;
wire [7:0] n0271;
wire [7:0] n0272;
wire [7:0] n0273;
wire [7:0] n0274;
wire [7:0] n0275;
wire [7:0] n0276;
wire [3:0] n0277;
wire [3:0] n0278;
wire [7:0] n0279;
wire [7:0] n0280;
wire n0281;
wire [7:0] n0282;
wire n0283;
wire [7:0] n0284;
wire n0285;
wire [7:0] n0286;
wire n0287;
wire [7:0] n0288;
wire n0289;
wire [7:0] n0290;
wire n0291;
wire [7:0] n0292;
wire n0293;
wire [7:0] n0294;
wire n0295;
wire [7:0] n0296;
wire n0297;
wire [7:0] n0298;
wire n0299;
wire [7:0] n0300;
wire n0301;
wire [7:0] n0302;
wire n0303;
wire [7:0] n0304;
wire n0305;
wire [7:0] n0306;
wire n0307;
wire [7:0] n0308;
wire n0309;
wire [7:0] n0310;
wire n0311;
wire [7:0] n0312;
wire n0313;
wire [7:0] n0314;
wire n0315;
wire [7:0] n0316;
wire n0317;
wire [7:0] n0318;
wire n0319;
wire [7:0] n0320;
wire n0321;
wire [7:0] n0322;
wire n0323;
wire [7:0] n0324;
wire n0325;
wire [7:0] n0326;
wire n0327;
wire [7:0] n0328;
wire n0329;
wire [7:0] n0330;
wire n0331;
wire [7:0] n0332;
wire n0333;
wire [7:0] n0334;
wire n0335;
wire [7:0] n0336;
wire n0337;
wire [7:0] n0338;
wire n0339;
wire [7:0] n0340;
wire n0341;
wire [7:0] n0342;
wire n0343;
wire [7:0] n0344;
wire n0345;
wire [7:0] n0346;
wire n0347;
wire [7:0] n0348;
wire n0349;
wire [7:0] n0350;
wire n0351;
wire [7:0] n0352;
wire n0353;
wire [7:0] n0354;
wire n0355;
wire [7:0] n0356;
wire n0357;
wire [7:0] n0358;
wire n0359;
wire [7:0] n0360;
wire n0361;
wire [7:0] n0362;
wire n0363;
wire [7:0] n0364;
wire n0365;
wire [7:0] n0366;
wire n0367;
wire [7:0] n0368;
wire n0369;
wire [7:0] n0370;
wire n0371;
wire [7:0] n0372;
wire n0373;
wire n0374;
wire n0375;
wire n0376;
wire n0377;
wire n0378;
wire n0379;
wire n0380;
wire [7:0] n0381;
wire n0382;
wire [7:0] n0383;
wire n0384;
wire [7:0] n0385;
wire n0386;
wire [7:0] n0387;
wire n0388;
wire [7:0] n0389;
wire n0390;
wire [7:0] n0391;
wire n0392;
wire n0393;
wire [7:0] n0394;
wire n0395;
wire [7:0] n0396;
wire n0397;
wire [7:0] n0398;
wire n0399;
wire [7:0] n0400;
wire n0401;
wire [7:0] n0402;
wire n0403;
wire [7:0] n0404;
wire n0405;
wire [7:0] n0406;
wire n0407;
wire [7:0] n0408;
wire n0409;
wire [7:0] n0410;
wire n0411;
wire [7:0] n0412;
wire n0413;
wire [7:0] n0414;
wire n0415;
wire [7:0] n0416;
wire n0417;
wire [7:0] n0418;
wire n0419;
wire [7:0] n0420;
wire n0421;
wire [7:0] n0422;
wire n0423;
wire [7:0] n0424;
wire n0425;
wire [7:0] n0426;
wire n0427;
wire [7:0] n0428;
wire n0429;
wire [7:0] n0430;
wire n0431;
wire [7:0] n0432;
wire n0433;
wire [7:0] n0434;
wire n0435;
wire [7:0] n0436;
wire n0437;
wire n0438;
wire [7:0] n0439;
wire n0440;
wire [7:0] n0441;
wire n0442;
wire [7:0] n0443;
wire n0444;
wire [7:0] n0445;
wire n0446;
wire [7:0] n0447;
wire n0448;
wire [7:0] n0449;
wire n0450;
wire [7:0] n0451;
wire n0452;
wire [7:0] n0453;
wire n0454;
wire [7:0] n0455;
wire n0456;
wire [7:0] n0457;
wire n0458;
wire [7:0] n0459;
wire n0460;
wire [7:0] n0461;
wire n0462;
wire [7:0] n0463;
wire n0464;
wire [7:0] n0465;
wire n0466;
wire [7:0] n0467;
wire n0468;
wire [7:0] n0469;
wire n0470;
wire [7:0] n0471;
wire n0472;
wire [7:0] n0473;
wire n0474;
wire [7:0] n0475;
wire n0476;
wire [7:0] n0477;
wire n0478;
wire [7:0] n0479;
wire n0480;
wire [7:0] n0481;
wire n0482;
wire [7:0] n0483;
wire n0484;
wire [7:0] n0485;
wire n0486;
wire [7:0] n0487;
wire n0488;

reg [7:0] IRAM[15:0];
reg [7:0] XRAM[65535:0];

// port: IRAM->RD_IRAM_0
// port: IRAM->RD_IRAM_1
// port: ROM->RD_ROM_0
// port: ROM->RD_ROM_1
// port: ROM->RD_ROM_2
// port: XRAM->RD_XRAM_0
// RD_IRAM_0_ADDR=(if (eq RD_ROM_0 (bv 75 8)) (concat (bv 0 3) (extract 4 3 PSW) (bv 3 3)) RD_IRAM_0_ABSTR_ADDR)
assign n0001 = 8'h4b;
assign n0002 = ( RD_ROM_0 == n0001 );
assign n0003 = 3'h0;
assign n0004 = PSW[4:3];
assign n0005 = 3'h3;
assign n0006 = { ( n0003 ), ( n0004 ), ( n0005 ) };
assign n0007 = ( n0002 ) ? ( n0006 ) : ( RD_IRAM_0_ABSTR_ADDR );
assign RD_IRAM_0_ADDR = n0007;
assign n0008 = n0007[3:0];
assign n0009 = IRAM[n0008];
assign RD_IRAM_0 = n0009;
// RD_IRAM_1_ADDR=RD_IRAM_1_ABSTR_ADDR
assign RD_IRAM_1_ADDR = RD_IRAM_1_ABSTR_ADDR;
assign n0010 = RD_IRAM_1_ABSTR_ADDR[3:0];
assign n0011 = IRAM[n0010];
assign RD_IRAM_1 = n0011;
// RD_ROM_0_ADDR=PC
assign RD_ROM_0_ADDR = PC;
// RD_ROM_1_ADDR=RD_ROM_1_ABSTR_ADDR
assign RD_ROM_1_ADDR = RD_ROM_1_ABSTR_ADDR;
// RD_ROM_2_ADDR=RD_ROM_2_ABSTR_ADDR
assign RD_ROM_2_ADDR = RD_ROM_2_ABSTR_ADDR;
// RD_XRAM_0_ADDR=RD_XRAM_0_ABSTR_ADDR
assign RD_XRAM_0_ADDR = RD_XRAM_0_ABSTR_ADDR;
assign n0012 = XRAM[RD_XRAM_0_ABSTR_ADDR];
assign RD_XRAM_0 = n0012;
// 
// ACC_00
// 
// 
// P1_00
// 
// 
// DPL_00
// 
// 
// DPH_00
// 
// 
// PC_00
// 
// 
// P2_00
// 
// 
// P3_00
// 
// 
// P0_00
// 
// 
// B_00
// 
// 
// SP_00
// 
// 
// PSW_00
// 
// 
// ACC_01
// 
// 
// P1_01
// 
// 
// DPL_01
// 
// 
// DPH_01
// 
// 
// PC_01
// 
// 
// P2_01
// 
// 
// P3_01
// 
// 
// P0_01
// 
// 
// B_01
// 
// 
// SP_01
// 
// 
// PSW_01
// 
// 
// ACC_02
// 
// 
// B_02
// 
// 
// DPL_02
// 
// 
// DPH_02
// 
// 
// PC_02
// 
// 
// P2_02
// 
// 
// P3_02
// 
// 
// P0_02
// 
// 
// P1_02
// 
// 
// SP_02
// 
// 
// PSW_02
// 
// 
// ACC_03
// 
// 
// B_03
// 
// 
// DPL_03
// 
// 
// DPH_03
// 
// 
// PC_03
// 
// 
// P2_03
// 
// 
// P3_03
// 
// 
// P0_03
// 
// 
// P1_03
// 
// 
// SP_03
// 
// 
// PSW_03
// 
// 
// ACC_04
// 
// 
// P1_04
// 
// 
// DPL_04
// 
// 
// DPH_04
// 
// 
// PC_04
// 
// 
// P2_04
// 
// 
// P3_04
// 
// 
// P0_04
// 
// 
// B_04
// 
// 
// SP_04
// 
// 
// PSW_04
// 
// 
// ACC_05
// 
// 
// P1_05
// 
// 
// DPL_05
// 
// 
// DPH_05
// 
// 
// PC_05
// 
// 
// P2_05
// 
// 
// P3_05
// 
// 
// P0_05
// 
// 
// B_05
// 
// 
// IRAM_05
// 
assign n0013 = RD_ROM_1[7:7];
assign n0014 = 1'h0;
assign n0015 = ( n0013 == n0014 );
assign n0016 = RD_ROM_1[3:0];
assign n0017 = 8'h80;
assign n0018 = ( RD_ROM_1 == n0017 );
assign n0019 = 8'h81;
assign n0020 = ( RD_ROM_1 == n0019 );
assign n0021 = 8'h82;
assign n0022 = ( RD_ROM_1 == n0021 );
assign n0023 = 8'h83;
assign n0024 = ( RD_ROM_1 == n0023 );
assign n0025 = 8'h87;
assign n0026 = ( RD_ROM_1 == n0025 );
assign n0027 = 8'h88;
assign n0028 = ( RD_ROM_1 == n0027 );
assign n0029 = 8'h89;
assign n0030 = ( RD_ROM_1 == n0029 );
assign n0031 = 8'h8a;
assign n0032 = ( RD_ROM_1 == n0031 );
assign n0033 = 8'h8c;
assign n0034 = ( RD_ROM_1 == n0033 );
assign n0035 = 8'h8b;
assign n0036 = ( RD_ROM_1 == n0035 );
assign n0037 = 8'h8d;
assign n0038 = ( RD_ROM_1 == n0037 );
assign n0039 = 8'h90;
assign n0040 = ( RD_ROM_1 == n0039 );
assign n0041 = 8'h98;
assign n0042 = ( RD_ROM_1 == n0041 );
assign n0043 = 8'h99;
assign n0044 = ( RD_ROM_1 == n0043 );
assign n0045 = 8'ha0;
assign n0046 = ( RD_ROM_1 == n0045 );
assign n0047 = 8'ha8;
assign n0048 = ( RD_ROM_1 == n0047 );
assign n0049 = 8'hb0;
assign n0050 = ( RD_ROM_1 == n0049 );
assign n0051 = 8'hb8;
assign n0052 = ( RD_ROM_1 == n0051 );
assign n0053 = 8'hd0;
assign n0054 = ( RD_ROM_1 == n0053 );
assign n0055 = 8'he0;
assign n0056 = ( RD_ROM_1 == n0055 );
assign n0057 = 8'hf0;
assign n0058 = ( RD_ROM_1 == n0057 );
assign n0059 = 8'h0;
assign n0060 = ( n0058 ) ? ( B ) : ( n0059 );
assign n0061 = ( n0056 ) ? ( ACC ) : ( n0060 );
assign n0062 = ( n0054 ) ? ( PSW ) : ( n0061 );
assign n0063 = ( n0052 ) ? ( IP ) : ( n0062 );
assign n0064 = ( n0050 ) ? ( P3 ) : ( n0063 );
assign n0065 = ( n0048 ) ? ( IE ) : ( n0064 );
assign n0066 = ( n0046 ) ? ( P2 ) : ( n0065 );
assign n0067 = ( n0044 ) ? ( SBUF ) : ( n0066 );
assign n0068 = ( n0042 ) ? ( SCON ) : ( n0067 );
assign n0069 = ( n0040 ) ? ( P1 ) : ( n0068 );
assign n0070 = ( n0038 ) ? ( TH1 ) : ( n0069 );
assign n0071 = ( n0036 ) ? ( TL1 ) : ( n0070 );
assign n0072 = ( n0034 ) ? ( TH0 ) : ( n0071 );
assign n0073 = ( n0032 ) ? ( TL0 ) : ( n0072 );
assign n0074 = ( n0030 ) ? ( TMOD ) : ( n0073 );
assign n0075 = ( n0028 ) ? ( TCON ) : ( n0074 );
assign n0076 = ( n0026 ) ? ( PCON ) : ( n0075 );
assign n0077 = ( n0024 ) ? ( DPH ) : ( n0076 );
assign n0078 = ( n0022 ) ? ( DPL ) : ( n0077 );
assign n0079 = ( n0020 ) ? ( SP ) : ( n0078 );
assign n0080 = ( n0018 ) ? ( P0 ) : ( n0079 );
assign n0081 = ( n0015 ) ? ( RD_IRAM_0 ) : ( n0080 );
assign n0082 = 8'h1;
assign n0083 = ( n0081 + n0082 );
// 
// SP_05
// 
// 
// PSW_05
// 
// 
// ACC_06
// 
// 
// B_06
// 
// 
// DPL_06
// 
// 
// DPH_06
// 
// 
// PC_06
// 
// 
// P2_06
// 
// 
// P3_06
// 
// 
// P0_06
// 
// 
// P1_06
// 
// 
// IRAM_06
// 
assign n0084 = RD_IRAM_0[3:0];
assign n0085 = ( RD_IRAM_1 + n0082 );
// 
// SP_06
// 
// 
// PSW_06
// 
// 
// ACC_07
// 
// 
// B_07
// 
// 
// DPL_07
// 
// 
// DPH_07
// 
// 
// PC_07
// 
// 
// P2_07
// 
// 
// P3_07
// 
// 
// P0_07
// 
// 
// P1_07
// 
// 
// IRAM_07
// 
// 
// SP_07
// 
// 
// PSW_07
// 
// 
// ACC_08
// 
// 
// B_08
// 
// 
// DPL_08
// 
// 
// DPH_08
// 
// 
// PC_08
// 
// 
// P2_08
// 
// 
// P3_08
// 
// 
// P0_08
// 
// 
// P1_08
// 
// 
// IRAM_08
// 
assign n0086 = { ( n0003 ), ( n0004 ), ( n0003 ) };
assign n0087 = n0086[3:0];
assign n0088 = ( RD_IRAM_0 + n0082 );
// 
// SP_08
// 
// 
// PSW_08
// 
// 
// ACC_09
// 
// 
// B_09
// 
// 
// DPL_09
// 
// 
// DPH_09
// 
// 
// PC_09
// 
// 
// P2_09
// 
// 
// P3_09
// 
// 
// P0_09
// 
// 
// P1_09
// 
// 
// IRAM_09
// 
assign n0089 = 3'h1;
assign n0090 = { ( n0003 ), ( n0004 ), ( n0089 ) };
assign n0091 = n0090[3:0];
// 
// SP_09
// 
// 
// PSW_09
// 
// 
// ACC_0a
// 
// 
// B_0a
// 
// 
// DPL_0a
// 
// 
// DPH_0a
// 
// 
// PC_0a
// 
// 
// P2_0a
// 
// 
// P3_0a
// 
// 
// P0_0a
// 
// 
// P1_0a
// 
// 
// IRAM_0a
// 
assign n0092 = 3'h2;
assign n0093 = { ( n0003 ), ( n0004 ), ( n0092 ) };
assign n0094 = n0093[3:0];
// 
// SP_0a
// 
// 
// PSW_0a
// 
// 
// ACC_0b
// 
// 
// P1_0b
// 
// 
// DPL_0b
// 
// 
// DPH_0b
// 
// 
// PC_0b
// 
// 
// P2_0b
// 
// 
// P3_0b
// 
// 
// P0_0b
// 
// 
// B_0b
// 
// 
// IRAM_0b
// 
assign n0095 = n0006[3:0];
// 
// SP_0b
// 
// 
// PSW_0b
// 
// 
// ACC_0c
// 
// 
// P1_0c
// 
// 
// DPL_0c
// 
// 
// DPH_0c
// 
// 
// PC_0c
// 
// 
// P2_0c
// 
// 
// P3_0c
// 
// 
// P0_0c
// 
// 
// B_0c
// 
// 
// IRAM_0c
// 
assign n0096 = 3'h4;
assign n0097 = { ( n0003 ), ( n0004 ), ( n0096 ) };
assign n0098 = n0097[3:0];
// 
// SP_0c
// 
// 
// PSW_0c
// 
// 
// ACC_0d
// 
// 
// B_0d
// 
// 
// DPL_0d
// 
// 
// DPH_0d
// 
// 
// PC_0d
// 
// 
// P2_0d
// 
// 
// P3_0d
// 
// 
// P0_0d
// 
// 
// P1_0d
// 
// 
// IRAM_0d
// 
assign n0099 = 3'h5;
assign n0100 = { ( n0003 ), ( n0004 ), ( n0099 ) };
assign n0101 = n0100[3:0];
// 
// SP_0d
// 
// 
// PSW_0d
// 
// 
// ACC_0e
// 
// 
// B_0e
// 
// 
// DPL_0e
// 
// 
// DPH_0e
// 
// 
// PC_0e
// 
// 
// P2_0e
// 
// 
// P3_0e
// 
// 
// P0_0e
// 
// 
// P1_0e
// 
// 
// IRAM_0e
// 
assign n0102 = 3'h6;
assign n0103 = { ( n0003 ), ( n0004 ), ( n0102 ) };
assign n0104 = n0103[3:0];
// 
// SP_0e
// 
// 
// PSW_0e
// 
// 
// ACC_0f
// 
// 
// P1_0f
// 
// 
// DPL_0f
// 
// 
// DPH_0f
// 
// 
// PC_0f
// 
// 
// P2_0f
// 
// 
// P3_0f
// 
// 
// P0_0f
// 
// 
// B_0f
// 
// 
// IRAM_0f
// 
assign n0105 = 3'h7;
assign n0106 = { ( n0003 ), ( n0004 ), ( n0105 ) };
assign n0107 = n0106[3:0];
// 
// SP_0f
// 
// 
// PSW_0f
// 
// 
// ACC_10
// 
// 
// P1_10
// 
// 
// DPL_10
// 
// 
// DPH_10
// 
// 
// PC_10
// 
// 
// P2_10
// 
// 
// P3_10
// 
// 
// P0_10
// 
// 
// B_10
// 
// 
// IRAM_10
// 
assign n0108 = 1'h1;
assign n0109 = ( n0013 == n0108 );
assign n0110 = RD_ROM_1[7:3];
assign n0111 = { ( n0110 ), ( n0003 ) };
assign n0112 = { 3'b0, n0110 };
assign n0113 = 8'h20;
assign n0114 = ( n0112 + n0113 );
assign n0115 = ( n0109 ) ? ( n0111 ) : ( n0114 );
assign n0116 = n0115[7:7];
assign n0117 = ( n0116 == n0014 );
assign n0118 = n0115[3:0];
assign n0119 = RD_ROM_1[2:0];
assign n0120 = { 5'b0, n0119 };
assign n0121 = ( n0082 << n0120 );
assign n0122 = ~( n0121 );
assign n0123 = ( n0115 == n0017 );
assign n0124 = ( n0115 == n0027 );
assign n0125 = ( n0115 == n0039 );
assign n0126 = ( n0115 == n0041 );
assign n0127 = ( n0115 == n0045 );
assign n0128 = ( n0115 == n0047 );
assign n0129 = ( n0115 == n0049 );
assign n0130 = ( n0115 == n0051 );
assign n0131 = ( n0115 == n0053 );
assign n0132 = ( n0115 == n0055 );
assign n0133 = ( n0115 == n0057 );
assign n0134 = ( n0133 ) ? ( B ) : ( n0059 );
assign n0135 = ( n0132 ) ? ( ACC ) : ( n0134 );
assign n0136 = ( n0131 ) ? ( PSW ) : ( n0135 );
assign n0137 = ( n0130 ) ? ( IP ) : ( n0136 );
assign n0138 = ( n0129 ) ? ( P3INREG ) : ( n0137 );
assign n0139 = ( n0128 ) ? ( IE ) : ( n0138 );
assign n0140 = ( n0127 ) ? ( P2INREG ) : ( n0139 );
assign n0141 = ( n0126 ) ? ( SCON ) : ( n0140 );
assign n0142 = ( n0125 ) ? ( P1INREG ) : ( n0141 );
assign n0143 = ( n0124 ) ? ( TCON ) : ( n0142 );
assign n0144 = ( n0123 ) ? ( P0INREG ) : ( n0143 );
assign n0145 = ( n0117 ) ? ( RD_IRAM_0 ) : ( n0144 );
assign n0146 = ( n0122 & n0145 );
assign n0147 = { 7'b0, n0014 };
assign n0148 = ( n0147 << n0120 );
assign n0149 = ( n0146 | n0148 );
// 
// SP_10
// 
// 
// PSW_10
// 
// 
// ACC_11
// 
// 
// B_11
// 
// 
// DPL_11
// 
// 
// DPH_11
// 
// 
// PC_11
// 
// 
// P2_11
// 
// 
// P3_11
// 
// 
// P0_11
// 
// 
// P1_11
// 
// 
// IRAM_11
// 
assign n0150 = ( SP + n0082 );
assign n0151 = n0150[3:0];
assign n0152 = 16'h2;
assign n0153 = ( PC + n0152 );
assign n0154 = n0153[7:0];
assign n0155 = ( n0150 + n0082 );
assign n0156 = n0155[3:0];
assign n0157 = n0153[15:8];
// 
// SP_11
// 
// 
// PSW_11
// 
// 
// ACC_12
// 
// 
// B_12
// 
// 
// DPL_12
// 
// 
// DPH_12
// 
// 
// PC_12
// 
// 
// P2_12
// 
// 
// P3_12
// 
// 
// P0_12
// 
// 
// P1_12
// 
// 
// IRAM_12
// 
assign n0158 = 16'h3;
assign n0159 = ( PC + n0158 );
assign n0160 = n0159[7:0];
assign n0161 = n0159[15:8];
// 
// SP_12
// 
// 
// PSW_12
// 
// 
// ACC_13
// 
// 
// B_13
// 
// 
// DPL_13
// 
// 
// DPH_13
// 
// 
// PC_13
// 
// 
// P2_13
// 
// 
// P3_13
// 
// 
// P0_13
// 
// 
// P1_13
// 
// 
// SP_13
// 
// 
// PSW_13
// 
// 
// ACC_14
// 
// 
// P1_14
// 
// 
// DPL_14
// 
// 
// DPH_14
// 
// 
// PC_14
// 
// 
// P2_14
// 
// 
// P3_14
// 
// 
// P0_14
// 
// 
// B_14
// 
// 
// SP_14
// 
// 
// PSW_14
// 
// 
// ACC_15
// 
// 
// P1_15
// 
// 
// DPL_15
// 
// 
// DPH_15
// 
// 
// PC_15
// 
// 
// P2_15
// 
// 
// P3_15
// 
// 
// P0_15
// 
// 
// B_15
// 
// 
// IRAM_15
// 
assign n0162 = ( n0081 - n0082 );
// 
// SP_15
// 
// 
// PSW_15
// 
// 
// ACC_16
// 
// 
// B_16
// 
// 
// DPL_16
// 
// 
// DPH_16
// 
// 
// PC_16
// 
// 
// P2_16
// 
// 
// P3_16
// 
// 
// P0_16
// 
// 
// P1_16
// 
// 
// IRAM_16
// 
assign n0163 = ( RD_IRAM_1 - n0082 );
// 
// SP_16
// 
// 
// PSW_16
// 
// 
// ACC_17
// 
// 
// B_17
// 
// 
// DPL_17
// 
// 
// DPH_17
// 
// 
// PC_17
// 
// 
// P2_17
// 
// 
// P3_17
// 
// 
// P0_17
// 
// 
// P1_17
// 
// 
// IRAM_17
// 
// 
// SP_17
// 
// 
// PSW_17
// 
// 
// ACC_18
// 
// 
// P1_18
// 
// 
// DPL_18
// 
// 
// DPH_18
// 
// 
// PC_18
// 
// 
// P2_18
// 
// 
// P3_18
// 
// 
// P0_18
// 
// 
// B_18
// 
// 
// IRAM_18
// 
assign n0164 = ( RD_IRAM_0 - n0082 );
// 
// SP_18
// 
// 
// PSW_18
// 
// 
// ACC_19
// 
// 
// P1_19
// 
// 
// DPL_19
// 
// 
// DPH_19
// 
// 
// PC_19
// 
// 
// P2_19
// 
// 
// P3_19
// 
// 
// P0_19
// 
// 
// B_19
// 
// 
// IRAM_19
// 
// 
// SP_19
// 
// 
// PSW_19
// 
// 
// ACC_1a
// 
// 
// P1_1a
// 
// 
// DPL_1a
// 
// 
// DPH_1a
// 
// 
// PC_1a
// 
// 
// P2_1a
// 
// 
// P3_1a
// 
// 
// P0_1a
// 
// 
// B_1a
// 
// 
// IRAM_1a
// 
// 
// SP_1a
// 
// 
// PSW_1a
// 
// 
// ACC_1b
// 
// 
// B_1b
// 
// 
// DPL_1b
// 
// 
// DPH_1b
// 
// 
// PC_1b
// 
// 
// P2_1b
// 
// 
// P3_1b
// 
// 
// P0_1b
// 
// 
// P1_1b
// 
// 
// IRAM_1b
// 
// 
// SP_1b
// 
// 
// PSW_1b
// 
// 
// ACC_1c
// 
// 
// B_1c
// 
// 
// DPL_1c
// 
// 
// DPH_1c
// 
// 
// PC_1c
// 
// 
// P2_1c
// 
// 
// P3_1c
// 
// 
// P0_1c
// 
// 
// P1_1c
// 
// 
// IRAM_1c
// 
// 
// SP_1c
// 
// 
// PSW_1c
// 
// 
// ACC_1d
// 
// 
// B_1d
// 
// 
// DPL_1d
// 
// 
// DPH_1d
// 
// 
// PC_1d
// 
// 
// P2_1d
// 
// 
// P3_1d
// 
// 
// P0_1d
// 
// 
// P1_1d
// 
// 
// IRAM_1d
// 
// 
// SP_1d
// 
// 
// PSW_1d
// 
// 
// ACC_1e
// 
// 
// P1_1e
// 
// 
// DPL_1e
// 
// 
// DPH_1e
// 
// 
// PC_1e
// 
// 
// P2_1e
// 
// 
// P3_1e
// 
// 
// P0_1e
// 
// 
// B_1e
// 
// 
// IRAM_1e
// 
// 
// SP_1e
// 
// 
// PSW_1e
// 
// 
// ACC_1f
// 
// 
// B_1f
// 
// 
// DPL_1f
// 
// 
// DPH_1f
// 
// 
// PC_1f
// 
// 
// P2_1f
// 
// 
// P3_1f
// 
// 
// P0_1f
// 
// 
// P1_1f
// 
// 
// IRAM_1f
// 
// 
// SP_1f
// 
// 
// PSW_1f
// 
// 
// ACC_20
// 
// 
// B_20
// 
// 
// DPL_20
// 
// 
// DPH_20
// 
// 
// PC_20
// 
// 
// P2_20
// 
// 
// P3_20
// 
// 
// P0_20
// 
// 
// P1_20
// 
// 
// SP_20
// 
// 
// PSW_20
// 
// 
// ACC_21
// 
// 
// B_21
// 
// 
// DPL_21
// 
// 
// DPH_21
// 
// 
// PC_21
// 
// 
// P2_21
// 
// 
// P3_21
// 
// 
// P0_21
// 
// 
// P1_21
// 
// 
// SP_21
// 
// 
// PSW_21
// 
// 
// ACC_22
// 
// 
// P1_22
// 
// 
// DPL_22
// 
// 
// DPH_22
// 
// 
// PC_22
// 
// 
// P2_22
// 
// 
// P3_22
// 
// 
// P0_22
// 
// 
// B_22
// 
// 
// SP_22
// 
// 
// PSW_22
// 
// 
// ACC_23
// 
// 
// B_23
// 
// 
// DPL_23
// 
// 
// DPH_23
// 
// 
// PC_23
// 
// 
// P2_23
// 
// 
// P3_23
// 
// 
// P0_23
// 
// 
// P1_23
// 
// 
// SP_23
// 
// 
// PSW_23
// 
// 
// ACC_24
// 
// 
// B_24
// 
// 
// DPL_24
// 
// 
// DPH_24
// 
// 
// PC_24
// 
// 
// P2_24
// 
// 
// P3_24
// 
// 
// P0_24
// 
// 
// P1_24
// 
// 
// SP_24
// 
// 
// PSW_24
// 
// 
// ACC_25
// 
// 
// P1_25
// 
// 
// DPL_25
// 
// 
// DPH_25
// 
// 
// PC_25
// 
// 
// P2_25
// 
// 
// P3_25
// 
// 
// P0_25
// 
// 
// B_25
// 
// 
// SP_25
// 
// 
// PSW_25
// 
// 
// ACC_26
// 
// 
// P1_26
// 
// 
// DPL_26
// 
// 
// DPH_26
// 
// 
// PC_26
// 
// 
// P2_26
// 
// 
// P3_26
// 
// 
// P0_26
// 
// 
// B_26
// 
// 
// SP_26
// 
// 
// PSW_26
// 
// 
// ACC_27
// 
// 
// B_27
// 
// 
// DPL_27
// 
// 
// DPH_27
// 
// 
// PC_27
// 
// 
// P2_27
// 
// 
// P3_27
// 
// 
// P0_27
// 
// 
// P1_27
// 
// 
// SP_27
// 
// 
// PSW_27
// 
// 
// ACC_28
// 
// 
// P1_28
// 
// 
// DPL_28
// 
// 
// DPH_28
// 
// 
// PC_28
// 
// 
// P2_28
// 
// 
// P3_28
// 
// 
// P0_28
// 
// 
// B_28
// 
// 
// SP_28
// 
// 
// PSW_28
// 
// 
// ACC_29
// 
// 
// P1_29
// 
// 
// DPL_29
// 
// 
// DPH_29
// 
// 
// PC_29
// 
// 
// P2_29
// 
// 
// P3_29
// 
// 
// P0_29
// 
// 
// B_29
// 
// 
// SP_29
// 
// 
// PSW_29
// 
// 
// ACC_2a
// 
// 
// B_2a
// 
// 
// DPL_2a
// 
// 
// DPH_2a
// 
// 
// PC_2a
// 
// 
// P2_2a
// 
// 
// P3_2a
// 
// 
// P0_2a
// 
// 
// P1_2a
// 
// 
// SP_2a
// 
// 
// PSW_2a
// 
// 
// ACC_2b
// 
// 
// B_2b
// 
// 
// DPL_2b
// 
// 
// DPH_2b
// 
// 
// PC_2b
// 
// 
// P2_2b
// 
// 
// P3_2b
// 
// 
// P0_2b
// 
// 
// P1_2b
// 
// 
// SP_2b
// 
// 
// PSW_2b
// 
// 
// ACC_2c
// 
// 
// B_2c
// 
// 
// DPL_2c
// 
// 
// DPH_2c
// 
// 
// PC_2c
// 
// 
// P2_2c
// 
// 
// P3_2c
// 
// 
// P0_2c
// 
// 
// P1_2c
// 
// 
// SP_2c
// 
// 
// PSW_2c
// 
// 
// ACC_2d
// 
// 
// P1_2d
// 
// 
// DPL_2d
// 
// 
// DPH_2d
// 
// 
// PC_2d
// 
// 
// P2_2d
// 
// 
// P3_2d
// 
// 
// P0_2d
// 
// 
// B_2d
// 
// 
// SP_2d
// 
// 
// PSW_2d
// 
// 
// ACC_2e
// 
// 
// B_2e
// 
// 
// DPL_2e
// 
// 
// DPH_2e
// 
// 
// PC_2e
// 
// 
// P2_2e
// 
// 
// P3_2e
// 
// 
// P0_2e
// 
// 
// P1_2e
// 
// 
// SP_2e
// 
// 
// PSW_2e
// 
// 
// ACC_2f
// 
// 
// P1_2f
// 
// 
// DPL_2f
// 
// 
// DPH_2f
// 
// 
// PC_2f
// 
// 
// P2_2f
// 
// 
// P3_2f
// 
// 
// P0_2f
// 
// 
// B_2f
// 
// 
// SP_2f
// 
// 
// PSW_2f
// 
// 
// ACC_30
// 
// 
// P1_30
// 
// 
// DPL_30
// 
// 
// DPH_30
// 
// 
// PC_30
// 
// 
// P2_30
// 
// 
// P3_30
// 
// 
// P0_30
// 
// 
// B_30
// 
// 
// SP_30
// 
// 
// PSW_30
// 
// 
// ACC_31
// 
// 
// B_31
// 
// 
// DPL_31
// 
// 
// DPH_31
// 
// 
// PC_31
// 
// 
// P2_31
// 
// 
// P3_31
// 
// 
// P0_31
// 
// 
// P1_31
// 
// 
// IRAM_31
// 
// 
// SP_31
// 
// 
// PSW_31
// 
// 
// ACC_32
// 
// 
// B_32
// 
// 
// DPL_32
// 
// 
// DPH_32
// 
// 
// PC_32
// 
// 
// P2_32
// 
// 
// P3_32
// 
// 
// P0_32
// 
// 
// P1_32
// 
// 
// SP_32
// 
// 
// PSW_32
// 
// 
// ACC_33
// 
// 
// B_33
// 
// 
// DPL_33
// 
// 
// DPH_33
// 
// 
// PC_33
// 
// 
// P2_33
// 
// 
// P3_33
// 
// 
// P0_33
// 
// 
// P1_33
// 
// 
// SP_33
// 
// 
// PSW_33
// 
// 
// ACC_34
// 
// 
// B_34
// 
// 
// DPL_34
// 
// 
// DPH_34
// 
// 
// PC_34
// 
// 
// P2_34
// 
// 
// P3_34
// 
// 
// P0_34
// 
// 
// P1_34
// 
// 
// SP_34
// 
// 
// PSW_34
// 
// 
// ACC_35
// 
// 
// B_35
// 
// 
// DPL_35
// 
// 
// DPH_35
// 
// 
// PC_35
// 
// 
// P2_35
// 
// 
// P3_35
// 
// 
// P0_35
// 
// 
// P1_35
// 
// 
// SP_35
// 
// 
// PSW_35
// 
// 
// ACC_36
// 
// 
// B_36
// 
// 
// DPL_36
// 
// 
// DPH_36
// 
// 
// PC_36
// 
// 
// P2_36
// 
// 
// P3_36
// 
// 
// P0_36
// 
// 
// P1_36
// 
// 
// SP_36
// 
// 
// PSW_36
// 
// 
// ACC_37
// 
// 
// B_37
// 
// 
// DPL_37
// 
// 
// DPH_37
// 
// 
// PC_37
// 
// 
// P2_37
// 
// 
// P3_37
// 
// 
// P0_37
// 
// 
// P1_37
// 
// 
// SP_37
// 
// 
// PSW_37
// 
// 
// ACC_38
// 
// 
// B_38
// 
// 
// DPL_38
// 
// 
// DPH_38
// 
// 
// PC_38
// 
// 
// P2_38
// 
// 
// P3_38
// 
// 
// P0_38
// 
// 
// P1_38
// 
// 
// SP_38
// 
// 
// PSW_38
// 
// 
// ACC_39
// 
// 
// P1_39
// 
// 
// DPL_39
// 
// 
// DPH_39
// 
// 
// PC_39
// 
// 
// P2_39
// 
// 
// P3_39
// 
// 
// P0_39
// 
// 
// B_39
// 
// 
// SP_39
// 
// 
// PSW_39
// 
// 
// ACC_3a
// 
// 
// P1_3a
// 
// 
// DPL_3a
// 
// 
// DPH_3a
// 
// 
// PC_3a
// 
// 
// P2_3a
// 
// 
// P3_3a
// 
// 
// P0_3a
// 
// 
// B_3a
// 
// 
// SP_3a
// 
// 
// PSW_3a
// 
// 
// ACC_3b
// 
// 
// B_3b
// 
// 
// DPL_3b
// 
// 
// DPH_3b
// 
// 
// PC_3b
// 
// 
// P2_3b
// 
// 
// P3_3b
// 
// 
// P0_3b
// 
// 
// P1_3b
// 
// 
// SP_3b
// 
// 
// PSW_3b
// 
// 
// ACC_3c
// 
// 
// P1_3c
// 
// 
// DPL_3c
// 
// 
// DPH_3c
// 
// 
// PC_3c
// 
// 
// P2_3c
// 
// 
// P3_3c
// 
// 
// P0_3c
// 
// 
// B_3c
// 
// 
// SP_3c
// 
// 
// PSW_3c
// 
// 
// ACC_3d
// 
// 
// B_3d
// 
// 
// DPL_3d
// 
// 
// DPH_3d
// 
// 
// PC_3d
// 
// 
// P2_3d
// 
// 
// P3_3d
// 
// 
// P0_3d
// 
// 
// P1_3d
// 
// 
// SP_3d
// 
// 
// PSW_3d
// 
// 
// ACC_3e
// 
// 
// B_3e
// 
// 
// DPL_3e
// 
// 
// DPH_3e
// 
// 
// PC_3e
// 
// 
// P2_3e
// 
// 
// P3_3e
// 
// 
// P0_3e
// 
// 
// P1_3e
// 
// 
// SP_3e
// 
// 
// PSW_3e
// 
// 
// ACC_3f
// 
// 
// P1_3f
// 
// 
// DPL_3f
// 
// 
// DPH_3f
// 
// 
// PC_3f
// 
// 
// P2_3f
// 
// 
// P3_3f
// 
// 
// P0_3f
// 
// 
// B_3f
// 
// 
// SP_3f
// 
// 
// PSW_3f
// 
// 
// ACC_40
// 
// 
// B_40
// 
// 
// DPL_40
// 
// 
// DPH_40
// 
// 
// PC_40
// 
// 
// P2_40
// 
// 
// P3_40
// 
// 
// P0_40
// 
// 
// P1_40
// 
// 
// SP_40
// 
// 
// PSW_40
// 
// 
// ACC_41
// 
// 
// B_41
// 
// 
// DPL_41
// 
// 
// DPH_41
// 
// 
// PC_41
// 
// 
// P2_41
// 
// 
// P3_41
// 
// 
// P0_41
// 
// 
// P1_41
// 
// 
// SP_41
// 
// 
// PSW_41
// 
// 
// ACC_42
// 
// 
// B_42
// 
// 
// DPL_42
// 
// 
// DPH_42
// 
// 
// PC_42
// 
// 
// P2_42
// 
// 
// P3_42
// 
// 
// P0_42
// 
// 
// P1_42
// 
// 
// IRAM_42
// 
assign n0165 = ( n0081 | ACC );
// 
// SP_42
// 
// 
// PSW_42
// 
// 
// ACC_43
// 
// 
// P1_43
// 
// 
// DPL_43
// 
// 
// DPH_43
// 
// 
// PC_43
// 
// 
// P2_43
// 
// 
// P3_43
// 
// 
// P0_43
// 
// 
// B_43
// 
// 
// IRAM_43
// 
assign n0166 = ( n0081 | RD_ROM_2 );
// 
// SP_43
// 
// 
// PSW_43
// 
// 
// ACC_44
// 
// 
// B_44
// 
// 
// DPL_44
// 
// 
// DPH_44
// 
// 
// PC_44
// 
// 
// P2_44
// 
// 
// P3_44
// 
// 
// P0_44
// 
// 
// P1_44
// 
// 
// SP_44
// 
// 
// PSW_44
// 
// 
// ACC_45
// 
// 
// P1_45
// 
// 
// DPL_45
// 
// 
// DPH_45
// 
// 
// PC_45
// 
// 
// P2_45
// 
// 
// P3_45
// 
// 
// P0_45
// 
// 
// B_45
// 
// 
// SP_45
// 
// 
// PSW_45
// 
// 
// ACC_46
// 
// 
// B_46
// 
// 
// DPL_46
// 
// 
// DPH_46
// 
// 
// PC_46
// 
// 
// P2_46
// 
// 
// P3_46
// 
// 
// P0_46
// 
// 
// P1_46
// 
// 
// SP_46
// 
// 
// PSW_46
// 
// 
// ACC_47
// 
// 
// P1_47
// 
// 
// DPL_47
// 
// 
// DPH_47
// 
// 
// PC_47
// 
// 
// P2_47
// 
// 
// P3_47
// 
// 
// P0_47
// 
// 
// B_47
// 
// 
// SP_47
// 
// 
// PSW_47
// 
// 
// ACC_48
// 
// 
// P1_48
// 
// 
// DPL_48
// 
// 
// DPH_48
// 
// 
// PC_48
// 
// 
// P2_48
// 
// 
// P3_48
// 
// 
// P0_48
// 
// 
// B_48
// 
// 
// SP_48
// 
// 
// PSW_48
// 
// 
// ACC_49
// 
// 
// B_49
// 
// 
// DPL_49
// 
// 
// DPH_49
// 
// 
// PC_49
// 
// 
// P2_49
// 
// 
// P3_49
// 
// 
// P0_49
// 
// 
// P1_49
// 
// 
// SP_49
// 
// 
// PSW_49
// 
// 
// ACC_4a
// 
// 
// P1_4a
// 
// 
// DPL_4a
// 
// 
// DPH_4a
// 
// 
// PC_4a
// 
// 
// P2_4a
// 
// 
// P3_4a
// 
// 
// P0_4a
// 
// 
// B_4a
// 
// 
// SP_4a
// 
// 
// PSW_4a
// 
// 
// ACC_4b
// 
assign n0167 = ( ACC | RD_IRAM_0 );
assign ACC_4b = n0167;
// 
// P1_4b
// 
assign P1_4b = P1;
// 
// DPL_4b
// 
assign DPL_4b = DPL;
// 
// DPH_4b
// 
assign DPH_4b = DPH;
// 
// PC_4b
// 
assign n0168 = 16'h1;
assign n0169 = ( PC + n0168 );
assign PC_4b = n0169;
// 
// P2_4b
// 
assign P2_4b = P2;
// 
// P3_4b
// 
assign P3_4b = P3;
// 
// P0_4b
// 
assign P0_4b = P0;
// 
// B_4b
// 
assign B_4b = B;
// 
// SP_4b
// 
assign SP_4b = SP;
// 
// PSW_4b
// 
assign n0170 = PSW[7:1];
assign n0171 = n0167[7:7];
assign n0172 = n0167[6:6];
assign n0173 = n0167[5:5];
assign n0174 = n0167[4:4];
assign n0175 = n0167[3:3];
assign n0176 = n0167[2:2];
assign n0177 = n0167[1:1];
assign n0178 = n0167[0:0];
assign n0179 = ( n0177 ^ n0178 );
assign n0180 = ( n0176 ^ n0179 );
assign n0181 = ( n0175 ^ n0180 );
assign n0182 = ( n0174 ^ n0181 );
assign n0183 = ( n0173 ^ n0182 );
assign n0184 = ( n0172 ^ n0183 );
assign n0185 = ( n0171 ^ n0184 );
assign n0186 = { ( n0170 ), ( n0185 ) };
assign PSW_4b = n0186;
// 
// ACC_4c
// 
// 
// P1_4c
// 
// 
// DPL_4c
// 
// 
// DPH_4c
// 
// 
// PC_4c
// 
// 
// P2_4c
// 
// 
// P3_4c
// 
// 
// P0_4c
// 
// 
// B_4c
// 
// 
// SP_4c
// 
// 
// PSW_4c
// 
// 
// ACC_4d
// 
// 
// B_4d
// 
// 
// DPL_4d
// 
// 
// DPH_4d
// 
// 
// PC_4d
// 
// 
// P2_4d
// 
// 
// P3_4d
// 
// 
// P0_4d
// 
// 
// P1_4d
// 
// 
// SP_4d
// 
// 
// PSW_4d
// 
// 
// ACC_4e
// 
// 
// P1_4e
// 
// 
// DPL_4e
// 
// 
// DPH_4e
// 
// 
// PC_4e
// 
// 
// P2_4e
// 
// 
// P3_4e
// 
// 
// P0_4e
// 
// 
// B_4e
// 
// 
// SP_4e
// 
// 
// PSW_4e
// 
// 
// ACC_4f
// 
// 
// P1_4f
// 
// 
// DPL_4f
// 
// 
// DPH_4f
// 
// 
// PC_4f
// 
// 
// P2_4f
// 
// 
// P3_4f
// 
// 
// P0_4f
// 
// 
// B_4f
// 
// 
// SP_4f
// 
// 
// PSW_4f
// 
// 
// ACC_50
// 
// 
// B_50
// 
// 
// DPL_50
// 
// 
// DPH_50
// 
// 
// PC_50
// 
// 
// P2_50
// 
// 
// P3_50
// 
// 
// P0_50
// 
// 
// P1_50
// 
// 
// SP_50
// 
// 
// PSW_50
// 
// 
// ACC_51
// 
// 
// B_51
// 
// 
// DPL_51
// 
// 
// DPH_51
// 
// 
// PC_51
// 
// 
// P2_51
// 
// 
// P3_51
// 
// 
// P0_51
// 
// 
// P1_51
// 
// 
// IRAM_51
// 
// 
// SP_51
// 
// 
// PSW_51
// 
// 
// ACC_52
// 
// 
// B_52
// 
// 
// DPL_52
// 
// 
// DPH_52
// 
// 
// PC_52
// 
// 
// P2_52
// 
// 
// P3_52
// 
// 
// P0_52
// 
// 
// P1_52
// 
// 
// IRAM_52
// 
assign n0187 = ( n0081 & ACC );
// 
// SP_52
// 
// 
// PSW_52
// 
// 
// ACC_53
// 
// 
// P1_53
// 
// 
// DPL_53
// 
// 
// DPH_53
// 
// 
// PC_53
// 
// 
// P2_53
// 
// 
// P3_53
// 
// 
// P0_53
// 
// 
// B_53
// 
// 
// IRAM_53
// 
assign n0188 = ( n0081 & RD_ROM_2 );
// 
// SP_53
// 
// 
// PSW_53
// 
// 
// ACC_54
// 
// 
// P1_54
// 
// 
// DPL_54
// 
// 
// DPH_54
// 
// 
// PC_54
// 
// 
// P2_54
// 
// 
// P3_54
// 
// 
// P0_54
// 
// 
// B_54
// 
// 
// SP_54
// 
// 
// PSW_54
// 
// 
// ACC_55
// 
// 
// B_55
// 
// 
// DPL_55
// 
// 
// DPH_55
// 
// 
// PC_55
// 
// 
// P2_55
// 
// 
// P3_55
// 
// 
// P0_55
// 
// 
// P1_55
// 
// 
// SP_55
// 
// 
// PSW_55
// 
// 
// ACC_56
// 
// 
// B_56
// 
// 
// DPL_56
// 
// 
// DPH_56
// 
// 
// PC_56
// 
// 
// P2_56
// 
// 
// P3_56
// 
// 
// P0_56
// 
// 
// P1_56
// 
// 
// SP_56
// 
// 
// PSW_56
// 
// 
// ACC_57
// 
// 
// B_57
// 
// 
// DPL_57
// 
// 
// DPH_57
// 
// 
// PC_57
// 
// 
// P2_57
// 
// 
// P3_57
// 
// 
// P0_57
// 
// 
// P1_57
// 
// 
// SP_57
// 
// 
// PSW_57
// 
// 
// ACC_58
// 
// 
// B_58
// 
// 
// DPL_58
// 
// 
// DPH_58
// 
// 
// PC_58
// 
// 
// P2_58
// 
// 
// P3_58
// 
// 
// P0_58
// 
// 
// P1_58
// 
// 
// SP_58
// 
// 
// PSW_58
// 
// 
// ACC_59
// 
// 
// P1_59
// 
// 
// DPL_59
// 
// 
// DPH_59
// 
// 
// PC_59
// 
// 
// P2_59
// 
// 
// P3_59
// 
// 
// P0_59
// 
// 
// B_59
// 
// 
// SP_59
// 
// 
// PSW_59
// 
// 
// ACC_5a
// 
// 
// B_5a
// 
// 
// DPL_5a
// 
// 
// DPH_5a
// 
// 
// PC_5a
// 
// 
// P2_5a
// 
// 
// P3_5a
// 
// 
// P0_5a
// 
// 
// P1_5a
// 
// 
// SP_5a
// 
// 
// PSW_5a
// 
// 
// ACC_5b
// 
// 
// B_5b
// 
// 
// DPL_5b
// 
// 
// DPH_5b
// 
// 
// PC_5b
// 
// 
// P2_5b
// 
// 
// P3_5b
// 
// 
// P0_5b
// 
// 
// P1_5b
// 
// 
// SP_5b
// 
// 
// PSW_5b
// 
// 
// ACC_5c
// 
// 
// B_5c
// 
// 
// DPL_5c
// 
// 
// DPH_5c
// 
// 
// PC_5c
// 
// 
// P2_5c
// 
// 
// P3_5c
// 
// 
// P0_5c
// 
// 
// P1_5c
// 
// 
// SP_5c
// 
// 
// PSW_5c
// 
// 
// ACC_5d
// 
// 
// P1_5d
// 
// 
// DPL_5d
// 
// 
// DPH_5d
// 
// 
// PC_5d
// 
// 
// P2_5d
// 
// 
// P3_5d
// 
// 
// P0_5d
// 
// 
// B_5d
// 
// 
// SP_5d
// 
// 
// PSW_5d
// 
// 
// ACC_5e
// 
// 
// B_5e
// 
// 
// DPL_5e
// 
// 
// DPH_5e
// 
// 
// PC_5e
// 
// 
// P2_5e
// 
// 
// P3_5e
// 
// 
// P0_5e
// 
// 
// P1_5e
// 
// 
// SP_5e
// 
// 
// PSW_5e
// 
// 
// ACC_5f
// 
// 
// B_5f
// 
// 
// DPL_5f
// 
// 
// DPH_5f
// 
// 
// PC_5f
// 
// 
// P2_5f
// 
// 
// P3_5f
// 
// 
// P0_5f
// 
// 
// P1_5f
// 
// 
// SP_5f
// 
// 
// PSW_5f
// 
// 
// ACC_60
// 
// 
// P1_60
// 
// 
// DPL_60
// 
// 
// DPH_60
// 
// 
// PC_60
// 
// 
// P2_60
// 
// 
// P3_60
// 
// 
// P0_60
// 
// 
// B_60
// 
// 
// SP_60
// 
// 
// PSW_60
// 
// 
// ACC_61
// 
// 
// P1_61
// 
// 
// DPL_61
// 
// 
// DPH_61
// 
// 
// PC_61
// 
// 
// P2_61
// 
// 
// P3_61
// 
// 
// P0_61
// 
// 
// B_61
// 
// 
// SP_61
// 
// 
// PSW_61
// 
// 
// ACC_62
// 
// 
// P1_62
// 
// 
// DPL_62
// 
// 
// DPH_62
// 
// 
// PC_62
// 
// 
// P2_62
// 
// 
// P3_62
// 
// 
// P0_62
// 
// 
// B_62
// 
// 
// IRAM_62
// 
assign n0189 = ( n0081 ^ ACC );
// 
// SP_62
// 
// 
// PSW_62
// 
// 
// ACC_63
// 
// 
// P1_63
// 
// 
// DPL_63
// 
// 
// DPH_63
// 
// 
// PC_63
// 
// 
// P2_63
// 
// 
// P3_63
// 
// 
// P0_63
// 
// 
// B_63
// 
// 
// IRAM_63
// 
assign n0190 = ( n0081 ^ RD_ROM_2 );
// 
// SP_63
// 
// 
// PSW_63
// 
// 
// ACC_64
// 
// 
// B_64
// 
// 
// DPL_64
// 
// 
// DPH_64
// 
// 
// PC_64
// 
// 
// P2_64
// 
// 
// P3_64
// 
// 
// P0_64
// 
// 
// P1_64
// 
// 
// SP_64
// 
// 
// PSW_64
// 
// 
// ACC_65
// 
// 
// B_65
// 
// 
// DPL_65
// 
// 
// DPH_65
// 
// 
// PC_65
// 
// 
// P2_65
// 
// 
// P3_65
// 
// 
// P0_65
// 
// 
// P1_65
// 
// 
// SP_65
// 
// 
// PSW_65
// 
// 
// ACC_66
// 
// 
// B_66
// 
// 
// DPL_66
// 
// 
// DPH_66
// 
// 
// PC_66
// 
// 
// P2_66
// 
// 
// P3_66
// 
// 
// P0_66
// 
// 
// P1_66
// 
// 
// SP_66
// 
// 
// PSW_66
// 
// 
// ACC_67
// 
// 
// P1_67
// 
// 
// DPL_67
// 
// 
// DPH_67
// 
// 
// PC_67
// 
// 
// P2_67
// 
// 
// P3_67
// 
// 
// P0_67
// 
// 
// B_67
// 
// 
// SP_67
// 
// 
// PSW_67
// 
// 
// ACC_68
// 
// 
// B_68
// 
// 
// DPL_68
// 
// 
// DPH_68
// 
// 
// PC_68
// 
// 
// P2_68
// 
// 
// P3_68
// 
// 
// P0_68
// 
// 
// P1_68
// 
// 
// SP_68
// 
// 
// PSW_68
// 
// 
// ACC_69
// 
// 
// B_69
// 
// 
// DPL_69
// 
// 
// DPH_69
// 
// 
// PC_69
// 
// 
// P2_69
// 
// 
// P3_69
// 
// 
// P0_69
// 
// 
// P1_69
// 
// 
// SP_69
// 
// 
// PSW_69
// 
// 
// ACC_6a
// 
// 
// B_6a
// 
// 
// DPL_6a
// 
// 
// DPH_6a
// 
// 
// PC_6a
// 
// 
// P2_6a
// 
// 
// P3_6a
// 
// 
// P0_6a
// 
// 
// P1_6a
// 
// 
// SP_6a
// 
// 
// PSW_6a
// 
// 
// ACC_6b
// 
// 
// P1_6b
// 
// 
// DPL_6b
// 
// 
// DPH_6b
// 
// 
// PC_6b
// 
// 
// P2_6b
// 
// 
// P3_6b
// 
// 
// P0_6b
// 
// 
// B_6b
// 
// 
// SP_6b
// 
// 
// PSW_6b
// 
// 
// ACC_6c
// 
// 
// B_6c
// 
// 
// DPL_6c
// 
// 
// DPH_6c
// 
// 
// PC_6c
// 
// 
// P2_6c
// 
// 
// P3_6c
// 
// 
// P0_6c
// 
// 
// P1_6c
// 
// 
// SP_6c
// 
// 
// PSW_6c
// 
// 
// ACC_6d
// 
// 
// B_6d
// 
// 
// DPL_6d
// 
// 
// DPH_6d
// 
// 
// PC_6d
// 
// 
// P2_6d
// 
// 
// P3_6d
// 
// 
// P0_6d
// 
// 
// P1_6d
// 
// 
// SP_6d
// 
// 
// PSW_6d
// 
// 
// ACC_6e
// 
// 
// P1_6e
// 
// 
// DPL_6e
// 
// 
// DPH_6e
// 
// 
// PC_6e
// 
// 
// P2_6e
// 
// 
// P3_6e
// 
// 
// P0_6e
// 
// 
// B_6e
// 
// 
// SP_6e
// 
// 
// PSW_6e
// 
// 
// ACC_6f
// 
// 
// B_6f
// 
// 
// DPL_6f
// 
// 
// DPH_6f
// 
// 
// PC_6f
// 
// 
// P2_6f
// 
// 
// P3_6f
// 
// 
// P0_6f
// 
// 
// P1_6f
// 
// 
// SP_6f
// 
// 
// PSW_6f
// 
// 
// ACC_70
// 
// 
// B_70
// 
// 
// DPL_70
// 
// 
// DPH_70
// 
// 
// PC_70
// 
// 
// P2_70
// 
// 
// P3_70
// 
// 
// P0_70
// 
// 
// P1_70
// 
// 
// SP_70
// 
// 
// PSW_70
// 
// 
// ACC_71
// 
// 
// P1_71
// 
// 
// DPL_71
// 
// 
// DPH_71
// 
// 
// PC_71
// 
// 
// P2_71
// 
// 
// P3_71
// 
// 
// P0_71
// 
// 
// B_71
// 
// 
// IRAM_71
// 
// 
// SP_71
// 
// 
// PSW_71
// 
// 
// ACC_72
// 
// 
// B_72
// 
// 
// DPL_72
// 
// 
// DPH_72
// 
// 
// PC_72
// 
// 
// P2_72
// 
// 
// P3_72
// 
// 
// P0_72
// 
// 
// P1_72
// 
// 
// SP_72
// 
// 
// PSW_72
// 
// 
// ACC_73
// 
// 
// B_73
// 
// 
// DPL_73
// 
// 
// DPH_73
// 
// 
// PC_73
// 
// 
// P2_73
// 
// 
// P3_73
// 
// 
// P0_73
// 
// 
// P1_73
// 
// 
// SP_73
// 
// 
// PSW_73
// 
// 
// ACC_74
// 
// 
// B_74
// 
// 
// DPL_74
// 
// 
// DPH_74
// 
// 
// PC_74
// 
// 
// P2_74
// 
// 
// P3_74
// 
// 
// P0_74
// 
// 
// P1_74
// 
// 
// SP_74
// 
// 
// PSW_74
// 
// 
// ACC_75
// 
// 
// P1_75
// 
// 
// DPL_75
// 
// 
// DPH_75
// 
// 
// PC_75
// 
// 
// P2_75
// 
// 
// P3_75
// 
// 
// P0_75
// 
// 
// B_75
// 
// 
// IRAM_75
// 
// 
// SP_75
// 
// 
// PSW_75
// 
// 
// ACC_76
// 
// 
// P1_76
// 
// 
// DPL_76
// 
// 
// DPH_76
// 
// 
// PC_76
// 
// 
// P2_76
// 
// 
// P3_76
// 
// 
// P0_76
// 
// 
// B_76
// 
// 
// IRAM_76
// 
// 
// SP_76
// 
// 
// PSW_76
// 
// 
// ACC_77
// 
// 
// P1_77
// 
// 
// DPL_77
// 
// 
// DPH_77
// 
// 
// PC_77
// 
// 
// P2_77
// 
// 
// P3_77
// 
// 
// P0_77
// 
// 
// B_77
// 
// 
// IRAM_77
// 
// 
// SP_77
// 
// 
// PSW_77
// 
// 
// ACC_78
// 
// 
// P1_78
// 
// 
// DPL_78
// 
// 
// DPH_78
// 
// 
// PC_78
// 
// 
// P2_78
// 
// 
// P3_78
// 
// 
// P0_78
// 
// 
// B_78
// 
// 
// IRAM_78
// 
// 
// SP_78
// 
// 
// PSW_78
// 
// 
// ACC_79
// 
// 
// B_79
// 
// 
// DPL_79
// 
// 
// DPH_79
// 
// 
// PC_79
// 
// 
// P2_79
// 
// 
// P3_79
// 
// 
// P0_79
// 
// 
// P1_79
// 
// 
// IRAM_79
// 
// 
// SP_79
// 
// 
// PSW_79
// 
// 
// ACC_7a
// 
// 
// P1_7a
// 
// 
// DPL_7a
// 
// 
// DPH_7a
// 
// 
// PC_7a
// 
// 
// P2_7a
// 
// 
// P3_7a
// 
// 
// P0_7a
// 
// 
// B_7a
// 
// 
// IRAM_7a
// 
// 
// SP_7a
// 
// 
// PSW_7a
// 
// 
// ACC_7b
// 
// 
// P1_7b
// 
// 
// DPL_7b
// 
// 
// DPH_7b
// 
// 
// PC_7b
// 
// 
// P2_7b
// 
// 
// P3_7b
// 
// 
// P0_7b
// 
// 
// B_7b
// 
// 
// IRAM_7b
// 
// 
// SP_7b
// 
// 
// PSW_7b
// 
// 
// ACC_7c
// 
// 
// P1_7c
// 
// 
// DPL_7c
// 
// 
// DPH_7c
// 
// 
// PC_7c
// 
// 
// P2_7c
// 
// 
// P3_7c
// 
// 
// P0_7c
// 
// 
// B_7c
// 
// 
// IRAM_7c
// 
// 
// SP_7c
// 
// 
// PSW_7c
// 
// 
// ACC_7d
// 
// 
// B_7d
// 
// 
// DPL_7d
// 
// 
// DPH_7d
// 
// 
// PC_7d
// 
// 
// P2_7d
// 
// 
// P3_7d
// 
// 
// P0_7d
// 
// 
// P1_7d
// 
// 
// IRAM_7d
// 
// 
// SP_7d
// 
// 
// PSW_7d
// 
// 
// ACC_7e
// 
// 
// B_7e
// 
// 
// DPL_7e
// 
// 
// DPH_7e
// 
// 
// PC_7e
// 
// 
// P2_7e
// 
// 
// P3_7e
// 
// 
// P0_7e
// 
// 
// P1_7e
// 
// 
// IRAM_7e
// 
// 
// SP_7e
// 
// 
// PSW_7e
// 
// 
// ACC_7f
// 
// 
// B_7f
// 
// 
// DPL_7f
// 
// 
// DPH_7f
// 
// 
// PC_7f
// 
// 
// P2_7f
// 
// 
// P3_7f
// 
// 
// P0_7f
// 
// 
// P1_7f
// 
// 
// IRAM_7f
// 
// 
// SP_7f
// 
// 
// PSW_7f
// 
// 
// ACC_80
// 
// 
// B_80
// 
// 
// DPL_80
// 
// 
// DPH_80
// 
// 
// PC_80
// 
// 
// P2_80
// 
// 
// P3_80
// 
// 
// P0_80
// 
// 
// P1_80
// 
// 
// SP_80
// 
// 
// PSW_80
// 
// 
// ACC_81
// 
// 
// B_81
// 
// 
// DPL_81
// 
// 
// DPH_81
// 
// 
// PC_81
// 
// 
// P2_81
// 
// 
// P3_81
// 
// 
// P0_81
// 
// 
// P1_81
// 
// 
// SP_81
// 
// 
// PSW_81
// 
// 
// ACC_82
// 
// 
// B_82
// 
// 
// DPL_82
// 
// 
// DPH_82
// 
// 
// PC_82
// 
// 
// P2_82
// 
// 
// P3_82
// 
// 
// P0_82
// 
// 
// P1_82
// 
// 
// SP_82
// 
// 
// PSW_82
// 
// 
// ACC_83
// 
// 
// P1_83
// 
// 
// DPL_83
// 
// 
// DPH_83
// 
// 
// PC_83
// 
// 
// P2_83
// 
// 
// P3_83
// 
// 
// P0_83
// 
// 
// B_83
// 
// 
// SP_83
// 
// 
// PSW_83
// 
// 
// ACC_84
// 
// 
// B_84
// 
// 
// DPL_84
// 
// 
// DPH_84
// 
// 
// PC_84
// 
// 
// P2_84
// 
// 
// P3_84
// 
// 
// P0_84
// 
// 
// P1_84
// 
// 
// SP_84
// 
// 
// PSW_84
// 
// 
// ACC_85
// 
// 
// B_85
// 
// 
// DPL_85
// 
// 
// DPH_85
// 
// 
// PC_85
// 
// 
// P2_85
// 
// 
// P3_85
// 
// 
// P0_85
// 
// 
// P1_85
// 
// 
// IRAM_85
// 
assign n0191 = RD_ROM_2[7:7];
assign n0192 = ( n0191 == n0014 );
assign n0193 = ( RD_ROM_2 == n0017 );
assign n0194 = ( RD_ROM_2 == n0019 );
assign n0195 = ( RD_ROM_2 == n0021 );
assign n0196 = ( RD_ROM_2 == n0023 );
assign n0197 = ( RD_ROM_2 == n0025 );
assign n0198 = ( RD_ROM_2 == n0027 );
assign n0199 = ( RD_ROM_2 == n0029 );
assign n0200 = ( RD_ROM_2 == n0031 );
assign n0201 = ( RD_ROM_2 == n0033 );
assign n0202 = ( RD_ROM_2 == n0035 );
assign n0203 = ( RD_ROM_2 == n0037 );
assign n0204 = ( RD_ROM_2 == n0039 );
assign n0205 = ( RD_ROM_2 == n0041 );
assign n0206 = ( RD_ROM_2 == n0043 );
assign n0207 = ( RD_ROM_2 == n0045 );
assign n0208 = ( RD_ROM_2 == n0047 );
assign n0209 = ( RD_ROM_2 == n0049 );
assign n0210 = ( RD_ROM_2 == n0051 );
assign n0211 = ( RD_ROM_2 == n0053 );
assign n0212 = ( RD_ROM_2 == n0055 );
assign n0213 = ( RD_ROM_2 == n0057 );
assign n0214 = ( n0213 ) ? ( B ) : ( n0059 );
assign n0215 = ( n0212 ) ? ( ACC ) : ( n0214 );
assign n0216 = ( n0211 ) ? ( PSW ) : ( n0215 );
assign n0217 = ( n0210 ) ? ( IP ) : ( n0216 );
assign n0218 = ( n0209 ) ? ( P3INREG ) : ( n0217 );
assign n0219 = ( n0208 ) ? ( IE ) : ( n0218 );
assign n0220 = ( n0207 ) ? ( P2INREG ) : ( n0219 );
assign n0221 = ( n0206 ) ? ( SBUF ) : ( n0220 );
assign n0222 = ( n0205 ) ? ( SCON ) : ( n0221 );
assign n0223 = ( n0204 ) ? ( P1INREG ) : ( n0222 );
assign n0224 = ( n0203 ) ? ( TH1 ) : ( n0223 );
assign n0225 = ( n0202 ) ? ( TL1 ) : ( n0224 );
assign n0226 = ( n0201 ) ? ( TH0 ) : ( n0225 );
assign n0227 = ( n0200 ) ? ( TL0 ) : ( n0226 );
assign n0228 = ( n0199 ) ? ( TMOD ) : ( n0227 );
assign n0229 = ( n0198 ) ? ( TCON ) : ( n0228 );
assign n0230 = ( n0197 ) ? ( PCON ) : ( n0229 );
assign n0231 = ( n0196 ) ? ( DPH ) : ( n0230 );
assign n0232 = ( n0195 ) ? ( DPL ) : ( n0231 );
assign n0233 = ( n0194 ) ? ( SP ) : ( n0232 );
assign n0234 = ( n0193 ) ? ( P0INREG ) : ( n0233 );
assign n0235 = ( n0192 ) ? ( RD_IRAM_0 ) : ( n0234 );
// 
// SP_85
// 
// 
// PSW_85
// 
// 
// ACC_86
// 
// 
// P1_86
// 
// 
// DPL_86
// 
// 
// DPH_86
// 
// 
// PC_86
// 
// 
// P2_86
// 
// 
// P3_86
// 
// 
// P0_86
// 
// 
// B_86
// 
// 
// IRAM_86
// 
// 
// SP_86
// 
// 
// PSW_86
// 
// 
// ACC_87
// 
// 
// B_87
// 
// 
// DPL_87
// 
// 
// DPH_87
// 
// 
// PC_87
// 
// 
// P2_87
// 
// 
// P3_87
// 
// 
// P0_87
// 
// 
// P1_87
// 
// 
// IRAM_87
// 
// 
// SP_87
// 
// 
// PSW_87
// 
// 
// ACC_88
// 
// 
// B_88
// 
// 
// DPL_88
// 
// 
// DPH_88
// 
// 
// PC_88
// 
// 
// P2_88
// 
// 
// P3_88
// 
// 
// P0_88
// 
// 
// P1_88
// 
// 
// IRAM_88
// 
// 
// SP_88
// 
// 
// PSW_88
// 
// 
// ACC_89
// 
// 
// B_89
// 
// 
// DPL_89
// 
// 
// DPH_89
// 
// 
// PC_89
// 
// 
// P2_89
// 
// 
// P3_89
// 
// 
// P0_89
// 
// 
// P1_89
// 
// 
// IRAM_89
// 
// 
// SP_89
// 
// 
// PSW_89
// 
// 
// ACC_8a
// 
// 
// P1_8a
// 
// 
// DPL_8a
// 
// 
// DPH_8a
// 
// 
// PC_8a
// 
// 
// P2_8a
// 
// 
// P3_8a
// 
// 
// P0_8a
// 
// 
// B_8a
// 
// 
// IRAM_8a
// 
// 
// SP_8a
// 
// 
// PSW_8a
// 
// 
// ACC_8b
// 
// 
// B_8b
// 
// 
// DPL_8b
// 
// 
// DPH_8b
// 
// 
// PC_8b
// 
// 
// P2_8b
// 
// 
// P3_8b
// 
// 
// P0_8b
// 
// 
// P1_8b
// 
// 
// IRAM_8b
// 
// 
// SP_8b
// 
// 
// PSW_8b
// 
// 
// ACC_8c
// 
// 
// B_8c
// 
// 
// DPL_8c
// 
// 
// DPH_8c
// 
// 
// PC_8c
// 
// 
// P2_8c
// 
// 
// P3_8c
// 
// 
// P0_8c
// 
// 
// P1_8c
// 
// 
// IRAM_8c
// 
// 
// SP_8c
// 
// 
// PSW_8c
// 
// 
// ACC_8d
// 
// 
// B_8d
// 
// 
// DPL_8d
// 
// 
// DPH_8d
// 
// 
// PC_8d
// 
// 
// P2_8d
// 
// 
// P3_8d
// 
// 
// P0_8d
// 
// 
// P1_8d
// 
// 
// IRAM_8d
// 
// 
// SP_8d
// 
// 
// PSW_8d
// 
// 
// ACC_8e
// 
// 
// B_8e
// 
// 
// DPL_8e
// 
// 
// DPH_8e
// 
// 
// PC_8e
// 
// 
// P2_8e
// 
// 
// P3_8e
// 
// 
// P0_8e
// 
// 
// P1_8e
// 
// 
// IRAM_8e
// 
// 
// SP_8e
// 
// 
// PSW_8e
// 
// 
// ACC_8f
// 
// 
// P1_8f
// 
// 
// DPL_8f
// 
// 
// DPH_8f
// 
// 
// PC_8f
// 
// 
// P2_8f
// 
// 
// P3_8f
// 
// 
// P0_8f
// 
// 
// B_8f
// 
// 
// IRAM_8f
// 
// 
// SP_8f
// 
// 
// PSW_8f
// 
// 
// ACC_90
// 
// 
// B_90
// 
// 
// DPL_90
// 
// 
// DPH_90
// 
// 
// PC_90
// 
// 
// P2_90
// 
// 
// P3_90
// 
// 
// P0_90
// 
// 
// P1_90
// 
// 
// SP_90
// 
// 
// PSW_90
// 
// 
// ACC_91
// 
// 
// P1_91
// 
// 
// DPL_91
// 
// 
// DPH_91
// 
// 
// PC_91
// 
// 
// P2_91
// 
// 
// P3_91
// 
// 
// P0_91
// 
// 
// B_91
// 
// 
// IRAM_91
// 
// 
// SP_91
// 
// 
// PSW_91
// 
// 
// ACC_92
// 
// 
// P1_92
// 
// 
// DPL_92
// 
// 
// DPH_92
// 
// 
// PC_92
// 
// 
// P2_92
// 
// 
// P3_92
// 
// 
// P0_92
// 
// 
// B_92
// 
// 
// IRAM_92
// 
assign n0236 = PSW[7:7];
assign n0237 = { 7'b0, n0236 };
assign n0238 = ( n0237 << n0120 );
assign n0239 = ( n0146 | n0238 );
// 
// SP_92
// 
// 
// PSW_92
// 
// 
// ACC_93
// 
// 
// B_93
// 
// 
// DPL_93
// 
// 
// DPH_93
// 
// 
// PC_93
// 
// 
// P2_93
// 
// 
// P3_93
// 
// 
// P0_93
// 
// 
// P1_93
// 
// 
// SP_93
// 
// 
// PSW_93
// 
// 
// ACC_94
// 
// 
// B_94
// 
// 
// DPL_94
// 
// 
// DPH_94
// 
// 
// PC_94
// 
// 
// P2_94
// 
// 
// P3_94
// 
// 
// P0_94
// 
// 
// P1_94
// 
// 
// SP_94
// 
// 
// PSW_94
// 
// 
// ACC_95
// 
// 
// B_95
// 
// 
// DPL_95
// 
// 
// DPH_95
// 
// 
// PC_95
// 
// 
// P2_95
// 
// 
// P3_95
// 
// 
// P0_95
// 
// 
// P1_95
// 
// 
// SP_95
// 
// 
// PSW_95
// 
// 
// ACC_96
// 
// 
// B_96
// 
// 
// DPL_96
// 
// 
// DPH_96
// 
// 
// PC_96
// 
// 
// P2_96
// 
// 
// P3_96
// 
// 
// P0_96
// 
// 
// P1_96
// 
// 
// SP_96
// 
// 
// PSW_96
// 
// 
// ACC_97
// 
// 
// P1_97
// 
// 
// DPL_97
// 
// 
// DPH_97
// 
// 
// PC_97
// 
// 
// P2_97
// 
// 
// P3_97
// 
// 
// P0_97
// 
// 
// B_97
// 
// 
// SP_97
// 
// 
// PSW_97
// 
// 
// ACC_98
// 
// 
// P1_98
// 
// 
// DPL_98
// 
// 
// DPH_98
// 
// 
// PC_98
// 
// 
// P2_98
// 
// 
// P3_98
// 
// 
// P0_98
// 
// 
// B_98
// 
// 
// SP_98
// 
// 
// PSW_98
// 
// 
// ACC_99
// 
// 
// B_99
// 
// 
// DPL_99
// 
// 
// DPH_99
// 
// 
// PC_99
// 
// 
// P2_99
// 
// 
// P3_99
// 
// 
// P0_99
// 
// 
// P1_99
// 
// 
// SP_99
// 
// 
// PSW_99
// 
// 
// ACC_9a
// 
// 
// B_9a
// 
// 
// DPL_9a
// 
// 
// DPH_9a
// 
// 
// PC_9a
// 
// 
// P2_9a
// 
// 
// P3_9a
// 
// 
// P0_9a
// 
// 
// P1_9a
// 
// 
// SP_9a
// 
// 
// PSW_9a
// 
// 
// ACC_9b
// 
// 
// B_9b
// 
// 
// DPL_9b
// 
// 
// DPH_9b
// 
// 
// PC_9b
// 
// 
// P2_9b
// 
// 
// P3_9b
// 
// 
// P0_9b
// 
// 
// P1_9b
// 
// 
// SP_9b
// 
// 
// PSW_9b
// 
// 
// ACC_9c
// 
// 
// B_9c
// 
// 
// DPL_9c
// 
// 
// DPH_9c
// 
// 
// PC_9c
// 
// 
// P2_9c
// 
// 
// P3_9c
// 
// 
// P0_9c
// 
// 
// P1_9c
// 
// 
// SP_9c
// 
// 
// PSW_9c
// 
// 
// ACC_9d
// 
// 
// B_9d
// 
// 
// DPL_9d
// 
// 
// DPH_9d
// 
// 
// PC_9d
// 
// 
// P2_9d
// 
// 
// P3_9d
// 
// 
// P0_9d
// 
// 
// P1_9d
// 
// 
// SP_9d
// 
// 
// PSW_9d
// 
// 
// ACC_9e
// 
// 
// B_9e
// 
// 
// DPL_9e
// 
// 
// DPH_9e
// 
// 
// PC_9e
// 
// 
// P2_9e
// 
// 
// P3_9e
// 
// 
// P0_9e
// 
// 
// P1_9e
// 
// 
// SP_9e
// 
// 
// PSW_9e
// 
// 
// ACC_9f
// 
// 
// B_9f
// 
// 
// DPL_9f
// 
// 
// DPH_9f
// 
// 
// PC_9f
// 
// 
// P2_9f
// 
// 
// P3_9f
// 
// 
// P0_9f
// 
// 
// P1_9f
// 
// 
// SP_9f
// 
// 
// PSW_9f
// 
// 
// ACC_a0
// 
// 
// B_a0
// 
// 
// DPL_a0
// 
// 
// DPH_a0
// 
// 
// PC_a0
// 
// 
// P2_a0
// 
// 
// P3_a0
// 
// 
// P0_a0
// 
// 
// P1_a0
// 
// 
// SP_a0
// 
// 
// PSW_a0
// 
// 
// ACC_a1
// 
// 
// B_a1
// 
// 
// DPL_a1
// 
// 
// DPH_a1
// 
// 
// PC_a1
// 
// 
// P2_a1
// 
// 
// P3_a1
// 
// 
// P0_a1
// 
// 
// P1_a1
// 
// 
// SP_a1
// 
// 
// PSW_a1
// 
// 
// ACC_a2
// 
// 
// P1_a2
// 
// 
// DPL_a2
// 
// 
// DPH_a2
// 
// 
// PC_a2
// 
// 
// P2_a2
// 
// 
// P3_a2
// 
// 
// P0_a2
// 
// 
// B_a2
// 
// 
// SP_a2
// 
// 
// PSW_a2
// 
// 
// ACC_a3
// 
// 
// P1_a3
// 
// 
// DPL_a3
// 
// 
// DPH_a3
// 
// 
// PC_a3
// 
// 
// P2_a3
// 
// 
// P3_a3
// 
// 
// P0_a3
// 
// 
// B_a3
// 
// 
// SP_a3
// 
// 
// PSW_a3
// 
// 
// ACC_a4
// 
// 
// P1_a4
// 
// 
// DPL_a4
// 
// 
// DPH_a4
// 
// 
// PC_a4
// 
// 
// P2_a4
// 
// 
// P3_a4
// 
// 
// P0_a4
// 
// 
// B_a4
// 
// 
// SP_a4
// 
// 
// PSW_a4
// 
// 
// ACC_a5
// 
// 
// P1_a5
// 
// 
// DPL_a5
// 
// 
// DPH_a5
// 
// 
// PC_a5
// 
// 
// P2_a5
// 
// 
// P3_a5
// 
// 
// P0_a5
// 
// 
// B_a5
// 
// 
// SP_a5
// 
// 
// PSW_a5
// 
// 
// ACC_a6
// 
// 
// B_a6
// 
// 
// DPL_a6
// 
// 
// DPH_a6
// 
// 
// PC_a6
// 
// 
// P2_a6
// 
// 
// P3_a6
// 
// 
// P0_a6
// 
// 
// P1_a6
// 
// 
// IRAM_a6
// 
assign n0240 = ( n0050 ) ? ( P3INREG ) : ( n0063 );
assign n0241 = ( n0048 ) ? ( IE ) : ( n0240 );
assign n0242 = ( n0046 ) ? ( P2INREG ) : ( n0241 );
assign n0243 = ( n0044 ) ? ( SBUF ) : ( n0242 );
assign n0244 = ( n0042 ) ? ( SCON ) : ( n0243 );
assign n0245 = ( n0040 ) ? ( P1INREG ) : ( n0244 );
assign n0246 = ( n0038 ) ? ( TH1 ) : ( n0245 );
assign n0247 = ( n0036 ) ? ( TL1 ) : ( n0246 );
assign n0248 = ( n0034 ) ? ( TH0 ) : ( n0247 );
assign n0249 = ( n0032 ) ? ( TL0 ) : ( n0248 );
assign n0250 = ( n0030 ) ? ( TMOD ) : ( n0249 );
assign n0251 = ( n0028 ) ? ( TCON ) : ( n0250 );
assign n0252 = ( n0026 ) ? ( PCON ) : ( n0251 );
assign n0253 = ( n0024 ) ? ( DPH ) : ( n0252 );
assign n0254 = ( n0022 ) ? ( DPL ) : ( n0253 );
assign n0255 = ( n0020 ) ? ( SP ) : ( n0254 );
assign n0256 = ( n0018 ) ? ( P0INREG ) : ( n0255 );
assign n0257 = ( n0015 ) ? ( RD_IRAM_1 ) : ( n0256 );
// 
// SP_a6
// 
// 
// PSW_a6
// 
// 
// ACC_a7
// 
// 
// B_a7
// 
// 
// DPL_a7
// 
// 
// DPH_a7
// 
// 
// PC_a7
// 
// 
// P2_a7
// 
// 
// P3_a7
// 
// 
// P0_a7
// 
// 
// P1_a7
// 
// 
// IRAM_a7
// 
// 
// SP_a7
// 
// 
// PSW_a7
// 
// 
// ACC_a8
// 
// 
// P1_a8
// 
// 
// DPL_a8
// 
// 
// DPH_a8
// 
// 
// PC_a8
// 
// 
// P2_a8
// 
// 
// P3_a8
// 
// 
// P0_a8
// 
// 
// B_a8
// 
// 
// IRAM_a8
// 
assign n0258 = ( n0015 ) ? ( RD_IRAM_0 ) : ( n0256 );
// 
// SP_a8
// 
// 
// PSW_a8
// 
// 
// ACC_a9
// 
// 
// B_a9
// 
// 
// DPL_a9
// 
// 
// DPH_a9
// 
// 
// PC_a9
// 
// 
// P2_a9
// 
// 
// P3_a9
// 
// 
// P0_a9
// 
// 
// P1_a9
// 
// 
// IRAM_a9
// 
// 
// SP_a9
// 
// 
// PSW_a9
// 
// 
// ACC_aa
// 
// 
// B_aa
// 
// 
// DPL_aa
// 
// 
// DPH_aa
// 
// 
// PC_aa
// 
// 
// P2_aa
// 
// 
// P3_aa
// 
// 
// P0_aa
// 
// 
// P1_aa
// 
// 
// IRAM_aa
// 
// 
// SP_aa
// 
// 
// PSW_aa
// 
// 
// ACC_ab
// 
// 
// P1_ab
// 
// 
// DPL_ab
// 
// 
// DPH_ab
// 
// 
// PC_ab
// 
// 
// P2_ab
// 
// 
// P3_ab
// 
// 
// P0_ab
// 
// 
// B_ab
// 
// 
// IRAM_ab
// 
// 
// SP_ab
// 
// 
// PSW_ab
// 
// 
// ACC_ac
// 
// 
// B_ac
// 
// 
// DPL_ac
// 
// 
// DPH_ac
// 
// 
// PC_ac
// 
// 
// P2_ac
// 
// 
// P3_ac
// 
// 
// P0_ac
// 
// 
// P1_ac
// 
// 
// IRAM_ac
// 
// 
// SP_ac
// 
// 
// PSW_ac
// 
// 
// ACC_ad
// 
// 
// B_ad
// 
// 
// DPL_ad
// 
// 
// DPH_ad
// 
// 
// PC_ad
// 
// 
// P2_ad
// 
// 
// P3_ad
// 
// 
// P0_ad
// 
// 
// P1_ad
// 
// 
// IRAM_ad
// 
// 
// SP_ad
// 
// 
// PSW_ad
// 
// 
// ACC_ae
// 
// 
// B_ae
// 
// 
// DPL_ae
// 
// 
// DPH_ae
// 
// 
// PC_ae
// 
// 
// P2_ae
// 
// 
// P3_ae
// 
// 
// P0_ae
// 
// 
// P1_ae
// 
// 
// IRAM_ae
// 
// 
// SP_ae
// 
// 
// PSW_ae
// 
// 
// ACC_af
// 
// 
// B_af
// 
// 
// DPL_af
// 
// 
// DPH_af
// 
// 
// PC_af
// 
// 
// P2_af
// 
// 
// P3_af
// 
// 
// P0_af
// 
// 
// P1_af
// 
// 
// IRAM_af
// 
// 
// SP_af
// 
// 
// PSW_af
// 
// 
// ACC_b0
// 
// 
// B_b0
// 
// 
// DPL_b0
// 
// 
// DPH_b0
// 
// 
// PC_b0
// 
// 
// P2_b0
// 
// 
// P3_b0
// 
// 
// P0_b0
// 
// 
// P1_b0
// 
// 
// SP_b0
// 
// 
// PSW_b0
// 
// 
// ACC_b1
// 
// 
// B_b1
// 
// 
// DPL_b1
// 
// 
// DPH_b1
// 
// 
// PC_b1
// 
// 
// P2_b1
// 
// 
// P3_b1
// 
// 
// P0_b1
// 
// 
// P1_b1
// 
// 
// IRAM_b1
// 
// 
// SP_b1
// 
// 
// PSW_b1
// 
// 
// ACC_b2
// 
// 
// P1_b2
// 
// 
// DPL_b2
// 
// 
// DPH_b2
// 
// 
// PC_b2
// 
// 
// P2_b2
// 
// 
// P3_b2
// 
// 
// P0_b2
// 
// 
// B_b2
// 
// 
// IRAM_b2
// 
assign n0259 = ( n0129 ) ? ( P3 ) : ( n0137 );
assign n0260 = ( n0128 ) ? ( IE ) : ( n0259 );
assign n0261 = ( n0127 ) ? ( P2 ) : ( n0260 );
assign n0262 = ( n0126 ) ? ( SCON ) : ( n0261 );
assign n0263 = ( n0125 ) ? ( P1 ) : ( n0262 );
assign n0264 = ( n0124 ) ? ( TCON ) : ( n0263 );
assign n0265 = ( n0123 ) ? ( P0 ) : ( n0264 );
assign n0266 = ( n0117 ) ? ( RD_IRAM_0 ) : ( n0265 );
assign n0267 = ( n0122 & n0266 );
assign n0268 = n0266[n0119];
assign n0269 = ~( n0268 );
assign n0270 = { 7'b0, n0269 };
assign n0271 = ( n0270 << n0120 );
assign n0272 = ( n0267 | n0271 );
// 
// SP_b2
// 
// 
// PSW_b2
// 
// 
// ACC_b3
// 
// 
// B_b3
// 
// 
// DPL_b3
// 
// 
// DPH_b3
// 
// 
// PC_b3
// 
// 
// P2_b3
// 
// 
// P3_b3
// 
// 
// P0_b3
// 
// 
// P1_b3
// 
// 
// SP_b3
// 
// 
// PSW_b3
// 
// 
// ACC_b4
// 
// 
// P1_b4
// 
// 
// DPL_b4
// 
// 
// DPH_b4
// 
// 
// PC_b4
// 
// 
// P2_b4
// 
// 
// P3_b4
// 
// 
// P0_b4
// 
// 
// B_b4
// 
// 
// SP_b4
// 
// 
// PSW_b4
// 
// 
// ACC_b5
// 
// 
// P1_b5
// 
// 
// DPL_b5
// 
// 
// DPH_b5
// 
// 
// PC_b5
// 
// 
// P2_b5
// 
// 
// P3_b5
// 
// 
// P0_b5
// 
// 
// B_b5
// 
// 
// SP_b5
// 
// 
// PSW_b5
// 
// 
// ACC_b6
// 
// 
// P1_b6
// 
// 
// DPL_b6
// 
// 
// DPH_b6
// 
// 
// PC_b6
// 
// 
// P2_b6
// 
// 
// P3_b6
// 
// 
// P0_b6
// 
// 
// B_b6
// 
// 
// SP_b6
// 
// 
// PSW_b6
// 
// 
// ACC_b7
// 
// 
// B_b7
// 
// 
// DPL_b7
// 
// 
// DPH_b7
// 
// 
// PC_b7
// 
// 
// P2_b7
// 
// 
// P3_b7
// 
// 
// P0_b7
// 
// 
// P1_b7
// 
// 
// SP_b7
// 
// 
// PSW_b7
// 
// 
// ACC_b8
// 
// 
// B_b8
// 
// 
// DPL_b8
// 
// 
// DPH_b8
// 
// 
// PC_b8
// 
// 
// P2_b8
// 
// 
// P3_b8
// 
// 
// P0_b8
// 
// 
// P1_b8
// 
// 
// SP_b8
// 
// 
// PSW_b8
// 
// 
// ACC_b9
// 
// 
// P1_b9
// 
// 
// DPL_b9
// 
// 
// DPH_b9
// 
// 
// PC_b9
// 
// 
// P2_b9
// 
// 
// P3_b9
// 
// 
// P0_b9
// 
// 
// B_b9
// 
// 
// SP_b9
// 
// 
// PSW_b9
// 
// 
// ACC_ba
// 
// 
// P1_ba
// 
// 
// DPL_ba
// 
// 
// DPH_ba
// 
// 
// PC_ba
// 
// 
// P2_ba
// 
// 
// P3_ba
// 
// 
// P0_ba
// 
// 
// B_ba
// 
// 
// SP_ba
// 
// 
// PSW_ba
// 
// 
// ACC_bb
// 
// 
// B_bb
// 
// 
// DPL_bb
// 
// 
// DPH_bb
// 
// 
// PC_bb
// 
// 
// P2_bb
// 
// 
// P3_bb
// 
// 
// P0_bb
// 
// 
// P1_bb
// 
// 
// SP_bb
// 
// 
// PSW_bb
// 
// 
// ACC_bc
// 
// 
// P1_bc
// 
// 
// DPL_bc
// 
// 
// DPH_bc
// 
// 
// PC_bc
// 
// 
// P2_bc
// 
// 
// P3_bc
// 
// 
// P0_bc
// 
// 
// B_bc
// 
// 
// SP_bc
// 
// 
// PSW_bc
// 
// 
// ACC_bd
// 
// 
// B_bd
// 
// 
// DPL_bd
// 
// 
// DPH_bd
// 
// 
// PC_bd
// 
// 
// P2_bd
// 
// 
// P3_bd
// 
// 
// P0_bd
// 
// 
// P1_bd
// 
// 
// SP_bd
// 
// 
// PSW_bd
// 
// 
// ACC_be
// 
// 
// B_be
// 
// 
// DPL_be
// 
// 
// DPH_be
// 
// 
// PC_be
// 
// 
// P2_be
// 
// 
// P3_be
// 
// 
// P0_be
// 
// 
// P1_be
// 
// 
// SP_be
// 
// 
// PSW_be
// 
// 
// ACC_bf
// 
// 
// B_bf
// 
// 
// DPL_bf
// 
// 
// DPH_bf
// 
// 
// PC_bf
// 
// 
// P2_bf
// 
// 
// P3_bf
// 
// 
// P0_bf
// 
// 
// P1_bf
// 
// 
// SP_bf
// 
// 
// PSW_bf
// 
// 
// ACC_c0
// 
// 
// B_c0
// 
// 
// DPL_c0
// 
// 
// DPH_c0
// 
// 
// PC_c0
// 
// 
// P2_c0
// 
// 
// P3_c0
// 
// 
// P0_c0
// 
// 
// P1_c0
// 
// 
// IRAM_c0
// 
// 
// SP_c0
// 
// 
// PSW_c0
// 
// 
// ACC_c1
// 
// 
// B_c1
// 
// 
// DPL_c1
// 
// 
// DPH_c1
// 
// 
// PC_c1
// 
// 
// P2_c1
// 
// 
// P3_c1
// 
// 
// P0_c1
// 
// 
// P1_c1
// 
// 
// SP_c1
// 
// 
// PSW_c1
// 
// 
// ACC_c2
// 
// 
// P1_c2
// 
// 
// DPL_c2
// 
// 
// DPH_c2
// 
// 
// PC_c2
// 
// 
// P2_c2
// 
// 
// P3_c2
// 
// 
// P0_c2
// 
// 
// B_c2
// 
// 
// IRAM_c2
// 
assign n0273 = ( n0267 | n0148 );
// 
// SP_c2
// 
// 
// PSW_c2
// 
// 
// ACC_c3
// 
// 
// B_c3
// 
// 
// DPL_c3
// 
// 
// DPH_c3
// 
// 
// PC_c3
// 
// 
// P2_c3
// 
// 
// P3_c3
// 
// 
// P0_c3
// 
// 
// P1_c3
// 
// 
// SP_c3
// 
// 
// PSW_c3
// 
// 
// ACC_c4
// 
// 
// P1_c4
// 
// 
// DPL_c4
// 
// 
// DPH_c4
// 
// 
// PC_c4
// 
// 
// P2_c4
// 
// 
// P3_c4
// 
// 
// P0_c4
// 
// 
// B_c4
// 
// 
// SP_c4
// 
// 
// PSW_c4
// 
// 
// ACC_c5
// 
// 
// P1_c5
// 
// 
// DPL_c5
// 
// 
// DPH_c5
// 
// 
// PC_c5
// 
// 
// P2_c5
// 
// 
// P3_c5
// 
// 
// P0_c5
// 
// 
// B_c5
// 
// 
// IRAM_c5
// 
// 
// SP_c5
// 
// 
// PSW_c5
// 
// 
// ACC_c6
// 
// 
// B_c6
// 
// 
// DPL_c6
// 
// 
// DPH_c6
// 
// 
// PC_c6
// 
// 
// P2_c6
// 
// 
// P3_c6
// 
// 
// P0_c6
// 
// 
// P1_c6
// 
// 
// IRAM_c6
// 
// 
// SP_c6
// 
// 
// PSW_c6
// 
// 
// ACC_c7
// 
// 
// P1_c7
// 
// 
// DPL_c7
// 
// 
// DPH_c7
// 
// 
// PC_c7
// 
// 
// P2_c7
// 
// 
// P3_c7
// 
// 
// P0_c7
// 
// 
// B_c7
// 
// 
// IRAM_c7
// 
// 
// SP_c7
// 
// 
// PSW_c7
// 
// 
// ACC_c8
// 
// 
// B_c8
// 
// 
// DPL_c8
// 
// 
// DPH_c8
// 
// 
// PC_c8
// 
// 
// P2_c8
// 
// 
// P3_c8
// 
// 
// P0_c8
// 
// 
// P1_c8
// 
// 
// IRAM_c8
// 
// 
// SP_c8
// 
// 
// PSW_c8
// 
// 
// ACC_c9
// 
// 
// B_c9
// 
// 
// DPL_c9
// 
// 
// DPH_c9
// 
// 
// PC_c9
// 
// 
// P2_c9
// 
// 
// P3_c9
// 
// 
// P0_c9
// 
// 
// P1_c9
// 
// 
// IRAM_c9
// 
// 
// SP_c9
// 
// 
// PSW_c9
// 
// 
// ACC_ca
// 
// 
// B_ca
// 
// 
// DPL_ca
// 
// 
// DPH_ca
// 
// 
// PC_ca
// 
// 
// P2_ca
// 
// 
// P3_ca
// 
// 
// P0_ca
// 
// 
// P1_ca
// 
// 
// IRAM_ca
// 
// 
// SP_ca
// 
// 
// PSW_ca
// 
// 
// ACC_cb
// 
// 
// P1_cb
// 
// 
// DPL_cb
// 
// 
// DPH_cb
// 
// 
// PC_cb
// 
// 
// P2_cb
// 
// 
// P3_cb
// 
// 
// P0_cb
// 
// 
// B_cb
// 
// 
// IRAM_cb
// 
// 
// SP_cb
// 
// 
// PSW_cb
// 
// 
// ACC_cc
// 
// 
// B_cc
// 
// 
// DPL_cc
// 
// 
// DPH_cc
// 
// 
// PC_cc
// 
// 
// P2_cc
// 
// 
// P3_cc
// 
// 
// P0_cc
// 
// 
// P1_cc
// 
// 
// IRAM_cc
// 
// 
// SP_cc
// 
// 
// PSW_cc
// 
// 
// ACC_cd
// 
// 
// B_cd
// 
// 
// DPL_cd
// 
// 
// DPH_cd
// 
// 
// PC_cd
// 
// 
// P2_cd
// 
// 
// P3_cd
// 
// 
// P0_cd
// 
// 
// P1_cd
// 
// 
// IRAM_cd
// 
// 
// SP_cd
// 
// 
// PSW_cd
// 
// 
// ACC_ce
// 
// 
// B_ce
// 
// 
// DPL_ce
// 
// 
// DPH_ce
// 
// 
// PC_ce
// 
// 
// P2_ce
// 
// 
// P3_ce
// 
// 
// P0_ce
// 
// 
// P1_ce
// 
// 
// IRAM_ce
// 
// 
// SP_ce
// 
// 
// PSW_ce
// 
// 
// ACC_cf
// 
// 
// B_cf
// 
// 
// DPL_cf
// 
// 
// DPH_cf
// 
// 
// PC_cf
// 
// 
// P2_cf
// 
// 
// P3_cf
// 
// 
// P0_cf
// 
// 
// P1_cf
// 
// 
// IRAM_cf
// 
// 
// SP_cf
// 
// 
// PSW_cf
// 
// 
// ACC_d0
// 
// 
// B_d0
// 
// 
// DPL_d0
// 
// 
// DPH_d0
// 
// 
// PC_d0
// 
// 
// P2_d0
// 
// 
// P3_d0
// 
// 
// P0_d0
// 
// 
// P1_d0
// 
// 
// IRAM_d0
// 
// 
// SP_d0
// 
// 
// PSW_d0
// 
// 
// ACC_d1
// 
// 
// B_d1
// 
// 
// DPL_d1
// 
// 
// DPH_d1
// 
// 
// PC_d1
// 
// 
// P2_d1
// 
// 
// P3_d1
// 
// 
// P0_d1
// 
// 
// P1_d1
// 
// 
// IRAM_d1
// 
// 
// SP_d1
// 
// 
// PSW_d1
// 
// 
// ACC_d2
// 
// 
// P1_d2
// 
// 
// DPL_d2
// 
// 
// DPH_d2
// 
// 
// PC_d2
// 
// 
// P2_d2
// 
// 
// P3_d2
// 
// 
// P0_d2
// 
// 
// B_d2
// 
// 
// IRAM_d2
// 
assign n0274 = { 7'b0, n0108 };
assign n0275 = ( n0274 << n0120 );
assign n0276 = ( n0267 | n0275 );
// 
// SP_d2
// 
// 
// PSW_d2
// 
// 
// ACC_d3
// 
// 
// B_d3
// 
// 
// DPL_d3
// 
// 
// DPH_d3
// 
// 
// PC_d3
// 
// 
// P2_d3
// 
// 
// P3_d3
// 
// 
// P0_d3
// 
// 
// P1_d3
// 
// 
// SP_d3
// 
// 
// PSW_d3
// 
// 
// ACC_d4
// 
// 
// P1_d4
// 
// 
// DPL_d4
// 
// 
// DPH_d4
// 
// 
// PC_d4
// 
// 
// P2_d4
// 
// 
// P3_d4
// 
// 
// P0_d4
// 
// 
// B_d4
// 
// 
// SP_d4
// 
// 
// PSW_d4
// 
// 
// ACC_d5
// 
// 
// B_d5
// 
// 
// DPL_d5
// 
// 
// DPH_d5
// 
// 
// PC_d5
// 
// 
// P2_d5
// 
// 
// P3_d5
// 
// 
// P0_d5
// 
// 
// P1_d5
// 
// 
// IRAM_d5
// 
// 
// SP_d5
// 
// 
// PSW_d5
// 
// 
// ACC_d6
// 
// 
// B_d6
// 
// 
// DPL_d6
// 
// 
// DPH_d6
// 
// 
// PC_d6
// 
// 
// P2_d6
// 
// 
// P3_d6
// 
// 
// P0_d6
// 
// 
// P1_d6
// 
// 
// IRAM_d6
// 
assign n0277 = RD_IRAM_1[7:4];
assign n0278 = ACC[3:0];
assign n0279 = { ( n0277 ), ( n0278 ) };
// 
// SP_d6
// 
// 
// PSW_d6
// 
// 
// ACC_d7
// 
// 
// P1_d7
// 
// 
// DPL_d7
// 
// 
// DPH_d7
// 
// 
// PC_d7
// 
// 
// P2_d7
// 
// 
// P3_d7
// 
// 
// P0_d7
// 
// 
// B_d7
// 
// 
// IRAM_d7
// 
// 
// SP_d7
// 
// 
// PSW_d7
// 
// 
// ACC_d8
// 
// 
// B_d8
// 
// 
// DPL_d8
// 
// 
// DPH_d8
// 
// 
// PC_d8
// 
// 
// P2_d8
// 
// 
// P3_d8
// 
// 
// P0_d8
// 
// 
// P1_d8
// 
// 
// IRAM_d8
// 
// 
// SP_d8
// 
// 
// PSW_d8
// 
// 
// ACC_d9
// 
// 
// P1_d9
// 
// 
// DPL_d9
// 
// 
// DPH_d9
// 
// 
// PC_d9
// 
// 
// P2_d9
// 
// 
// P3_d9
// 
// 
// P0_d9
// 
// 
// B_d9
// 
// 
// IRAM_d9
// 
// 
// SP_d9
// 
// 
// PSW_d9
// 
// 
// ACC_da
// 
// 
// B_da
// 
// 
// DPL_da
// 
// 
// DPH_da
// 
// 
// PC_da
// 
// 
// P2_da
// 
// 
// P3_da
// 
// 
// P0_da
// 
// 
// P1_da
// 
// 
// IRAM_da
// 
// 
// SP_da
// 
// 
// PSW_da
// 
// 
// ACC_db
// 
// 
// B_db
// 
// 
// DPL_db
// 
// 
// DPH_db
// 
// 
// PC_db
// 
// 
// P2_db
// 
// 
// P3_db
// 
// 
// P0_db
// 
// 
// P1_db
// 
// 
// IRAM_db
// 
// 
// SP_db
// 
// 
// PSW_db
// 
// 
// ACC_dc
// 
// 
// P1_dc
// 
// 
// DPL_dc
// 
// 
// DPH_dc
// 
// 
// PC_dc
// 
// 
// P2_dc
// 
// 
// P3_dc
// 
// 
// P0_dc
// 
// 
// B_dc
// 
// 
// IRAM_dc
// 
// 
// SP_dc
// 
// 
// PSW_dc
// 
// 
// ACC_dd
// 
// 
// P1_dd
// 
// 
// DPL_dd
// 
// 
// DPH_dd
// 
// 
// PC_dd
// 
// 
// P2_dd
// 
// 
// P3_dd
// 
// 
// P0_dd
// 
// 
// B_dd
// 
// 
// IRAM_dd
// 
// 
// SP_dd
// 
// 
// PSW_dd
// 
// 
// ACC_de
// 
// 
// B_de
// 
// 
// DPL_de
// 
// 
// DPH_de
// 
// 
// PC_de
// 
// 
// P2_de
// 
// 
// P3_de
// 
// 
// P0_de
// 
// 
// P1_de
// 
// 
// IRAM_de
// 
// 
// SP_de
// 
// 
// PSW_de
// 
// 
// ACC_df
// 
// 
// B_df
// 
// 
// DPL_df
// 
// 
// DPH_df
// 
// 
// PC_df
// 
// 
// P2_df
// 
// 
// P3_df
// 
// 
// P0_df
// 
// 
// P1_df
// 
// 
// IRAM_df
// 
// 
// SP_df
// 
// 
// PSW_df
// 
// 
// ACC_e1
// 
// 
// P1_e1
// 
// 
// DPL_e1
// 
// 
// DPH_e1
// 
// 
// PC_e1
// 
// 
// P2_e1
// 
// 
// P3_e1
// 
// 
// P0_e1
// 
// 
// B_e1
// 
// 
// SP_e1
// 
// 
// PSW_e1
// 
// 
// ACC_e4
// 
// 
// P1_e4
// 
// 
// DPL_e4
// 
// 
// DPH_e4
// 
// 
// PC_e4
// 
// 
// P2_e4
// 
// 
// P3_e4
// 
// 
// P0_e4
// 
// 
// B_e4
// 
// 
// SP_e4
// 
// 
// PSW_e4
// 
// 
// ACC_e5
// 
// 
// P1_e5
// 
// 
// DPL_e5
// 
// 
// DPH_e5
// 
// 
// PC_e5
// 
// 
// P2_e5
// 
// 
// P3_e5
// 
// 
// P0_e5
// 
// 
// B_e5
// 
// 
// SP_e5
// 
// 
// PSW_e5
// 
// 
// ACC_e6
// 
// 
// P1_e6
// 
// 
// DPL_e6
// 
// 
// DPH_e6
// 
// 
// PC_e6
// 
// 
// P2_e6
// 
// 
// P3_e6
// 
// 
// P0_e6
// 
// 
// B_e6
// 
// 
// SP_e6
// 
// 
// PSW_e6
// 
// 
// ACC_e7
// 
// 
// B_e7
// 
// 
// DPL_e7
// 
// 
// DPH_e7
// 
// 
// PC_e7
// 
// 
// P2_e7
// 
// 
// P3_e7
// 
// 
// P0_e7
// 
// 
// P1_e7
// 
// 
// SP_e7
// 
// 
// PSW_e7
// 
// 
// ACC_e8
// 
// 
// B_e8
// 
// 
// DPL_e8
// 
// 
// DPH_e8
// 
// 
// PC_e8
// 
// 
// P2_e8
// 
// 
// P3_e8
// 
// 
// P0_e8
// 
// 
// P1_e8
// 
// 
// SP_e8
// 
// 
// PSW_e8
// 
// 
// ACC_e9
// 
// 
// B_e9
// 
// 
// DPL_e9
// 
// 
// DPH_e9
// 
// 
// PC_e9
// 
// 
// P2_e9
// 
// 
// P3_e9
// 
// 
// P0_e9
// 
// 
// P1_e9
// 
// 
// SP_e9
// 
// 
// PSW_e9
// 
// 
// ACC_ea
// 
// 
// B_ea
// 
// 
// DPL_ea
// 
// 
// DPH_ea
// 
// 
// PC_ea
// 
// 
// P2_ea
// 
// 
// P3_ea
// 
// 
// P0_ea
// 
// 
// P1_ea
// 
// 
// SP_ea
// 
// 
// PSW_ea
// 
// 
// ACC_eb
// 
// 
// P1_eb
// 
// 
// DPL_eb
// 
// 
// DPH_eb
// 
// 
// PC_eb
// 
// 
// P2_eb
// 
// 
// P3_eb
// 
// 
// P0_eb
// 
// 
// B_eb
// 
// 
// SP_eb
// 
// 
// PSW_eb
// 
// 
// ACC_ec
// 
// 
// B_ec
// 
// 
// DPL_ec
// 
// 
// DPH_ec
// 
// 
// PC_ec
// 
// 
// P2_ec
// 
// 
// P3_ec
// 
// 
// P0_ec
// 
// 
// P1_ec
// 
// 
// SP_ec
// 
// 
// PSW_ec
// 
// 
// ACC_ed
// 
// 
// B_ed
// 
// 
// DPL_ed
// 
// 
// DPH_ed
// 
// 
// PC_ed
// 
// 
// P2_ed
// 
// 
// P3_ed
// 
// 
// P0_ed
// 
// 
// P1_ed
// 
// 
// SP_ed
// 
// 
// PSW_ed
// 
// 
// ACC_ee
// 
// 
// P1_ee
// 
// 
// DPL_ee
// 
// 
// DPH_ee
// 
// 
// PC_ee
// 
// 
// P2_ee
// 
// 
// P3_ee
// 
// 
// P0_ee
// 
// 
// B_ee
// 
// 
// SP_ee
// 
// 
// PSW_ee
// 
// 
// ACC_ef
// 
// 
// P1_ef
// 
// 
// DPL_ef
// 
// 
// DPH_ef
// 
// 
// PC_ef
// 
// 
// P2_ef
// 
// 
// P3_ef
// 
// 
// P0_ef
// 
// 
// B_ef
// 
// 
// SP_ef
// 
// 
// PSW_ef
// 
// 
// ACC_f1
// 
// 
// P1_f1
// 
// 
// DPL_f1
// 
// 
// DPH_f1
// 
// 
// PC_f1
// 
// 
// P2_f1
// 
// 
// P3_f1
// 
// 
// P0_f1
// 
// 
// B_f1
// 
// 
// IRAM_f1
// 
// 
// SP_f1
// 
// 
// PSW_f1
// 
// 
// ACC_f4
// 
// 
// B_f4
// 
// 
// DPL_f4
// 
// 
// DPH_f4
// 
// 
// PC_f4
// 
// 
// P2_f4
// 
// 
// P3_f4
// 
// 
// P0_f4
// 
// 
// P1_f4
// 
// 
// SP_f4
// 
// 
// PSW_f4
// 
// 
// ACC_f5
// 
// 
// P1_f5
// 
// 
// DPL_f5
// 
// 
// DPH_f5
// 
// 
// PC_f5
// 
// 
// P2_f5
// 
// 
// P3_f5
// 
// 
// P0_f5
// 
// 
// B_f5
// 
// 
// IRAM_f5
// 
// 
// SP_f5
// 
// 
// PSW_f5
// 
// 
// ACC_f6
// 
// 
// P1_f6
// 
// 
// DPL_f6
// 
// 
// DPH_f6
// 
// 
// PC_f6
// 
// 
// P2_f6
// 
// 
// P3_f6
// 
// 
// P0_f6
// 
// 
// B_f6
// 
// 
// IRAM_f6
// 
// 
// SP_f6
// 
// 
// PSW_f6
// 
// 
// ACC_f7
// 
// 
// P1_f7
// 
// 
// DPL_f7
// 
// 
// DPH_f7
// 
// 
// PC_f7
// 
// 
// P2_f7
// 
// 
// P3_f7
// 
// 
// P0_f7
// 
// 
// B_f7
// 
// 
// IRAM_f7
// 
// 
// SP_f7
// 
// 
// PSW_f7
// 
// 
// ACC_f8
// 
// 
// B_f8
// 
// 
// DPL_f8
// 
// 
// DPH_f8
// 
// 
// PC_f8
// 
// 
// P2_f8
// 
// 
// P3_f8
// 
// 
// P0_f8
// 
// 
// P1_f8
// 
// 
// IRAM_f8
// 
// 
// SP_f8
// 
// 
// PSW_f8
// 
// 
// ACC_f9
// 
// 
// B_f9
// 
// 
// DPL_f9
// 
// 
// DPH_f9
// 
// 
// PC_f9
// 
// 
// P2_f9
// 
// 
// P3_f9
// 
// 
// P0_f9
// 
// 
// P1_f9
// 
// 
// IRAM_f9
// 
// 
// SP_f9
// 
// 
// PSW_f9
// 
// 
// ACC_fa
// 
// 
// B_fa
// 
// 
// DPL_fa
// 
// 
// DPH_fa
// 
// 
// PC_fa
// 
// 
// P2_fa
// 
// 
// P3_fa
// 
// 
// P0_fa
// 
// 
// P1_fa
// 
// 
// IRAM_fa
// 
// 
// SP_fa
// 
// 
// PSW_fa
// 
// 
// ACC_fb
// 
// 
// B_fb
// 
// 
// DPL_fb
// 
// 
// DPH_fb
// 
// 
// PC_fb
// 
// 
// P2_fb
// 
// 
// P3_fb
// 
// 
// P0_fb
// 
// 
// P1_fb
// 
// 
// IRAM_fb
// 
// 
// SP_fb
// 
// 
// PSW_fb
// 
// 
// ACC_fc
// 
// 
// B_fc
// 
// 
// DPL_fc
// 
// 
// DPH_fc
// 
// 
// PC_fc
// 
// 
// P2_fc
// 
// 
// P3_fc
// 
// 
// P0_fc
// 
// 
// P1_fc
// 
// 
// IRAM_fc
// 
// 
// SP_fc
// 
// 
// PSW_fc
// 
// 
// ACC_fd
// 
// 
// B_fd
// 
// 
// DPL_fd
// 
// 
// DPH_fd
// 
// 
// PC_fd
// 
// 
// P2_fd
// 
// 
// P3_fd
// 
// 
// P0_fd
// 
// 
// P1_fd
// 
// 
// IRAM_fd
// 
// 
// SP_fd
// 
// 
// PSW_fd
// 
// 
// ACC_fe
// 
// 
// B_fe
// 
// 
// DPL_fe
// 
// 
// DPH_fe
// 
// 
// PC_fe
// 
// 
// P2_fe
// 
// 
// P3_fe
// 
// 
// P0_fe
// 
// 
// P1_fe
// 
// 
// IRAM_fe
// 
// 
// SP_fe
// 
// 
// PSW_fe
// 
// 
// ACC_ff
// 
// 
// B_ff
// 
// 
// DPL_ff
// 
// 
// DPH_ff
// 
// 
// PC_ff
// 
// 
// P2_ff
// 
// 
// P3_ff
// 
// 
// P0_ff
// 
// 
// P1_ff
// 
// 
// IRAM_ff
// 
// 
// SP_ff
// 
// 
// PSW_ff
// 
assign ACC_next =   ( n0002 ) ? ( ACC_4b ) :  ( ACC_abstr );
assign P2_next =   ( n0002 ) ? ( P2_4b ) :  ( P2_abstr );
assign P0_next =   ( n0002 ) ? ( P0_4b ) :  ( P0_abstr );
assign P1_next =   ( n0002 ) ? ( P1_4b ) :  ( P1_abstr );
assign P3_next =   ( n0002 ) ? ( P3_4b ) :  ( P3_abstr );
assign SP_next =   ( n0002 ) ? ( SP_4b ) :  ( SP_abstr );
assign PC_next =   ( n0002 ) ? ( PC_4b ) :  ( PC_abstr );
assign B_next =   ( n0002 ) ? ( B_4b ) :  ( B_abstr );
assign DPL_next =   ( n0002 ) ? ( DPL_4b ) :  ( DPL_abstr );
assign PSW_next =   ( n0002 ) ? ( PSW_4b ) :  ( PSW_abstr );
assign DPH_next =   ( n0002 ) ? ( DPH_4b ) :  ( DPH_abstr );
assign n0280 = 8'h5;
assign n0281 = ( RD_ROM_0 == n0280 );
assign n0282 = 8'h6;
assign n0283 = ( RD_ROM_0 == n0282 );
assign n0284 = 8'h7;
assign n0285 = ( RD_ROM_0 == n0284 );
assign n0286 = 8'h8;
assign n0287 = ( RD_ROM_0 == n0286 );
assign n0288 = 8'h9;
assign n0289 = ( RD_ROM_0 == n0288 );
assign n0290 = 8'ha;
assign n0291 = ( RD_ROM_0 == n0290 );
assign n0292 = 8'hb;
assign n0293 = ( RD_ROM_0 == n0292 );
assign n0294 = 8'hc;
assign n0295 = ( RD_ROM_0 == n0294 );
assign n0296 = 8'hd;
assign n0297 = ( RD_ROM_0 == n0296 );
assign n0298 = 8'he;
assign n0299 = ( RD_ROM_0 == n0298 );
assign n0300 = 8'hf;
assign n0301 = ( RD_ROM_0 == n0300 );
assign n0302 = 8'h10;
assign n0303 = ( RD_ROM_0 == n0302 );
assign n0304 = 8'h11;
assign n0305 = ( RD_ROM_0 == n0304 );
assign n0306 = 8'h12;
assign n0307 = ( RD_ROM_0 == n0306 );
assign n0308 = 8'h15;
assign n0309 = ( RD_ROM_0 == n0308 );
assign n0310 = 8'h16;
assign n0311 = ( RD_ROM_0 == n0310 );
assign n0312 = 8'h17;
assign n0313 = ( RD_ROM_0 == n0312 );
assign n0314 = 8'h18;
assign n0315 = ( RD_ROM_0 == n0314 );
assign n0316 = 8'h19;
assign n0317 = ( RD_ROM_0 == n0316 );
assign n0318 = 8'h1a;
assign n0319 = ( RD_ROM_0 == n0318 );
assign n0320 = 8'h1b;
assign n0321 = ( RD_ROM_0 == n0320 );
assign n0322 = 8'h1c;
assign n0323 = ( RD_ROM_0 == n0322 );
assign n0324 = 8'h1d;
assign n0325 = ( RD_ROM_0 == n0324 );
assign n0326 = 8'h1e;
assign n0327 = ( RD_ROM_0 == n0326 );
assign n0328 = 8'h1f;
assign n0329 = ( RD_ROM_0 == n0328 );
assign n0330 = 8'h31;
assign n0331 = ( RD_ROM_0 == n0330 );
assign n0332 = 8'h42;
assign n0333 = ( RD_ROM_0 == n0332 );
assign n0334 = 8'h43;
assign n0335 = ( RD_ROM_0 == n0334 );
assign n0336 = 8'h51;
assign n0337 = ( RD_ROM_0 == n0336 );
assign n0338 = 8'h52;
assign n0339 = ( RD_ROM_0 == n0338 );
assign n0340 = 8'h53;
assign n0341 = ( RD_ROM_0 == n0340 );
assign n0342 = 8'h62;
assign n0343 = ( RD_ROM_0 == n0342 );
assign n0344 = 8'h63;
assign n0345 = ( RD_ROM_0 == n0344 );
assign n0346 = 8'h71;
assign n0347 = ( RD_ROM_0 == n0346 );
assign n0348 = 8'h75;
assign n0349 = ( RD_ROM_0 == n0348 );
assign n0350 = 8'h76;
assign n0351 = ( RD_ROM_0 == n0350 );
assign n0352 = 8'h77;
assign n0353 = ( RD_ROM_0 == n0352 );
assign n0354 = 8'h78;
assign n0355 = ( RD_ROM_0 == n0354 );
assign n0356 = 8'h79;
assign n0357 = ( RD_ROM_0 == n0356 );
assign n0358 = 8'h7a;
assign n0359 = ( RD_ROM_0 == n0358 );
assign n0360 = 8'h7b;
assign n0361 = ( RD_ROM_0 == n0360 );
assign n0362 = 8'h7c;
assign n0363 = ( RD_ROM_0 == n0362 );
assign n0364 = 8'h7d;
assign n0365 = ( RD_ROM_0 == n0364 );
assign n0366 = 8'h7e;
assign n0367 = ( RD_ROM_0 == n0366 );
assign n0368 = 8'h7f;
assign n0369 = ( RD_ROM_0 == n0368 );
assign n0370 = 8'h85;
assign n0371 = ( RD_ROM_0 == n0370 );
assign n0372 = 8'h86;
assign n0373 = ( RD_ROM_0 == n0372 );
assign n0374 = ( RD_ROM_0 == n0025 );
assign n0375 = ( RD_ROM_0 == n0027 );
assign n0376 = ( RD_ROM_0 == n0029 );
assign n0377 = ( RD_ROM_0 == n0031 );
assign n0378 = ( RD_ROM_0 == n0035 );
assign n0379 = ( RD_ROM_0 == n0033 );
assign n0380 = ( RD_ROM_0 == n0037 );
assign n0381 = 8'h8e;
assign n0382 = ( RD_ROM_0 == n0381 );
assign n0383 = 8'h8f;
assign n0384 = ( RD_ROM_0 == n0383 );
assign n0385 = 8'h91;
assign n0386 = ( RD_ROM_0 == n0385 );
assign n0387 = 8'h92;
assign n0388 = ( RD_ROM_0 == n0387 );
assign n0389 = 8'ha6;
assign n0390 = ( RD_ROM_0 == n0389 );
assign n0391 = 8'ha7;
assign n0392 = ( RD_ROM_0 == n0391 );
assign n0393 = ( RD_ROM_0 == n0047 );
assign n0394 = 8'ha9;
assign n0395 = ( RD_ROM_0 == n0394 );
assign n0396 = 8'haa;
assign n0397 = ( RD_ROM_0 == n0396 );
assign n0398 = 8'hab;
assign n0399 = ( RD_ROM_0 == n0398 );
assign n0400 = 8'hac;
assign n0401 = ( RD_ROM_0 == n0400 );
assign n0402 = 8'had;
assign n0403 = ( RD_ROM_0 == n0402 );
assign n0404 = 8'hae;
assign n0405 = ( RD_ROM_0 == n0404 );
assign n0406 = 8'haf;
assign n0407 = ( RD_ROM_0 == n0406 );
assign n0408 = 8'hb1;
assign n0409 = ( RD_ROM_0 == n0408 );
assign n0410 = 8'hb2;
assign n0411 = ( RD_ROM_0 == n0410 );
assign n0412 = 8'hc0;
assign n0413 = ( RD_ROM_0 == n0412 );
assign n0414 = 8'hc2;
assign n0415 = ( RD_ROM_0 == n0414 );
assign n0416 = 8'hc5;
assign n0417 = ( RD_ROM_0 == n0416 );
assign n0418 = 8'hc6;
assign n0419 = ( RD_ROM_0 == n0418 );
assign n0420 = 8'hc7;
assign n0421 = ( RD_ROM_0 == n0420 );
assign n0422 = 8'hc8;
assign n0423 = ( RD_ROM_0 == n0422 );
assign n0424 = 8'hc9;
assign n0425 = ( RD_ROM_0 == n0424 );
assign n0426 = 8'hca;
assign n0427 = ( RD_ROM_0 == n0426 );
assign n0428 = 8'hcb;
assign n0429 = ( RD_ROM_0 == n0428 );
assign n0430 = 8'hcc;
assign n0431 = ( RD_ROM_0 == n0430 );
assign n0432 = 8'hcd;
assign n0433 = ( RD_ROM_0 == n0432 );
assign n0434 = 8'hce;
assign n0435 = ( RD_ROM_0 == n0434 );
assign n0436 = 8'hcf;
assign n0437 = ( RD_ROM_0 == n0436 );
assign n0438 = ( RD_ROM_0 == n0053 );
assign n0439 = 8'hd1;
assign n0440 = ( RD_ROM_0 == n0439 );
assign n0441 = 8'hd2;
assign n0442 = ( RD_ROM_0 == n0441 );
assign n0443 = 8'hd5;
assign n0444 = ( RD_ROM_0 == n0443 );
assign n0445 = 8'hd6;
assign n0446 = ( RD_ROM_0 == n0445 );
assign n0447 = 8'hd7;
assign n0448 = ( RD_ROM_0 == n0447 );
assign n0449 = 8'hd8;
assign n0450 = ( RD_ROM_0 == n0449 );
assign n0451 = 8'hd9;
assign n0452 = ( RD_ROM_0 == n0451 );
assign n0453 = 8'hda;
assign n0454 = ( RD_ROM_0 == n0453 );
assign n0455 = 8'hdb;
assign n0456 = ( RD_ROM_0 == n0455 );
assign n0457 = 8'hdc;
assign n0458 = ( RD_ROM_0 == n0457 );
assign n0459 = 8'hdd;
assign n0460 = ( RD_ROM_0 == n0459 );
assign n0461 = 8'hde;
assign n0462 = ( RD_ROM_0 == n0461 );
assign n0463 = 8'hdf;
assign n0464 = ( RD_ROM_0 == n0463 );
assign n0465 = 8'hf1;
assign n0466 = ( RD_ROM_0 == n0465 );
assign n0467 = 8'hf5;
assign n0468 = ( RD_ROM_0 == n0467 );
assign n0469 = 8'hf6;
assign n0470 = ( RD_ROM_0 == n0469 );
assign n0471 = 8'hf7;
assign n0472 = ( RD_ROM_0 == n0471 );
assign n0473 = 8'hf8;
assign n0474 = ( RD_ROM_0 == n0473 );
assign n0475 = 8'hf9;
assign n0476 = ( RD_ROM_0 == n0475 );
assign n0477 = 8'hfa;
assign n0478 = ( RD_ROM_0 == n0477 );
assign n0479 = 8'hfb;
assign n0480 = ( RD_ROM_0 == n0479 );
assign n0481 = 8'hfc;
assign n0482 = ( RD_ROM_0 == n0481 );
assign n0483 = 8'hfd;
assign n0484 = ( RD_ROM_0 == n0483 );
assign n0485 = 8'hfe;
assign n0486 = ( RD_ROM_0 == n0485 );
assign n0487 = 8'hff;
assign n0488 = ( RD_ROM_0 == n0487 );
assign WR_ADDR_0_IRAM = WR_ADDR_ABSTR_IRAM_0;
assign WR_DATA_0_IRAM = WR_DATA_ABSTR_IRAM_0;
assign WR_COND_0_IRAM = ((WR_COND_ABSTR_IRAM_0 && !(n0002)));
assign WR_ADDR_1_IRAM = WR_ADDR_ABSTR_IRAM_1;
assign WR_DATA_1_IRAM = WR_DATA_ABSTR_IRAM_1;
assign WR_COND_1_IRAM = ((WR_COND_ABSTR_IRAM_1 && !(n0002)));
assign IRAM_full = {IRAM[15], IRAM[14], IRAM[13], IRAM[12], IRAM[11], IRAM[10], IRAM[9], IRAM[8], IRAM[7], IRAM[6], IRAM[5], IRAM[4], IRAM[3], IRAM[2], IRAM[1], IRAM[0]} ;
assign SBUF_next = SBUF;
assign SCON_next = SCON;
assign PCON_next = PCON;
assign TCON_next = TCON;
assign TL0_next = TL0;
assign TL1_next = TL1;
assign TH0_next = TH0;
assign TH1_next = TH1;
assign TMOD_next = TMOD;
assign IE_next = IE;
assign IP_next = IP;

always @(posedge clk) begin
  if (rst) begin
    ACC <= 8'h0;
    B <= 8'h0;
    DPH <= 8'h0;
    DPL <= 8'h0;
    IE <= 8'h0;
    IP <= 8'h0;
    P0 <= 8'hff;
    P0INREG <= 8'h0;
    P1 <= 8'hff;
    P1INREG <= 8'h0;
    P2 <= 8'hff;
    P2INREG <= 8'h0;
    P3 <= 8'hff;
    P3INREG <= 8'h0;
    PC <= 16'h0;
    PCON <= 8'h0;
    PSW <= 8'h0;
    SBUF <= 8'h0;
    SCON <= 8'h0;
    SP <= 8'h7;
    TCON <= 8'h0;
    TH0 <= 8'h0;
    TH1 <= 8'h0;
    TL0 <= 8'h0;
    TL1 <= 8'h0;
    TMOD <= 8'h0;
`ifdef OC8051_SIMULATION
    IRAM[0] = 8'b0;
    IRAM[1] = 8'b0;
    IRAM[2] = 8'b0;
    IRAM[3] = 8'b0;
    IRAM[4] = 8'b0;
    IRAM[5] = 8'b0;
    IRAM[6] = 8'b0;
    IRAM[7] = 8'b0;
    IRAM[8] = 8'b0;
    IRAM[9] = 8'b0;
    IRAM[10] = 8'b0;
    IRAM[11] = 8'b0;
    IRAM[12] = 8'b0;
    IRAM[13] = 8'b0;
    IRAM[14] = 8'b0;
    IRAM[15] = 8'b0;
`endif
`ifdef OC8051_SIMULATION
    XRAM[0] = 8'b0;
    XRAM[1] = 8'b0;
    XRAM[2] = 8'b0;
    XRAM[3] = 8'b0;
    XRAM[4] = 8'b0;
    XRAM[5] = 8'b0;
    XRAM[6] = 8'b0;
    XRAM[7] = 8'b0;
    XRAM[8] = 8'b0;
    XRAM[9] = 8'b0;
    XRAM[10] = 8'b0;
    XRAM[11] = 8'b0;
    XRAM[12] = 8'b0;
    XRAM[13] = 8'b0;
    XRAM[14] = 8'b0;
    XRAM[15] = 8'b0;
    XRAM[16] = 8'b0;
    XRAM[17] = 8'b0;
    XRAM[18] = 8'b0;
    XRAM[19] = 8'b0;
    XRAM[20] = 8'b0;
    XRAM[21] = 8'b0;
    XRAM[22] = 8'b0;
    XRAM[23] = 8'b0;
    XRAM[24] = 8'b0;
    XRAM[25] = 8'b0;
    XRAM[26] = 8'b0;
    XRAM[27] = 8'b0;
    XRAM[28] = 8'b0;
    XRAM[29] = 8'b0;
    XRAM[30] = 8'b0;
    XRAM[31] = 8'b0;
    XRAM[32] = 8'b0;
    XRAM[33] = 8'b0;
    XRAM[34] = 8'b0;
    XRAM[35] = 8'b0;
    XRAM[36] = 8'b0;
    XRAM[37] = 8'b0;
    XRAM[38] = 8'b0;
    XRAM[39] = 8'b0;
    XRAM[40] = 8'b0;
    XRAM[41] = 8'b0;
    XRAM[42] = 8'b0;
    XRAM[43] = 8'b0;
    XRAM[44] = 8'b0;
    XRAM[45] = 8'b0;
    XRAM[46] = 8'b0;
    XRAM[47] = 8'b0;
    XRAM[48] = 8'b0;
    XRAM[49] = 8'b0;
    XRAM[50] = 8'b0;
    XRAM[51] = 8'b0;
    XRAM[52] = 8'b0;
    XRAM[53] = 8'b0;
    XRAM[54] = 8'b0;
    XRAM[55] = 8'b0;
    XRAM[56] = 8'b0;
    XRAM[57] = 8'b0;
    XRAM[58] = 8'b0;
    XRAM[59] = 8'b0;
    XRAM[60] = 8'b0;
    XRAM[61] = 8'b0;
    XRAM[62] = 8'b0;
    XRAM[63] = 8'b0;
    XRAM[64] = 8'b0;
    XRAM[65] = 8'b0;
    XRAM[66] = 8'b0;
    XRAM[67] = 8'b0;
    XRAM[68] = 8'b0;
    XRAM[69] = 8'b0;
    XRAM[70] = 8'b0;
    XRAM[71] = 8'b0;
    XRAM[72] = 8'b0;
    XRAM[73] = 8'b0;
    XRAM[74] = 8'b0;
    XRAM[75] = 8'b0;
    XRAM[76] = 8'b0;
    XRAM[77] = 8'b0;
    XRAM[78] = 8'b0;
    XRAM[79] = 8'b0;
    XRAM[80] = 8'b0;
    XRAM[81] = 8'b0;
    XRAM[82] = 8'b0;
    XRAM[83] = 8'b0;
    XRAM[84] = 8'b0;
    XRAM[85] = 8'b0;
    XRAM[86] = 8'b0;
    XRAM[87] = 8'b0;
    XRAM[88] = 8'b0;
    XRAM[89] = 8'b0;
    XRAM[90] = 8'b0;
    XRAM[91] = 8'b0;
    XRAM[92] = 8'b0;
    XRAM[93] = 8'b0;
    XRAM[94] = 8'b0;
    XRAM[95] = 8'b0;
    XRAM[96] = 8'b0;
    XRAM[97] = 8'b0;
    XRAM[98] = 8'b0;
    XRAM[99] = 8'b0;
    XRAM[100] = 8'b0;
    XRAM[101] = 8'b0;
    XRAM[102] = 8'b0;
    XRAM[103] = 8'b0;
    XRAM[104] = 8'b0;
    XRAM[105] = 8'b0;
    XRAM[106] = 8'b0;
    XRAM[107] = 8'b0;
    XRAM[108] = 8'b0;
    XRAM[109] = 8'b0;
    XRAM[110] = 8'b0;
    XRAM[111] = 8'b0;
    XRAM[112] = 8'b0;
    XRAM[113] = 8'b0;
    XRAM[114] = 8'b0;
    XRAM[115] = 8'b0;
    XRAM[116] = 8'b0;
    XRAM[117] = 8'b0;
    XRAM[118] = 8'b0;
    XRAM[119] = 8'b0;
    XRAM[120] = 8'b0;
    XRAM[121] = 8'b0;
    XRAM[122] = 8'b0;
    XRAM[123] = 8'b0;
    XRAM[124] = 8'b0;
    XRAM[125] = 8'b0;
    XRAM[126] = 8'b0;
    XRAM[127] = 8'b0;
    XRAM[128] = 8'b0;
    XRAM[129] = 8'b0;
    XRAM[130] = 8'b0;
    XRAM[131] = 8'b0;
    XRAM[132] = 8'b0;
    XRAM[133] = 8'b0;
    XRAM[134] = 8'b0;
    XRAM[135] = 8'b0;
    XRAM[136] = 8'b0;
    XRAM[137] = 8'b0;
    XRAM[138] = 8'b0;
    XRAM[139] = 8'b0;
    XRAM[140] = 8'b0;
    XRAM[141] = 8'b0;
    XRAM[142] = 8'b0;
    XRAM[143] = 8'b0;
    XRAM[144] = 8'b0;
    XRAM[145] = 8'b0;
    XRAM[146] = 8'b0;
    XRAM[147] = 8'b0;
    XRAM[148] = 8'b0;
    XRAM[149] = 8'b0;
    XRAM[150] = 8'b0;
    XRAM[151] = 8'b0;
    XRAM[152] = 8'b0;
    XRAM[153] = 8'b0;
    XRAM[154] = 8'b0;
    XRAM[155] = 8'b0;
    XRAM[156] = 8'b0;
    XRAM[157] = 8'b0;
    XRAM[158] = 8'b0;
    XRAM[159] = 8'b0;
    XRAM[160] = 8'b0;
    XRAM[161] = 8'b0;
    XRAM[162] = 8'b0;
    XRAM[163] = 8'b0;
    XRAM[164] = 8'b0;
    XRAM[165] = 8'b0;
    XRAM[166] = 8'b0;
    XRAM[167] = 8'b0;
    XRAM[168] = 8'b0;
    XRAM[169] = 8'b0;
    XRAM[170] = 8'b0;
    XRAM[171] = 8'b0;
    XRAM[172] = 8'b0;
    XRAM[173] = 8'b0;
    XRAM[174] = 8'b0;
    XRAM[175] = 8'b0;
    XRAM[176] = 8'b0;
    XRAM[177] = 8'b0;
    XRAM[178] = 8'b0;
    XRAM[179] = 8'b0;
    XRAM[180] = 8'b0;
    XRAM[181] = 8'b0;
    XRAM[182] = 8'b0;
    XRAM[183] = 8'b0;
    XRAM[184] = 8'b0;
    XRAM[185] = 8'b0;
    XRAM[186] = 8'b0;
    XRAM[187] = 8'b0;
    XRAM[188] = 8'b0;
    XRAM[189] = 8'b0;
    XRAM[190] = 8'b0;
    XRAM[191] = 8'b0;
    XRAM[192] = 8'b0;
    XRAM[193] = 8'b0;
    XRAM[194] = 8'b0;
    XRAM[195] = 8'b0;
    XRAM[196] = 8'b0;
    XRAM[197] = 8'b0;
    XRAM[198] = 8'b0;
    XRAM[199] = 8'b0;
    XRAM[200] = 8'b0;
    XRAM[201] = 8'b0;
    XRAM[202] = 8'b0;
    XRAM[203] = 8'b0;
    XRAM[204] = 8'b0;
    XRAM[205] = 8'b0;
    XRAM[206] = 8'b0;
    XRAM[207] = 8'b0;
    XRAM[208] = 8'b0;
    XRAM[209] = 8'b0;
    XRAM[210] = 8'b0;
    XRAM[211] = 8'b0;
    XRAM[212] = 8'b0;
    XRAM[213] = 8'b0;
    XRAM[214] = 8'b0;
    XRAM[215] = 8'b0;
    XRAM[216] = 8'b0;
    XRAM[217] = 8'b0;
    XRAM[218] = 8'b0;
    XRAM[219] = 8'b0;
    XRAM[220] = 8'b0;
    XRAM[221] = 8'b0;
    XRAM[222] = 8'b0;
    XRAM[223] = 8'b0;
    XRAM[224] = 8'b0;
    XRAM[225] = 8'b0;
    XRAM[226] = 8'b0;
    XRAM[227] = 8'b0;
    XRAM[228] = 8'b0;
    XRAM[229] = 8'b0;
    XRAM[230] = 8'b0;
    XRAM[231] = 8'b0;
    XRAM[232] = 8'b0;
    XRAM[233] = 8'b0;
    XRAM[234] = 8'b0;
    XRAM[235] = 8'b0;
    XRAM[236] = 8'b0;
    XRAM[237] = 8'b0;
    XRAM[238] = 8'b0;
    XRAM[239] = 8'b0;
    XRAM[240] = 8'b0;
    XRAM[241] = 8'b0;
    XRAM[242] = 8'b0;
    XRAM[243] = 8'b0;
    XRAM[244] = 8'b0;
    XRAM[245] = 8'b0;
    XRAM[246] = 8'b0;
    XRAM[247] = 8'b0;
    XRAM[248] = 8'b0;
    XRAM[249] = 8'b0;
    XRAM[250] = 8'b0;
    XRAM[251] = 8'b0;
    XRAM[252] = 8'b0;
    XRAM[253] = 8'b0;
    XRAM[254] = 8'b0;
    XRAM[255] = 8'b0;
    XRAM[256] = 8'b0;
    XRAM[257] = 8'b0;
    XRAM[258] = 8'b0;
    XRAM[259] = 8'b0;
    XRAM[260] = 8'b0;
    XRAM[261] = 8'b0;
    XRAM[262] = 8'b0;
    XRAM[263] = 8'b0;
    XRAM[264] = 8'b0;
    XRAM[265] = 8'b0;
    XRAM[266] = 8'b0;
    XRAM[267] = 8'b0;
    XRAM[268] = 8'b0;
    XRAM[269] = 8'b0;
    XRAM[270] = 8'b0;
    XRAM[271] = 8'b0;
    XRAM[272] = 8'b0;
    XRAM[273] = 8'b0;
    XRAM[274] = 8'b0;
    XRAM[275] = 8'b0;
    XRAM[276] = 8'b0;
    XRAM[277] = 8'b0;
    XRAM[278] = 8'b0;
    XRAM[279] = 8'b0;
    XRAM[280] = 8'b0;
    XRAM[281] = 8'b0;
    XRAM[282] = 8'b0;
    XRAM[283] = 8'b0;
    XRAM[284] = 8'b0;
    XRAM[285] = 8'b0;
    XRAM[286] = 8'b0;
    XRAM[287] = 8'b0;
    XRAM[288] = 8'b0;
    XRAM[289] = 8'b0;
    XRAM[290] = 8'b0;
    XRAM[291] = 8'b0;
    XRAM[292] = 8'b0;
    XRAM[293] = 8'b0;
    XRAM[294] = 8'b0;
    XRAM[295] = 8'b0;
    XRAM[296] = 8'b0;
    XRAM[297] = 8'b0;
    XRAM[298] = 8'b0;
    XRAM[299] = 8'b0;
    XRAM[300] = 8'b0;
    XRAM[301] = 8'b0;
    XRAM[302] = 8'b0;
    XRAM[303] = 8'b0;
    XRAM[304] = 8'b0;
    XRAM[305] = 8'b0;
    XRAM[306] = 8'b0;
    XRAM[307] = 8'b0;
    XRAM[308] = 8'b0;
    XRAM[309] = 8'b0;
    XRAM[310] = 8'b0;
    XRAM[311] = 8'b0;
    XRAM[312] = 8'b0;
    XRAM[313] = 8'b0;
    XRAM[314] = 8'b0;
    XRAM[315] = 8'b0;
    XRAM[316] = 8'b0;
    XRAM[317] = 8'b0;
    XRAM[318] = 8'b0;
    XRAM[319] = 8'b0;
    XRAM[320] = 8'b0;
    XRAM[321] = 8'b0;
    XRAM[322] = 8'b0;
    XRAM[323] = 8'b0;
    XRAM[324] = 8'b0;
    XRAM[325] = 8'b0;
    XRAM[326] = 8'b0;
    XRAM[327] = 8'b0;
    XRAM[328] = 8'b0;
    XRAM[329] = 8'b0;
    XRAM[330] = 8'b0;
    XRAM[331] = 8'b0;
    XRAM[332] = 8'b0;
    XRAM[333] = 8'b0;
    XRAM[334] = 8'b0;
    XRAM[335] = 8'b0;
    XRAM[336] = 8'b0;
    XRAM[337] = 8'b0;
    XRAM[338] = 8'b0;
    XRAM[339] = 8'b0;
    XRAM[340] = 8'b0;
    XRAM[341] = 8'b0;
    XRAM[342] = 8'b0;
    XRAM[343] = 8'b0;
    XRAM[344] = 8'b0;
    XRAM[345] = 8'b0;
    XRAM[346] = 8'b0;
    XRAM[347] = 8'b0;
    XRAM[348] = 8'b0;
    XRAM[349] = 8'b0;
    XRAM[350] = 8'b0;
    XRAM[351] = 8'b0;
    XRAM[352] = 8'b0;
    XRAM[353] = 8'b0;
    XRAM[354] = 8'b0;
    XRAM[355] = 8'b0;
    XRAM[356] = 8'b0;
    XRAM[357] = 8'b0;
    XRAM[358] = 8'b0;
    XRAM[359] = 8'b0;
    XRAM[360] = 8'b0;
    XRAM[361] = 8'b0;
    XRAM[362] = 8'b0;
    XRAM[363] = 8'b0;
    XRAM[364] = 8'b0;
    XRAM[365] = 8'b0;
    XRAM[366] = 8'b0;
    XRAM[367] = 8'b0;
    XRAM[368] = 8'b0;
    XRAM[369] = 8'b0;
    XRAM[370] = 8'b0;
    XRAM[371] = 8'b0;
    XRAM[372] = 8'b0;
    XRAM[373] = 8'b0;
    XRAM[374] = 8'b0;
    XRAM[375] = 8'b0;
    XRAM[376] = 8'b0;
    XRAM[377] = 8'b0;
    XRAM[378] = 8'b0;
    XRAM[379] = 8'b0;
    XRAM[380] = 8'b0;
    XRAM[381] = 8'b0;
    XRAM[382] = 8'b0;
    XRAM[383] = 8'b0;
    XRAM[384] = 8'b0;
    XRAM[385] = 8'b0;
    XRAM[386] = 8'b0;
    XRAM[387] = 8'b0;
    XRAM[388] = 8'b0;
    XRAM[389] = 8'b0;
    XRAM[390] = 8'b0;
    XRAM[391] = 8'b0;
    XRAM[392] = 8'b0;
    XRAM[393] = 8'b0;
    XRAM[394] = 8'b0;
    XRAM[395] = 8'b0;
    XRAM[396] = 8'b0;
    XRAM[397] = 8'b0;
    XRAM[398] = 8'b0;
    XRAM[399] = 8'b0;
    XRAM[400] = 8'b0;
    XRAM[401] = 8'b0;
    XRAM[402] = 8'b0;
    XRAM[403] = 8'b0;
    XRAM[404] = 8'b0;
    XRAM[405] = 8'b0;
    XRAM[406] = 8'b0;
    XRAM[407] = 8'b0;
    XRAM[408] = 8'b0;
    XRAM[409] = 8'b0;
    XRAM[410] = 8'b0;
    XRAM[411] = 8'b0;
    XRAM[412] = 8'b0;
    XRAM[413] = 8'b0;
    XRAM[414] = 8'b0;
    XRAM[415] = 8'b0;
    XRAM[416] = 8'b0;
    XRAM[417] = 8'b0;
    XRAM[418] = 8'b0;
    XRAM[419] = 8'b0;
    XRAM[420] = 8'b0;
    XRAM[421] = 8'b0;
    XRAM[422] = 8'b0;
    XRAM[423] = 8'b0;
    XRAM[424] = 8'b0;
    XRAM[425] = 8'b0;
    XRAM[426] = 8'b0;
    XRAM[427] = 8'b0;
    XRAM[428] = 8'b0;
    XRAM[429] = 8'b0;
    XRAM[430] = 8'b0;
    XRAM[431] = 8'b0;
    XRAM[432] = 8'b0;
    XRAM[433] = 8'b0;
    XRAM[434] = 8'b0;
    XRAM[435] = 8'b0;
    XRAM[436] = 8'b0;
    XRAM[437] = 8'b0;
    XRAM[438] = 8'b0;
    XRAM[439] = 8'b0;
    XRAM[440] = 8'b0;
    XRAM[441] = 8'b0;
    XRAM[442] = 8'b0;
    XRAM[443] = 8'b0;
    XRAM[444] = 8'b0;
    XRAM[445] = 8'b0;
    XRAM[446] = 8'b0;
    XRAM[447] = 8'b0;
    XRAM[448] = 8'b0;
    XRAM[449] = 8'b0;
    XRAM[450] = 8'b0;
    XRAM[451] = 8'b0;
    XRAM[452] = 8'b0;
    XRAM[453] = 8'b0;
    XRAM[454] = 8'b0;
    XRAM[455] = 8'b0;
    XRAM[456] = 8'b0;
    XRAM[457] = 8'b0;
    XRAM[458] = 8'b0;
    XRAM[459] = 8'b0;
    XRAM[460] = 8'b0;
    XRAM[461] = 8'b0;
    XRAM[462] = 8'b0;
    XRAM[463] = 8'b0;
    XRAM[464] = 8'b0;
    XRAM[465] = 8'b0;
    XRAM[466] = 8'b0;
    XRAM[467] = 8'b0;
    XRAM[468] = 8'b0;
    XRAM[469] = 8'b0;
    XRAM[470] = 8'b0;
    XRAM[471] = 8'b0;
    XRAM[472] = 8'b0;
    XRAM[473] = 8'b0;
    XRAM[474] = 8'b0;
    XRAM[475] = 8'b0;
    XRAM[476] = 8'b0;
    XRAM[477] = 8'b0;
    XRAM[478] = 8'b0;
    XRAM[479] = 8'b0;
    XRAM[480] = 8'b0;
    XRAM[481] = 8'b0;
    XRAM[482] = 8'b0;
    XRAM[483] = 8'b0;
    XRAM[484] = 8'b0;
    XRAM[485] = 8'b0;
    XRAM[486] = 8'b0;
    XRAM[487] = 8'b0;
    XRAM[488] = 8'b0;
    XRAM[489] = 8'b0;
    XRAM[490] = 8'b0;
    XRAM[491] = 8'b0;
    XRAM[492] = 8'b0;
    XRAM[493] = 8'b0;
    XRAM[494] = 8'b0;
    XRAM[495] = 8'b0;
    XRAM[496] = 8'b0;
    XRAM[497] = 8'b0;
    XRAM[498] = 8'b0;
    XRAM[499] = 8'b0;
    XRAM[500] = 8'b0;
    XRAM[501] = 8'b0;
    XRAM[502] = 8'b0;
    XRAM[503] = 8'b0;
    XRAM[504] = 8'b0;
    XRAM[505] = 8'b0;
    XRAM[506] = 8'b0;
    XRAM[507] = 8'b0;
    XRAM[508] = 8'b0;
    XRAM[509] = 8'b0;
    XRAM[510] = 8'b0;
    XRAM[511] = 8'b0;
    XRAM[512] = 8'b0;
    XRAM[513] = 8'b0;
    XRAM[514] = 8'b0;
    XRAM[515] = 8'b0;
    XRAM[516] = 8'b0;
    XRAM[517] = 8'b0;
    XRAM[518] = 8'b0;
    XRAM[519] = 8'b0;
    XRAM[520] = 8'b0;
    XRAM[521] = 8'b0;
    XRAM[522] = 8'b0;
    XRAM[523] = 8'b0;
    XRAM[524] = 8'b0;
    XRAM[525] = 8'b0;
    XRAM[526] = 8'b0;
    XRAM[527] = 8'b0;
    XRAM[528] = 8'b0;
    XRAM[529] = 8'b0;
    XRAM[530] = 8'b0;
    XRAM[531] = 8'b0;
    XRAM[532] = 8'b0;
    XRAM[533] = 8'b0;
    XRAM[534] = 8'b0;
    XRAM[535] = 8'b0;
    XRAM[536] = 8'b0;
    XRAM[537] = 8'b0;
    XRAM[538] = 8'b0;
    XRAM[539] = 8'b0;
    XRAM[540] = 8'b0;
    XRAM[541] = 8'b0;
    XRAM[542] = 8'b0;
    XRAM[543] = 8'b0;
    XRAM[544] = 8'b0;
    XRAM[545] = 8'b0;
    XRAM[546] = 8'b0;
    XRAM[547] = 8'b0;
    XRAM[548] = 8'b0;
    XRAM[549] = 8'b0;
    XRAM[550] = 8'b0;
    XRAM[551] = 8'b0;
    XRAM[552] = 8'b0;
    XRAM[553] = 8'b0;
    XRAM[554] = 8'b0;
    XRAM[555] = 8'b0;
    XRAM[556] = 8'b0;
    XRAM[557] = 8'b0;
    XRAM[558] = 8'b0;
    XRAM[559] = 8'b0;
    XRAM[560] = 8'b0;
    XRAM[561] = 8'b0;
    XRAM[562] = 8'b0;
    XRAM[563] = 8'b0;
    XRAM[564] = 8'b0;
    XRAM[565] = 8'b0;
    XRAM[566] = 8'b0;
    XRAM[567] = 8'b0;
    XRAM[568] = 8'b0;
    XRAM[569] = 8'b0;
    XRAM[570] = 8'b0;
    XRAM[571] = 8'b0;
    XRAM[572] = 8'b0;
    XRAM[573] = 8'b0;
    XRAM[574] = 8'b0;
    XRAM[575] = 8'b0;
    XRAM[576] = 8'b0;
    XRAM[577] = 8'b0;
    XRAM[578] = 8'b0;
    XRAM[579] = 8'b0;
    XRAM[580] = 8'b0;
    XRAM[581] = 8'b0;
    XRAM[582] = 8'b0;
    XRAM[583] = 8'b0;
    XRAM[584] = 8'b0;
    XRAM[585] = 8'b0;
    XRAM[586] = 8'b0;
    XRAM[587] = 8'b0;
    XRAM[588] = 8'b0;
    XRAM[589] = 8'b0;
    XRAM[590] = 8'b0;
    XRAM[591] = 8'b0;
    XRAM[592] = 8'b0;
    XRAM[593] = 8'b0;
    XRAM[594] = 8'b0;
    XRAM[595] = 8'b0;
    XRAM[596] = 8'b0;
    XRAM[597] = 8'b0;
    XRAM[598] = 8'b0;
    XRAM[599] = 8'b0;
    XRAM[600] = 8'b0;
    XRAM[601] = 8'b0;
    XRAM[602] = 8'b0;
    XRAM[603] = 8'b0;
    XRAM[604] = 8'b0;
    XRAM[605] = 8'b0;
    XRAM[606] = 8'b0;
    XRAM[607] = 8'b0;
    XRAM[608] = 8'b0;
    XRAM[609] = 8'b0;
    XRAM[610] = 8'b0;
    XRAM[611] = 8'b0;
    XRAM[612] = 8'b0;
    XRAM[613] = 8'b0;
    XRAM[614] = 8'b0;
    XRAM[615] = 8'b0;
    XRAM[616] = 8'b0;
    XRAM[617] = 8'b0;
    XRAM[618] = 8'b0;
    XRAM[619] = 8'b0;
    XRAM[620] = 8'b0;
    XRAM[621] = 8'b0;
    XRAM[622] = 8'b0;
    XRAM[623] = 8'b0;
    XRAM[624] = 8'b0;
    XRAM[625] = 8'b0;
    XRAM[626] = 8'b0;
    XRAM[627] = 8'b0;
    XRAM[628] = 8'b0;
    XRAM[629] = 8'b0;
    XRAM[630] = 8'b0;
    XRAM[631] = 8'b0;
    XRAM[632] = 8'b0;
    XRAM[633] = 8'b0;
    XRAM[634] = 8'b0;
    XRAM[635] = 8'b0;
    XRAM[636] = 8'b0;
    XRAM[637] = 8'b0;
    XRAM[638] = 8'b0;
    XRAM[639] = 8'b0;
    XRAM[640] = 8'b0;
    XRAM[641] = 8'b0;
    XRAM[642] = 8'b0;
    XRAM[643] = 8'b0;
    XRAM[644] = 8'b0;
    XRAM[645] = 8'b0;
    XRAM[646] = 8'b0;
    XRAM[647] = 8'b0;
    XRAM[648] = 8'b0;
    XRAM[649] = 8'b0;
    XRAM[650] = 8'b0;
    XRAM[651] = 8'b0;
    XRAM[652] = 8'b0;
    XRAM[653] = 8'b0;
    XRAM[654] = 8'b0;
    XRAM[655] = 8'b0;
    XRAM[656] = 8'b0;
    XRAM[657] = 8'b0;
    XRAM[658] = 8'b0;
    XRAM[659] = 8'b0;
    XRAM[660] = 8'b0;
    XRAM[661] = 8'b0;
    XRAM[662] = 8'b0;
    XRAM[663] = 8'b0;
    XRAM[664] = 8'b0;
    XRAM[665] = 8'b0;
    XRAM[666] = 8'b0;
    XRAM[667] = 8'b0;
    XRAM[668] = 8'b0;
    XRAM[669] = 8'b0;
    XRAM[670] = 8'b0;
    XRAM[671] = 8'b0;
    XRAM[672] = 8'b0;
    XRAM[673] = 8'b0;
    XRAM[674] = 8'b0;
    XRAM[675] = 8'b0;
    XRAM[676] = 8'b0;
    XRAM[677] = 8'b0;
    XRAM[678] = 8'b0;
    XRAM[679] = 8'b0;
    XRAM[680] = 8'b0;
    XRAM[681] = 8'b0;
    XRAM[682] = 8'b0;
    XRAM[683] = 8'b0;
    XRAM[684] = 8'b0;
    XRAM[685] = 8'b0;
    XRAM[686] = 8'b0;
    XRAM[687] = 8'b0;
    XRAM[688] = 8'b0;
    XRAM[689] = 8'b0;
    XRAM[690] = 8'b0;
    XRAM[691] = 8'b0;
    XRAM[692] = 8'b0;
    XRAM[693] = 8'b0;
    XRAM[694] = 8'b0;
    XRAM[695] = 8'b0;
    XRAM[696] = 8'b0;
    XRAM[697] = 8'b0;
    XRAM[698] = 8'b0;
    XRAM[699] = 8'b0;
    XRAM[700] = 8'b0;
    XRAM[701] = 8'b0;
    XRAM[702] = 8'b0;
    XRAM[703] = 8'b0;
    XRAM[704] = 8'b0;
    XRAM[705] = 8'b0;
    XRAM[706] = 8'b0;
    XRAM[707] = 8'b0;
    XRAM[708] = 8'b0;
    XRAM[709] = 8'b0;
    XRAM[710] = 8'b0;
    XRAM[711] = 8'b0;
    XRAM[712] = 8'b0;
    XRAM[713] = 8'b0;
    XRAM[714] = 8'b0;
    XRAM[715] = 8'b0;
    XRAM[716] = 8'b0;
    XRAM[717] = 8'b0;
    XRAM[718] = 8'b0;
    XRAM[719] = 8'b0;
    XRAM[720] = 8'b0;
    XRAM[721] = 8'b0;
    XRAM[722] = 8'b0;
    XRAM[723] = 8'b0;
    XRAM[724] = 8'b0;
    XRAM[725] = 8'b0;
    XRAM[726] = 8'b0;
    XRAM[727] = 8'b0;
    XRAM[728] = 8'b0;
    XRAM[729] = 8'b0;
    XRAM[730] = 8'b0;
    XRAM[731] = 8'b0;
    XRAM[732] = 8'b0;
    XRAM[733] = 8'b0;
    XRAM[734] = 8'b0;
    XRAM[735] = 8'b0;
    XRAM[736] = 8'b0;
    XRAM[737] = 8'b0;
    XRAM[738] = 8'b0;
    XRAM[739] = 8'b0;
    XRAM[740] = 8'b0;
    XRAM[741] = 8'b0;
    XRAM[742] = 8'b0;
    XRAM[743] = 8'b0;
    XRAM[744] = 8'b0;
    XRAM[745] = 8'b0;
    XRAM[746] = 8'b0;
    XRAM[747] = 8'b0;
    XRAM[748] = 8'b0;
    XRAM[749] = 8'b0;
    XRAM[750] = 8'b0;
    XRAM[751] = 8'b0;
    XRAM[752] = 8'b0;
    XRAM[753] = 8'b0;
    XRAM[754] = 8'b0;
    XRAM[755] = 8'b0;
    XRAM[756] = 8'b0;
    XRAM[757] = 8'b0;
    XRAM[758] = 8'b0;
    XRAM[759] = 8'b0;
    XRAM[760] = 8'b0;
    XRAM[761] = 8'b0;
    XRAM[762] = 8'b0;
    XRAM[763] = 8'b0;
    XRAM[764] = 8'b0;
    XRAM[765] = 8'b0;
    XRAM[766] = 8'b0;
    XRAM[767] = 8'b0;
    XRAM[768] = 8'b0;
    XRAM[769] = 8'b0;
    XRAM[770] = 8'b0;
    XRAM[771] = 8'b0;
    XRAM[772] = 8'b0;
    XRAM[773] = 8'b0;
    XRAM[774] = 8'b0;
    XRAM[775] = 8'b0;
    XRAM[776] = 8'b0;
    XRAM[777] = 8'b0;
    XRAM[778] = 8'b0;
    XRAM[779] = 8'b0;
    XRAM[780] = 8'b0;
    XRAM[781] = 8'b0;
    XRAM[782] = 8'b0;
    XRAM[783] = 8'b0;
    XRAM[784] = 8'b0;
    XRAM[785] = 8'b0;
    XRAM[786] = 8'b0;
    XRAM[787] = 8'b0;
    XRAM[788] = 8'b0;
    XRAM[789] = 8'b0;
    XRAM[790] = 8'b0;
    XRAM[791] = 8'b0;
    XRAM[792] = 8'b0;
    XRAM[793] = 8'b0;
    XRAM[794] = 8'b0;
    XRAM[795] = 8'b0;
    XRAM[796] = 8'b0;
    XRAM[797] = 8'b0;
    XRAM[798] = 8'b0;
    XRAM[799] = 8'b0;
    XRAM[800] = 8'b0;
    XRAM[801] = 8'b0;
    XRAM[802] = 8'b0;
    XRAM[803] = 8'b0;
    XRAM[804] = 8'b0;
    XRAM[805] = 8'b0;
    XRAM[806] = 8'b0;
    XRAM[807] = 8'b0;
    XRAM[808] = 8'b0;
    XRAM[809] = 8'b0;
    XRAM[810] = 8'b0;
    XRAM[811] = 8'b0;
    XRAM[812] = 8'b0;
    XRAM[813] = 8'b0;
    XRAM[814] = 8'b0;
    XRAM[815] = 8'b0;
    XRAM[816] = 8'b0;
    XRAM[817] = 8'b0;
    XRAM[818] = 8'b0;
    XRAM[819] = 8'b0;
    XRAM[820] = 8'b0;
    XRAM[821] = 8'b0;
    XRAM[822] = 8'b0;
    XRAM[823] = 8'b0;
    XRAM[824] = 8'b0;
    XRAM[825] = 8'b0;
    XRAM[826] = 8'b0;
    XRAM[827] = 8'b0;
    XRAM[828] = 8'b0;
    XRAM[829] = 8'b0;
    XRAM[830] = 8'b0;
    XRAM[831] = 8'b0;
    XRAM[832] = 8'b0;
    XRAM[833] = 8'b0;
    XRAM[834] = 8'b0;
    XRAM[835] = 8'b0;
    XRAM[836] = 8'b0;
    XRAM[837] = 8'b0;
    XRAM[838] = 8'b0;
    XRAM[839] = 8'b0;
    XRAM[840] = 8'b0;
    XRAM[841] = 8'b0;
    XRAM[842] = 8'b0;
    XRAM[843] = 8'b0;
    XRAM[844] = 8'b0;
    XRAM[845] = 8'b0;
    XRAM[846] = 8'b0;
    XRAM[847] = 8'b0;
    XRAM[848] = 8'b0;
    XRAM[849] = 8'b0;
    XRAM[850] = 8'b0;
    XRAM[851] = 8'b0;
    XRAM[852] = 8'b0;
    XRAM[853] = 8'b0;
    XRAM[854] = 8'b0;
    XRAM[855] = 8'b0;
    XRAM[856] = 8'b0;
    XRAM[857] = 8'b0;
    XRAM[858] = 8'b0;
    XRAM[859] = 8'b0;
    XRAM[860] = 8'b0;
    XRAM[861] = 8'b0;
    XRAM[862] = 8'b0;
    XRAM[863] = 8'b0;
    XRAM[864] = 8'b0;
    XRAM[865] = 8'b0;
    XRAM[866] = 8'b0;
    XRAM[867] = 8'b0;
    XRAM[868] = 8'b0;
    XRAM[869] = 8'b0;
    XRAM[870] = 8'b0;
    XRAM[871] = 8'b0;
    XRAM[872] = 8'b0;
    XRAM[873] = 8'b0;
    XRAM[874] = 8'b0;
    XRAM[875] = 8'b0;
    XRAM[876] = 8'b0;
    XRAM[877] = 8'b0;
    XRAM[878] = 8'b0;
    XRAM[879] = 8'b0;
    XRAM[880] = 8'b0;
    XRAM[881] = 8'b0;
    XRAM[882] = 8'b0;
    XRAM[883] = 8'b0;
    XRAM[884] = 8'b0;
    XRAM[885] = 8'b0;
    XRAM[886] = 8'b0;
    XRAM[887] = 8'b0;
    XRAM[888] = 8'b0;
    XRAM[889] = 8'b0;
    XRAM[890] = 8'b0;
    XRAM[891] = 8'b0;
    XRAM[892] = 8'b0;
    XRAM[893] = 8'b0;
    XRAM[894] = 8'b0;
    XRAM[895] = 8'b0;
    XRAM[896] = 8'b0;
    XRAM[897] = 8'b0;
    XRAM[898] = 8'b0;
    XRAM[899] = 8'b0;
    XRAM[900] = 8'b0;
    XRAM[901] = 8'b0;
    XRAM[902] = 8'b0;
    XRAM[903] = 8'b0;
    XRAM[904] = 8'b0;
    XRAM[905] = 8'b0;
    XRAM[906] = 8'b0;
    XRAM[907] = 8'b0;
    XRAM[908] = 8'b0;
    XRAM[909] = 8'b0;
    XRAM[910] = 8'b0;
    XRAM[911] = 8'b0;
    XRAM[912] = 8'b0;
    XRAM[913] = 8'b0;
    XRAM[914] = 8'b0;
    XRAM[915] = 8'b0;
    XRAM[916] = 8'b0;
    XRAM[917] = 8'b0;
    XRAM[918] = 8'b0;
    XRAM[919] = 8'b0;
    XRAM[920] = 8'b0;
    XRAM[921] = 8'b0;
    XRAM[922] = 8'b0;
    XRAM[923] = 8'b0;
    XRAM[924] = 8'b0;
    XRAM[925] = 8'b0;
    XRAM[926] = 8'b0;
    XRAM[927] = 8'b0;
    XRAM[928] = 8'b0;
    XRAM[929] = 8'b0;
    XRAM[930] = 8'b0;
    XRAM[931] = 8'b0;
    XRAM[932] = 8'b0;
    XRAM[933] = 8'b0;
    XRAM[934] = 8'b0;
    XRAM[935] = 8'b0;
    XRAM[936] = 8'b0;
    XRAM[937] = 8'b0;
    XRAM[938] = 8'b0;
    XRAM[939] = 8'b0;
    XRAM[940] = 8'b0;
    XRAM[941] = 8'b0;
    XRAM[942] = 8'b0;
    XRAM[943] = 8'b0;
    XRAM[944] = 8'b0;
    XRAM[945] = 8'b0;
    XRAM[946] = 8'b0;
    XRAM[947] = 8'b0;
    XRAM[948] = 8'b0;
    XRAM[949] = 8'b0;
    XRAM[950] = 8'b0;
    XRAM[951] = 8'b0;
    XRAM[952] = 8'b0;
    XRAM[953] = 8'b0;
    XRAM[954] = 8'b0;
    XRAM[955] = 8'b0;
    XRAM[956] = 8'b0;
    XRAM[957] = 8'b0;
    XRAM[958] = 8'b0;
    XRAM[959] = 8'b0;
    XRAM[960] = 8'b0;
    XRAM[961] = 8'b0;
    XRAM[962] = 8'b0;
    XRAM[963] = 8'b0;
    XRAM[964] = 8'b0;
    XRAM[965] = 8'b0;
    XRAM[966] = 8'b0;
    XRAM[967] = 8'b0;
    XRAM[968] = 8'b0;
    XRAM[969] = 8'b0;
    XRAM[970] = 8'b0;
    XRAM[971] = 8'b0;
    XRAM[972] = 8'b0;
    XRAM[973] = 8'b0;
    XRAM[974] = 8'b0;
    XRAM[975] = 8'b0;
    XRAM[976] = 8'b0;
    XRAM[977] = 8'b0;
    XRAM[978] = 8'b0;
    XRAM[979] = 8'b0;
    XRAM[980] = 8'b0;
    XRAM[981] = 8'b0;
    XRAM[982] = 8'b0;
    XRAM[983] = 8'b0;
    XRAM[984] = 8'b0;
    XRAM[985] = 8'b0;
    XRAM[986] = 8'b0;
    XRAM[987] = 8'b0;
    XRAM[988] = 8'b0;
    XRAM[989] = 8'b0;
    XRAM[990] = 8'b0;
    XRAM[991] = 8'b0;
    XRAM[992] = 8'b0;
    XRAM[993] = 8'b0;
    XRAM[994] = 8'b0;
    XRAM[995] = 8'b0;
    XRAM[996] = 8'b0;
    XRAM[997] = 8'b0;
    XRAM[998] = 8'b0;
    XRAM[999] = 8'b0;
    XRAM[1000] = 8'b0;
    XRAM[1001] = 8'b0;
    XRAM[1002] = 8'b0;
    XRAM[1003] = 8'b0;
    XRAM[1004] = 8'b0;
    XRAM[1005] = 8'b0;
    XRAM[1006] = 8'b0;
    XRAM[1007] = 8'b0;
    XRAM[1008] = 8'b0;
    XRAM[1009] = 8'b0;
    XRAM[1010] = 8'b0;
    XRAM[1011] = 8'b0;
    XRAM[1012] = 8'b0;
    XRAM[1013] = 8'b0;
    XRAM[1014] = 8'b0;
    XRAM[1015] = 8'b0;
    XRAM[1016] = 8'b0;
    XRAM[1017] = 8'b0;
    XRAM[1018] = 8'b0;
    XRAM[1019] = 8'b0;
    XRAM[1020] = 8'b0;
    XRAM[1021] = 8'b0;
    XRAM[1022] = 8'b0;
    XRAM[1023] = 8'b0;
    XRAM[1024] = 8'b0;
    XRAM[1025] = 8'b0;
    XRAM[1026] = 8'b0;
    XRAM[1027] = 8'b0;
    XRAM[1028] = 8'b0;
    XRAM[1029] = 8'b0;
    XRAM[1030] = 8'b0;
    XRAM[1031] = 8'b0;
    XRAM[1032] = 8'b0;
    XRAM[1033] = 8'b0;
    XRAM[1034] = 8'b0;
    XRAM[1035] = 8'b0;
    XRAM[1036] = 8'b0;
    XRAM[1037] = 8'b0;
    XRAM[1038] = 8'b0;
    XRAM[1039] = 8'b0;
    XRAM[1040] = 8'b0;
    XRAM[1041] = 8'b0;
    XRAM[1042] = 8'b0;
    XRAM[1043] = 8'b0;
    XRAM[1044] = 8'b0;
    XRAM[1045] = 8'b0;
    XRAM[1046] = 8'b0;
    XRAM[1047] = 8'b0;
    XRAM[1048] = 8'b0;
    XRAM[1049] = 8'b0;
    XRAM[1050] = 8'b0;
    XRAM[1051] = 8'b0;
    XRAM[1052] = 8'b0;
    XRAM[1053] = 8'b0;
    XRAM[1054] = 8'b0;
    XRAM[1055] = 8'b0;
    XRAM[1056] = 8'b0;
    XRAM[1057] = 8'b0;
    XRAM[1058] = 8'b0;
    XRAM[1059] = 8'b0;
    XRAM[1060] = 8'b0;
    XRAM[1061] = 8'b0;
    XRAM[1062] = 8'b0;
    XRAM[1063] = 8'b0;
    XRAM[1064] = 8'b0;
    XRAM[1065] = 8'b0;
    XRAM[1066] = 8'b0;
    XRAM[1067] = 8'b0;
    XRAM[1068] = 8'b0;
    XRAM[1069] = 8'b0;
    XRAM[1070] = 8'b0;
    XRAM[1071] = 8'b0;
    XRAM[1072] = 8'b0;
    XRAM[1073] = 8'b0;
    XRAM[1074] = 8'b0;
    XRAM[1075] = 8'b0;
    XRAM[1076] = 8'b0;
    XRAM[1077] = 8'b0;
    XRAM[1078] = 8'b0;
    XRAM[1079] = 8'b0;
    XRAM[1080] = 8'b0;
    XRAM[1081] = 8'b0;
    XRAM[1082] = 8'b0;
    XRAM[1083] = 8'b0;
    XRAM[1084] = 8'b0;
    XRAM[1085] = 8'b0;
    XRAM[1086] = 8'b0;
    XRAM[1087] = 8'b0;
    XRAM[1088] = 8'b0;
    XRAM[1089] = 8'b0;
    XRAM[1090] = 8'b0;
    XRAM[1091] = 8'b0;
    XRAM[1092] = 8'b0;
    XRAM[1093] = 8'b0;
    XRAM[1094] = 8'b0;
    XRAM[1095] = 8'b0;
    XRAM[1096] = 8'b0;
    XRAM[1097] = 8'b0;
    XRAM[1098] = 8'b0;
    XRAM[1099] = 8'b0;
    XRAM[1100] = 8'b0;
    XRAM[1101] = 8'b0;
    XRAM[1102] = 8'b0;
    XRAM[1103] = 8'b0;
    XRAM[1104] = 8'b0;
    XRAM[1105] = 8'b0;
    XRAM[1106] = 8'b0;
    XRAM[1107] = 8'b0;
    XRAM[1108] = 8'b0;
    XRAM[1109] = 8'b0;
    XRAM[1110] = 8'b0;
    XRAM[1111] = 8'b0;
    XRAM[1112] = 8'b0;
    XRAM[1113] = 8'b0;
    XRAM[1114] = 8'b0;
    XRAM[1115] = 8'b0;
    XRAM[1116] = 8'b0;
    XRAM[1117] = 8'b0;
    XRAM[1118] = 8'b0;
    XRAM[1119] = 8'b0;
    XRAM[1120] = 8'b0;
    XRAM[1121] = 8'b0;
    XRAM[1122] = 8'b0;
    XRAM[1123] = 8'b0;
    XRAM[1124] = 8'b0;
    XRAM[1125] = 8'b0;
    XRAM[1126] = 8'b0;
    XRAM[1127] = 8'b0;
    XRAM[1128] = 8'b0;
    XRAM[1129] = 8'b0;
    XRAM[1130] = 8'b0;
    XRAM[1131] = 8'b0;
    XRAM[1132] = 8'b0;
    XRAM[1133] = 8'b0;
    XRAM[1134] = 8'b0;
    XRAM[1135] = 8'b0;
    XRAM[1136] = 8'b0;
    XRAM[1137] = 8'b0;
    XRAM[1138] = 8'b0;
    XRAM[1139] = 8'b0;
    XRAM[1140] = 8'b0;
    XRAM[1141] = 8'b0;
    XRAM[1142] = 8'b0;
    XRAM[1143] = 8'b0;
    XRAM[1144] = 8'b0;
    XRAM[1145] = 8'b0;
    XRAM[1146] = 8'b0;
    XRAM[1147] = 8'b0;
    XRAM[1148] = 8'b0;
    XRAM[1149] = 8'b0;
    XRAM[1150] = 8'b0;
    XRAM[1151] = 8'b0;
    XRAM[1152] = 8'b0;
    XRAM[1153] = 8'b0;
    XRAM[1154] = 8'b0;
    XRAM[1155] = 8'b0;
    XRAM[1156] = 8'b0;
    XRAM[1157] = 8'b0;
    XRAM[1158] = 8'b0;
    XRAM[1159] = 8'b0;
    XRAM[1160] = 8'b0;
    XRAM[1161] = 8'b0;
    XRAM[1162] = 8'b0;
    XRAM[1163] = 8'b0;
    XRAM[1164] = 8'b0;
    XRAM[1165] = 8'b0;
    XRAM[1166] = 8'b0;
    XRAM[1167] = 8'b0;
    XRAM[1168] = 8'b0;
    XRAM[1169] = 8'b0;
    XRAM[1170] = 8'b0;
    XRAM[1171] = 8'b0;
    XRAM[1172] = 8'b0;
    XRAM[1173] = 8'b0;
    XRAM[1174] = 8'b0;
    XRAM[1175] = 8'b0;
    XRAM[1176] = 8'b0;
    XRAM[1177] = 8'b0;
    XRAM[1178] = 8'b0;
    XRAM[1179] = 8'b0;
    XRAM[1180] = 8'b0;
    XRAM[1181] = 8'b0;
    XRAM[1182] = 8'b0;
    XRAM[1183] = 8'b0;
    XRAM[1184] = 8'b0;
    XRAM[1185] = 8'b0;
    XRAM[1186] = 8'b0;
    XRAM[1187] = 8'b0;
    XRAM[1188] = 8'b0;
    XRAM[1189] = 8'b0;
    XRAM[1190] = 8'b0;
    XRAM[1191] = 8'b0;
    XRAM[1192] = 8'b0;
    XRAM[1193] = 8'b0;
    XRAM[1194] = 8'b0;
    XRAM[1195] = 8'b0;
    XRAM[1196] = 8'b0;
    XRAM[1197] = 8'b0;
    XRAM[1198] = 8'b0;
    XRAM[1199] = 8'b0;
    XRAM[1200] = 8'b0;
    XRAM[1201] = 8'b0;
    XRAM[1202] = 8'b0;
    XRAM[1203] = 8'b0;
    XRAM[1204] = 8'b0;
    XRAM[1205] = 8'b0;
    XRAM[1206] = 8'b0;
    XRAM[1207] = 8'b0;
    XRAM[1208] = 8'b0;
    XRAM[1209] = 8'b0;
    XRAM[1210] = 8'b0;
    XRAM[1211] = 8'b0;
    XRAM[1212] = 8'b0;
    XRAM[1213] = 8'b0;
    XRAM[1214] = 8'b0;
    XRAM[1215] = 8'b0;
    XRAM[1216] = 8'b0;
    XRAM[1217] = 8'b0;
    XRAM[1218] = 8'b0;
    XRAM[1219] = 8'b0;
    XRAM[1220] = 8'b0;
    XRAM[1221] = 8'b0;
    XRAM[1222] = 8'b0;
    XRAM[1223] = 8'b0;
    XRAM[1224] = 8'b0;
    XRAM[1225] = 8'b0;
    XRAM[1226] = 8'b0;
    XRAM[1227] = 8'b0;
    XRAM[1228] = 8'b0;
    XRAM[1229] = 8'b0;
    XRAM[1230] = 8'b0;
    XRAM[1231] = 8'b0;
    XRAM[1232] = 8'b0;
    XRAM[1233] = 8'b0;
    XRAM[1234] = 8'b0;
    XRAM[1235] = 8'b0;
    XRAM[1236] = 8'b0;
    XRAM[1237] = 8'b0;
    XRAM[1238] = 8'b0;
    XRAM[1239] = 8'b0;
    XRAM[1240] = 8'b0;
    XRAM[1241] = 8'b0;
    XRAM[1242] = 8'b0;
    XRAM[1243] = 8'b0;
    XRAM[1244] = 8'b0;
    XRAM[1245] = 8'b0;
    XRAM[1246] = 8'b0;
    XRAM[1247] = 8'b0;
    XRAM[1248] = 8'b0;
    XRAM[1249] = 8'b0;
    XRAM[1250] = 8'b0;
    XRAM[1251] = 8'b0;
    XRAM[1252] = 8'b0;
    XRAM[1253] = 8'b0;
    XRAM[1254] = 8'b0;
    XRAM[1255] = 8'b0;
    XRAM[1256] = 8'b0;
    XRAM[1257] = 8'b0;
    XRAM[1258] = 8'b0;
    XRAM[1259] = 8'b0;
    XRAM[1260] = 8'b0;
    XRAM[1261] = 8'b0;
    XRAM[1262] = 8'b0;
    XRAM[1263] = 8'b0;
    XRAM[1264] = 8'b0;
    XRAM[1265] = 8'b0;
    XRAM[1266] = 8'b0;
    XRAM[1267] = 8'b0;
    XRAM[1268] = 8'b0;
    XRAM[1269] = 8'b0;
    XRAM[1270] = 8'b0;
    XRAM[1271] = 8'b0;
    XRAM[1272] = 8'b0;
    XRAM[1273] = 8'b0;
    XRAM[1274] = 8'b0;
    XRAM[1275] = 8'b0;
    XRAM[1276] = 8'b0;
    XRAM[1277] = 8'b0;
    XRAM[1278] = 8'b0;
    XRAM[1279] = 8'b0;
    XRAM[1280] = 8'b0;
    XRAM[1281] = 8'b0;
    XRAM[1282] = 8'b0;
    XRAM[1283] = 8'b0;
    XRAM[1284] = 8'b0;
    XRAM[1285] = 8'b0;
    XRAM[1286] = 8'b0;
    XRAM[1287] = 8'b0;
    XRAM[1288] = 8'b0;
    XRAM[1289] = 8'b0;
    XRAM[1290] = 8'b0;
    XRAM[1291] = 8'b0;
    XRAM[1292] = 8'b0;
    XRAM[1293] = 8'b0;
    XRAM[1294] = 8'b0;
    XRAM[1295] = 8'b0;
    XRAM[1296] = 8'b0;
    XRAM[1297] = 8'b0;
    XRAM[1298] = 8'b0;
    XRAM[1299] = 8'b0;
    XRAM[1300] = 8'b0;
    XRAM[1301] = 8'b0;
    XRAM[1302] = 8'b0;
    XRAM[1303] = 8'b0;
    XRAM[1304] = 8'b0;
    XRAM[1305] = 8'b0;
    XRAM[1306] = 8'b0;
    XRAM[1307] = 8'b0;
    XRAM[1308] = 8'b0;
    XRAM[1309] = 8'b0;
    XRAM[1310] = 8'b0;
    XRAM[1311] = 8'b0;
    XRAM[1312] = 8'b0;
    XRAM[1313] = 8'b0;
    XRAM[1314] = 8'b0;
    XRAM[1315] = 8'b0;
    XRAM[1316] = 8'b0;
    XRAM[1317] = 8'b0;
    XRAM[1318] = 8'b0;
    XRAM[1319] = 8'b0;
    XRAM[1320] = 8'b0;
    XRAM[1321] = 8'b0;
    XRAM[1322] = 8'b0;
    XRAM[1323] = 8'b0;
    XRAM[1324] = 8'b0;
    XRAM[1325] = 8'b0;
    XRAM[1326] = 8'b0;
    XRAM[1327] = 8'b0;
    XRAM[1328] = 8'b0;
    XRAM[1329] = 8'b0;
    XRAM[1330] = 8'b0;
    XRAM[1331] = 8'b0;
    XRAM[1332] = 8'b0;
    XRAM[1333] = 8'b0;
    XRAM[1334] = 8'b0;
    XRAM[1335] = 8'b0;
    XRAM[1336] = 8'b0;
    XRAM[1337] = 8'b0;
    XRAM[1338] = 8'b0;
    XRAM[1339] = 8'b0;
    XRAM[1340] = 8'b0;
    XRAM[1341] = 8'b0;
    XRAM[1342] = 8'b0;
    XRAM[1343] = 8'b0;
    XRAM[1344] = 8'b0;
    XRAM[1345] = 8'b0;
    XRAM[1346] = 8'b0;
    XRAM[1347] = 8'b0;
    XRAM[1348] = 8'b0;
    XRAM[1349] = 8'b0;
    XRAM[1350] = 8'b0;
    XRAM[1351] = 8'b0;
    XRAM[1352] = 8'b0;
    XRAM[1353] = 8'b0;
    XRAM[1354] = 8'b0;
    XRAM[1355] = 8'b0;
    XRAM[1356] = 8'b0;
    XRAM[1357] = 8'b0;
    XRAM[1358] = 8'b0;
    XRAM[1359] = 8'b0;
    XRAM[1360] = 8'b0;
    XRAM[1361] = 8'b0;
    XRAM[1362] = 8'b0;
    XRAM[1363] = 8'b0;
    XRAM[1364] = 8'b0;
    XRAM[1365] = 8'b0;
    XRAM[1366] = 8'b0;
    XRAM[1367] = 8'b0;
    XRAM[1368] = 8'b0;
    XRAM[1369] = 8'b0;
    XRAM[1370] = 8'b0;
    XRAM[1371] = 8'b0;
    XRAM[1372] = 8'b0;
    XRAM[1373] = 8'b0;
    XRAM[1374] = 8'b0;
    XRAM[1375] = 8'b0;
    XRAM[1376] = 8'b0;
    XRAM[1377] = 8'b0;
    XRAM[1378] = 8'b0;
    XRAM[1379] = 8'b0;
    XRAM[1380] = 8'b0;
    XRAM[1381] = 8'b0;
    XRAM[1382] = 8'b0;
    XRAM[1383] = 8'b0;
    XRAM[1384] = 8'b0;
    XRAM[1385] = 8'b0;
    XRAM[1386] = 8'b0;
    XRAM[1387] = 8'b0;
    XRAM[1388] = 8'b0;
    XRAM[1389] = 8'b0;
    XRAM[1390] = 8'b0;
    XRAM[1391] = 8'b0;
    XRAM[1392] = 8'b0;
    XRAM[1393] = 8'b0;
    XRAM[1394] = 8'b0;
    XRAM[1395] = 8'b0;
    XRAM[1396] = 8'b0;
    XRAM[1397] = 8'b0;
    XRAM[1398] = 8'b0;
    XRAM[1399] = 8'b0;
    XRAM[1400] = 8'b0;
    XRAM[1401] = 8'b0;
    XRAM[1402] = 8'b0;
    XRAM[1403] = 8'b0;
    XRAM[1404] = 8'b0;
    XRAM[1405] = 8'b0;
    XRAM[1406] = 8'b0;
    XRAM[1407] = 8'b0;
    XRAM[1408] = 8'b0;
    XRAM[1409] = 8'b0;
    XRAM[1410] = 8'b0;
    XRAM[1411] = 8'b0;
    XRAM[1412] = 8'b0;
    XRAM[1413] = 8'b0;
    XRAM[1414] = 8'b0;
    XRAM[1415] = 8'b0;
    XRAM[1416] = 8'b0;
    XRAM[1417] = 8'b0;
    XRAM[1418] = 8'b0;
    XRAM[1419] = 8'b0;
    XRAM[1420] = 8'b0;
    XRAM[1421] = 8'b0;
    XRAM[1422] = 8'b0;
    XRAM[1423] = 8'b0;
    XRAM[1424] = 8'b0;
    XRAM[1425] = 8'b0;
    XRAM[1426] = 8'b0;
    XRAM[1427] = 8'b0;
    XRAM[1428] = 8'b0;
    XRAM[1429] = 8'b0;
    XRAM[1430] = 8'b0;
    XRAM[1431] = 8'b0;
    XRAM[1432] = 8'b0;
    XRAM[1433] = 8'b0;
    XRAM[1434] = 8'b0;
    XRAM[1435] = 8'b0;
    XRAM[1436] = 8'b0;
    XRAM[1437] = 8'b0;
    XRAM[1438] = 8'b0;
    XRAM[1439] = 8'b0;
    XRAM[1440] = 8'b0;
    XRAM[1441] = 8'b0;
    XRAM[1442] = 8'b0;
    XRAM[1443] = 8'b0;
    XRAM[1444] = 8'b0;
    XRAM[1445] = 8'b0;
    XRAM[1446] = 8'b0;
    XRAM[1447] = 8'b0;
    XRAM[1448] = 8'b0;
    XRAM[1449] = 8'b0;
    XRAM[1450] = 8'b0;
    XRAM[1451] = 8'b0;
    XRAM[1452] = 8'b0;
    XRAM[1453] = 8'b0;
    XRAM[1454] = 8'b0;
    XRAM[1455] = 8'b0;
    XRAM[1456] = 8'b0;
    XRAM[1457] = 8'b0;
    XRAM[1458] = 8'b0;
    XRAM[1459] = 8'b0;
    XRAM[1460] = 8'b0;
    XRAM[1461] = 8'b0;
    XRAM[1462] = 8'b0;
    XRAM[1463] = 8'b0;
    XRAM[1464] = 8'b0;
    XRAM[1465] = 8'b0;
    XRAM[1466] = 8'b0;
    XRAM[1467] = 8'b0;
    XRAM[1468] = 8'b0;
    XRAM[1469] = 8'b0;
    XRAM[1470] = 8'b0;
    XRAM[1471] = 8'b0;
    XRAM[1472] = 8'b0;
    XRAM[1473] = 8'b0;
    XRAM[1474] = 8'b0;
    XRAM[1475] = 8'b0;
    XRAM[1476] = 8'b0;
    XRAM[1477] = 8'b0;
    XRAM[1478] = 8'b0;
    XRAM[1479] = 8'b0;
    XRAM[1480] = 8'b0;
    XRAM[1481] = 8'b0;
    XRAM[1482] = 8'b0;
    XRAM[1483] = 8'b0;
    XRAM[1484] = 8'b0;
    XRAM[1485] = 8'b0;
    XRAM[1486] = 8'b0;
    XRAM[1487] = 8'b0;
    XRAM[1488] = 8'b0;
    XRAM[1489] = 8'b0;
    XRAM[1490] = 8'b0;
    XRAM[1491] = 8'b0;
    XRAM[1492] = 8'b0;
    XRAM[1493] = 8'b0;
    XRAM[1494] = 8'b0;
    XRAM[1495] = 8'b0;
    XRAM[1496] = 8'b0;
    XRAM[1497] = 8'b0;
    XRAM[1498] = 8'b0;
    XRAM[1499] = 8'b0;
    XRAM[1500] = 8'b0;
    XRAM[1501] = 8'b0;
    XRAM[1502] = 8'b0;
    XRAM[1503] = 8'b0;
    XRAM[1504] = 8'b0;
    XRAM[1505] = 8'b0;
    XRAM[1506] = 8'b0;
    XRAM[1507] = 8'b0;
    XRAM[1508] = 8'b0;
    XRAM[1509] = 8'b0;
    XRAM[1510] = 8'b0;
    XRAM[1511] = 8'b0;
    XRAM[1512] = 8'b0;
    XRAM[1513] = 8'b0;
    XRAM[1514] = 8'b0;
    XRAM[1515] = 8'b0;
    XRAM[1516] = 8'b0;
    XRAM[1517] = 8'b0;
    XRAM[1518] = 8'b0;
    XRAM[1519] = 8'b0;
    XRAM[1520] = 8'b0;
    XRAM[1521] = 8'b0;
    XRAM[1522] = 8'b0;
    XRAM[1523] = 8'b0;
    XRAM[1524] = 8'b0;
    XRAM[1525] = 8'b0;
    XRAM[1526] = 8'b0;
    XRAM[1527] = 8'b0;
    XRAM[1528] = 8'b0;
    XRAM[1529] = 8'b0;
    XRAM[1530] = 8'b0;
    XRAM[1531] = 8'b0;
    XRAM[1532] = 8'b0;
    XRAM[1533] = 8'b0;
    XRAM[1534] = 8'b0;
    XRAM[1535] = 8'b0;
    XRAM[1536] = 8'b0;
    XRAM[1537] = 8'b0;
    XRAM[1538] = 8'b0;
    XRAM[1539] = 8'b0;
    XRAM[1540] = 8'b0;
    XRAM[1541] = 8'b0;
    XRAM[1542] = 8'b0;
    XRAM[1543] = 8'b0;
    XRAM[1544] = 8'b0;
    XRAM[1545] = 8'b0;
    XRAM[1546] = 8'b0;
    XRAM[1547] = 8'b0;
    XRAM[1548] = 8'b0;
    XRAM[1549] = 8'b0;
    XRAM[1550] = 8'b0;
    XRAM[1551] = 8'b0;
    XRAM[1552] = 8'b0;
    XRAM[1553] = 8'b0;
    XRAM[1554] = 8'b0;
    XRAM[1555] = 8'b0;
    XRAM[1556] = 8'b0;
    XRAM[1557] = 8'b0;
    XRAM[1558] = 8'b0;
    XRAM[1559] = 8'b0;
    XRAM[1560] = 8'b0;
    XRAM[1561] = 8'b0;
    XRAM[1562] = 8'b0;
    XRAM[1563] = 8'b0;
    XRAM[1564] = 8'b0;
    XRAM[1565] = 8'b0;
    XRAM[1566] = 8'b0;
    XRAM[1567] = 8'b0;
    XRAM[1568] = 8'b0;
    XRAM[1569] = 8'b0;
    XRAM[1570] = 8'b0;
    XRAM[1571] = 8'b0;
    XRAM[1572] = 8'b0;
    XRAM[1573] = 8'b0;
    XRAM[1574] = 8'b0;
    XRAM[1575] = 8'b0;
    XRAM[1576] = 8'b0;
    XRAM[1577] = 8'b0;
    XRAM[1578] = 8'b0;
    XRAM[1579] = 8'b0;
    XRAM[1580] = 8'b0;
    XRAM[1581] = 8'b0;
    XRAM[1582] = 8'b0;
    XRAM[1583] = 8'b0;
    XRAM[1584] = 8'b0;
    XRAM[1585] = 8'b0;
    XRAM[1586] = 8'b0;
    XRAM[1587] = 8'b0;
    XRAM[1588] = 8'b0;
    XRAM[1589] = 8'b0;
    XRAM[1590] = 8'b0;
    XRAM[1591] = 8'b0;
    XRAM[1592] = 8'b0;
    XRAM[1593] = 8'b0;
    XRAM[1594] = 8'b0;
    XRAM[1595] = 8'b0;
    XRAM[1596] = 8'b0;
    XRAM[1597] = 8'b0;
    XRAM[1598] = 8'b0;
    XRAM[1599] = 8'b0;
    XRAM[1600] = 8'b0;
    XRAM[1601] = 8'b0;
    XRAM[1602] = 8'b0;
    XRAM[1603] = 8'b0;
    XRAM[1604] = 8'b0;
    XRAM[1605] = 8'b0;
    XRAM[1606] = 8'b0;
    XRAM[1607] = 8'b0;
    XRAM[1608] = 8'b0;
    XRAM[1609] = 8'b0;
    XRAM[1610] = 8'b0;
    XRAM[1611] = 8'b0;
    XRAM[1612] = 8'b0;
    XRAM[1613] = 8'b0;
    XRAM[1614] = 8'b0;
    XRAM[1615] = 8'b0;
    XRAM[1616] = 8'b0;
    XRAM[1617] = 8'b0;
    XRAM[1618] = 8'b0;
    XRAM[1619] = 8'b0;
    XRAM[1620] = 8'b0;
    XRAM[1621] = 8'b0;
    XRAM[1622] = 8'b0;
    XRAM[1623] = 8'b0;
    XRAM[1624] = 8'b0;
    XRAM[1625] = 8'b0;
    XRAM[1626] = 8'b0;
    XRAM[1627] = 8'b0;
    XRAM[1628] = 8'b0;
    XRAM[1629] = 8'b0;
    XRAM[1630] = 8'b0;
    XRAM[1631] = 8'b0;
    XRAM[1632] = 8'b0;
    XRAM[1633] = 8'b0;
    XRAM[1634] = 8'b0;
    XRAM[1635] = 8'b0;
    XRAM[1636] = 8'b0;
    XRAM[1637] = 8'b0;
    XRAM[1638] = 8'b0;
    XRAM[1639] = 8'b0;
    XRAM[1640] = 8'b0;
    XRAM[1641] = 8'b0;
    XRAM[1642] = 8'b0;
    XRAM[1643] = 8'b0;
    XRAM[1644] = 8'b0;
    XRAM[1645] = 8'b0;
    XRAM[1646] = 8'b0;
    XRAM[1647] = 8'b0;
    XRAM[1648] = 8'b0;
    XRAM[1649] = 8'b0;
    XRAM[1650] = 8'b0;
    XRAM[1651] = 8'b0;
    XRAM[1652] = 8'b0;
    XRAM[1653] = 8'b0;
    XRAM[1654] = 8'b0;
    XRAM[1655] = 8'b0;
    XRAM[1656] = 8'b0;
    XRAM[1657] = 8'b0;
    XRAM[1658] = 8'b0;
    XRAM[1659] = 8'b0;
    XRAM[1660] = 8'b0;
    XRAM[1661] = 8'b0;
    XRAM[1662] = 8'b0;
    XRAM[1663] = 8'b0;
    XRAM[1664] = 8'b0;
    XRAM[1665] = 8'b0;
    XRAM[1666] = 8'b0;
    XRAM[1667] = 8'b0;
    XRAM[1668] = 8'b0;
    XRAM[1669] = 8'b0;
    XRAM[1670] = 8'b0;
    XRAM[1671] = 8'b0;
    XRAM[1672] = 8'b0;
    XRAM[1673] = 8'b0;
    XRAM[1674] = 8'b0;
    XRAM[1675] = 8'b0;
    XRAM[1676] = 8'b0;
    XRAM[1677] = 8'b0;
    XRAM[1678] = 8'b0;
    XRAM[1679] = 8'b0;
    XRAM[1680] = 8'b0;
    XRAM[1681] = 8'b0;
    XRAM[1682] = 8'b0;
    XRAM[1683] = 8'b0;
    XRAM[1684] = 8'b0;
    XRAM[1685] = 8'b0;
    XRAM[1686] = 8'b0;
    XRAM[1687] = 8'b0;
    XRAM[1688] = 8'b0;
    XRAM[1689] = 8'b0;
    XRAM[1690] = 8'b0;
    XRAM[1691] = 8'b0;
    XRAM[1692] = 8'b0;
    XRAM[1693] = 8'b0;
    XRAM[1694] = 8'b0;
    XRAM[1695] = 8'b0;
    XRAM[1696] = 8'b0;
    XRAM[1697] = 8'b0;
    XRAM[1698] = 8'b0;
    XRAM[1699] = 8'b0;
    XRAM[1700] = 8'b0;
    XRAM[1701] = 8'b0;
    XRAM[1702] = 8'b0;
    XRAM[1703] = 8'b0;
    XRAM[1704] = 8'b0;
    XRAM[1705] = 8'b0;
    XRAM[1706] = 8'b0;
    XRAM[1707] = 8'b0;
    XRAM[1708] = 8'b0;
    XRAM[1709] = 8'b0;
    XRAM[1710] = 8'b0;
    XRAM[1711] = 8'b0;
    XRAM[1712] = 8'b0;
    XRAM[1713] = 8'b0;
    XRAM[1714] = 8'b0;
    XRAM[1715] = 8'b0;
    XRAM[1716] = 8'b0;
    XRAM[1717] = 8'b0;
    XRAM[1718] = 8'b0;
    XRAM[1719] = 8'b0;
    XRAM[1720] = 8'b0;
    XRAM[1721] = 8'b0;
    XRAM[1722] = 8'b0;
    XRAM[1723] = 8'b0;
    XRAM[1724] = 8'b0;
    XRAM[1725] = 8'b0;
    XRAM[1726] = 8'b0;
    XRAM[1727] = 8'b0;
    XRAM[1728] = 8'b0;
    XRAM[1729] = 8'b0;
    XRAM[1730] = 8'b0;
    XRAM[1731] = 8'b0;
    XRAM[1732] = 8'b0;
    XRAM[1733] = 8'b0;
    XRAM[1734] = 8'b0;
    XRAM[1735] = 8'b0;
    XRAM[1736] = 8'b0;
    XRAM[1737] = 8'b0;
    XRAM[1738] = 8'b0;
    XRAM[1739] = 8'b0;
    XRAM[1740] = 8'b0;
    XRAM[1741] = 8'b0;
    XRAM[1742] = 8'b0;
    XRAM[1743] = 8'b0;
    XRAM[1744] = 8'b0;
    XRAM[1745] = 8'b0;
    XRAM[1746] = 8'b0;
    XRAM[1747] = 8'b0;
    XRAM[1748] = 8'b0;
    XRAM[1749] = 8'b0;
    XRAM[1750] = 8'b0;
    XRAM[1751] = 8'b0;
    XRAM[1752] = 8'b0;
    XRAM[1753] = 8'b0;
    XRAM[1754] = 8'b0;
    XRAM[1755] = 8'b0;
    XRAM[1756] = 8'b0;
    XRAM[1757] = 8'b0;
    XRAM[1758] = 8'b0;
    XRAM[1759] = 8'b0;
    XRAM[1760] = 8'b0;
    XRAM[1761] = 8'b0;
    XRAM[1762] = 8'b0;
    XRAM[1763] = 8'b0;
    XRAM[1764] = 8'b0;
    XRAM[1765] = 8'b0;
    XRAM[1766] = 8'b0;
    XRAM[1767] = 8'b0;
    XRAM[1768] = 8'b0;
    XRAM[1769] = 8'b0;
    XRAM[1770] = 8'b0;
    XRAM[1771] = 8'b0;
    XRAM[1772] = 8'b0;
    XRAM[1773] = 8'b0;
    XRAM[1774] = 8'b0;
    XRAM[1775] = 8'b0;
    XRAM[1776] = 8'b0;
    XRAM[1777] = 8'b0;
    XRAM[1778] = 8'b0;
    XRAM[1779] = 8'b0;
    XRAM[1780] = 8'b0;
    XRAM[1781] = 8'b0;
    XRAM[1782] = 8'b0;
    XRAM[1783] = 8'b0;
    XRAM[1784] = 8'b0;
    XRAM[1785] = 8'b0;
    XRAM[1786] = 8'b0;
    XRAM[1787] = 8'b0;
    XRAM[1788] = 8'b0;
    XRAM[1789] = 8'b0;
    XRAM[1790] = 8'b0;
    XRAM[1791] = 8'b0;
    XRAM[1792] = 8'b0;
    XRAM[1793] = 8'b0;
    XRAM[1794] = 8'b0;
    XRAM[1795] = 8'b0;
    XRAM[1796] = 8'b0;
    XRAM[1797] = 8'b0;
    XRAM[1798] = 8'b0;
    XRAM[1799] = 8'b0;
    XRAM[1800] = 8'b0;
    XRAM[1801] = 8'b0;
    XRAM[1802] = 8'b0;
    XRAM[1803] = 8'b0;
    XRAM[1804] = 8'b0;
    XRAM[1805] = 8'b0;
    XRAM[1806] = 8'b0;
    XRAM[1807] = 8'b0;
    XRAM[1808] = 8'b0;
    XRAM[1809] = 8'b0;
    XRAM[1810] = 8'b0;
    XRAM[1811] = 8'b0;
    XRAM[1812] = 8'b0;
    XRAM[1813] = 8'b0;
    XRAM[1814] = 8'b0;
    XRAM[1815] = 8'b0;
    XRAM[1816] = 8'b0;
    XRAM[1817] = 8'b0;
    XRAM[1818] = 8'b0;
    XRAM[1819] = 8'b0;
    XRAM[1820] = 8'b0;
    XRAM[1821] = 8'b0;
    XRAM[1822] = 8'b0;
    XRAM[1823] = 8'b0;
    XRAM[1824] = 8'b0;
    XRAM[1825] = 8'b0;
    XRAM[1826] = 8'b0;
    XRAM[1827] = 8'b0;
    XRAM[1828] = 8'b0;
    XRAM[1829] = 8'b0;
    XRAM[1830] = 8'b0;
    XRAM[1831] = 8'b0;
    XRAM[1832] = 8'b0;
    XRAM[1833] = 8'b0;
    XRAM[1834] = 8'b0;
    XRAM[1835] = 8'b0;
    XRAM[1836] = 8'b0;
    XRAM[1837] = 8'b0;
    XRAM[1838] = 8'b0;
    XRAM[1839] = 8'b0;
    XRAM[1840] = 8'b0;
    XRAM[1841] = 8'b0;
    XRAM[1842] = 8'b0;
    XRAM[1843] = 8'b0;
    XRAM[1844] = 8'b0;
    XRAM[1845] = 8'b0;
    XRAM[1846] = 8'b0;
    XRAM[1847] = 8'b0;
    XRAM[1848] = 8'b0;
    XRAM[1849] = 8'b0;
    XRAM[1850] = 8'b0;
    XRAM[1851] = 8'b0;
    XRAM[1852] = 8'b0;
    XRAM[1853] = 8'b0;
    XRAM[1854] = 8'b0;
    XRAM[1855] = 8'b0;
    XRAM[1856] = 8'b0;
    XRAM[1857] = 8'b0;
    XRAM[1858] = 8'b0;
    XRAM[1859] = 8'b0;
    XRAM[1860] = 8'b0;
    XRAM[1861] = 8'b0;
    XRAM[1862] = 8'b0;
    XRAM[1863] = 8'b0;
    XRAM[1864] = 8'b0;
    XRAM[1865] = 8'b0;
    XRAM[1866] = 8'b0;
    XRAM[1867] = 8'b0;
    XRAM[1868] = 8'b0;
    XRAM[1869] = 8'b0;
    XRAM[1870] = 8'b0;
    XRAM[1871] = 8'b0;
    XRAM[1872] = 8'b0;
    XRAM[1873] = 8'b0;
    XRAM[1874] = 8'b0;
    XRAM[1875] = 8'b0;
    XRAM[1876] = 8'b0;
    XRAM[1877] = 8'b0;
    XRAM[1878] = 8'b0;
    XRAM[1879] = 8'b0;
    XRAM[1880] = 8'b0;
    XRAM[1881] = 8'b0;
    XRAM[1882] = 8'b0;
    XRAM[1883] = 8'b0;
    XRAM[1884] = 8'b0;
    XRAM[1885] = 8'b0;
    XRAM[1886] = 8'b0;
    XRAM[1887] = 8'b0;
    XRAM[1888] = 8'b0;
    XRAM[1889] = 8'b0;
    XRAM[1890] = 8'b0;
    XRAM[1891] = 8'b0;
    XRAM[1892] = 8'b0;
    XRAM[1893] = 8'b0;
    XRAM[1894] = 8'b0;
    XRAM[1895] = 8'b0;
    XRAM[1896] = 8'b0;
    XRAM[1897] = 8'b0;
    XRAM[1898] = 8'b0;
    XRAM[1899] = 8'b0;
    XRAM[1900] = 8'b0;
    XRAM[1901] = 8'b0;
    XRAM[1902] = 8'b0;
    XRAM[1903] = 8'b0;
    XRAM[1904] = 8'b0;
    XRAM[1905] = 8'b0;
    XRAM[1906] = 8'b0;
    XRAM[1907] = 8'b0;
    XRAM[1908] = 8'b0;
    XRAM[1909] = 8'b0;
    XRAM[1910] = 8'b0;
    XRAM[1911] = 8'b0;
    XRAM[1912] = 8'b0;
    XRAM[1913] = 8'b0;
    XRAM[1914] = 8'b0;
    XRAM[1915] = 8'b0;
    XRAM[1916] = 8'b0;
    XRAM[1917] = 8'b0;
    XRAM[1918] = 8'b0;
    XRAM[1919] = 8'b0;
    XRAM[1920] = 8'b0;
    XRAM[1921] = 8'b0;
    XRAM[1922] = 8'b0;
    XRAM[1923] = 8'b0;
    XRAM[1924] = 8'b0;
    XRAM[1925] = 8'b0;
    XRAM[1926] = 8'b0;
    XRAM[1927] = 8'b0;
    XRAM[1928] = 8'b0;
    XRAM[1929] = 8'b0;
    XRAM[1930] = 8'b0;
    XRAM[1931] = 8'b0;
    XRAM[1932] = 8'b0;
    XRAM[1933] = 8'b0;
    XRAM[1934] = 8'b0;
    XRAM[1935] = 8'b0;
    XRAM[1936] = 8'b0;
    XRAM[1937] = 8'b0;
    XRAM[1938] = 8'b0;
    XRAM[1939] = 8'b0;
    XRAM[1940] = 8'b0;
    XRAM[1941] = 8'b0;
    XRAM[1942] = 8'b0;
    XRAM[1943] = 8'b0;
    XRAM[1944] = 8'b0;
    XRAM[1945] = 8'b0;
    XRAM[1946] = 8'b0;
    XRAM[1947] = 8'b0;
    XRAM[1948] = 8'b0;
    XRAM[1949] = 8'b0;
    XRAM[1950] = 8'b0;
    XRAM[1951] = 8'b0;
    XRAM[1952] = 8'b0;
    XRAM[1953] = 8'b0;
    XRAM[1954] = 8'b0;
    XRAM[1955] = 8'b0;
    XRAM[1956] = 8'b0;
    XRAM[1957] = 8'b0;
    XRAM[1958] = 8'b0;
    XRAM[1959] = 8'b0;
    XRAM[1960] = 8'b0;
    XRAM[1961] = 8'b0;
    XRAM[1962] = 8'b0;
    XRAM[1963] = 8'b0;
    XRAM[1964] = 8'b0;
    XRAM[1965] = 8'b0;
    XRAM[1966] = 8'b0;
    XRAM[1967] = 8'b0;
    XRAM[1968] = 8'b0;
    XRAM[1969] = 8'b0;
    XRAM[1970] = 8'b0;
    XRAM[1971] = 8'b0;
    XRAM[1972] = 8'b0;
    XRAM[1973] = 8'b0;
    XRAM[1974] = 8'b0;
    XRAM[1975] = 8'b0;
    XRAM[1976] = 8'b0;
    XRAM[1977] = 8'b0;
    XRAM[1978] = 8'b0;
    XRAM[1979] = 8'b0;
    XRAM[1980] = 8'b0;
    XRAM[1981] = 8'b0;
    XRAM[1982] = 8'b0;
    XRAM[1983] = 8'b0;
    XRAM[1984] = 8'b0;
    XRAM[1985] = 8'b0;
    XRAM[1986] = 8'b0;
    XRAM[1987] = 8'b0;
    XRAM[1988] = 8'b0;
    XRAM[1989] = 8'b0;
    XRAM[1990] = 8'b0;
    XRAM[1991] = 8'b0;
    XRAM[1992] = 8'b0;
    XRAM[1993] = 8'b0;
    XRAM[1994] = 8'b0;
    XRAM[1995] = 8'b0;
    XRAM[1996] = 8'b0;
    XRAM[1997] = 8'b0;
    XRAM[1998] = 8'b0;
    XRAM[1999] = 8'b0;
    XRAM[2000] = 8'b0;
    XRAM[2001] = 8'b0;
    XRAM[2002] = 8'b0;
    XRAM[2003] = 8'b0;
    XRAM[2004] = 8'b0;
    XRAM[2005] = 8'b0;
    XRAM[2006] = 8'b0;
    XRAM[2007] = 8'b0;
    XRAM[2008] = 8'b0;
    XRAM[2009] = 8'b0;
    XRAM[2010] = 8'b0;
    XRAM[2011] = 8'b0;
    XRAM[2012] = 8'b0;
    XRAM[2013] = 8'b0;
    XRAM[2014] = 8'b0;
    XRAM[2015] = 8'b0;
    XRAM[2016] = 8'b0;
    XRAM[2017] = 8'b0;
    XRAM[2018] = 8'b0;
    XRAM[2019] = 8'b0;
    XRAM[2020] = 8'b0;
    XRAM[2021] = 8'b0;
    XRAM[2022] = 8'b0;
    XRAM[2023] = 8'b0;
    XRAM[2024] = 8'b0;
    XRAM[2025] = 8'b0;
    XRAM[2026] = 8'b0;
    XRAM[2027] = 8'b0;
    XRAM[2028] = 8'b0;
    XRAM[2029] = 8'b0;
    XRAM[2030] = 8'b0;
    XRAM[2031] = 8'b0;
    XRAM[2032] = 8'b0;
    XRAM[2033] = 8'b0;
    XRAM[2034] = 8'b0;
    XRAM[2035] = 8'b0;
    XRAM[2036] = 8'b0;
    XRAM[2037] = 8'b0;
    XRAM[2038] = 8'b0;
    XRAM[2039] = 8'b0;
    XRAM[2040] = 8'b0;
    XRAM[2041] = 8'b0;
    XRAM[2042] = 8'b0;
    XRAM[2043] = 8'b0;
    XRAM[2044] = 8'b0;
    XRAM[2045] = 8'b0;
    XRAM[2046] = 8'b0;
    XRAM[2047] = 8'b0;
    XRAM[2048] = 8'b0;
    XRAM[2049] = 8'b0;
    XRAM[2050] = 8'b0;
    XRAM[2051] = 8'b0;
    XRAM[2052] = 8'b0;
    XRAM[2053] = 8'b0;
    XRAM[2054] = 8'b0;
    XRAM[2055] = 8'b0;
    XRAM[2056] = 8'b0;
    XRAM[2057] = 8'b0;
    XRAM[2058] = 8'b0;
    XRAM[2059] = 8'b0;
    XRAM[2060] = 8'b0;
    XRAM[2061] = 8'b0;
    XRAM[2062] = 8'b0;
    XRAM[2063] = 8'b0;
    XRAM[2064] = 8'b0;
    XRAM[2065] = 8'b0;
    XRAM[2066] = 8'b0;
    XRAM[2067] = 8'b0;
    XRAM[2068] = 8'b0;
    XRAM[2069] = 8'b0;
    XRAM[2070] = 8'b0;
    XRAM[2071] = 8'b0;
    XRAM[2072] = 8'b0;
    XRAM[2073] = 8'b0;
    XRAM[2074] = 8'b0;
    XRAM[2075] = 8'b0;
    XRAM[2076] = 8'b0;
    XRAM[2077] = 8'b0;
    XRAM[2078] = 8'b0;
    XRAM[2079] = 8'b0;
    XRAM[2080] = 8'b0;
    XRAM[2081] = 8'b0;
    XRAM[2082] = 8'b0;
    XRAM[2083] = 8'b0;
    XRAM[2084] = 8'b0;
    XRAM[2085] = 8'b0;
    XRAM[2086] = 8'b0;
    XRAM[2087] = 8'b0;
    XRAM[2088] = 8'b0;
    XRAM[2089] = 8'b0;
    XRAM[2090] = 8'b0;
    XRAM[2091] = 8'b0;
    XRAM[2092] = 8'b0;
    XRAM[2093] = 8'b0;
    XRAM[2094] = 8'b0;
    XRAM[2095] = 8'b0;
    XRAM[2096] = 8'b0;
    XRAM[2097] = 8'b0;
    XRAM[2098] = 8'b0;
    XRAM[2099] = 8'b0;
    XRAM[2100] = 8'b0;
    XRAM[2101] = 8'b0;
    XRAM[2102] = 8'b0;
    XRAM[2103] = 8'b0;
    XRAM[2104] = 8'b0;
    XRAM[2105] = 8'b0;
    XRAM[2106] = 8'b0;
    XRAM[2107] = 8'b0;
    XRAM[2108] = 8'b0;
    XRAM[2109] = 8'b0;
    XRAM[2110] = 8'b0;
    XRAM[2111] = 8'b0;
    XRAM[2112] = 8'b0;
    XRAM[2113] = 8'b0;
    XRAM[2114] = 8'b0;
    XRAM[2115] = 8'b0;
    XRAM[2116] = 8'b0;
    XRAM[2117] = 8'b0;
    XRAM[2118] = 8'b0;
    XRAM[2119] = 8'b0;
    XRAM[2120] = 8'b0;
    XRAM[2121] = 8'b0;
    XRAM[2122] = 8'b0;
    XRAM[2123] = 8'b0;
    XRAM[2124] = 8'b0;
    XRAM[2125] = 8'b0;
    XRAM[2126] = 8'b0;
    XRAM[2127] = 8'b0;
    XRAM[2128] = 8'b0;
    XRAM[2129] = 8'b0;
    XRAM[2130] = 8'b0;
    XRAM[2131] = 8'b0;
    XRAM[2132] = 8'b0;
    XRAM[2133] = 8'b0;
    XRAM[2134] = 8'b0;
    XRAM[2135] = 8'b0;
    XRAM[2136] = 8'b0;
    XRAM[2137] = 8'b0;
    XRAM[2138] = 8'b0;
    XRAM[2139] = 8'b0;
    XRAM[2140] = 8'b0;
    XRAM[2141] = 8'b0;
    XRAM[2142] = 8'b0;
    XRAM[2143] = 8'b0;
    XRAM[2144] = 8'b0;
    XRAM[2145] = 8'b0;
    XRAM[2146] = 8'b0;
    XRAM[2147] = 8'b0;
    XRAM[2148] = 8'b0;
    XRAM[2149] = 8'b0;
    XRAM[2150] = 8'b0;
    XRAM[2151] = 8'b0;
    XRAM[2152] = 8'b0;
    XRAM[2153] = 8'b0;
    XRAM[2154] = 8'b0;
    XRAM[2155] = 8'b0;
    XRAM[2156] = 8'b0;
    XRAM[2157] = 8'b0;
    XRAM[2158] = 8'b0;
    XRAM[2159] = 8'b0;
    XRAM[2160] = 8'b0;
    XRAM[2161] = 8'b0;
    XRAM[2162] = 8'b0;
    XRAM[2163] = 8'b0;
    XRAM[2164] = 8'b0;
    XRAM[2165] = 8'b0;
    XRAM[2166] = 8'b0;
    XRAM[2167] = 8'b0;
    XRAM[2168] = 8'b0;
    XRAM[2169] = 8'b0;
    XRAM[2170] = 8'b0;
    XRAM[2171] = 8'b0;
    XRAM[2172] = 8'b0;
    XRAM[2173] = 8'b0;
    XRAM[2174] = 8'b0;
    XRAM[2175] = 8'b0;
    XRAM[2176] = 8'b0;
    XRAM[2177] = 8'b0;
    XRAM[2178] = 8'b0;
    XRAM[2179] = 8'b0;
    XRAM[2180] = 8'b0;
    XRAM[2181] = 8'b0;
    XRAM[2182] = 8'b0;
    XRAM[2183] = 8'b0;
    XRAM[2184] = 8'b0;
    XRAM[2185] = 8'b0;
    XRAM[2186] = 8'b0;
    XRAM[2187] = 8'b0;
    XRAM[2188] = 8'b0;
    XRAM[2189] = 8'b0;
    XRAM[2190] = 8'b0;
    XRAM[2191] = 8'b0;
    XRAM[2192] = 8'b0;
    XRAM[2193] = 8'b0;
    XRAM[2194] = 8'b0;
    XRAM[2195] = 8'b0;
    XRAM[2196] = 8'b0;
    XRAM[2197] = 8'b0;
    XRAM[2198] = 8'b0;
    XRAM[2199] = 8'b0;
    XRAM[2200] = 8'b0;
    XRAM[2201] = 8'b0;
    XRAM[2202] = 8'b0;
    XRAM[2203] = 8'b0;
    XRAM[2204] = 8'b0;
    XRAM[2205] = 8'b0;
    XRAM[2206] = 8'b0;
    XRAM[2207] = 8'b0;
    XRAM[2208] = 8'b0;
    XRAM[2209] = 8'b0;
    XRAM[2210] = 8'b0;
    XRAM[2211] = 8'b0;
    XRAM[2212] = 8'b0;
    XRAM[2213] = 8'b0;
    XRAM[2214] = 8'b0;
    XRAM[2215] = 8'b0;
    XRAM[2216] = 8'b0;
    XRAM[2217] = 8'b0;
    XRAM[2218] = 8'b0;
    XRAM[2219] = 8'b0;
    XRAM[2220] = 8'b0;
    XRAM[2221] = 8'b0;
    XRAM[2222] = 8'b0;
    XRAM[2223] = 8'b0;
    XRAM[2224] = 8'b0;
    XRAM[2225] = 8'b0;
    XRAM[2226] = 8'b0;
    XRAM[2227] = 8'b0;
    XRAM[2228] = 8'b0;
    XRAM[2229] = 8'b0;
    XRAM[2230] = 8'b0;
    XRAM[2231] = 8'b0;
    XRAM[2232] = 8'b0;
    XRAM[2233] = 8'b0;
    XRAM[2234] = 8'b0;
    XRAM[2235] = 8'b0;
    XRAM[2236] = 8'b0;
    XRAM[2237] = 8'b0;
    XRAM[2238] = 8'b0;
    XRAM[2239] = 8'b0;
    XRAM[2240] = 8'b0;
    XRAM[2241] = 8'b0;
    XRAM[2242] = 8'b0;
    XRAM[2243] = 8'b0;
    XRAM[2244] = 8'b0;
    XRAM[2245] = 8'b0;
    XRAM[2246] = 8'b0;
    XRAM[2247] = 8'b0;
    XRAM[2248] = 8'b0;
    XRAM[2249] = 8'b0;
    XRAM[2250] = 8'b0;
    XRAM[2251] = 8'b0;
    XRAM[2252] = 8'b0;
    XRAM[2253] = 8'b0;
    XRAM[2254] = 8'b0;
    XRAM[2255] = 8'b0;
    XRAM[2256] = 8'b0;
    XRAM[2257] = 8'b0;
    XRAM[2258] = 8'b0;
    XRAM[2259] = 8'b0;
    XRAM[2260] = 8'b0;
    XRAM[2261] = 8'b0;
    XRAM[2262] = 8'b0;
    XRAM[2263] = 8'b0;
    XRAM[2264] = 8'b0;
    XRAM[2265] = 8'b0;
    XRAM[2266] = 8'b0;
    XRAM[2267] = 8'b0;
    XRAM[2268] = 8'b0;
    XRAM[2269] = 8'b0;
    XRAM[2270] = 8'b0;
    XRAM[2271] = 8'b0;
    XRAM[2272] = 8'b0;
    XRAM[2273] = 8'b0;
    XRAM[2274] = 8'b0;
    XRAM[2275] = 8'b0;
    XRAM[2276] = 8'b0;
    XRAM[2277] = 8'b0;
    XRAM[2278] = 8'b0;
    XRAM[2279] = 8'b0;
    XRAM[2280] = 8'b0;
    XRAM[2281] = 8'b0;
    XRAM[2282] = 8'b0;
    XRAM[2283] = 8'b0;
    XRAM[2284] = 8'b0;
    XRAM[2285] = 8'b0;
    XRAM[2286] = 8'b0;
    XRAM[2287] = 8'b0;
    XRAM[2288] = 8'b0;
    XRAM[2289] = 8'b0;
    XRAM[2290] = 8'b0;
    XRAM[2291] = 8'b0;
    XRAM[2292] = 8'b0;
    XRAM[2293] = 8'b0;
    XRAM[2294] = 8'b0;
    XRAM[2295] = 8'b0;
    XRAM[2296] = 8'b0;
    XRAM[2297] = 8'b0;
    XRAM[2298] = 8'b0;
    XRAM[2299] = 8'b0;
    XRAM[2300] = 8'b0;
    XRAM[2301] = 8'b0;
    XRAM[2302] = 8'b0;
    XRAM[2303] = 8'b0;
    XRAM[2304] = 8'b0;
    XRAM[2305] = 8'b0;
    XRAM[2306] = 8'b0;
    XRAM[2307] = 8'b0;
    XRAM[2308] = 8'b0;
    XRAM[2309] = 8'b0;
    XRAM[2310] = 8'b0;
    XRAM[2311] = 8'b0;
    XRAM[2312] = 8'b0;
    XRAM[2313] = 8'b0;
    XRAM[2314] = 8'b0;
    XRAM[2315] = 8'b0;
    XRAM[2316] = 8'b0;
    XRAM[2317] = 8'b0;
    XRAM[2318] = 8'b0;
    XRAM[2319] = 8'b0;
    XRAM[2320] = 8'b0;
    XRAM[2321] = 8'b0;
    XRAM[2322] = 8'b0;
    XRAM[2323] = 8'b0;
    XRAM[2324] = 8'b0;
    XRAM[2325] = 8'b0;
    XRAM[2326] = 8'b0;
    XRAM[2327] = 8'b0;
    XRAM[2328] = 8'b0;
    XRAM[2329] = 8'b0;
    XRAM[2330] = 8'b0;
    XRAM[2331] = 8'b0;
    XRAM[2332] = 8'b0;
    XRAM[2333] = 8'b0;
    XRAM[2334] = 8'b0;
    XRAM[2335] = 8'b0;
    XRAM[2336] = 8'b0;
    XRAM[2337] = 8'b0;
    XRAM[2338] = 8'b0;
    XRAM[2339] = 8'b0;
    XRAM[2340] = 8'b0;
    XRAM[2341] = 8'b0;
    XRAM[2342] = 8'b0;
    XRAM[2343] = 8'b0;
    XRAM[2344] = 8'b0;
    XRAM[2345] = 8'b0;
    XRAM[2346] = 8'b0;
    XRAM[2347] = 8'b0;
    XRAM[2348] = 8'b0;
    XRAM[2349] = 8'b0;
    XRAM[2350] = 8'b0;
    XRAM[2351] = 8'b0;
    XRAM[2352] = 8'b0;
    XRAM[2353] = 8'b0;
    XRAM[2354] = 8'b0;
    XRAM[2355] = 8'b0;
    XRAM[2356] = 8'b0;
    XRAM[2357] = 8'b0;
    XRAM[2358] = 8'b0;
    XRAM[2359] = 8'b0;
    XRAM[2360] = 8'b0;
    XRAM[2361] = 8'b0;
    XRAM[2362] = 8'b0;
    XRAM[2363] = 8'b0;
    XRAM[2364] = 8'b0;
    XRAM[2365] = 8'b0;
    XRAM[2366] = 8'b0;
    XRAM[2367] = 8'b0;
    XRAM[2368] = 8'b0;
    XRAM[2369] = 8'b0;
    XRAM[2370] = 8'b0;
    XRAM[2371] = 8'b0;
    XRAM[2372] = 8'b0;
    XRAM[2373] = 8'b0;
    XRAM[2374] = 8'b0;
    XRAM[2375] = 8'b0;
    XRAM[2376] = 8'b0;
    XRAM[2377] = 8'b0;
    XRAM[2378] = 8'b0;
    XRAM[2379] = 8'b0;
    XRAM[2380] = 8'b0;
    XRAM[2381] = 8'b0;
    XRAM[2382] = 8'b0;
    XRAM[2383] = 8'b0;
    XRAM[2384] = 8'b0;
    XRAM[2385] = 8'b0;
    XRAM[2386] = 8'b0;
    XRAM[2387] = 8'b0;
    XRAM[2388] = 8'b0;
    XRAM[2389] = 8'b0;
    XRAM[2390] = 8'b0;
    XRAM[2391] = 8'b0;
    XRAM[2392] = 8'b0;
    XRAM[2393] = 8'b0;
    XRAM[2394] = 8'b0;
    XRAM[2395] = 8'b0;
    XRAM[2396] = 8'b0;
    XRAM[2397] = 8'b0;
    XRAM[2398] = 8'b0;
    XRAM[2399] = 8'b0;
    XRAM[2400] = 8'b0;
    XRAM[2401] = 8'b0;
    XRAM[2402] = 8'b0;
    XRAM[2403] = 8'b0;
    XRAM[2404] = 8'b0;
    XRAM[2405] = 8'b0;
    XRAM[2406] = 8'b0;
    XRAM[2407] = 8'b0;
    XRAM[2408] = 8'b0;
    XRAM[2409] = 8'b0;
    XRAM[2410] = 8'b0;
    XRAM[2411] = 8'b0;
    XRAM[2412] = 8'b0;
    XRAM[2413] = 8'b0;
    XRAM[2414] = 8'b0;
    XRAM[2415] = 8'b0;
    XRAM[2416] = 8'b0;
    XRAM[2417] = 8'b0;
    XRAM[2418] = 8'b0;
    XRAM[2419] = 8'b0;
    XRAM[2420] = 8'b0;
    XRAM[2421] = 8'b0;
    XRAM[2422] = 8'b0;
    XRAM[2423] = 8'b0;
    XRAM[2424] = 8'b0;
    XRAM[2425] = 8'b0;
    XRAM[2426] = 8'b0;
    XRAM[2427] = 8'b0;
    XRAM[2428] = 8'b0;
    XRAM[2429] = 8'b0;
    XRAM[2430] = 8'b0;
    XRAM[2431] = 8'b0;
    XRAM[2432] = 8'b0;
    XRAM[2433] = 8'b0;
    XRAM[2434] = 8'b0;
    XRAM[2435] = 8'b0;
    XRAM[2436] = 8'b0;
    XRAM[2437] = 8'b0;
    XRAM[2438] = 8'b0;
    XRAM[2439] = 8'b0;
    XRAM[2440] = 8'b0;
    XRAM[2441] = 8'b0;
    XRAM[2442] = 8'b0;
    XRAM[2443] = 8'b0;
    XRAM[2444] = 8'b0;
    XRAM[2445] = 8'b0;
    XRAM[2446] = 8'b0;
    XRAM[2447] = 8'b0;
    XRAM[2448] = 8'b0;
    XRAM[2449] = 8'b0;
    XRAM[2450] = 8'b0;
    XRAM[2451] = 8'b0;
    XRAM[2452] = 8'b0;
    XRAM[2453] = 8'b0;
    XRAM[2454] = 8'b0;
    XRAM[2455] = 8'b0;
    XRAM[2456] = 8'b0;
    XRAM[2457] = 8'b0;
    XRAM[2458] = 8'b0;
    XRAM[2459] = 8'b0;
    XRAM[2460] = 8'b0;
    XRAM[2461] = 8'b0;
    XRAM[2462] = 8'b0;
    XRAM[2463] = 8'b0;
    XRAM[2464] = 8'b0;
    XRAM[2465] = 8'b0;
    XRAM[2466] = 8'b0;
    XRAM[2467] = 8'b0;
    XRAM[2468] = 8'b0;
    XRAM[2469] = 8'b0;
    XRAM[2470] = 8'b0;
    XRAM[2471] = 8'b0;
    XRAM[2472] = 8'b0;
    XRAM[2473] = 8'b0;
    XRAM[2474] = 8'b0;
    XRAM[2475] = 8'b0;
    XRAM[2476] = 8'b0;
    XRAM[2477] = 8'b0;
    XRAM[2478] = 8'b0;
    XRAM[2479] = 8'b0;
    XRAM[2480] = 8'b0;
    XRAM[2481] = 8'b0;
    XRAM[2482] = 8'b0;
    XRAM[2483] = 8'b0;
    XRAM[2484] = 8'b0;
    XRAM[2485] = 8'b0;
    XRAM[2486] = 8'b0;
    XRAM[2487] = 8'b0;
    XRAM[2488] = 8'b0;
    XRAM[2489] = 8'b0;
    XRAM[2490] = 8'b0;
    XRAM[2491] = 8'b0;
    XRAM[2492] = 8'b0;
    XRAM[2493] = 8'b0;
    XRAM[2494] = 8'b0;
    XRAM[2495] = 8'b0;
    XRAM[2496] = 8'b0;
    XRAM[2497] = 8'b0;
    XRAM[2498] = 8'b0;
    XRAM[2499] = 8'b0;
    XRAM[2500] = 8'b0;
    XRAM[2501] = 8'b0;
    XRAM[2502] = 8'b0;
    XRAM[2503] = 8'b0;
    XRAM[2504] = 8'b0;
    XRAM[2505] = 8'b0;
    XRAM[2506] = 8'b0;
    XRAM[2507] = 8'b0;
    XRAM[2508] = 8'b0;
    XRAM[2509] = 8'b0;
    XRAM[2510] = 8'b0;
    XRAM[2511] = 8'b0;
    XRAM[2512] = 8'b0;
    XRAM[2513] = 8'b0;
    XRAM[2514] = 8'b0;
    XRAM[2515] = 8'b0;
    XRAM[2516] = 8'b0;
    XRAM[2517] = 8'b0;
    XRAM[2518] = 8'b0;
    XRAM[2519] = 8'b0;
    XRAM[2520] = 8'b0;
    XRAM[2521] = 8'b0;
    XRAM[2522] = 8'b0;
    XRAM[2523] = 8'b0;
    XRAM[2524] = 8'b0;
    XRAM[2525] = 8'b0;
    XRAM[2526] = 8'b0;
    XRAM[2527] = 8'b0;
    XRAM[2528] = 8'b0;
    XRAM[2529] = 8'b0;
    XRAM[2530] = 8'b0;
    XRAM[2531] = 8'b0;
    XRAM[2532] = 8'b0;
    XRAM[2533] = 8'b0;
    XRAM[2534] = 8'b0;
    XRAM[2535] = 8'b0;
    XRAM[2536] = 8'b0;
    XRAM[2537] = 8'b0;
    XRAM[2538] = 8'b0;
    XRAM[2539] = 8'b0;
    XRAM[2540] = 8'b0;
    XRAM[2541] = 8'b0;
    XRAM[2542] = 8'b0;
    XRAM[2543] = 8'b0;
    XRAM[2544] = 8'b0;
    XRAM[2545] = 8'b0;
    XRAM[2546] = 8'b0;
    XRAM[2547] = 8'b0;
    XRAM[2548] = 8'b0;
    XRAM[2549] = 8'b0;
    XRAM[2550] = 8'b0;
    XRAM[2551] = 8'b0;
    XRAM[2552] = 8'b0;
    XRAM[2553] = 8'b0;
    XRAM[2554] = 8'b0;
    XRAM[2555] = 8'b0;
    XRAM[2556] = 8'b0;
    XRAM[2557] = 8'b0;
    XRAM[2558] = 8'b0;
    XRAM[2559] = 8'b0;
    XRAM[2560] = 8'b0;
    XRAM[2561] = 8'b0;
    XRAM[2562] = 8'b0;
    XRAM[2563] = 8'b0;
    XRAM[2564] = 8'b0;
    XRAM[2565] = 8'b0;
    XRAM[2566] = 8'b0;
    XRAM[2567] = 8'b0;
    XRAM[2568] = 8'b0;
    XRAM[2569] = 8'b0;
    XRAM[2570] = 8'b0;
    XRAM[2571] = 8'b0;
    XRAM[2572] = 8'b0;
    XRAM[2573] = 8'b0;
    XRAM[2574] = 8'b0;
    XRAM[2575] = 8'b0;
    XRAM[2576] = 8'b0;
    XRAM[2577] = 8'b0;
    XRAM[2578] = 8'b0;
    XRAM[2579] = 8'b0;
    XRAM[2580] = 8'b0;
    XRAM[2581] = 8'b0;
    XRAM[2582] = 8'b0;
    XRAM[2583] = 8'b0;
    XRAM[2584] = 8'b0;
    XRAM[2585] = 8'b0;
    XRAM[2586] = 8'b0;
    XRAM[2587] = 8'b0;
    XRAM[2588] = 8'b0;
    XRAM[2589] = 8'b0;
    XRAM[2590] = 8'b0;
    XRAM[2591] = 8'b0;
    XRAM[2592] = 8'b0;
    XRAM[2593] = 8'b0;
    XRAM[2594] = 8'b0;
    XRAM[2595] = 8'b0;
    XRAM[2596] = 8'b0;
    XRAM[2597] = 8'b0;
    XRAM[2598] = 8'b0;
    XRAM[2599] = 8'b0;
    XRAM[2600] = 8'b0;
    XRAM[2601] = 8'b0;
    XRAM[2602] = 8'b0;
    XRAM[2603] = 8'b0;
    XRAM[2604] = 8'b0;
    XRAM[2605] = 8'b0;
    XRAM[2606] = 8'b0;
    XRAM[2607] = 8'b0;
    XRAM[2608] = 8'b0;
    XRAM[2609] = 8'b0;
    XRAM[2610] = 8'b0;
    XRAM[2611] = 8'b0;
    XRAM[2612] = 8'b0;
    XRAM[2613] = 8'b0;
    XRAM[2614] = 8'b0;
    XRAM[2615] = 8'b0;
    XRAM[2616] = 8'b0;
    XRAM[2617] = 8'b0;
    XRAM[2618] = 8'b0;
    XRAM[2619] = 8'b0;
    XRAM[2620] = 8'b0;
    XRAM[2621] = 8'b0;
    XRAM[2622] = 8'b0;
    XRAM[2623] = 8'b0;
    XRAM[2624] = 8'b0;
    XRAM[2625] = 8'b0;
    XRAM[2626] = 8'b0;
    XRAM[2627] = 8'b0;
    XRAM[2628] = 8'b0;
    XRAM[2629] = 8'b0;
    XRAM[2630] = 8'b0;
    XRAM[2631] = 8'b0;
    XRAM[2632] = 8'b0;
    XRAM[2633] = 8'b0;
    XRAM[2634] = 8'b0;
    XRAM[2635] = 8'b0;
    XRAM[2636] = 8'b0;
    XRAM[2637] = 8'b0;
    XRAM[2638] = 8'b0;
    XRAM[2639] = 8'b0;
    XRAM[2640] = 8'b0;
    XRAM[2641] = 8'b0;
    XRAM[2642] = 8'b0;
    XRAM[2643] = 8'b0;
    XRAM[2644] = 8'b0;
    XRAM[2645] = 8'b0;
    XRAM[2646] = 8'b0;
    XRAM[2647] = 8'b0;
    XRAM[2648] = 8'b0;
    XRAM[2649] = 8'b0;
    XRAM[2650] = 8'b0;
    XRAM[2651] = 8'b0;
    XRAM[2652] = 8'b0;
    XRAM[2653] = 8'b0;
    XRAM[2654] = 8'b0;
    XRAM[2655] = 8'b0;
    XRAM[2656] = 8'b0;
    XRAM[2657] = 8'b0;
    XRAM[2658] = 8'b0;
    XRAM[2659] = 8'b0;
    XRAM[2660] = 8'b0;
    XRAM[2661] = 8'b0;
    XRAM[2662] = 8'b0;
    XRAM[2663] = 8'b0;
    XRAM[2664] = 8'b0;
    XRAM[2665] = 8'b0;
    XRAM[2666] = 8'b0;
    XRAM[2667] = 8'b0;
    XRAM[2668] = 8'b0;
    XRAM[2669] = 8'b0;
    XRAM[2670] = 8'b0;
    XRAM[2671] = 8'b0;
    XRAM[2672] = 8'b0;
    XRAM[2673] = 8'b0;
    XRAM[2674] = 8'b0;
    XRAM[2675] = 8'b0;
    XRAM[2676] = 8'b0;
    XRAM[2677] = 8'b0;
    XRAM[2678] = 8'b0;
    XRAM[2679] = 8'b0;
    XRAM[2680] = 8'b0;
    XRAM[2681] = 8'b0;
    XRAM[2682] = 8'b0;
    XRAM[2683] = 8'b0;
    XRAM[2684] = 8'b0;
    XRAM[2685] = 8'b0;
    XRAM[2686] = 8'b0;
    XRAM[2687] = 8'b0;
    XRAM[2688] = 8'b0;
    XRAM[2689] = 8'b0;
    XRAM[2690] = 8'b0;
    XRAM[2691] = 8'b0;
    XRAM[2692] = 8'b0;
    XRAM[2693] = 8'b0;
    XRAM[2694] = 8'b0;
    XRAM[2695] = 8'b0;
    XRAM[2696] = 8'b0;
    XRAM[2697] = 8'b0;
    XRAM[2698] = 8'b0;
    XRAM[2699] = 8'b0;
    XRAM[2700] = 8'b0;
    XRAM[2701] = 8'b0;
    XRAM[2702] = 8'b0;
    XRAM[2703] = 8'b0;
    XRAM[2704] = 8'b0;
    XRAM[2705] = 8'b0;
    XRAM[2706] = 8'b0;
    XRAM[2707] = 8'b0;
    XRAM[2708] = 8'b0;
    XRAM[2709] = 8'b0;
    XRAM[2710] = 8'b0;
    XRAM[2711] = 8'b0;
    XRAM[2712] = 8'b0;
    XRAM[2713] = 8'b0;
    XRAM[2714] = 8'b0;
    XRAM[2715] = 8'b0;
    XRAM[2716] = 8'b0;
    XRAM[2717] = 8'b0;
    XRAM[2718] = 8'b0;
    XRAM[2719] = 8'b0;
    XRAM[2720] = 8'b0;
    XRAM[2721] = 8'b0;
    XRAM[2722] = 8'b0;
    XRAM[2723] = 8'b0;
    XRAM[2724] = 8'b0;
    XRAM[2725] = 8'b0;
    XRAM[2726] = 8'b0;
    XRAM[2727] = 8'b0;
    XRAM[2728] = 8'b0;
    XRAM[2729] = 8'b0;
    XRAM[2730] = 8'b0;
    XRAM[2731] = 8'b0;
    XRAM[2732] = 8'b0;
    XRAM[2733] = 8'b0;
    XRAM[2734] = 8'b0;
    XRAM[2735] = 8'b0;
    XRAM[2736] = 8'b0;
    XRAM[2737] = 8'b0;
    XRAM[2738] = 8'b0;
    XRAM[2739] = 8'b0;
    XRAM[2740] = 8'b0;
    XRAM[2741] = 8'b0;
    XRAM[2742] = 8'b0;
    XRAM[2743] = 8'b0;
    XRAM[2744] = 8'b0;
    XRAM[2745] = 8'b0;
    XRAM[2746] = 8'b0;
    XRAM[2747] = 8'b0;
    XRAM[2748] = 8'b0;
    XRAM[2749] = 8'b0;
    XRAM[2750] = 8'b0;
    XRAM[2751] = 8'b0;
    XRAM[2752] = 8'b0;
    XRAM[2753] = 8'b0;
    XRAM[2754] = 8'b0;
    XRAM[2755] = 8'b0;
    XRAM[2756] = 8'b0;
    XRAM[2757] = 8'b0;
    XRAM[2758] = 8'b0;
    XRAM[2759] = 8'b0;
    XRAM[2760] = 8'b0;
    XRAM[2761] = 8'b0;
    XRAM[2762] = 8'b0;
    XRAM[2763] = 8'b0;
    XRAM[2764] = 8'b0;
    XRAM[2765] = 8'b0;
    XRAM[2766] = 8'b0;
    XRAM[2767] = 8'b0;
    XRAM[2768] = 8'b0;
    XRAM[2769] = 8'b0;
    XRAM[2770] = 8'b0;
    XRAM[2771] = 8'b0;
    XRAM[2772] = 8'b0;
    XRAM[2773] = 8'b0;
    XRAM[2774] = 8'b0;
    XRAM[2775] = 8'b0;
    XRAM[2776] = 8'b0;
    XRAM[2777] = 8'b0;
    XRAM[2778] = 8'b0;
    XRAM[2779] = 8'b0;
    XRAM[2780] = 8'b0;
    XRAM[2781] = 8'b0;
    XRAM[2782] = 8'b0;
    XRAM[2783] = 8'b0;
    XRAM[2784] = 8'b0;
    XRAM[2785] = 8'b0;
    XRAM[2786] = 8'b0;
    XRAM[2787] = 8'b0;
    XRAM[2788] = 8'b0;
    XRAM[2789] = 8'b0;
    XRAM[2790] = 8'b0;
    XRAM[2791] = 8'b0;
    XRAM[2792] = 8'b0;
    XRAM[2793] = 8'b0;
    XRAM[2794] = 8'b0;
    XRAM[2795] = 8'b0;
    XRAM[2796] = 8'b0;
    XRAM[2797] = 8'b0;
    XRAM[2798] = 8'b0;
    XRAM[2799] = 8'b0;
    XRAM[2800] = 8'b0;
    XRAM[2801] = 8'b0;
    XRAM[2802] = 8'b0;
    XRAM[2803] = 8'b0;
    XRAM[2804] = 8'b0;
    XRAM[2805] = 8'b0;
    XRAM[2806] = 8'b0;
    XRAM[2807] = 8'b0;
    XRAM[2808] = 8'b0;
    XRAM[2809] = 8'b0;
    XRAM[2810] = 8'b0;
    XRAM[2811] = 8'b0;
    XRAM[2812] = 8'b0;
    XRAM[2813] = 8'b0;
    XRAM[2814] = 8'b0;
    XRAM[2815] = 8'b0;
    XRAM[2816] = 8'b0;
    XRAM[2817] = 8'b0;
    XRAM[2818] = 8'b0;
    XRAM[2819] = 8'b0;
    XRAM[2820] = 8'b0;
    XRAM[2821] = 8'b0;
    XRAM[2822] = 8'b0;
    XRAM[2823] = 8'b0;
    XRAM[2824] = 8'b0;
    XRAM[2825] = 8'b0;
    XRAM[2826] = 8'b0;
    XRAM[2827] = 8'b0;
    XRAM[2828] = 8'b0;
    XRAM[2829] = 8'b0;
    XRAM[2830] = 8'b0;
    XRAM[2831] = 8'b0;
    XRAM[2832] = 8'b0;
    XRAM[2833] = 8'b0;
    XRAM[2834] = 8'b0;
    XRAM[2835] = 8'b0;
    XRAM[2836] = 8'b0;
    XRAM[2837] = 8'b0;
    XRAM[2838] = 8'b0;
    XRAM[2839] = 8'b0;
    XRAM[2840] = 8'b0;
    XRAM[2841] = 8'b0;
    XRAM[2842] = 8'b0;
    XRAM[2843] = 8'b0;
    XRAM[2844] = 8'b0;
    XRAM[2845] = 8'b0;
    XRAM[2846] = 8'b0;
    XRAM[2847] = 8'b0;
    XRAM[2848] = 8'b0;
    XRAM[2849] = 8'b0;
    XRAM[2850] = 8'b0;
    XRAM[2851] = 8'b0;
    XRAM[2852] = 8'b0;
    XRAM[2853] = 8'b0;
    XRAM[2854] = 8'b0;
    XRAM[2855] = 8'b0;
    XRAM[2856] = 8'b0;
    XRAM[2857] = 8'b0;
    XRAM[2858] = 8'b0;
    XRAM[2859] = 8'b0;
    XRAM[2860] = 8'b0;
    XRAM[2861] = 8'b0;
    XRAM[2862] = 8'b0;
    XRAM[2863] = 8'b0;
    XRAM[2864] = 8'b0;
    XRAM[2865] = 8'b0;
    XRAM[2866] = 8'b0;
    XRAM[2867] = 8'b0;
    XRAM[2868] = 8'b0;
    XRAM[2869] = 8'b0;
    XRAM[2870] = 8'b0;
    XRAM[2871] = 8'b0;
    XRAM[2872] = 8'b0;
    XRAM[2873] = 8'b0;
    XRAM[2874] = 8'b0;
    XRAM[2875] = 8'b0;
    XRAM[2876] = 8'b0;
    XRAM[2877] = 8'b0;
    XRAM[2878] = 8'b0;
    XRAM[2879] = 8'b0;
    XRAM[2880] = 8'b0;
    XRAM[2881] = 8'b0;
    XRAM[2882] = 8'b0;
    XRAM[2883] = 8'b0;
    XRAM[2884] = 8'b0;
    XRAM[2885] = 8'b0;
    XRAM[2886] = 8'b0;
    XRAM[2887] = 8'b0;
    XRAM[2888] = 8'b0;
    XRAM[2889] = 8'b0;
    XRAM[2890] = 8'b0;
    XRAM[2891] = 8'b0;
    XRAM[2892] = 8'b0;
    XRAM[2893] = 8'b0;
    XRAM[2894] = 8'b0;
    XRAM[2895] = 8'b0;
    XRAM[2896] = 8'b0;
    XRAM[2897] = 8'b0;
    XRAM[2898] = 8'b0;
    XRAM[2899] = 8'b0;
    XRAM[2900] = 8'b0;
    XRAM[2901] = 8'b0;
    XRAM[2902] = 8'b0;
    XRAM[2903] = 8'b0;
    XRAM[2904] = 8'b0;
    XRAM[2905] = 8'b0;
    XRAM[2906] = 8'b0;
    XRAM[2907] = 8'b0;
    XRAM[2908] = 8'b0;
    XRAM[2909] = 8'b0;
    XRAM[2910] = 8'b0;
    XRAM[2911] = 8'b0;
    XRAM[2912] = 8'b0;
    XRAM[2913] = 8'b0;
    XRAM[2914] = 8'b0;
    XRAM[2915] = 8'b0;
    XRAM[2916] = 8'b0;
    XRAM[2917] = 8'b0;
    XRAM[2918] = 8'b0;
    XRAM[2919] = 8'b0;
    XRAM[2920] = 8'b0;
    XRAM[2921] = 8'b0;
    XRAM[2922] = 8'b0;
    XRAM[2923] = 8'b0;
    XRAM[2924] = 8'b0;
    XRAM[2925] = 8'b0;
    XRAM[2926] = 8'b0;
    XRAM[2927] = 8'b0;
    XRAM[2928] = 8'b0;
    XRAM[2929] = 8'b0;
    XRAM[2930] = 8'b0;
    XRAM[2931] = 8'b0;
    XRAM[2932] = 8'b0;
    XRAM[2933] = 8'b0;
    XRAM[2934] = 8'b0;
    XRAM[2935] = 8'b0;
    XRAM[2936] = 8'b0;
    XRAM[2937] = 8'b0;
    XRAM[2938] = 8'b0;
    XRAM[2939] = 8'b0;
    XRAM[2940] = 8'b0;
    XRAM[2941] = 8'b0;
    XRAM[2942] = 8'b0;
    XRAM[2943] = 8'b0;
    XRAM[2944] = 8'b0;
    XRAM[2945] = 8'b0;
    XRAM[2946] = 8'b0;
    XRAM[2947] = 8'b0;
    XRAM[2948] = 8'b0;
    XRAM[2949] = 8'b0;
    XRAM[2950] = 8'b0;
    XRAM[2951] = 8'b0;
    XRAM[2952] = 8'b0;
    XRAM[2953] = 8'b0;
    XRAM[2954] = 8'b0;
    XRAM[2955] = 8'b0;
    XRAM[2956] = 8'b0;
    XRAM[2957] = 8'b0;
    XRAM[2958] = 8'b0;
    XRAM[2959] = 8'b0;
    XRAM[2960] = 8'b0;
    XRAM[2961] = 8'b0;
    XRAM[2962] = 8'b0;
    XRAM[2963] = 8'b0;
    XRAM[2964] = 8'b0;
    XRAM[2965] = 8'b0;
    XRAM[2966] = 8'b0;
    XRAM[2967] = 8'b0;
    XRAM[2968] = 8'b0;
    XRAM[2969] = 8'b0;
    XRAM[2970] = 8'b0;
    XRAM[2971] = 8'b0;
    XRAM[2972] = 8'b0;
    XRAM[2973] = 8'b0;
    XRAM[2974] = 8'b0;
    XRAM[2975] = 8'b0;
    XRAM[2976] = 8'b0;
    XRAM[2977] = 8'b0;
    XRAM[2978] = 8'b0;
    XRAM[2979] = 8'b0;
    XRAM[2980] = 8'b0;
    XRAM[2981] = 8'b0;
    XRAM[2982] = 8'b0;
    XRAM[2983] = 8'b0;
    XRAM[2984] = 8'b0;
    XRAM[2985] = 8'b0;
    XRAM[2986] = 8'b0;
    XRAM[2987] = 8'b0;
    XRAM[2988] = 8'b0;
    XRAM[2989] = 8'b0;
    XRAM[2990] = 8'b0;
    XRAM[2991] = 8'b0;
    XRAM[2992] = 8'b0;
    XRAM[2993] = 8'b0;
    XRAM[2994] = 8'b0;
    XRAM[2995] = 8'b0;
    XRAM[2996] = 8'b0;
    XRAM[2997] = 8'b0;
    XRAM[2998] = 8'b0;
    XRAM[2999] = 8'b0;
    XRAM[3000] = 8'b0;
    XRAM[3001] = 8'b0;
    XRAM[3002] = 8'b0;
    XRAM[3003] = 8'b0;
    XRAM[3004] = 8'b0;
    XRAM[3005] = 8'b0;
    XRAM[3006] = 8'b0;
    XRAM[3007] = 8'b0;
    XRAM[3008] = 8'b0;
    XRAM[3009] = 8'b0;
    XRAM[3010] = 8'b0;
    XRAM[3011] = 8'b0;
    XRAM[3012] = 8'b0;
    XRAM[3013] = 8'b0;
    XRAM[3014] = 8'b0;
    XRAM[3015] = 8'b0;
    XRAM[3016] = 8'b0;
    XRAM[3017] = 8'b0;
    XRAM[3018] = 8'b0;
    XRAM[3019] = 8'b0;
    XRAM[3020] = 8'b0;
    XRAM[3021] = 8'b0;
    XRAM[3022] = 8'b0;
    XRAM[3023] = 8'b0;
    XRAM[3024] = 8'b0;
    XRAM[3025] = 8'b0;
    XRAM[3026] = 8'b0;
    XRAM[3027] = 8'b0;
    XRAM[3028] = 8'b0;
    XRAM[3029] = 8'b0;
    XRAM[3030] = 8'b0;
    XRAM[3031] = 8'b0;
    XRAM[3032] = 8'b0;
    XRAM[3033] = 8'b0;
    XRAM[3034] = 8'b0;
    XRAM[3035] = 8'b0;
    XRAM[3036] = 8'b0;
    XRAM[3037] = 8'b0;
    XRAM[3038] = 8'b0;
    XRAM[3039] = 8'b0;
    XRAM[3040] = 8'b0;
    XRAM[3041] = 8'b0;
    XRAM[3042] = 8'b0;
    XRAM[3043] = 8'b0;
    XRAM[3044] = 8'b0;
    XRAM[3045] = 8'b0;
    XRAM[3046] = 8'b0;
    XRAM[3047] = 8'b0;
    XRAM[3048] = 8'b0;
    XRAM[3049] = 8'b0;
    XRAM[3050] = 8'b0;
    XRAM[3051] = 8'b0;
    XRAM[3052] = 8'b0;
    XRAM[3053] = 8'b0;
    XRAM[3054] = 8'b0;
    XRAM[3055] = 8'b0;
    XRAM[3056] = 8'b0;
    XRAM[3057] = 8'b0;
    XRAM[3058] = 8'b0;
    XRAM[3059] = 8'b0;
    XRAM[3060] = 8'b0;
    XRAM[3061] = 8'b0;
    XRAM[3062] = 8'b0;
    XRAM[3063] = 8'b0;
    XRAM[3064] = 8'b0;
    XRAM[3065] = 8'b0;
    XRAM[3066] = 8'b0;
    XRAM[3067] = 8'b0;
    XRAM[3068] = 8'b0;
    XRAM[3069] = 8'b0;
    XRAM[3070] = 8'b0;
    XRAM[3071] = 8'b0;
    XRAM[3072] = 8'b0;
    XRAM[3073] = 8'b0;
    XRAM[3074] = 8'b0;
    XRAM[3075] = 8'b0;
    XRAM[3076] = 8'b0;
    XRAM[3077] = 8'b0;
    XRAM[3078] = 8'b0;
    XRAM[3079] = 8'b0;
    XRAM[3080] = 8'b0;
    XRAM[3081] = 8'b0;
    XRAM[3082] = 8'b0;
    XRAM[3083] = 8'b0;
    XRAM[3084] = 8'b0;
    XRAM[3085] = 8'b0;
    XRAM[3086] = 8'b0;
    XRAM[3087] = 8'b0;
    XRAM[3088] = 8'b0;
    XRAM[3089] = 8'b0;
    XRAM[3090] = 8'b0;
    XRAM[3091] = 8'b0;
    XRAM[3092] = 8'b0;
    XRAM[3093] = 8'b0;
    XRAM[3094] = 8'b0;
    XRAM[3095] = 8'b0;
    XRAM[3096] = 8'b0;
    XRAM[3097] = 8'b0;
    XRAM[3098] = 8'b0;
    XRAM[3099] = 8'b0;
    XRAM[3100] = 8'b0;
    XRAM[3101] = 8'b0;
    XRAM[3102] = 8'b0;
    XRAM[3103] = 8'b0;
    XRAM[3104] = 8'b0;
    XRAM[3105] = 8'b0;
    XRAM[3106] = 8'b0;
    XRAM[3107] = 8'b0;
    XRAM[3108] = 8'b0;
    XRAM[3109] = 8'b0;
    XRAM[3110] = 8'b0;
    XRAM[3111] = 8'b0;
    XRAM[3112] = 8'b0;
    XRAM[3113] = 8'b0;
    XRAM[3114] = 8'b0;
    XRAM[3115] = 8'b0;
    XRAM[3116] = 8'b0;
    XRAM[3117] = 8'b0;
    XRAM[3118] = 8'b0;
    XRAM[3119] = 8'b0;
    XRAM[3120] = 8'b0;
    XRAM[3121] = 8'b0;
    XRAM[3122] = 8'b0;
    XRAM[3123] = 8'b0;
    XRAM[3124] = 8'b0;
    XRAM[3125] = 8'b0;
    XRAM[3126] = 8'b0;
    XRAM[3127] = 8'b0;
    XRAM[3128] = 8'b0;
    XRAM[3129] = 8'b0;
    XRAM[3130] = 8'b0;
    XRAM[3131] = 8'b0;
    XRAM[3132] = 8'b0;
    XRAM[3133] = 8'b0;
    XRAM[3134] = 8'b0;
    XRAM[3135] = 8'b0;
    XRAM[3136] = 8'b0;
    XRAM[3137] = 8'b0;
    XRAM[3138] = 8'b0;
    XRAM[3139] = 8'b0;
    XRAM[3140] = 8'b0;
    XRAM[3141] = 8'b0;
    XRAM[3142] = 8'b0;
    XRAM[3143] = 8'b0;
    XRAM[3144] = 8'b0;
    XRAM[3145] = 8'b0;
    XRAM[3146] = 8'b0;
    XRAM[3147] = 8'b0;
    XRAM[3148] = 8'b0;
    XRAM[3149] = 8'b0;
    XRAM[3150] = 8'b0;
    XRAM[3151] = 8'b0;
    XRAM[3152] = 8'b0;
    XRAM[3153] = 8'b0;
    XRAM[3154] = 8'b0;
    XRAM[3155] = 8'b0;
    XRAM[3156] = 8'b0;
    XRAM[3157] = 8'b0;
    XRAM[3158] = 8'b0;
    XRAM[3159] = 8'b0;
    XRAM[3160] = 8'b0;
    XRAM[3161] = 8'b0;
    XRAM[3162] = 8'b0;
    XRAM[3163] = 8'b0;
    XRAM[3164] = 8'b0;
    XRAM[3165] = 8'b0;
    XRAM[3166] = 8'b0;
    XRAM[3167] = 8'b0;
    XRAM[3168] = 8'b0;
    XRAM[3169] = 8'b0;
    XRAM[3170] = 8'b0;
    XRAM[3171] = 8'b0;
    XRAM[3172] = 8'b0;
    XRAM[3173] = 8'b0;
    XRAM[3174] = 8'b0;
    XRAM[3175] = 8'b0;
    XRAM[3176] = 8'b0;
    XRAM[3177] = 8'b0;
    XRAM[3178] = 8'b0;
    XRAM[3179] = 8'b0;
    XRAM[3180] = 8'b0;
    XRAM[3181] = 8'b0;
    XRAM[3182] = 8'b0;
    XRAM[3183] = 8'b0;
    XRAM[3184] = 8'b0;
    XRAM[3185] = 8'b0;
    XRAM[3186] = 8'b0;
    XRAM[3187] = 8'b0;
    XRAM[3188] = 8'b0;
    XRAM[3189] = 8'b0;
    XRAM[3190] = 8'b0;
    XRAM[3191] = 8'b0;
    XRAM[3192] = 8'b0;
    XRAM[3193] = 8'b0;
    XRAM[3194] = 8'b0;
    XRAM[3195] = 8'b0;
    XRAM[3196] = 8'b0;
    XRAM[3197] = 8'b0;
    XRAM[3198] = 8'b0;
    XRAM[3199] = 8'b0;
    XRAM[3200] = 8'b0;
    XRAM[3201] = 8'b0;
    XRAM[3202] = 8'b0;
    XRAM[3203] = 8'b0;
    XRAM[3204] = 8'b0;
    XRAM[3205] = 8'b0;
    XRAM[3206] = 8'b0;
    XRAM[3207] = 8'b0;
    XRAM[3208] = 8'b0;
    XRAM[3209] = 8'b0;
    XRAM[3210] = 8'b0;
    XRAM[3211] = 8'b0;
    XRAM[3212] = 8'b0;
    XRAM[3213] = 8'b0;
    XRAM[3214] = 8'b0;
    XRAM[3215] = 8'b0;
    XRAM[3216] = 8'b0;
    XRAM[3217] = 8'b0;
    XRAM[3218] = 8'b0;
    XRAM[3219] = 8'b0;
    XRAM[3220] = 8'b0;
    XRAM[3221] = 8'b0;
    XRAM[3222] = 8'b0;
    XRAM[3223] = 8'b0;
    XRAM[3224] = 8'b0;
    XRAM[3225] = 8'b0;
    XRAM[3226] = 8'b0;
    XRAM[3227] = 8'b0;
    XRAM[3228] = 8'b0;
    XRAM[3229] = 8'b0;
    XRAM[3230] = 8'b0;
    XRAM[3231] = 8'b0;
    XRAM[3232] = 8'b0;
    XRAM[3233] = 8'b0;
    XRAM[3234] = 8'b0;
    XRAM[3235] = 8'b0;
    XRAM[3236] = 8'b0;
    XRAM[3237] = 8'b0;
    XRAM[3238] = 8'b0;
    XRAM[3239] = 8'b0;
    XRAM[3240] = 8'b0;
    XRAM[3241] = 8'b0;
    XRAM[3242] = 8'b0;
    XRAM[3243] = 8'b0;
    XRAM[3244] = 8'b0;
    XRAM[3245] = 8'b0;
    XRAM[3246] = 8'b0;
    XRAM[3247] = 8'b0;
    XRAM[3248] = 8'b0;
    XRAM[3249] = 8'b0;
    XRAM[3250] = 8'b0;
    XRAM[3251] = 8'b0;
    XRAM[3252] = 8'b0;
    XRAM[3253] = 8'b0;
    XRAM[3254] = 8'b0;
    XRAM[3255] = 8'b0;
    XRAM[3256] = 8'b0;
    XRAM[3257] = 8'b0;
    XRAM[3258] = 8'b0;
    XRAM[3259] = 8'b0;
    XRAM[3260] = 8'b0;
    XRAM[3261] = 8'b0;
    XRAM[3262] = 8'b0;
    XRAM[3263] = 8'b0;
    XRAM[3264] = 8'b0;
    XRAM[3265] = 8'b0;
    XRAM[3266] = 8'b0;
    XRAM[3267] = 8'b0;
    XRAM[3268] = 8'b0;
    XRAM[3269] = 8'b0;
    XRAM[3270] = 8'b0;
    XRAM[3271] = 8'b0;
    XRAM[3272] = 8'b0;
    XRAM[3273] = 8'b0;
    XRAM[3274] = 8'b0;
    XRAM[3275] = 8'b0;
    XRAM[3276] = 8'b0;
    XRAM[3277] = 8'b0;
    XRAM[3278] = 8'b0;
    XRAM[3279] = 8'b0;
    XRAM[3280] = 8'b0;
    XRAM[3281] = 8'b0;
    XRAM[3282] = 8'b0;
    XRAM[3283] = 8'b0;
    XRAM[3284] = 8'b0;
    XRAM[3285] = 8'b0;
    XRAM[3286] = 8'b0;
    XRAM[3287] = 8'b0;
    XRAM[3288] = 8'b0;
    XRAM[3289] = 8'b0;
    XRAM[3290] = 8'b0;
    XRAM[3291] = 8'b0;
    XRAM[3292] = 8'b0;
    XRAM[3293] = 8'b0;
    XRAM[3294] = 8'b0;
    XRAM[3295] = 8'b0;
    XRAM[3296] = 8'b0;
    XRAM[3297] = 8'b0;
    XRAM[3298] = 8'b0;
    XRAM[3299] = 8'b0;
    XRAM[3300] = 8'b0;
    XRAM[3301] = 8'b0;
    XRAM[3302] = 8'b0;
    XRAM[3303] = 8'b0;
    XRAM[3304] = 8'b0;
    XRAM[3305] = 8'b0;
    XRAM[3306] = 8'b0;
    XRAM[3307] = 8'b0;
    XRAM[3308] = 8'b0;
    XRAM[3309] = 8'b0;
    XRAM[3310] = 8'b0;
    XRAM[3311] = 8'b0;
    XRAM[3312] = 8'b0;
    XRAM[3313] = 8'b0;
    XRAM[3314] = 8'b0;
    XRAM[3315] = 8'b0;
    XRAM[3316] = 8'b0;
    XRAM[3317] = 8'b0;
    XRAM[3318] = 8'b0;
    XRAM[3319] = 8'b0;
    XRAM[3320] = 8'b0;
    XRAM[3321] = 8'b0;
    XRAM[3322] = 8'b0;
    XRAM[3323] = 8'b0;
    XRAM[3324] = 8'b0;
    XRAM[3325] = 8'b0;
    XRAM[3326] = 8'b0;
    XRAM[3327] = 8'b0;
    XRAM[3328] = 8'b0;
    XRAM[3329] = 8'b0;
    XRAM[3330] = 8'b0;
    XRAM[3331] = 8'b0;
    XRAM[3332] = 8'b0;
    XRAM[3333] = 8'b0;
    XRAM[3334] = 8'b0;
    XRAM[3335] = 8'b0;
    XRAM[3336] = 8'b0;
    XRAM[3337] = 8'b0;
    XRAM[3338] = 8'b0;
    XRAM[3339] = 8'b0;
    XRAM[3340] = 8'b0;
    XRAM[3341] = 8'b0;
    XRAM[3342] = 8'b0;
    XRAM[3343] = 8'b0;
    XRAM[3344] = 8'b0;
    XRAM[3345] = 8'b0;
    XRAM[3346] = 8'b0;
    XRAM[3347] = 8'b0;
    XRAM[3348] = 8'b0;
    XRAM[3349] = 8'b0;
    XRAM[3350] = 8'b0;
    XRAM[3351] = 8'b0;
    XRAM[3352] = 8'b0;
    XRAM[3353] = 8'b0;
    XRAM[3354] = 8'b0;
    XRAM[3355] = 8'b0;
    XRAM[3356] = 8'b0;
    XRAM[3357] = 8'b0;
    XRAM[3358] = 8'b0;
    XRAM[3359] = 8'b0;
    XRAM[3360] = 8'b0;
    XRAM[3361] = 8'b0;
    XRAM[3362] = 8'b0;
    XRAM[3363] = 8'b0;
    XRAM[3364] = 8'b0;
    XRAM[3365] = 8'b0;
    XRAM[3366] = 8'b0;
    XRAM[3367] = 8'b0;
    XRAM[3368] = 8'b0;
    XRAM[3369] = 8'b0;
    XRAM[3370] = 8'b0;
    XRAM[3371] = 8'b0;
    XRAM[3372] = 8'b0;
    XRAM[3373] = 8'b0;
    XRAM[3374] = 8'b0;
    XRAM[3375] = 8'b0;
    XRAM[3376] = 8'b0;
    XRAM[3377] = 8'b0;
    XRAM[3378] = 8'b0;
    XRAM[3379] = 8'b0;
    XRAM[3380] = 8'b0;
    XRAM[3381] = 8'b0;
    XRAM[3382] = 8'b0;
    XRAM[3383] = 8'b0;
    XRAM[3384] = 8'b0;
    XRAM[3385] = 8'b0;
    XRAM[3386] = 8'b0;
    XRAM[3387] = 8'b0;
    XRAM[3388] = 8'b0;
    XRAM[3389] = 8'b0;
    XRAM[3390] = 8'b0;
    XRAM[3391] = 8'b0;
    XRAM[3392] = 8'b0;
    XRAM[3393] = 8'b0;
    XRAM[3394] = 8'b0;
    XRAM[3395] = 8'b0;
    XRAM[3396] = 8'b0;
    XRAM[3397] = 8'b0;
    XRAM[3398] = 8'b0;
    XRAM[3399] = 8'b0;
    XRAM[3400] = 8'b0;
    XRAM[3401] = 8'b0;
    XRAM[3402] = 8'b0;
    XRAM[3403] = 8'b0;
    XRAM[3404] = 8'b0;
    XRAM[3405] = 8'b0;
    XRAM[3406] = 8'b0;
    XRAM[3407] = 8'b0;
    XRAM[3408] = 8'b0;
    XRAM[3409] = 8'b0;
    XRAM[3410] = 8'b0;
    XRAM[3411] = 8'b0;
    XRAM[3412] = 8'b0;
    XRAM[3413] = 8'b0;
    XRAM[3414] = 8'b0;
    XRAM[3415] = 8'b0;
    XRAM[3416] = 8'b0;
    XRAM[3417] = 8'b0;
    XRAM[3418] = 8'b0;
    XRAM[3419] = 8'b0;
    XRAM[3420] = 8'b0;
    XRAM[3421] = 8'b0;
    XRAM[3422] = 8'b0;
    XRAM[3423] = 8'b0;
    XRAM[3424] = 8'b0;
    XRAM[3425] = 8'b0;
    XRAM[3426] = 8'b0;
    XRAM[3427] = 8'b0;
    XRAM[3428] = 8'b0;
    XRAM[3429] = 8'b0;
    XRAM[3430] = 8'b0;
    XRAM[3431] = 8'b0;
    XRAM[3432] = 8'b0;
    XRAM[3433] = 8'b0;
    XRAM[3434] = 8'b0;
    XRAM[3435] = 8'b0;
    XRAM[3436] = 8'b0;
    XRAM[3437] = 8'b0;
    XRAM[3438] = 8'b0;
    XRAM[3439] = 8'b0;
    XRAM[3440] = 8'b0;
    XRAM[3441] = 8'b0;
    XRAM[3442] = 8'b0;
    XRAM[3443] = 8'b0;
    XRAM[3444] = 8'b0;
    XRAM[3445] = 8'b0;
    XRAM[3446] = 8'b0;
    XRAM[3447] = 8'b0;
    XRAM[3448] = 8'b0;
    XRAM[3449] = 8'b0;
    XRAM[3450] = 8'b0;
    XRAM[3451] = 8'b0;
    XRAM[3452] = 8'b0;
    XRAM[3453] = 8'b0;
    XRAM[3454] = 8'b0;
    XRAM[3455] = 8'b0;
    XRAM[3456] = 8'b0;
    XRAM[3457] = 8'b0;
    XRAM[3458] = 8'b0;
    XRAM[3459] = 8'b0;
    XRAM[3460] = 8'b0;
    XRAM[3461] = 8'b0;
    XRAM[3462] = 8'b0;
    XRAM[3463] = 8'b0;
    XRAM[3464] = 8'b0;
    XRAM[3465] = 8'b0;
    XRAM[3466] = 8'b0;
    XRAM[3467] = 8'b0;
    XRAM[3468] = 8'b0;
    XRAM[3469] = 8'b0;
    XRAM[3470] = 8'b0;
    XRAM[3471] = 8'b0;
    XRAM[3472] = 8'b0;
    XRAM[3473] = 8'b0;
    XRAM[3474] = 8'b0;
    XRAM[3475] = 8'b0;
    XRAM[3476] = 8'b0;
    XRAM[3477] = 8'b0;
    XRAM[3478] = 8'b0;
    XRAM[3479] = 8'b0;
    XRAM[3480] = 8'b0;
    XRAM[3481] = 8'b0;
    XRAM[3482] = 8'b0;
    XRAM[3483] = 8'b0;
    XRAM[3484] = 8'b0;
    XRAM[3485] = 8'b0;
    XRAM[3486] = 8'b0;
    XRAM[3487] = 8'b0;
    XRAM[3488] = 8'b0;
    XRAM[3489] = 8'b0;
    XRAM[3490] = 8'b0;
    XRAM[3491] = 8'b0;
    XRAM[3492] = 8'b0;
    XRAM[3493] = 8'b0;
    XRAM[3494] = 8'b0;
    XRAM[3495] = 8'b0;
    XRAM[3496] = 8'b0;
    XRAM[3497] = 8'b0;
    XRAM[3498] = 8'b0;
    XRAM[3499] = 8'b0;
    XRAM[3500] = 8'b0;
    XRAM[3501] = 8'b0;
    XRAM[3502] = 8'b0;
    XRAM[3503] = 8'b0;
    XRAM[3504] = 8'b0;
    XRAM[3505] = 8'b0;
    XRAM[3506] = 8'b0;
    XRAM[3507] = 8'b0;
    XRAM[3508] = 8'b0;
    XRAM[3509] = 8'b0;
    XRAM[3510] = 8'b0;
    XRAM[3511] = 8'b0;
    XRAM[3512] = 8'b0;
    XRAM[3513] = 8'b0;
    XRAM[3514] = 8'b0;
    XRAM[3515] = 8'b0;
    XRAM[3516] = 8'b0;
    XRAM[3517] = 8'b0;
    XRAM[3518] = 8'b0;
    XRAM[3519] = 8'b0;
    XRAM[3520] = 8'b0;
    XRAM[3521] = 8'b0;
    XRAM[3522] = 8'b0;
    XRAM[3523] = 8'b0;
    XRAM[3524] = 8'b0;
    XRAM[3525] = 8'b0;
    XRAM[3526] = 8'b0;
    XRAM[3527] = 8'b0;
    XRAM[3528] = 8'b0;
    XRAM[3529] = 8'b0;
    XRAM[3530] = 8'b0;
    XRAM[3531] = 8'b0;
    XRAM[3532] = 8'b0;
    XRAM[3533] = 8'b0;
    XRAM[3534] = 8'b0;
    XRAM[3535] = 8'b0;
    XRAM[3536] = 8'b0;
    XRAM[3537] = 8'b0;
    XRAM[3538] = 8'b0;
    XRAM[3539] = 8'b0;
    XRAM[3540] = 8'b0;
    XRAM[3541] = 8'b0;
    XRAM[3542] = 8'b0;
    XRAM[3543] = 8'b0;
    XRAM[3544] = 8'b0;
    XRAM[3545] = 8'b0;
    XRAM[3546] = 8'b0;
    XRAM[3547] = 8'b0;
    XRAM[3548] = 8'b0;
    XRAM[3549] = 8'b0;
    XRAM[3550] = 8'b0;
    XRAM[3551] = 8'b0;
    XRAM[3552] = 8'b0;
    XRAM[3553] = 8'b0;
    XRAM[3554] = 8'b0;
    XRAM[3555] = 8'b0;
    XRAM[3556] = 8'b0;
    XRAM[3557] = 8'b0;
    XRAM[3558] = 8'b0;
    XRAM[3559] = 8'b0;
    XRAM[3560] = 8'b0;
    XRAM[3561] = 8'b0;
    XRAM[3562] = 8'b0;
    XRAM[3563] = 8'b0;
    XRAM[3564] = 8'b0;
    XRAM[3565] = 8'b0;
    XRAM[3566] = 8'b0;
    XRAM[3567] = 8'b0;
    XRAM[3568] = 8'b0;
    XRAM[3569] = 8'b0;
    XRAM[3570] = 8'b0;
    XRAM[3571] = 8'b0;
    XRAM[3572] = 8'b0;
    XRAM[3573] = 8'b0;
    XRAM[3574] = 8'b0;
    XRAM[3575] = 8'b0;
    XRAM[3576] = 8'b0;
    XRAM[3577] = 8'b0;
    XRAM[3578] = 8'b0;
    XRAM[3579] = 8'b0;
    XRAM[3580] = 8'b0;
    XRAM[3581] = 8'b0;
    XRAM[3582] = 8'b0;
    XRAM[3583] = 8'b0;
    XRAM[3584] = 8'b0;
    XRAM[3585] = 8'b0;
    XRAM[3586] = 8'b0;
    XRAM[3587] = 8'b0;
    XRAM[3588] = 8'b0;
    XRAM[3589] = 8'b0;
    XRAM[3590] = 8'b0;
    XRAM[3591] = 8'b0;
    XRAM[3592] = 8'b0;
    XRAM[3593] = 8'b0;
    XRAM[3594] = 8'b0;
    XRAM[3595] = 8'b0;
    XRAM[3596] = 8'b0;
    XRAM[3597] = 8'b0;
    XRAM[3598] = 8'b0;
    XRAM[3599] = 8'b0;
    XRAM[3600] = 8'b0;
    XRAM[3601] = 8'b0;
    XRAM[3602] = 8'b0;
    XRAM[3603] = 8'b0;
    XRAM[3604] = 8'b0;
    XRAM[3605] = 8'b0;
    XRAM[3606] = 8'b0;
    XRAM[3607] = 8'b0;
    XRAM[3608] = 8'b0;
    XRAM[3609] = 8'b0;
    XRAM[3610] = 8'b0;
    XRAM[3611] = 8'b0;
    XRAM[3612] = 8'b0;
    XRAM[3613] = 8'b0;
    XRAM[3614] = 8'b0;
    XRAM[3615] = 8'b0;
    XRAM[3616] = 8'b0;
    XRAM[3617] = 8'b0;
    XRAM[3618] = 8'b0;
    XRAM[3619] = 8'b0;
    XRAM[3620] = 8'b0;
    XRAM[3621] = 8'b0;
    XRAM[3622] = 8'b0;
    XRAM[3623] = 8'b0;
    XRAM[3624] = 8'b0;
    XRAM[3625] = 8'b0;
    XRAM[3626] = 8'b0;
    XRAM[3627] = 8'b0;
    XRAM[3628] = 8'b0;
    XRAM[3629] = 8'b0;
    XRAM[3630] = 8'b0;
    XRAM[3631] = 8'b0;
    XRAM[3632] = 8'b0;
    XRAM[3633] = 8'b0;
    XRAM[3634] = 8'b0;
    XRAM[3635] = 8'b0;
    XRAM[3636] = 8'b0;
    XRAM[3637] = 8'b0;
    XRAM[3638] = 8'b0;
    XRAM[3639] = 8'b0;
    XRAM[3640] = 8'b0;
    XRAM[3641] = 8'b0;
    XRAM[3642] = 8'b0;
    XRAM[3643] = 8'b0;
    XRAM[3644] = 8'b0;
    XRAM[3645] = 8'b0;
    XRAM[3646] = 8'b0;
    XRAM[3647] = 8'b0;
    XRAM[3648] = 8'b0;
    XRAM[3649] = 8'b0;
    XRAM[3650] = 8'b0;
    XRAM[3651] = 8'b0;
    XRAM[3652] = 8'b0;
    XRAM[3653] = 8'b0;
    XRAM[3654] = 8'b0;
    XRAM[3655] = 8'b0;
    XRAM[3656] = 8'b0;
    XRAM[3657] = 8'b0;
    XRAM[3658] = 8'b0;
    XRAM[3659] = 8'b0;
    XRAM[3660] = 8'b0;
    XRAM[3661] = 8'b0;
    XRAM[3662] = 8'b0;
    XRAM[3663] = 8'b0;
    XRAM[3664] = 8'b0;
    XRAM[3665] = 8'b0;
    XRAM[3666] = 8'b0;
    XRAM[3667] = 8'b0;
    XRAM[3668] = 8'b0;
    XRAM[3669] = 8'b0;
    XRAM[3670] = 8'b0;
    XRAM[3671] = 8'b0;
    XRAM[3672] = 8'b0;
    XRAM[3673] = 8'b0;
    XRAM[3674] = 8'b0;
    XRAM[3675] = 8'b0;
    XRAM[3676] = 8'b0;
    XRAM[3677] = 8'b0;
    XRAM[3678] = 8'b0;
    XRAM[3679] = 8'b0;
    XRAM[3680] = 8'b0;
    XRAM[3681] = 8'b0;
    XRAM[3682] = 8'b0;
    XRAM[3683] = 8'b0;
    XRAM[3684] = 8'b0;
    XRAM[3685] = 8'b0;
    XRAM[3686] = 8'b0;
    XRAM[3687] = 8'b0;
    XRAM[3688] = 8'b0;
    XRAM[3689] = 8'b0;
    XRAM[3690] = 8'b0;
    XRAM[3691] = 8'b0;
    XRAM[3692] = 8'b0;
    XRAM[3693] = 8'b0;
    XRAM[3694] = 8'b0;
    XRAM[3695] = 8'b0;
    XRAM[3696] = 8'b0;
    XRAM[3697] = 8'b0;
    XRAM[3698] = 8'b0;
    XRAM[3699] = 8'b0;
    XRAM[3700] = 8'b0;
    XRAM[3701] = 8'b0;
    XRAM[3702] = 8'b0;
    XRAM[3703] = 8'b0;
    XRAM[3704] = 8'b0;
    XRAM[3705] = 8'b0;
    XRAM[3706] = 8'b0;
    XRAM[3707] = 8'b0;
    XRAM[3708] = 8'b0;
    XRAM[3709] = 8'b0;
    XRAM[3710] = 8'b0;
    XRAM[3711] = 8'b0;
    XRAM[3712] = 8'b0;
    XRAM[3713] = 8'b0;
    XRAM[3714] = 8'b0;
    XRAM[3715] = 8'b0;
    XRAM[3716] = 8'b0;
    XRAM[3717] = 8'b0;
    XRAM[3718] = 8'b0;
    XRAM[3719] = 8'b0;
    XRAM[3720] = 8'b0;
    XRAM[3721] = 8'b0;
    XRAM[3722] = 8'b0;
    XRAM[3723] = 8'b0;
    XRAM[3724] = 8'b0;
    XRAM[3725] = 8'b0;
    XRAM[3726] = 8'b0;
    XRAM[3727] = 8'b0;
    XRAM[3728] = 8'b0;
    XRAM[3729] = 8'b0;
    XRAM[3730] = 8'b0;
    XRAM[3731] = 8'b0;
    XRAM[3732] = 8'b0;
    XRAM[3733] = 8'b0;
    XRAM[3734] = 8'b0;
    XRAM[3735] = 8'b0;
    XRAM[3736] = 8'b0;
    XRAM[3737] = 8'b0;
    XRAM[3738] = 8'b0;
    XRAM[3739] = 8'b0;
    XRAM[3740] = 8'b0;
    XRAM[3741] = 8'b0;
    XRAM[3742] = 8'b0;
    XRAM[3743] = 8'b0;
    XRAM[3744] = 8'b0;
    XRAM[3745] = 8'b0;
    XRAM[3746] = 8'b0;
    XRAM[3747] = 8'b0;
    XRAM[3748] = 8'b0;
    XRAM[3749] = 8'b0;
    XRAM[3750] = 8'b0;
    XRAM[3751] = 8'b0;
    XRAM[3752] = 8'b0;
    XRAM[3753] = 8'b0;
    XRAM[3754] = 8'b0;
    XRAM[3755] = 8'b0;
    XRAM[3756] = 8'b0;
    XRAM[3757] = 8'b0;
    XRAM[3758] = 8'b0;
    XRAM[3759] = 8'b0;
    XRAM[3760] = 8'b0;
    XRAM[3761] = 8'b0;
    XRAM[3762] = 8'b0;
    XRAM[3763] = 8'b0;
    XRAM[3764] = 8'b0;
    XRAM[3765] = 8'b0;
    XRAM[3766] = 8'b0;
    XRAM[3767] = 8'b0;
    XRAM[3768] = 8'b0;
    XRAM[3769] = 8'b0;
    XRAM[3770] = 8'b0;
    XRAM[3771] = 8'b0;
    XRAM[3772] = 8'b0;
    XRAM[3773] = 8'b0;
    XRAM[3774] = 8'b0;
    XRAM[3775] = 8'b0;
    XRAM[3776] = 8'b0;
    XRAM[3777] = 8'b0;
    XRAM[3778] = 8'b0;
    XRAM[3779] = 8'b0;
    XRAM[3780] = 8'b0;
    XRAM[3781] = 8'b0;
    XRAM[3782] = 8'b0;
    XRAM[3783] = 8'b0;
    XRAM[3784] = 8'b0;
    XRAM[3785] = 8'b0;
    XRAM[3786] = 8'b0;
    XRAM[3787] = 8'b0;
    XRAM[3788] = 8'b0;
    XRAM[3789] = 8'b0;
    XRAM[3790] = 8'b0;
    XRAM[3791] = 8'b0;
    XRAM[3792] = 8'b0;
    XRAM[3793] = 8'b0;
    XRAM[3794] = 8'b0;
    XRAM[3795] = 8'b0;
    XRAM[3796] = 8'b0;
    XRAM[3797] = 8'b0;
    XRAM[3798] = 8'b0;
    XRAM[3799] = 8'b0;
    XRAM[3800] = 8'b0;
    XRAM[3801] = 8'b0;
    XRAM[3802] = 8'b0;
    XRAM[3803] = 8'b0;
    XRAM[3804] = 8'b0;
    XRAM[3805] = 8'b0;
    XRAM[3806] = 8'b0;
    XRAM[3807] = 8'b0;
    XRAM[3808] = 8'b0;
    XRAM[3809] = 8'b0;
    XRAM[3810] = 8'b0;
    XRAM[3811] = 8'b0;
    XRAM[3812] = 8'b0;
    XRAM[3813] = 8'b0;
    XRAM[3814] = 8'b0;
    XRAM[3815] = 8'b0;
    XRAM[3816] = 8'b0;
    XRAM[3817] = 8'b0;
    XRAM[3818] = 8'b0;
    XRAM[3819] = 8'b0;
    XRAM[3820] = 8'b0;
    XRAM[3821] = 8'b0;
    XRAM[3822] = 8'b0;
    XRAM[3823] = 8'b0;
    XRAM[3824] = 8'b0;
    XRAM[3825] = 8'b0;
    XRAM[3826] = 8'b0;
    XRAM[3827] = 8'b0;
    XRAM[3828] = 8'b0;
    XRAM[3829] = 8'b0;
    XRAM[3830] = 8'b0;
    XRAM[3831] = 8'b0;
    XRAM[3832] = 8'b0;
    XRAM[3833] = 8'b0;
    XRAM[3834] = 8'b0;
    XRAM[3835] = 8'b0;
    XRAM[3836] = 8'b0;
    XRAM[3837] = 8'b0;
    XRAM[3838] = 8'b0;
    XRAM[3839] = 8'b0;
    XRAM[3840] = 8'b0;
    XRAM[3841] = 8'b0;
    XRAM[3842] = 8'b0;
    XRAM[3843] = 8'b0;
    XRAM[3844] = 8'b0;
    XRAM[3845] = 8'b0;
    XRAM[3846] = 8'b0;
    XRAM[3847] = 8'b0;
    XRAM[3848] = 8'b0;
    XRAM[3849] = 8'b0;
    XRAM[3850] = 8'b0;
    XRAM[3851] = 8'b0;
    XRAM[3852] = 8'b0;
    XRAM[3853] = 8'b0;
    XRAM[3854] = 8'b0;
    XRAM[3855] = 8'b0;
    XRAM[3856] = 8'b0;
    XRAM[3857] = 8'b0;
    XRAM[3858] = 8'b0;
    XRAM[3859] = 8'b0;
    XRAM[3860] = 8'b0;
    XRAM[3861] = 8'b0;
    XRAM[3862] = 8'b0;
    XRAM[3863] = 8'b0;
    XRAM[3864] = 8'b0;
    XRAM[3865] = 8'b0;
    XRAM[3866] = 8'b0;
    XRAM[3867] = 8'b0;
    XRAM[3868] = 8'b0;
    XRAM[3869] = 8'b0;
    XRAM[3870] = 8'b0;
    XRAM[3871] = 8'b0;
    XRAM[3872] = 8'b0;
    XRAM[3873] = 8'b0;
    XRAM[3874] = 8'b0;
    XRAM[3875] = 8'b0;
    XRAM[3876] = 8'b0;
    XRAM[3877] = 8'b0;
    XRAM[3878] = 8'b0;
    XRAM[3879] = 8'b0;
    XRAM[3880] = 8'b0;
    XRAM[3881] = 8'b0;
    XRAM[3882] = 8'b0;
    XRAM[3883] = 8'b0;
    XRAM[3884] = 8'b0;
    XRAM[3885] = 8'b0;
    XRAM[3886] = 8'b0;
    XRAM[3887] = 8'b0;
    XRAM[3888] = 8'b0;
    XRAM[3889] = 8'b0;
    XRAM[3890] = 8'b0;
    XRAM[3891] = 8'b0;
    XRAM[3892] = 8'b0;
    XRAM[3893] = 8'b0;
    XRAM[3894] = 8'b0;
    XRAM[3895] = 8'b0;
    XRAM[3896] = 8'b0;
    XRAM[3897] = 8'b0;
    XRAM[3898] = 8'b0;
    XRAM[3899] = 8'b0;
    XRAM[3900] = 8'b0;
    XRAM[3901] = 8'b0;
    XRAM[3902] = 8'b0;
    XRAM[3903] = 8'b0;
    XRAM[3904] = 8'b0;
    XRAM[3905] = 8'b0;
    XRAM[3906] = 8'b0;
    XRAM[3907] = 8'b0;
    XRAM[3908] = 8'b0;
    XRAM[3909] = 8'b0;
    XRAM[3910] = 8'b0;
    XRAM[3911] = 8'b0;
    XRAM[3912] = 8'b0;
    XRAM[3913] = 8'b0;
    XRAM[3914] = 8'b0;
    XRAM[3915] = 8'b0;
    XRAM[3916] = 8'b0;
    XRAM[3917] = 8'b0;
    XRAM[3918] = 8'b0;
    XRAM[3919] = 8'b0;
    XRAM[3920] = 8'b0;
    XRAM[3921] = 8'b0;
    XRAM[3922] = 8'b0;
    XRAM[3923] = 8'b0;
    XRAM[3924] = 8'b0;
    XRAM[3925] = 8'b0;
    XRAM[3926] = 8'b0;
    XRAM[3927] = 8'b0;
    XRAM[3928] = 8'b0;
    XRAM[3929] = 8'b0;
    XRAM[3930] = 8'b0;
    XRAM[3931] = 8'b0;
    XRAM[3932] = 8'b0;
    XRAM[3933] = 8'b0;
    XRAM[3934] = 8'b0;
    XRAM[3935] = 8'b0;
    XRAM[3936] = 8'b0;
    XRAM[3937] = 8'b0;
    XRAM[3938] = 8'b0;
    XRAM[3939] = 8'b0;
    XRAM[3940] = 8'b0;
    XRAM[3941] = 8'b0;
    XRAM[3942] = 8'b0;
    XRAM[3943] = 8'b0;
    XRAM[3944] = 8'b0;
    XRAM[3945] = 8'b0;
    XRAM[3946] = 8'b0;
    XRAM[3947] = 8'b0;
    XRAM[3948] = 8'b0;
    XRAM[3949] = 8'b0;
    XRAM[3950] = 8'b0;
    XRAM[3951] = 8'b0;
    XRAM[3952] = 8'b0;
    XRAM[3953] = 8'b0;
    XRAM[3954] = 8'b0;
    XRAM[3955] = 8'b0;
    XRAM[3956] = 8'b0;
    XRAM[3957] = 8'b0;
    XRAM[3958] = 8'b0;
    XRAM[3959] = 8'b0;
    XRAM[3960] = 8'b0;
    XRAM[3961] = 8'b0;
    XRAM[3962] = 8'b0;
    XRAM[3963] = 8'b0;
    XRAM[3964] = 8'b0;
    XRAM[3965] = 8'b0;
    XRAM[3966] = 8'b0;
    XRAM[3967] = 8'b0;
    XRAM[3968] = 8'b0;
    XRAM[3969] = 8'b0;
    XRAM[3970] = 8'b0;
    XRAM[3971] = 8'b0;
    XRAM[3972] = 8'b0;
    XRAM[3973] = 8'b0;
    XRAM[3974] = 8'b0;
    XRAM[3975] = 8'b0;
    XRAM[3976] = 8'b0;
    XRAM[3977] = 8'b0;
    XRAM[3978] = 8'b0;
    XRAM[3979] = 8'b0;
    XRAM[3980] = 8'b0;
    XRAM[3981] = 8'b0;
    XRAM[3982] = 8'b0;
    XRAM[3983] = 8'b0;
    XRAM[3984] = 8'b0;
    XRAM[3985] = 8'b0;
    XRAM[3986] = 8'b0;
    XRAM[3987] = 8'b0;
    XRAM[3988] = 8'b0;
    XRAM[3989] = 8'b0;
    XRAM[3990] = 8'b0;
    XRAM[3991] = 8'b0;
    XRAM[3992] = 8'b0;
    XRAM[3993] = 8'b0;
    XRAM[3994] = 8'b0;
    XRAM[3995] = 8'b0;
    XRAM[3996] = 8'b0;
    XRAM[3997] = 8'b0;
    XRAM[3998] = 8'b0;
    XRAM[3999] = 8'b0;
    XRAM[4000] = 8'b0;
    XRAM[4001] = 8'b0;
    XRAM[4002] = 8'b0;
    XRAM[4003] = 8'b0;
    XRAM[4004] = 8'b0;
    XRAM[4005] = 8'b0;
    XRAM[4006] = 8'b0;
    XRAM[4007] = 8'b0;
    XRAM[4008] = 8'b0;
    XRAM[4009] = 8'b0;
    XRAM[4010] = 8'b0;
    XRAM[4011] = 8'b0;
    XRAM[4012] = 8'b0;
    XRAM[4013] = 8'b0;
    XRAM[4014] = 8'b0;
    XRAM[4015] = 8'b0;
    XRAM[4016] = 8'b0;
    XRAM[4017] = 8'b0;
    XRAM[4018] = 8'b0;
    XRAM[4019] = 8'b0;
    XRAM[4020] = 8'b0;
    XRAM[4021] = 8'b0;
    XRAM[4022] = 8'b0;
    XRAM[4023] = 8'b0;
    XRAM[4024] = 8'b0;
    XRAM[4025] = 8'b0;
    XRAM[4026] = 8'b0;
    XRAM[4027] = 8'b0;
    XRAM[4028] = 8'b0;
    XRAM[4029] = 8'b0;
    XRAM[4030] = 8'b0;
    XRAM[4031] = 8'b0;
    XRAM[4032] = 8'b0;
    XRAM[4033] = 8'b0;
    XRAM[4034] = 8'b0;
    XRAM[4035] = 8'b0;
    XRAM[4036] = 8'b0;
    XRAM[4037] = 8'b0;
    XRAM[4038] = 8'b0;
    XRAM[4039] = 8'b0;
    XRAM[4040] = 8'b0;
    XRAM[4041] = 8'b0;
    XRAM[4042] = 8'b0;
    XRAM[4043] = 8'b0;
    XRAM[4044] = 8'b0;
    XRAM[4045] = 8'b0;
    XRAM[4046] = 8'b0;
    XRAM[4047] = 8'b0;
    XRAM[4048] = 8'b0;
    XRAM[4049] = 8'b0;
    XRAM[4050] = 8'b0;
    XRAM[4051] = 8'b0;
    XRAM[4052] = 8'b0;
    XRAM[4053] = 8'b0;
    XRAM[4054] = 8'b0;
    XRAM[4055] = 8'b0;
    XRAM[4056] = 8'b0;
    XRAM[4057] = 8'b0;
    XRAM[4058] = 8'b0;
    XRAM[4059] = 8'b0;
    XRAM[4060] = 8'b0;
    XRAM[4061] = 8'b0;
    XRAM[4062] = 8'b0;
    XRAM[4063] = 8'b0;
    XRAM[4064] = 8'b0;
    XRAM[4065] = 8'b0;
    XRAM[4066] = 8'b0;
    XRAM[4067] = 8'b0;
    XRAM[4068] = 8'b0;
    XRAM[4069] = 8'b0;
    XRAM[4070] = 8'b0;
    XRAM[4071] = 8'b0;
    XRAM[4072] = 8'b0;
    XRAM[4073] = 8'b0;
    XRAM[4074] = 8'b0;
    XRAM[4075] = 8'b0;
    XRAM[4076] = 8'b0;
    XRAM[4077] = 8'b0;
    XRAM[4078] = 8'b0;
    XRAM[4079] = 8'b0;
    XRAM[4080] = 8'b0;
    XRAM[4081] = 8'b0;
    XRAM[4082] = 8'b0;
    XRAM[4083] = 8'b0;
    XRAM[4084] = 8'b0;
    XRAM[4085] = 8'b0;
    XRAM[4086] = 8'b0;
    XRAM[4087] = 8'b0;
    XRAM[4088] = 8'b0;
    XRAM[4089] = 8'b0;
    XRAM[4090] = 8'b0;
    XRAM[4091] = 8'b0;
    XRAM[4092] = 8'b0;
    XRAM[4093] = 8'b0;
    XRAM[4094] = 8'b0;
    XRAM[4095] = 8'b0;
    XRAM[4096] = 8'b0;
    XRAM[4097] = 8'b0;
    XRAM[4098] = 8'b0;
    XRAM[4099] = 8'b0;
    XRAM[4100] = 8'b0;
    XRAM[4101] = 8'b0;
    XRAM[4102] = 8'b0;
    XRAM[4103] = 8'b0;
    XRAM[4104] = 8'b0;
    XRAM[4105] = 8'b0;
    XRAM[4106] = 8'b0;
    XRAM[4107] = 8'b0;
    XRAM[4108] = 8'b0;
    XRAM[4109] = 8'b0;
    XRAM[4110] = 8'b0;
    XRAM[4111] = 8'b0;
    XRAM[4112] = 8'b0;
    XRAM[4113] = 8'b0;
    XRAM[4114] = 8'b0;
    XRAM[4115] = 8'b0;
    XRAM[4116] = 8'b0;
    XRAM[4117] = 8'b0;
    XRAM[4118] = 8'b0;
    XRAM[4119] = 8'b0;
    XRAM[4120] = 8'b0;
    XRAM[4121] = 8'b0;
    XRAM[4122] = 8'b0;
    XRAM[4123] = 8'b0;
    XRAM[4124] = 8'b0;
    XRAM[4125] = 8'b0;
    XRAM[4126] = 8'b0;
    XRAM[4127] = 8'b0;
    XRAM[4128] = 8'b0;
    XRAM[4129] = 8'b0;
    XRAM[4130] = 8'b0;
    XRAM[4131] = 8'b0;
    XRAM[4132] = 8'b0;
    XRAM[4133] = 8'b0;
    XRAM[4134] = 8'b0;
    XRAM[4135] = 8'b0;
    XRAM[4136] = 8'b0;
    XRAM[4137] = 8'b0;
    XRAM[4138] = 8'b0;
    XRAM[4139] = 8'b0;
    XRAM[4140] = 8'b0;
    XRAM[4141] = 8'b0;
    XRAM[4142] = 8'b0;
    XRAM[4143] = 8'b0;
    XRAM[4144] = 8'b0;
    XRAM[4145] = 8'b0;
    XRAM[4146] = 8'b0;
    XRAM[4147] = 8'b0;
    XRAM[4148] = 8'b0;
    XRAM[4149] = 8'b0;
    XRAM[4150] = 8'b0;
    XRAM[4151] = 8'b0;
    XRAM[4152] = 8'b0;
    XRAM[4153] = 8'b0;
    XRAM[4154] = 8'b0;
    XRAM[4155] = 8'b0;
    XRAM[4156] = 8'b0;
    XRAM[4157] = 8'b0;
    XRAM[4158] = 8'b0;
    XRAM[4159] = 8'b0;
    XRAM[4160] = 8'b0;
    XRAM[4161] = 8'b0;
    XRAM[4162] = 8'b0;
    XRAM[4163] = 8'b0;
    XRAM[4164] = 8'b0;
    XRAM[4165] = 8'b0;
    XRAM[4166] = 8'b0;
    XRAM[4167] = 8'b0;
    XRAM[4168] = 8'b0;
    XRAM[4169] = 8'b0;
    XRAM[4170] = 8'b0;
    XRAM[4171] = 8'b0;
    XRAM[4172] = 8'b0;
    XRAM[4173] = 8'b0;
    XRAM[4174] = 8'b0;
    XRAM[4175] = 8'b0;
    XRAM[4176] = 8'b0;
    XRAM[4177] = 8'b0;
    XRAM[4178] = 8'b0;
    XRAM[4179] = 8'b0;
    XRAM[4180] = 8'b0;
    XRAM[4181] = 8'b0;
    XRAM[4182] = 8'b0;
    XRAM[4183] = 8'b0;
    XRAM[4184] = 8'b0;
    XRAM[4185] = 8'b0;
    XRAM[4186] = 8'b0;
    XRAM[4187] = 8'b0;
    XRAM[4188] = 8'b0;
    XRAM[4189] = 8'b0;
    XRAM[4190] = 8'b0;
    XRAM[4191] = 8'b0;
    XRAM[4192] = 8'b0;
    XRAM[4193] = 8'b0;
    XRAM[4194] = 8'b0;
    XRAM[4195] = 8'b0;
    XRAM[4196] = 8'b0;
    XRAM[4197] = 8'b0;
    XRAM[4198] = 8'b0;
    XRAM[4199] = 8'b0;
    XRAM[4200] = 8'b0;
    XRAM[4201] = 8'b0;
    XRAM[4202] = 8'b0;
    XRAM[4203] = 8'b0;
    XRAM[4204] = 8'b0;
    XRAM[4205] = 8'b0;
    XRAM[4206] = 8'b0;
    XRAM[4207] = 8'b0;
    XRAM[4208] = 8'b0;
    XRAM[4209] = 8'b0;
    XRAM[4210] = 8'b0;
    XRAM[4211] = 8'b0;
    XRAM[4212] = 8'b0;
    XRAM[4213] = 8'b0;
    XRAM[4214] = 8'b0;
    XRAM[4215] = 8'b0;
    XRAM[4216] = 8'b0;
    XRAM[4217] = 8'b0;
    XRAM[4218] = 8'b0;
    XRAM[4219] = 8'b0;
    XRAM[4220] = 8'b0;
    XRAM[4221] = 8'b0;
    XRAM[4222] = 8'b0;
    XRAM[4223] = 8'b0;
    XRAM[4224] = 8'b0;
    XRAM[4225] = 8'b0;
    XRAM[4226] = 8'b0;
    XRAM[4227] = 8'b0;
    XRAM[4228] = 8'b0;
    XRAM[4229] = 8'b0;
    XRAM[4230] = 8'b0;
    XRAM[4231] = 8'b0;
    XRAM[4232] = 8'b0;
    XRAM[4233] = 8'b0;
    XRAM[4234] = 8'b0;
    XRAM[4235] = 8'b0;
    XRAM[4236] = 8'b0;
    XRAM[4237] = 8'b0;
    XRAM[4238] = 8'b0;
    XRAM[4239] = 8'b0;
    XRAM[4240] = 8'b0;
    XRAM[4241] = 8'b0;
    XRAM[4242] = 8'b0;
    XRAM[4243] = 8'b0;
    XRAM[4244] = 8'b0;
    XRAM[4245] = 8'b0;
    XRAM[4246] = 8'b0;
    XRAM[4247] = 8'b0;
    XRAM[4248] = 8'b0;
    XRAM[4249] = 8'b0;
    XRAM[4250] = 8'b0;
    XRAM[4251] = 8'b0;
    XRAM[4252] = 8'b0;
    XRAM[4253] = 8'b0;
    XRAM[4254] = 8'b0;
    XRAM[4255] = 8'b0;
    XRAM[4256] = 8'b0;
    XRAM[4257] = 8'b0;
    XRAM[4258] = 8'b0;
    XRAM[4259] = 8'b0;
    XRAM[4260] = 8'b0;
    XRAM[4261] = 8'b0;
    XRAM[4262] = 8'b0;
    XRAM[4263] = 8'b0;
    XRAM[4264] = 8'b0;
    XRAM[4265] = 8'b0;
    XRAM[4266] = 8'b0;
    XRAM[4267] = 8'b0;
    XRAM[4268] = 8'b0;
    XRAM[4269] = 8'b0;
    XRAM[4270] = 8'b0;
    XRAM[4271] = 8'b0;
    XRAM[4272] = 8'b0;
    XRAM[4273] = 8'b0;
    XRAM[4274] = 8'b0;
    XRAM[4275] = 8'b0;
    XRAM[4276] = 8'b0;
    XRAM[4277] = 8'b0;
    XRAM[4278] = 8'b0;
    XRAM[4279] = 8'b0;
    XRAM[4280] = 8'b0;
    XRAM[4281] = 8'b0;
    XRAM[4282] = 8'b0;
    XRAM[4283] = 8'b0;
    XRAM[4284] = 8'b0;
    XRAM[4285] = 8'b0;
    XRAM[4286] = 8'b0;
    XRAM[4287] = 8'b0;
    XRAM[4288] = 8'b0;
    XRAM[4289] = 8'b0;
    XRAM[4290] = 8'b0;
    XRAM[4291] = 8'b0;
    XRAM[4292] = 8'b0;
    XRAM[4293] = 8'b0;
    XRAM[4294] = 8'b0;
    XRAM[4295] = 8'b0;
    XRAM[4296] = 8'b0;
    XRAM[4297] = 8'b0;
    XRAM[4298] = 8'b0;
    XRAM[4299] = 8'b0;
    XRAM[4300] = 8'b0;
    XRAM[4301] = 8'b0;
    XRAM[4302] = 8'b0;
    XRAM[4303] = 8'b0;
    XRAM[4304] = 8'b0;
    XRAM[4305] = 8'b0;
    XRAM[4306] = 8'b0;
    XRAM[4307] = 8'b0;
    XRAM[4308] = 8'b0;
    XRAM[4309] = 8'b0;
    XRAM[4310] = 8'b0;
    XRAM[4311] = 8'b0;
    XRAM[4312] = 8'b0;
    XRAM[4313] = 8'b0;
    XRAM[4314] = 8'b0;
    XRAM[4315] = 8'b0;
    XRAM[4316] = 8'b0;
    XRAM[4317] = 8'b0;
    XRAM[4318] = 8'b0;
    XRAM[4319] = 8'b0;
    XRAM[4320] = 8'b0;
    XRAM[4321] = 8'b0;
    XRAM[4322] = 8'b0;
    XRAM[4323] = 8'b0;
    XRAM[4324] = 8'b0;
    XRAM[4325] = 8'b0;
    XRAM[4326] = 8'b0;
    XRAM[4327] = 8'b0;
    XRAM[4328] = 8'b0;
    XRAM[4329] = 8'b0;
    XRAM[4330] = 8'b0;
    XRAM[4331] = 8'b0;
    XRAM[4332] = 8'b0;
    XRAM[4333] = 8'b0;
    XRAM[4334] = 8'b0;
    XRAM[4335] = 8'b0;
    XRAM[4336] = 8'b0;
    XRAM[4337] = 8'b0;
    XRAM[4338] = 8'b0;
    XRAM[4339] = 8'b0;
    XRAM[4340] = 8'b0;
    XRAM[4341] = 8'b0;
    XRAM[4342] = 8'b0;
    XRAM[4343] = 8'b0;
    XRAM[4344] = 8'b0;
    XRAM[4345] = 8'b0;
    XRAM[4346] = 8'b0;
    XRAM[4347] = 8'b0;
    XRAM[4348] = 8'b0;
    XRAM[4349] = 8'b0;
    XRAM[4350] = 8'b0;
    XRAM[4351] = 8'b0;
    XRAM[4352] = 8'b0;
    XRAM[4353] = 8'b0;
    XRAM[4354] = 8'b0;
    XRAM[4355] = 8'b0;
    XRAM[4356] = 8'b0;
    XRAM[4357] = 8'b0;
    XRAM[4358] = 8'b0;
    XRAM[4359] = 8'b0;
    XRAM[4360] = 8'b0;
    XRAM[4361] = 8'b0;
    XRAM[4362] = 8'b0;
    XRAM[4363] = 8'b0;
    XRAM[4364] = 8'b0;
    XRAM[4365] = 8'b0;
    XRAM[4366] = 8'b0;
    XRAM[4367] = 8'b0;
    XRAM[4368] = 8'b0;
    XRAM[4369] = 8'b0;
    XRAM[4370] = 8'b0;
    XRAM[4371] = 8'b0;
    XRAM[4372] = 8'b0;
    XRAM[4373] = 8'b0;
    XRAM[4374] = 8'b0;
    XRAM[4375] = 8'b0;
    XRAM[4376] = 8'b0;
    XRAM[4377] = 8'b0;
    XRAM[4378] = 8'b0;
    XRAM[4379] = 8'b0;
    XRAM[4380] = 8'b0;
    XRAM[4381] = 8'b0;
    XRAM[4382] = 8'b0;
    XRAM[4383] = 8'b0;
    XRAM[4384] = 8'b0;
    XRAM[4385] = 8'b0;
    XRAM[4386] = 8'b0;
    XRAM[4387] = 8'b0;
    XRAM[4388] = 8'b0;
    XRAM[4389] = 8'b0;
    XRAM[4390] = 8'b0;
    XRAM[4391] = 8'b0;
    XRAM[4392] = 8'b0;
    XRAM[4393] = 8'b0;
    XRAM[4394] = 8'b0;
    XRAM[4395] = 8'b0;
    XRAM[4396] = 8'b0;
    XRAM[4397] = 8'b0;
    XRAM[4398] = 8'b0;
    XRAM[4399] = 8'b0;
    XRAM[4400] = 8'b0;
    XRAM[4401] = 8'b0;
    XRAM[4402] = 8'b0;
    XRAM[4403] = 8'b0;
    XRAM[4404] = 8'b0;
    XRAM[4405] = 8'b0;
    XRAM[4406] = 8'b0;
    XRAM[4407] = 8'b0;
    XRAM[4408] = 8'b0;
    XRAM[4409] = 8'b0;
    XRAM[4410] = 8'b0;
    XRAM[4411] = 8'b0;
    XRAM[4412] = 8'b0;
    XRAM[4413] = 8'b0;
    XRAM[4414] = 8'b0;
    XRAM[4415] = 8'b0;
    XRAM[4416] = 8'b0;
    XRAM[4417] = 8'b0;
    XRAM[4418] = 8'b0;
    XRAM[4419] = 8'b0;
    XRAM[4420] = 8'b0;
    XRAM[4421] = 8'b0;
    XRAM[4422] = 8'b0;
    XRAM[4423] = 8'b0;
    XRAM[4424] = 8'b0;
    XRAM[4425] = 8'b0;
    XRAM[4426] = 8'b0;
    XRAM[4427] = 8'b0;
    XRAM[4428] = 8'b0;
    XRAM[4429] = 8'b0;
    XRAM[4430] = 8'b0;
    XRAM[4431] = 8'b0;
    XRAM[4432] = 8'b0;
    XRAM[4433] = 8'b0;
    XRAM[4434] = 8'b0;
    XRAM[4435] = 8'b0;
    XRAM[4436] = 8'b0;
    XRAM[4437] = 8'b0;
    XRAM[4438] = 8'b0;
    XRAM[4439] = 8'b0;
    XRAM[4440] = 8'b0;
    XRAM[4441] = 8'b0;
    XRAM[4442] = 8'b0;
    XRAM[4443] = 8'b0;
    XRAM[4444] = 8'b0;
    XRAM[4445] = 8'b0;
    XRAM[4446] = 8'b0;
    XRAM[4447] = 8'b0;
    XRAM[4448] = 8'b0;
    XRAM[4449] = 8'b0;
    XRAM[4450] = 8'b0;
    XRAM[4451] = 8'b0;
    XRAM[4452] = 8'b0;
    XRAM[4453] = 8'b0;
    XRAM[4454] = 8'b0;
    XRAM[4455] = 8'b0;
    XRAM[4456] = 8'b0;
    XRAM[4457] = 8'b0;
    XRAM[4458] = 8'b0;
    XRAM[4459] = 8'b0;
    XRAM[4460] = 8'b0;
    XRAM[4461] = 8'b0;
    XRAM[4462] = 8'b0;
    XRAM[4463] = 8'b0;
    XRAM[4464] = 8'b0;
    XRAM[4465] = 8'b0;
    XRAM[4466] = 8'b0;
    XRAM[4467] = 8'b0;
    XRAM[4468] = 8'b0;
    XRAM[4469] = 8'b0;
    XRAM[4470] = 8'b0;
    XRAM[4471] = 8'b0;
    XRAM[4472] = 8'b0;
    XRAM[4473] = 8'b0;
    XRAM[4474] = 8'b0;
    XRAM[4475] = 8'b0;
    XRAM[4476] = 8'b0;
    XRAM[4477] = 8'b0;
    XRAM[4478] = 8'b0;
    XRAM[4479] = 8'b0;
    XRAM[4480] = 8'b0;
    XRAM[4481] = 8'b0;
    XRAM[4482] = 8'b0;
    XRAM[4483] = 8'b0;
    XRAM[4484] = 8'b0;
    XRAM[4485] = 8'b0;
    XRAM[4486] = 8'b0;
    XRAM[4487] = 8'b0;
    XRAM[4488] = 8'b0;
    XRAM[4489] = 8'b0;
    XRAM[4490] = 8'b0;
    XRAM[4491] = 8'b0;
    XRAM[4492] = 8'b0;
    XRAM[4493] = 8'b0;
    XRAM[4494] = 8'b0;
    XRAM[4495] = 8'b0;
    XRAM[4496] = 8'b0;
    XRAM[4497] = 8'b0;
    XRAM[4498] = 8'b0;
    XRAM[4499] = 8'b0;
    XRAM[4500] = 8'b0;
    XRAM[4501] = 8'b0;
    XRAM[4502] = 8'b0;
    XRAM[4503] = 8'b0;
    XRAM[4504] = 8'b0;
    XRAM[4505] = 8'b0;
    XRAM[4506] = 8'b0;
    XRAM[4507] = 8'b0;
    XRAM[4508] = 8'b0;
    XRAM[4509] = 8'b0;
    XRAM[4510] = 8'b0;
    XRAM[4511] = 8'b0;
    XRAM[4512] = 8'b0;
    XRAM[4513] = 8'b0;
    XRAM[4514] = 8'b0;
    XRAM[4515] = 8'b0;
    XRAM[4516] = 8'b0;
    XRAM[4517] = 8'b0;
    XRAM[4518] = 8'b0;
    XRAM[4519] = 8'b0;
    XRAM[4520] = 8'b0;
    XRAM[4521] = 8'b0;
    XRAM[4522] = 8'b0;
    XRAM[4523] = 8'b0;
    XRAM[4524] = 8'b0;
    XRAM[4525] = 8'b0;
    XRAM[4526] = 8'b0;
    XRAM[4527] = 8'b0;
    XRAM[4528] = 8'b0;
    XRAM[4529] = 8'b0;
    XRAM[4530] = 8'b0;
    XRAM[4531] = 8'b0;
    XRAM[4532] = 8'b0;
    XRAM[4533] = 8'b0;
    XRAM[4534] = 8'b0;
    XRAM[4535] = 8'b0;
    XRAM[4536] = 8'b0;
    XRAM[4537] = 8'b0;
    XRAM[4538] = 8'b0;
    XRAM[4539] = 8'b0;
    XRAM[4540] = 8'b0;
    XRAM[4541] = 8'b0;
    XRAM[4542] = 8'b0;
    XRAM[4543] = 8'b0;
    XRAM[4544] = 8'b0;
    XRAM[4545] = 8'b0;
    XRAM[4546] = 8'b0;
    XRAM[4547] = 8'b0;
    XRAM[4548] = 8'b0;
    XRAM[4549] = 8'b0;
    XRAM[4550] = 8'b0;
    XRAM[4551] = 8'b0;
    XRAM[4552] = 8'b0;
    XRAM[4553] = 8'b0;
    XRAM[4554] = 8'b0;
    XRAM[4555] = 8'b0;
    XRAM[4556] = 8'b0;
    XRAM[4557] = 8'b0;
    XRAM[4558] = 8'b0;
    XRAM[4559] = 8'b0;
    XRAM[4560] = 8'b0;
    XRAM[4561] = 8'b0;
    XRAM[4562] = 8'b0;
    XRAM[4563] = 8'b0;
    XRAM[4564] = 8'b0;
    XRAM[4565] = 8'b0;
    XRAM[4566] = 8'b0;
    XRAM[4567] = 8'b0;
    XRAM[4568] = 8'b0;
    XRAM[4569] = 8'b0;
    XRAM[4570] = 8'b0;
    XRAM[4571] = 8'b0;
    XRAM[4572] = 8'b0;
    XRAM[4573] = 8'b0;
    XRAM[4574] = 8'b0;
    XRAM[4575] = 8'b0;
    XRAM[4576] = 8'b0;
    XRAM[4577] = 8'b0;
    XRAM[4578] = 8'b0;
    XRAM[4579] = 8'b0;
    XRAM[4580] = 8'b0;
    XRAM[4581] = 8'b0;
    XRAM[4582] = 8'b0;
    XRAM[4583] = 8'b0;
    XRAM[4584] = 8'b0;
    XRAM[4585] = 8'b0;
    XRAM[4586] = 8'b0;
    XRAM[4587] = 8'b0;
    XRAM[4588] = 8'b0;
    XRAM[4589] = 8'b0;
    XRAM[4590] = 8'b0;
    XRAM[4591] = 8'b0;
    XRAM[4592] = 8'b0;
    XRAM[4593] = 8'b0;
    XRAM[4594] = 8'b0;
    XRAM[4595] = 8'b0;
    XRAM[4596] = 8'b0;
    XRAM[4597] = 8'b0;
    XRAM[4598] = 8'b0;
    XRAM[4599] = 8'b0;
    XRAM[4600] = 8'b0;
    XRAM[4601] = 8'b0;
    XRAM[4602] = 8'b0;
    XRAM[4603] = 8'b0;
    XRAM[4604] = 8'b0;
    XRAM[4605] = 8'b0;
    XRAM[4606] = 8'b0;
    XRAM[4607] = 8'b0;
    XRAM[4608] = 8'b0;
    XRAM[4609] = 8'b0;
    XRAM[4610] = 8'b0;
    XRAM[4611] = 8'b0;
    XRAM[4612] = 8'b0;
    XRAM[4613] = 8'b0;
    XRAM[4614] = 8'b0;
    XRAM[4615] = 8'b0;
    XRAM[4616] = 8'b0;
    XRAM[4617] = 8'b0;
    XRAM[4618] = 8'b0;
    XRAM[4619] = 8'b0;
    XRAM[4620] = 8'b0;
    XRAM[4621] = 8'b0;
    XRAM[4622] = 8'b0;
    XRAM[4623] = 8'b0;
    XRAM[4624] = 8'b0;
    XRAM[4625] = 8'b0;
    XRAM[4626] = 8'b0;
    XRAM[4627] = 8'b0;
    XRAM[4628] = 8'b0;
    XRAM[4629] = 8'b0;
    XRAM[4630] = 8'b0;
    XRAM[4631] = 8'b0;
    XRAM[4632] = 8'b0;
    XRAM[4633] = 8'b0;
    XRAM[4634] = 8'b0;
    XRAM[4635] = 8'b0;
    XRAM[4636] = 8'b0;
    XRAM[4637] = 8'b0;
    XRAM[4638] = 8'b0;
    XRAM[4639] = 8'b0;
    XRAM[4640] = 8'b0;
    XRAM[4641] = 8'b0;
    XRAM[4642] = 8'b0;
    XRAM[4643] = 8'b0;
    XRAM[4644] = 8'b0;
    XRAM[4645] = 8'b0;
    XRAM[4646] = 8'b0;
    XRAM[4647] = 8'b0;
    XRAM[4648] = 8'b0;
    XRAM[4649] = 8'b0;
    XRAM[4650] = 8'b0;
    XRAM[4651] = 8'b0;
    XRAM[4652] = 8'b0;
    XRAM[4653] = 8'b0;
    XRAM[4654] = 8'b0;
    XRAM[4655] = 8'b0;
    XRAM[4656] = 8'b0;
    XRAM[4657] = 8'b0;
    XRAM[4658] = 8'b0;
    XRAM[4659] = 8'b0;
    XRAM[4660] = 8'b0;
    XRAM[4661] = 8'b0;
    XRAM[4662] = 8'b0;
    XRAM[4663] = 8'b0;
    XRAM[4664] = 8'b0;
    XRAM[4665] = 8'b0;
    XRAM[4666] = 8'b0;
    XRAM[4667] = 8'b0;
    XRAM[4668] = 8'b0;
    XRAM[4669] = 8'b0;
    XRAM[4670] = 8'b0;
    XRAM[4671] = 8'b0;
    XRAM[4672] = 8'b0;
    XRAM[4673] = 8'b0;
    XRAM[4674] = 8'b0;
    XRAM[4675] = 8'b0;
    XRAM[4676] = 8'b0;
    XRAM[4677] = 8'b0;
    XRAM[4678] = 8'b0;
    XRAM[4679] = 8'b0;
    XRAM[4680] = 8'b0;
    XRAM[4681] = 8'b0;
    XRAM[4682] = 8'b0;
    XRAM[4683] = 8'b0;
    XRAM[4684] = 8'b0;
    XRAM[4685] = 8'b0;
    XRAM[4686] = 8'b0;
    XRAM[4687] = 8'b0;
    XRAM[4688] = 8'b0;
    XRAM[4689] = 8'b0;
    XRAM[4690] = 8'b0;
    XRAM[4691] = 8'b0;
    XRAM[4692] = 8'b0;
    XRAM[4693] = 8'b0;
    XRAM[4694] = 8'b0;
    XRAM[4695] = 8'b0;
    XRAM[4696] = 8'b0;
    XRAM[4697] = 8'b0;
    XRAM[4698] = 8'b0;
    XRAM[4699] = 8'b0;
    XRAM[4700] = 8'b0;
    XRAM[4701] = 8'b0;
    XRAM[4702] = 8'b0;
    XRAM[4703] = 8'b0;
    XRAM[4704] = 8'b0;
    XRAM[4705] = 8'b0;
    XRAM[4706] = 8'b0;
    XRAM[4707] = 8'b0;
    XRAM[4708] = 8'b0;
    XRAM[4709] = 8'b0;
    XRAM[4710] = 8'b0;
    XRAM[4711] = 8'b0;
    XRAM[4712] = 8'b0;
    XRAM[4713] = 8'b0;
    XRAM[4714] = 8'b0;
    XRAM[4715] = 8'b0;
    XRAM[4716] = 8'b0;
    XRAM[4717] = 8'b0;
    XRAM[4718] = 8'b0;
    XRAM[4719] = 8'b0;
    XRAM[4720] = 8'b0;
    XRAM[4721] = 8'b0;
    XRAM[4722] = 8'b0;
    XRAM[4723] = 8'b0;
    XRAM[4724] = 8'b0;
    XRAM[4725] = 8'b0;
    XRAM[4726] = 8'b0;
    XRAM[4727] = 8'b0;
    XRAM[4728] = 8'b0;
    XRAM[4729] = 8'b0;
    XRAM[4730] = 8'b0;
    XRAM[4731] = 8'b0;
    XRAM[4732] = 8'b0;
    XRAM[4733] = 8'b0;
    XRAM[4734] = 8'b0;
    XRAM[4735] = 8'b0;
    XRAM[4736] = 8'b0;
    XRAM[4737] = 8'b0;
    XRAM[4738] = 8'b0;
    XRAM[4739] = 8'b0;
    XRAM[4740] = 8'b0;
    XRAM[4741] = 8'b0;
    XRAM[4742] = 8'b0;
    XRAM[4743] = 8'b0;
    XRAM[4744] = 8'b0;
    XRAM[4745] = 8'b0;
    XRAM[4746] = 8'b0;
    XRAM[4747] = 8'b0;
    XRAM[4748] = 8'b0;
    XRAM[4749] = 8'b0;
    XRAM[4750] = 8'b0;
    XRAM[4751] = 8'b0;
    XRAM[4752] = 8'b0;
    XRAM[4753] = 8'b0;
    XRAM[4754] = 8'b0;
    XRAM[4755] = 8'b0;
    XRAM[4756] = 8'b0;
    XRAM[4757] = 8'b0;
    XRAM[4758] = 8'b0;
    XRAM[4759] = 8'b0;
    XRAM[4760] = 8'b0;
    XRAM[4761] = 8'b0;
    XRAM[4762] = 8'b0;
    XRAM[4763] = 8'b0;
    XRAM[4764] = 8'b0;
    XRAM[4765] = 8'b0;
    XRAM[4766] = 8'b0;
    XRAM[4767] = 8'b0;
    XRAM[4768] = 8'b0;
    XRAM[4769] = 8'b0;
    XRAM[4770] = 8'b0;
    XRAM[4771] = 8'b0;
    XRAM[4772] = 8'b0;
    XRAM[4773] = 8'b0;
    XRAM[4774] = 8'b0;
    XRAM[4775] = 8'b0;
    XRAM[4776] = 8'b0;
    XRAM[4777] = 8'b0;
    XRAM[4778] = 8'b0;
    XRAM[4779] = 8'b0;
    XRAM[4780] = 8'b0;
    XRAM[4781] = 8'b0;
    XRAM[4782] = 8'b0;
    XRAM[4783] = 8'b0;
    XRAM[4784] = 8'b0;
    XRAM[4785] = 8'b0;
    XRAM[4786] = 8'b0;
    XRAM[4787] = 8'b0;
    XRAM[4788] = 8'b0;
    XRAM[4789] = 8'b0;
    XRAM[4790] = 8'b0;
    XRAM[4791] = 8'b0;
    XRAM[4792] = 8'b0;
    XRAM[4793] = 8'b0;
    XRAM[4794] = 8'b0;
    XRAM[4795] = 8'b0;
    XRAM[4796] = 8'b0;
    XRAM[4797] = 8'b0;
    XRAM[4798] = 8'b0;
    XRAM[4799] = 8'b0;
    XRAM[4800] = 8'b0;
    XRAM[4801] = 8'b0;
    XRAM[4802] = 8'b0;
    XRAM[4803] = 8'b0;
    XRAM[4804] = 8'b0;
    XRAM[4805] = 8'b0;
    XRAM[4806] = 8'b0;
    XRAM[4807] = 8'b0;
    XRAM[4808] = 8'b0;
    XRAM[4809] = 8'b0;
    XRAM[4810] = 8'b0;
    XRAM[4811] = 8'b0;
    XRAM[4812] = 8'b0;
    XRAM[4813] = 8'b0;
    XRAM[4814] = 8'b0;
    XRAM[4815] = 8'b0;
    XRAM[4816] = 8'b0;
    XRAM[4817] = 8'b0;
    XRAM[4818] = 8'b0;
    XRAM[4819] = 8'b0;
    XRAM[4820] = 8'b0;
    XRAM[4821] = 8'b0;
    XRAM[4822] = 8'b0;
    XRAM[4823] = 8'b0;
    XRAM[4824] = 8'b0;
    XRAM[4825] = 8'b0;
    XRAM[4826] = 8'b0;
    XRAM[4827] = 8'b0;
    XRAM[4828] = 8'b0;
    XRAM[4829] = 8'b0;
    XRAM[4830] = 8'b0;
    XRAM[4831] = 8'b0;
    XRAM[4832] = 8'b0;
    XRAM[4833] = 8'b0;
    XRAM[4834] = 8'b0;
    XRAM[4835] = 8'b0;
    XRAM[4836] = 8'b0;
    XRAM[4837] = 8'b0;
    XRAM[4838] = 8'b0;
    XRAM[4839] = 8'b0;
    XRAM[4840] = 8'b0;
    XRAM[4841] = 8'b0;
    XRAM[4842] = 8'b0;
    XRAM[4843] = 8'b0;
    XRAM[4844] = 8'b0;
    XRAM[4845] = 8'b0;
    XRAM[4846] = 8'b0;
    XRAM[4847] = 8'b0;
    XRAM[4848] = 8'b0;
    XRAM[4849] = 8'b0;
    XRAM[4850] = 8'b0;
    XRAM[4851] = 8'b0;
    XRAM[4852] = 8'b0;
    XRAM[4853] = 8'b0;
    XRAM[4854] = 8'b0;
    XRAM[4855] = 8'b0;
    XRAM[4856] = 8'b0;
    XRAM[4857] = 8'b0;
    XRAM[4858] = 8'b0;
    XRAM[4859] = 8'b0;
    XRAM[4860] = 8'b0;
    XRAM[4861] = 8'b0;
    XRAM[4862] = 8'b0;
    XRAM[4863] = 8'b0;
    XRAM[4864] = 8'b0;
    XRAM[4865] = 8'b0;
    XRAM[4866] = 8'b0;
    XRAM[4867] = 8'b0;
    XRAM[4868] = 8'b0;
    XRAM[4869] = 8'b0;
    XRAM[4870] = 8'b0;
    XRAM[4871] = 8'b0;
    XRAM[4872] = 8'b0;
    XRAM[4873] = 8'b0;
    XRAM[4874] = 8'b0;
    XRAM[4875] = 8'b0;
    XRAM[4876] = 8'b0;
    XRAM[4877] = 8'b0;
    XRAM[4878] = 8'b0;
    XRAM[4879] = 8'b0;
    XRAM[4880] = 8'b0;
    XRAM[4881] = 8'b0;
    XRAM[4882] = 8'b0;
    XRAM[4883] = 8'b0;
    XRAM[4884] = 8'b0;
    XRAM[4885] = 8'b0;
    XRAM[4886] = 8'b0;
    XRAM[4887] = 8'b0;
    XRAM[4888] = 8'b0;
    XRAM[4889] = 8'b0;
    XRAM[4890] = 8'b0;
    XRAM[4891] = 8'b0;
    XRAM[4892] = 8'b0;
    XRAM[4893] = 8'b0;
    XRAM[4894] = 8'b0;
    XRAM[4895] = 8'b0;
    XRAM[4896] = 8'b0;
    XRAM[4897] = 8'b0;
    XRAM[4898] = 8'b0;
    XRAM[4899] = 8'b0;
    XRAM[4900] = 8'b0;
    XRAM[4901] = 8'b0;
    XRAM[4902] = 8'b0;
    XRAM[4903] = 8'b0;
    XRAM[4904] = 8'b0;
    XRAM[4905] = 8'b0;
    XRAM[4906] = 8'b0;
    XRAM[4907] = 8'b0;
    XRAM[4908] = 8'b0;
    XRAM[4909] = 8'b0;
    XRAM[4910] = 8'b0;
    XRAM[4911] = 8'b0;
    XRAM[4912] = 8'b0;
    XRAM[4913] = 8'b0;
    XRAM[4914] = 8'b0;
    XRAM[4915] = 8'b0;
    XRAM[4916] = 8'b0;
    XRAM[4917] = 8'b0;
    XRAM[4918] = 8'b0;
    XRAM[4919] = 8'b0;
    XRAM[4920] = 8'b0;
    XRAM[4921] = 8'b0;
    XRAM[4922] = 8'b0;
    XRAM[4923] = 8'b0;
    XRAM[4924] = 8'b0;
    XRAM[4925] = 8'b0;
    XRAM[4926] = 8'b0;
    XRAM[4927] = 8'b0;
    XRAM[4928] = 8'b0;
    XRAM[4929] = 8'b0;
    XRAM[4930] = 8'b0;
    XRAM[4931] = 8'b0;
    XRAM[4932] = 8'b0;
    XRAM[4933] = 8'b0;
    XRAM[4934] = 8'b0;
    XRAM[4935] = 8'b0;
    XRAM[4936] = 8'b0;
    XRAM[4937] = 8'b0;
    XRAM[4938] = 8'b0;
    XRAM[4939] = 8'b0;
    XRAM[4940] = 8'b0;
    XRAM[4941] = 8'b0;
    XRAM[4942] = 8'b0;
    XRAM[4943] = 8'b0;
    XRAM[4944] = 8'b0;
    XRAM[4945] = 8'b0;
    XRAM[4946] = 8'b0;
    XRAM[4947] = 8'b0;
    XRAM[4948] = 8'b0;
    XRAM[4949] = 8'b0;
    XRAM[4950] = 8'b0;
    XRAM[4951] = 8'b0;
    XRAM[4952] = 8'b0;
    XRAM[4953] = 8'b0;
    XRAM[4954] = 8'b0;
    XRAM[4955] = 8'b0;
    XRAM[4956] = 8'b0;
    XRAM[4957] = 8'b0;
    XRAM[4958] = 8'b0;
    XRAM[4959] = 8'b0;
    XRAM[4960] = 8'b0;
    XRAM[4961] = 8'b0;
    XRAM[4962] = 8'b0;
    XRAM[4963] = 8'b0;
    XRAM[4964] = 8'b0;
    XRAM[4965] = 8'b0;
    XRAM[4966] = 8'b0;
    XRAM[4967] = 8'b0;
    XRAM[4968] = 8'b0;
    XRAM[4969] = 8'b0;
    XRAM[4970] = 8'b0;
    XRAM[4971] = 8'b0;
    XRAM[4972] = 8'b0;
    XRAM[4973] = 8'b0;
    XRAM[4974] = 8'b0;
    XRAM[4975] = 8'b0;
    XRAM[4976] = 8'b0;
    XRAM[4977] = 8'b0;
    XRAM[4978] = 8'b0;
    XRAM[4979] = 8'b0;
    XRAM[4980] = 8'b0;
    XRAM[4981] = 8'b0;
    XRAM[4982] = 8'b0;
    XRAM[4983] = 8'b0;
    XRAM[4984] = 8'b0;
    XRAM[4985] = 8'b0;
    XRAM[4986] = 8'b0;
    XRAM[4987] = 8'b0;
    XRAM[4988] = 8'b0;
    XRAM[4989] = 8'b0;
    XRAM[4990] = 8'b0;
    XRAM[4991] = 8'b0;
    XRAM[4992] = 8'b0;
    XRAM[4993] = 8'b0;
    XRAM[4994] = 8'b0;
    XRAM[4995] = 8'b0;
    XRAM[4996] = 8'b0;
    XRAM[4997] = 8'b0;
    XRAM[4998] = 8'b0;
    XRAM[4999] = 8'b0;
    XRAM[5000] = 8'b0;
    XRAM[5001] = 8'b0;
    XRAM[5002] = 8'b0;
    XRAM[5003] = 8'b0;
    XRAM[5004] = 8'b0;
    XRAM[5005] = 8'b0;
    XRAM[5006] = 8'b0;
    XRAM[5007] = 8'b0;
    XRAM[5008] = 8'b0;
    XRAM[5009] = 8'b0;
    XRAM[5010] = 8'b0;
    XRAM[5011] = 8'b0;
    XRAM[5012] = 8'b0;
    XRAM[5013] = 8'b0;
    XRAM[5014] = 8'b0;
    XRAM[5015] = 8'b0;
    XRAM[5016] = 8'b0;
    XRAM[5017] = 8'b0;
    XRAM[5018] = 8'b0;
    XRAM[5019] = 8'b0;
    XRAM[5020] = 8'b0;
    XRAM[5021] = 8'b0;
    XRAM[5022] = 8'b0;
    XRAM[5023] = 8'b0;
    XRAM[5024] = 8'b0;
    XRAM[5025] = 8'b0;
    XRAM[5026] = 8'b0;
    XRAM[5027] = 8'b0;
    XRAM[5028] = 8'b0;
    XRAM[5029] = 8'b0;
    XRAM[5030] = 8'b0;
    XRAM[5031] = 8'b0;
    XRAM[5032] = 8'b0;
    XRAM[5033] = 8'b0;
    XRAM[5034] = 8'b0;
    XRAM[5035] = 8'b0;
    XRAM[5036] = 8'b0;
    XRAM[5037] = 8'b0;
    XRAM[5038] = 8'b0;
    XRAM[5039] = 8'b0;
    XRAM[5040] = 8'b0;
    XRAM[5041] = 8'b0;
    XRAM[5042] = 8'b0;
    XRAM[5043] = 8'b0;
    XRAM[5044] = 8'b0;
    XRAM[5045] = 8'b0;
    XRAM[5046] = 8'b0;
    XRAM[5047] = 8'b0;
    XRAM[5048] = 8'b0;
    XRAM[5049] = 8'b0;
    XRAM[5050] = 8'b0;
    XRAM[5051] = 8'b0;
    XRAM[5052] = 8'b0;
    XRAM[5053] = 8'b0;
    XRAM[5054] = 8'b0;
    XRAM[5055] = 8'b0;
    XRAM[5056] = 8'b0;
    XRAM[5057] = 8'b0;
    XRAM[5058] = 8'b0;
    XRAM[5059] = 8'b0;
    XRAM[5060] = 8'b0;
    XRAM[5061] = 8'b0;
    XRAM[5062] = 8'b0;
    XRAM[5063] = 8'b0;
    XRAM[5064] = 8'b0;
    XRAM[5065] = 8'b0;
    XRAM[5066] = 8'b0;
    XRAM[5067] = 8'b0;
    XRAM[5068] = 8'b0;
    XRAM[5069] = 8'b0;
    XRAM[5070] = 8'b0;
    XRAM[5071] = 8'b0;
    XRAM[5072] = 8'b0;
    XRAM[5073] = 8'b0;
    XRAM[5074] = 8'b0;
    XRAM[5075] = 8'b0;
    XRAM[5076] = 8'b0;
    XRAM[5077] = 8'b0;
    XRAM[5078] = 8'b0;
    XRAM[5079] = 8'b0;
    XRAM[5080] = 8'b0;
    XRAM[5081] = 8'b0;
    XRAM[5082] = 8'b0;
    XRAM[5083] = 8'b0;
    XRAM[5084] = 8'b0;
    XRAM[5085] = 8'b0;
    XRAM[5086] = 8'b0;
    XRAM[5087] = 8'b0;
    XRAM[5088] = 8'b0;
    XRAM[5089] = 8'b0;
    XRAM[5090] = 8'b0;
    XRAM[5091] = 8'b0;
    XRAM[5092] = 8'b0;
    XRAM[5093] = 8'b0;
    XRAM[5094] = 8'b0;
    XRAM[5095] = 8'b0;
    XRAM[5096] = 8'b0;
    XRAM[5097] = 8'b0;
    XRAM[5098] = 8'b0;
    XRAM[5099] = 8'b0;
    XRAM[5100] = 8'b0;
    XRAM[5101] = 8'b0;
    XRAM[5102] = 8'b0;
    XRAM[5103] = 8'b0;
    XRAM[5104] = 8'b0;
    XRAM[5105] = 8'b0;
    XRAM[5106] = 8'b0;
    XRAM[5107] = 8'b0;
    XRAM[5108] = 8'b0;
    XRAM[5109] = 8'b0;
    XRAM[5110] = 8'b0;
    XRAM[5111] = 8'b0;
    XRAM[5112] = 8'b0;
    XRAM[5113] = 8'b0;
    XRAM[5114] = 8'b0;
    XRAM[5115] = 8'b0;
    XRAM[5116] = 8'b0;
    XRAM[5117] = 8'b0;
    XRAM[5118] = 8'b0;
    XRAM[5119] = 8'b0;
    XRAM[5120] = 8'b0;
    XRAM[5121] = 8'b0;
    XRAM[5122] = 8'b0;
    XRAM[5123] = 8'b0;
    XRAM[5124] = 8'b0;
    XRAM[5125] = 8'b0;
    XRAM[5126] = 8'b0;
    XRAM[5127] = 8'b0;
    XRAM[5128] = 8'b0;
    XRAM[5129] = 8'b0;
    XRAM[5130] = 8'b0;
    XRAM[5131] = 8'b0;
    XRAM[5132] = 8'b0;
    XRAM[5133] = 8'b0;
    XRAM[5134] = 8'b0;
    XRAM[5135] = 8'b0;
    XRAM[5136] = 8'b0;
    XRAM[5137] = 8'b0;
    XRAM[5138] = 8'b0;
    XRAM[5139] = 8'b0;
    XRAM[5140] = 8'b0;
    XRAM[5141] = 8'b0;
    XRAM[5142] = 8'b0;
    XRAM[5143] = 8'b0;
    XRAM[5144] = 8'b0;
    XRAM[5145] = 8'b0;
    XRAM[5146] = 8'b0;
    XRAM[5147] = 8'b0;
    XRAM[5148] = 8'b0;
    XRAM[5149] = 8'b0;
    XRAM[5150] = 8'b0;
    XRAM[5151] = 8'b0;
    XRAM[5152] = 8'b0;
    XRAM[5153] = 8'b0;
    XRAM[5154] = 8'b0;
    XRAM[5155] = 8'b0;
    XRAM[5156] = 8'b0;
    XRAM[5157] = 8'b0;
    XRAM[5158] = 8'b0;
    XRAM[5159] = 8'b0;
    XRAM[5160] = 8'b0;
    XRAM[5161] = 8'b0;
    XRAM[5162] = 8'b0;
    XRAM[5163] = 8'b0;
    XRAM[5164] = 8'b0;
    XRAM[5165] = 8'b0;
    XRAM[5166] = 8'b0;
    XRAM[5167] = 8'b0;
    XRAM[5168] = 8'b0;
    XRAM[5169] = 8'b0;
    XRAM[5170] = 8'b0;
    XRAM[5171] = 8'b0;
    XRAM[5172] = 8'b0;
    XRAM[5173] = 8'b0;
    XRAM[5174] = 8'b0;
    XRAM[5175] = 8'b0;
    XRAM[5176] = 8'b0;
    XRAM[5177] = 8'b0;
    XRAM[5178] = 8'b0;
    XRAM[5179] = 8'b0;
    XRAM[5180] = 8'b0;
    XRAM[5181] = 8'b0;
    XRAM[5182] = 8'b0;
    XRAM[5183] = 8'b0;
    XRAM[5184] = 8'b0;
    XRAM[5185] = 8'b0;
    XRAM[5186] = 8'b0;
    XRAM[5187] = 8'b0;
    XRAM[5188] = 8'b0;
    XRAM[5189] = 8'b0;
    XRAM[5190] = 8'b0;
    XRAM[5191] = 8'b0;
    XRAM[5192] = 8'b0;
    XRAM[5193] = 8'b0;
    XRAM[5194] = 8'b0;
    XRAM[5195] = 8'b0;
    XRAM[5196] = 8'b0;
    XRAM[5197] = 8'b0;
    XRAM[5198] = 8'b0;
    XRAM[5199] = 8'b0;
    XRAM[5200] = 8'b0;
    XRAM[5201] = 8'b0;
    XRAM[5202] = 8'b0;
    XRAM[5203] = 8'b0;
    XRAM[5204] = 8'b0;
    XRAM[5205] = 8'b0;
    XRAM[5206] = 8'b0;
    XRAM[5207] = 8'b0;
    XRAM[5208] = 8'b0;
    XRAM[5209] = 8'b0;
    XRAM[5210] = 8'b0;
    XRAM[5211] = 8'b0;
    XRAM[5212] = 8'b0;
    XRAM[5213] = 8'b0;
    XRAM[5214] = 8'b0;
    XRAM[5215] = 8'b0;
    XRAM[5216] = 8'b0;
    XRAM[5217] = 8'b0;
    XRAM[5218] = 8'b0;
    XRAM[5219] = 8'b0;
    XRAM[5220] = 8'b0;
    XRAM[5221] = 8'b0;
    XRAM[5222] = 8'b0;
    XRAM[5223] = 8'b0;
    XRAM[5224] = 8'b0;
    XRAM[5225] = 8'b0;
    XRAM[5226] = 8'b0;
    XRAM[5227] = 8'b0;
    XRAM[5228] = 8'b0;
    XRAM[5229] = 8'b0;
    XRAM[5230] = 8'b0;
    XRAM[5231] = 8'b0;
    XRAM[5232] = 8'b0;
    XRAM[5233] = 8'b0;
    XRAM[5234] = 8'b0;
    XRAM[5235] = 8'b0;
    XRAM[5236] = 8'b0;
    XRAM[5237] = 8'b0;
    XRAM[5238] = 8'b0;
    XRAM[5239] = 8'b0;
    XRAM[5240] = 8'b0;
    XRAM[5241] = 8'b0;
    XRAM[5242] = 8'b0;
    XRAM[5243] = 8'b0;
    XRAM[5244] = 8'b0;
    XRAM[5245] = 8'b0;
    XRAM[5246] = 8'b0;
    XRAM[5247] = 8'b0;
    XRAM[5248] = 8'b0;
    XRAM[5249] = 8'b0;
    XRAM[5250] = 8'b0;
    XRAM[5251] = 8'b0;
    XRAM[5252] = 8'b0;
    XRAM[5253] = 8'b0;
    XRAM[5254] = 8'b0;
    XRAM[5255] = 8'b0;
    XRAM[5256] = 8'b0;
    XRAM[5257] = 8'b0;
    XRAM[5258] = 8'b0;
    XRAM[5259] = 8'b0;
    XRAM[5260] = 8'b0;
    XRAM[5261] = 8'b0;
    XRAM[5262] = 8'b0;
    XRAM[5263] = 8'b0;
    XRAM[5264] = 8'b0;
    XRAM[5265] = 8'b0;
    XRAM[5266] = 8'b0;
    XRAM[5267] = 8'b0;
    XRAM[5268] = 8'b0;
    XRAM[5269] = 8'b0;
    XRAM[5270] = 8'b0;
    XRAM[5271] = 8'b0;
    XRAM[5272] = 8'b0;
    XRAM[5273] = 8'b0;
    XRAM[5274] = 8'b0;
    XRAM[5275] = 8'b0;
    XRAM[5276] = 8'b0;
    XRAM[5277] = 8'b0;
    XRAM[5278] = 8'b0;
    XRAM[5279] = 8'b0;
    XRAM[5280] = 8'b0;
    XRAM[5281] = 8'b0;
    XRAM[5282] = 8'b0;
    XRAM[5283] = 8'b0;
    XRAM[5284] = 8'b0;
    XRAM[5285] = 8'b0;
    XRAM[5286] = 8'b0;
    XRAM[5287] = 8'b0;
    XRAM[5288] = 8'b0;
    XRAM[5289] = 8'b0;
    XRAM[5290] = 8'b0;
    XRAM[5291] = 8'b0;
    XRAM[5292] = 8'b0;
    XRAM[5293] = 8'b0;
    XRAM[5294] = 8'b0;
    XRAM[5295] = 8'b0;
    XRAM[5296] = 8'b0;
    XRAM[5297] = 8'b0;
    XRAM[5298] = 8'b0;
    XRAM[5299] = 8'b0;
    XRAM[5300] = 8'b0;
    XRAM[5301] = 8'b0;
    XRAM[5302] = 8'b0;
    XRAM[5303] = 8'b0;
    XRAM[5304] = 8'b0;
    XRAM[5305] = 8'b0;
    XRAM[5306] = 8'b0;
    XRAM[5307] = 8'b0;
    XRAM[5308] = 8'b0;
    XRAM[5309] = 8'b0;
    XRAM[5310] = 8'b0;
    XRAM[5311] = 8'b0;
    XRAM[5312] = 8'b0;
    XRAM[5313] = 8'b0;
    XRAM[5314] = 8'b0;
    XRAM[5315] = 8'b0;
    XRAM[5316] = 8'b0;
    XRAM[5317] = 8'b0;
    XRAM[5318] = 8'b0;
    XRAM[5319] = 8'b0;
    XRAM[5320] = 8'b0;
    XRAM[5321] = 8'b0;
    XRAM[5322] = 8'b0;
    XRAM[5323] = 8'b0;
    XRAM[5324] = 8'b0;
    XRAM[5325] = 8'b0;
    XRAM[5326] = 8'b0;
    XRAM[5327] = 8'b0;
    XRAM[5328] = 8'b0;
    XRAM[5329] = 8'b0;
    XRAM[5330] = 8'b0;
    XRAM[5331] = 8'b0;
    XRAM[5332] = 8'b0;
    XRAM[5333] = 8'b0;
    XRAM[5334] = 8'b0;
    XRAM[5335] = 8'b0;
    XRAM[5336] = 8'b0;
    XRAM[5337] = 8'b0;
    XRAM[5338] = 8'b0;
    XRAM[5339] = 8'b0;
    XRAM[5340] = 8'b0;
    XRAM[5341] = 8'b0;
    XRAM[5342] = 8'b0;
    XRAM[5343] = 8'b0;
    XRAM[5344] = 8'b0;
    XRAM[5345] = 8'b0;
    XRAM[5346] = 8'b0;
    XRAM[5347] = 8'b0;
    XRAM[5348] = 8'b0;
    XRAM[5349] = 8'b0;
    XRAM[5350] = 8'b0;
    XRAM[5351] = 8'b0;
    XRAM[5352] = 8'b0;
    XRAM[5353] = 8'b0;
    XRAM[5354] = 8'b0;
    XRAM[5355] = 8'b0;
    XRAM[5356] = 8'b0;
    XRAM[5357] = 8'b0;
    XRAM[5358] = 8'b0;
    XRAM[5359] = 8'b0;
    XRAM[5360] = 8'b0;
    XRAM[5361] = 8'b0;
    XRAM[5362] = 8'b0;
    XRAM[5363] = 8'b0;
    XRAM[5364] = 8'b0;
    XRAM[5365] = 8'b0;
    XRAM[5366] = 8'b0;
    XRAM[5367] = 8'b0;
    XRAM[5368] = 8'b0;
    XRAM[5369] = 8'b0;
    XRAM[5370] = 8'b0;
    XRAM[5371] = 8'b0;
    XRAM[5372] = 8'b0;
    XRAM[5373] = 8'b0;
    XRAM[5374] = 8'b0;
    XRAM[5375] = 8'b0;
    XRAM[5376] = 8'b0;
    XRAM[5377] = 8'b0;
    XRAM[5378] = 8'b0;
    XRAM[5379] = 8'b0;
    XRAM[5380] = 8'b0;
    XRAM[5381] = 8'b0;
    XRAM[5382] = 8'b0;
    XRAM[5383] = 8'b0;
    XRAM[5384] = 8'b0;
    XRAM[5385] = 8'b0;
    XRAM[5386] = 8'b0;
    XRAM[5387] = 8'b0;
    XRAM[5388] = 8'b0;
    XRAM[5389] = 8'b0;
    XRAM[5390] = 8'b0;
    XRAM[5391] = 8'b0;
    XRAM[5392] = 8'b0;
    XRAM[5393] = 8'b0;
    XRAM[5394] = 8'b0;
    XRAM[5395] = 8'b0;
    XRAM[5396] = 8'b0;
    XRAM[5397] = 8'b0;
    XRAM[5398] = 8'b0;
    XRAM[5399] = 8'b0;
    XRAM[5400] = 8'b0;
    XRAM[5401] = 8'b0;
    XRAM[5402] = 8'b0;
    XRAM[5403] = 8'b0;
    XRAM[5404] = 8'b0;
    XRAM[5405] = 8'b0;
    XRAM[5406] = 8'b0;
    XRAM[5407] = 8'b0;
    XRAM[5408] = 8'b0;
    XRAM[5409] = 8'b0;
    XRAM[5410] = 8'b0;
    XRAM[5411] = 8'b0;
    XRAM[5412] = 8'b0;
    XRAM[5413] = 8'b0;
    XRAM[5414] = 8'b0;
    XRAM[5415] = 8'b0;
    XRAM[5416] = 8'b0;
    XRAM[5417] = 8'b0;
    XRAM[5418] = 8'b0;
    XRAM[5419] = 8'b0;
    XRAM[5420] = 8'b0;
    XRAM[5421] = 8'b0;
    XRAM[5422] = 8'b0;
    XRAM[5423] = 8'b0;
    XRAM[5424] = 8'b0;
    XRAM[5425] = 8'b0;
    XRAM[5426] = 8'b0;
    XRAM[5427] = 8'b0;
    XRAM[5428] = 8'b0;
    XRAM[5429] = 8'b0;
    XRAM[5430] = 8'b0;
    XRAM[5431] = 8'b0;
    XRAM[5432] = 8'b0;
    XRAM[5433] = 8'b0;
    XRAM[5434] = 8'b0;
    XRAM[5435] = 8'b0;
    XRAM[5436] = 8'b0;
    XRAM[5437] = 8'b0;
    XRAM[5438] = 8'b0;
    XRAM[5439] = 8'b0;
    XRAM[5440] = 8'b0;
    XRAM[5441] = 8'b0;
    XRAM[5442] = 8'b0;
    XRAM[5443] = 8'b0;
    XRAM[5444] = 8'b0;
    XRAM[5445] = 8'b0;
    XRAM[5446] = 8'b0;
    XRAM[5447] = 8'b0;
    XRAM[5448] = 8'b0;
    XRAM[5449] = 8'b0;
    XRAM[5450] = 8'b0;
    XRAM[5451] = 8'b0;
    XRAM[5452] = 8'b0;
    XRAM[5453] = 8'b0;
    XRAM[5454] = 8'b0;
    XRAM[5455] = 8'b0;
    XRAM[5456] = 8'b0;
    XRAM[5457] = 8'b0;
    XRAM[5458] = 8'b0;
    XRAM[5459] = 8'b0;
    XRAM[5460] = 8'b0;
    XRAM[5461] = 8'b0;
    XRAM[5462] = 8'b0;
    XRAM[5463] = 8'b0;
    XRAM[5464] = 8'b0;
    XRAM[5465] = 8'b0;
    XRAM[5466] = 8'b0;
    XRAM[5467] = 8'b0;
    XRAM[5468] = 8'b0;
    XRAM[5469] = 8'b0;
    XRAM[5470] = 8'b0;
    XRAM[5471] = 8'b0;
    XRAM[5472] = 8'b0;
    XRAM[5473] = 8'b0;
    XRAM[5474] = 8'b0;
    XRAM[5475] = 8'b0;
    XRAM[5476] = 8'b0;
    XRAM[5477] = 8'b0;
    XRAM[5478] = 8'b0;
    XRAM[5479] = 8'b0;
    XRAM[5480] = 8'b0;
    XRAM[5481] = 8'b0;
    XRAM[5482] = 8'b0;
    XRAM[5483] = 8'b0;
    XRAM[5484] = 8'b0;
    XRAM[5485] = 8'b0;
    XRAM[5486] = 8'b0;
    XRAM[5487] = 8'b0;
    XRAM[5488] = 8'b0;
    XRAM[5489] = 8'b0;
    XRAM[5490] = 8'b0;
    XRAM[5491] = 8'b0;
    XRAM[5492] = 8'b0;
    XRAM[5493] = 8'b0;
    XRAM[5494] = 8'b0;
    XRAM[5495] = 8'b0;
    XRAM[5496] = 8'b0;
    XRAM[5497] = 8'b0;
    XRAM[5498] = 8'b0;
    XRAM[5499] = 8'b0;
    XRAM[5500] = 8'b0;
    XRAM[5501] = 8'b0;
    XRAM[5502] = 8'b0;
    XRAM[5503] = 8'b0;
    XRAM[5504] = 8'b0;
    XRAM[5505] = 8'b0;
    XRAM[5506] = 8'b0;
    XRAM[5507] = 8'b0;
    XRAM[5508] = 8'b0;
    XRAM[5509] = 8'b0;
    XRAM[5510] = 8'b0;
    XRAM[5511] = 8'b0;
    XRAM[5512] = 8'b0;
    XRAM[5513] = 8'b0;
    XRAM[5514] = 8'b0;
    XRAM[5515] = 8'b0;
    XRAM[5516] = 8'b0;
    XRAM[5517] = 8'b0;
    XRAM[5518] = 8'b0;
    XRAM[5519] = 8'b0;
    XRAM[5520] = 8'b0;
    XRAM[5521] = 8'b0;
    XRAM[5522] = 8'b0;
    XRAM[5523] = 8'b0;
    XRAM[5524] = 8'b0;
    XRAM[5525] = 8'b0;
    XRAM[5526] = 8'b0;
    XRAM[5527] = 8'b0;
    XRAM[5528] = 8'b0;
    XRAM[5529] = 8'b0;
    XRAM[5530] = 8'b0;
    XRAM[5531] = 8'b0;
    XRAM[5532] = 8'b0;
    XRAM[5533] = 8'b0;
    XRAM[5534] = 8'b0;
    XRAM[5535] = 8'b0;
    XRAM[5536] = 8'b0;
    XRAM[5537] = 8'b0;
    XRAM[5538] = 8'b0;
    XRAM[5539] = 8'b0;
    XRAM[5540] = 8'b0;
    XRAM[5541] = 8'b0;
    XRAM[5542] = 8'b0;
    XRAM[5543] = 8'b0;
    XRAM[5544] = 8'b0;
    XRAM[5545] = 8'b0;
    XRAM[5546] = 8'b0;
    XRAM[5547] = 8'b0;
    XRAM[5548] = 8'b0;
    XRAM[5549] = 8'b0;
    XRAM[5550] = 8'b0;
    XRAM[5551] = 8'b0;
    XRAM[5552] = 8'b0;
    XRAM[5553] = 8'b0;
    XRAM[5554] = 8'b0;
    XRAM[5555] = 8'b0;
    XRAM[5556] = 8'b0;
    XRAM[5557] = 8'b0;
    XRAM[5558] = 8'b0;
    XRAM[5559] = 8'b0;
    XRAM[5560] = 8'b0;
    XRAM[5561] = 8'b0;
    XRAM[5562] = 8'b0;
    XRAM[5563] = 8'b0;
    XRAM[5564] = 8'b0;
    XRAM[5565] = 8'b0;
    XRAM[5566] = 8'b0;
    XRAM[5567] = 8'b0;
    XRAM[5568] = 8'b0;
    XRAM[5569] = 8'b0;
    XRAM[5570] = 8'b0;
    XRAM[5571] = 8'b0;
    XRAM[5572] = 8'b0;
    XRAM[5573] = 8'b0;
    XRAM[5574] = 8'b0;
    XRAM[5575] = 8'b0;
    XRAM[5576] = 8'b0;
    XRAM[5577] = 8'b0;
    XRAM[5578] = 8'b0;
    XRAM[5579] = 8'b0;
    XRAM[5580] = 8'b0;
    XRAM[5581] = 8'b0;
    XRAM[5582] = 8'b0;
    XRAM[5583] = 8'b0;
    XRAM[5584] = 8'b0;
    XRAM[5585] = 8'b0;
    XRAM[5586] = 8'b0;
    XRAM[5587] = 8'b0;
    XRAM[5588] = 8'b0;
    XRAM[5589] = 8'b0;
    XRAM[5590] = 8'b0;
    XRAM[5591] = 8'b0;
    XRAM[5592] = 8'b0;
    XRAM[5593] = 8'b0;
    XRAM[5594] = 8'b0;
    XRAM[5595] = 8'b0;
    XRAM[5596] = 8'b0;
    XRAM[5597] = 8'b0;
    XRAM[5598] = 8'b0;
    XRAM[5599] = 8'b0;
    XRAM[5600] = 8'b0;
    XRAM[5601] = 8'b0;
    XRAM[5602] = 8'b0;
    XRAM[5603] = 8'b0;
    XRAM[5604] = 8'b0;
    XRAM[5605] = 8'b0;
    XRAM[5606] = 8'b0;
    XRAM[5607] = 8'b0;
    XRAM[5608] = 8'b0;
    XRAM[5609] = 8'b0;
    XRAM[5610] = 8'b0;
    XRAM[5611] = 8'b0;
    XRAM[5612] = 8'b0;
    XRAM[5613] = 8'b0;
    XRAM[5614] = 8'b0;
    XRAM[5615] = 8'b0;
    XRAM[5616] = 8'b0;
    XRAM[5617] = 8'b0;
    XRAM[5618] = 8'b0;
    XRAM[5619] = 8'b0;
    XRAM[5620] = 8'b0;
    XRAM[5621] = 8'b0;
    XRAM[5622] = 8'b0;
    XRAM[5623] = 8'b0;
    XRAM[5624] = 8'b0;
    XRAM[5625] = 8'b0;
    XRAM[5626] = 8'b0;
    XRAM[5627] = 8'b0;
    XRAM[5628] = 8'b0;
    XRAM[5629] = 8'b0;
    XRAM[5630] = 8'b0;
    XRAM[5631] = 8'b0;
    XRAM[5632] = 8'b0;
    XRAM[5633] = 8'b0;
    XRAM[5634] = 8'b0;
    XRAM[5635] = 8'b0;
    XRAM[5636] = 8'b0;
    XRAM[5637] = 8'b0;
    XRAM[5638] = 8'b0;
    XRAM[5639] = 8'b0;
    XRAM[5640] = 8'b0;
    XRAM[5641] = 8'b0;
    XRAM[5642] = 8'b0;
    XRAM[5643] = 8'b0;
    XRAM[5644] = 8'b0;
    XRAM[5645] = 8'b0;
    XRAM[5646] = 8'b0;
    XRAM[5647] = 8'b0;
    XRAM[5648] = 8'b0;
    XRAM[5649] = 8'b0;
    XRAM[5650] = 8'b0;
    XRAM[5651] = 8'b0;
    XRAM[5652] = 8'b0;
    XRAM[5653] = 8'b0;
    XRAM[5654] = 8'b0;
    XRAM[5655] = 8'b0;
    XRAM[5656] = 8'b0;
    XRAM[5657] = 8'b0;
    XRAM[5658] = 8'b0;
    XRAM[5659] = 8'b0;
    XRAM[5660] = 8'b0;
    XRAM[5661] = 8'b0;
    XRAM[5662] = 8'b0;
    XRAM[5663] = 8'b0;
    XRAM[5664] = 8'b0;
    XRAM[5665] = 8'b0;
    XRAM[5666] = 8'b0;
    XRAM[5667] = 8'b0;
    XRAM[5668] = 8'b0;
    XRAM[5669] = 8'b0;
    XRAM[5670] = 8'b0;
    XRAM[5671] = 8'b0;
    XRAM[5672] = 8'b0;
    XRAM[5673] = 8'b0;
    XRAM[5674] = 8'b0;
    XRAM[5675] = 8'b0;
    XRAM[5676] = 8'b0;
    XRAM[5677] = 8'b0;
    XRAM[5678] = 8'b0;
    XRAM[5679] = 8'b0;
    XRAM[5680] = 8'b0;
    XRAM[5681] = 8'b0;
    XRAM[5682] = 8'b0;
    XRAM[5683] = 8'b0;
    XRAM[5684] = 8'b0;
    XRAM[5685] = 8'b0;
    XRAM[5686] = 8'b0;
    XRAM[5687] = 8'b0;
    XRAM[5688] = 8'b0;
    XRAM[5689] = 8'b0;
    XRAM[5690] = 8'b0;
    XRAM[5691] = 8'b0;
    XRAM[5692] = 8'b0;
    XRAM[5693] = 8'b0;
    XRAM[5694] = 8'b0;
    XRAM[5695] = 8'b0;
    XRAM[5696] = 8'b0;
    XRAM[5697] = 8'b0;
    XRAM[5698] = 8'b0;
    XRAM[5699] = 8'b0;
    XRAM[5700] = 8'b0;
    XRAM[5701] = 8'b0;
    XRAM[5702] = 8'b0;
    XRAM[5703] = 8'b0;
    XRAM[5704] = 8'b0;
    XRAM[5705] = 8'b0;
    XRAM[5706] = 8'b0;
    XRAM[5707] = 8'b0;
    XRAM[5708] = 8'b0;
    XRAM[5709] = 8'b0;
    XRAM[5710] = 8'b0;
    XRAM[5711] = 8'b0;
    XRAM[5712] = 8'b0;
    XRAM[5713] = 8'b0;
    XRAM[5714] = 8'b0;
    XRAM[5715] = 8'b0;
    XRAM[5716] = 8'b0;
    XRAM[5717] = 8'b0;
    XRAM[5718] = 8'b0;
    XRAM[5719] = 8'b0;
    XRAM[5720] = 8'b0;
    XRAM[5721] = 8'b0;
    XRAM[5722] = 8'b0;
    XRAM[5723] = 8'b0;
    XRAM[5724] = 8'b0;
    XRAM[5725] = 8'b0;
    XRAM[5726] = 8'b0;
    XRAM[5727] = 8'b0;
    XRAM[5728] = 8'b0;
    XRAM[5729] = 8'b0;
    XRAM[5730] = 8'b0;
    XRAM[5731] = 8'b0;
    XRAM[5732] = 8'b0;
    XRAM[5733] = 8'b0;
    XRAM[5734] = 8'b0;
    XRAM[5735] = 8'b0;
    XRAM[5736] = 8'b0;
    XRAM[5737] = 8'b0;
    XRAM[5738] = 8'b0;
    XRAM[5739] = 8'b0;
    XRAM[5740] = 8'b0;
    XRAM[5741] = 8'b0;
    XRAM[5742] = 8'b0;
    XRAM[5743] = 8'b0;
    XRAM[5744] = 8'b0;
    XRAM[5745] = 8'b0;
    XRAM[5746] = 8'b0;
    XRAM[5747] = 8'b0;
    XRAM[5748] = 8'b0;
    XRAM[5749] = 8'b0;
    XRAM[5750] = 8'b0;
    XRAM[5751] = 8'b0;
    XRAM[5752] = 8'b0;
    XRAM[5753] = 8'b0;
    XRAM[5754] = 8'b0;
    XRAM[5755] = 8'b0;
    XRAM[5756] = 8'b0;
    XRAM[5757] = 8'b0;
    XRAM[5758] = 8'b0;
    XRAM[5759] = 8'b0;
    XRAM[5760] = 8'b0;
    XRAM[5761] = 8'b0;
    XRAM[5762] = 8'b0;
    XRAM[5763] = 8'b0;
    XRAM[5764] = 8'b0;
    XRAM[5765] = 8'b0;
    XRAM[5766] = 8'b0;
    XRAM[5767] = 8'b0;
    XRAM[5768] = 8'b0;
    XRAM[5769] = 8'b0;
    XRAM[5770] = 8'b0;
    XRAM[5771] = 8'b0;
    XRAM[5772] = 8'b0;
    XRAM[5773] = 8'b0;
    XRAM[5774] = 8'b0;
    XRAM[5775] = 8'b0;
    XRAM[5776] = 8'b0;
    XRAM[5777] = 8'b0;
    XRAM[5778] = 8'b0;
    XRAM[5779] = 8'b0;
    XRAM[5780] = 8'b0;
    XRAM[5781] = 8'b0;
    XRAM[5782] = 8'b0;
    XRAM[5783] = 8'b0;
    XRAM[5784] = 8'b0;
    XRAM[5785] = 8'b0;
    XRAM[5786] = 8'b0;
    XRAM[5787] = 8'b0;
    XRAM[5788] = 8'b0;
    XRAM[5789] = 8'b0;
    XRAM[5790] = 8'b0;
    XRAM[5791] = 8'b0;
    XRAM[5792] = 8'b0;
    XRAM[5793] = 8'b0;
    XRAM[5794] = 8'b0;
    XRAM[5795] = 8'b0;
    XRAM[5796] = 8'b0;
    XRAM[5797] = 8'b0;
    XRAM[5798] = 8'b0;
    XRAM[5799] = 8'b0;
    XRAM[5800] = 8'b0;
    XRAM[5801] = 8'b0;
    XRAM[5802] = 8'b0;
    XRAM[5803] = 8'b0;
    XRAM[5804] = 8'b0;
    XRAM[5805] = 8'b0;
    XRAM[5806] = 8'b0;
    XRAM[5807] = 8'b0;
    XRAM[5808] = 8'b0;
    XRAM[5809] = 8'b0;
    XRAM[5810] = 8'b0;
    XRAM[5811] = 8'b0;
    XRAM[5812] = 8'b0;
    XRAM[5813] = 8'b0;
    XRAM[5814] = 8'b0;
    XRAM[5815] = 8'b0;
    XRAM[5816] = 8'b0;
    XRAM[5817] = 8'b0;
    XRAM[5818] = 8'b0;
    XRAM[5819] = 8'b0;
    XRAM[5820] = 8'b0;
    XRAM[5821] = 8'b0;
    XRAM[5822] = 8'b0;
    XRAM[5823] = 8'b0;
    XRAM[5824] = 8'b0;
    XRAM[5825] = 8'b0;
    XRAM[5826] = 8'b0;
    XRAM[5827] = 8'b0;
    XRAM[5828] = 8'b0;
    XRAM[5829] = 8'b0;
    XRAM[5830] = 8'b0;
    XRAM[5831] = 8'b0;
    XRAM[5832] = 8'b0;
    XRAM[5833] = 8'b0;
    XRAM[5834] = 8'b0;
    XRAM[5835] = 8'b0;
    XRAM[5836] = 8'b0;
    XRAM[5837] = 8'b0;
    XRAM[5838] = 8'b0;
    XRAM[5839] = 8'b0;
    XRAM[5840] = 8'b0;
    XRAM[5841] = 8'b0;
    XRAM[5842] = 8'b0;
    XRAM[5843] = 8'b0;
    XRAM[5844] = 8'b0;
    XRAM[5845] = 8'b0;
    XRAM[5846] = 8'b0;
    XRAM[5847] = 8'b0;
    XRAM[5848] = 8'b0;
    XRAM[5849] = 8'b0;
    XRAM[5850] = 8'b0;
    XRAM[5851] = 8'b0;
    XRAM[5852] = 8'b0;
    XRAM[5853] = 8'b0;
    XRAM[5854] = 8'b0;
    XRAM[5855] = 8'b0;
    XRAM[5856] = 8'b0;
    XRAM[5857] = 8'b0;
    XRAM[5858] = 8'b0;
    XRAM[5859] = 8'b0;
    XRAM[5860] = 8'b0;
    XRAM[5861] = 8'b0;
    XRAM[5862] = 8'b0;
    XRAM[5863] = 8'b0;
    XRAM[5864] = 8'b0;
    XRAM[5865] = 8'b0;
    XRAM[5866] = 8'b0;
    XRAM[5867] = 8'b0;
    XRAM[5868] = 8'b0;
    XRAM[5869] = 8'b0;
    XRAM[5870] = 8'b0;
    XRAM[5871] = 8'b0;
    XRAM[5872] = 8'b0;
    XRAM[5873] = 8'b0;
    XRAM[5874] = 8'b0;
    XRAM[5875] = 8'b0;
    XRAM[5876] = 8'b0;
    XRAM[5877] = 8'b0;
    XRAM[5878] = 8'b0;
    XRAM[5879] = 8'b0;
    XRAM[5880] = 8'b0;
    XRAM[5881] = 8'b0;
    XRAM[5882] = 8'b0;
    XRAM[5883] = 8'b0;
    XRAM[5884] = 8'b0;
    XRAM[5885] = 8'b0;
    XRAM[5886] = 8'b0;
    XRAM[5887] = 8'b0;
    XRAM[5888] = 8'b0;
    XRAM[5889] = 8'b0;
    XRAM[5890] = 8'b0;
    XRAM[5891] = 8'b0;
    XRAM[5892] = 8'b0;
    XRAM[5893] = 8'b0;
    XRAM[5894] = 8'b0;
    XRAM[5895] = 8'b0;
    XRAM[5896] = 8'b0;
    XRAM[5897] = 8'b0;
    XRAM[5898] = 8'b0;
    XRAM[5899] = 8'b0;
    XRAM[5900] = 8'b0;
    XRAM[5901] = 8'b0;
    XRAM[5902] = 8'b0;
    XRAM[5903] = 8'b0;
    XRAM[5904] = 8'b0;
    XRAM[5905] = 8'b0;
    XRAM[5906] = 8'b0;
    XRAM[5907] = 8'b0;
    XRAM[5908] = 8'b0;
    XRAM[5909] = 8'b0;
    XRAM[5910] = 8'b0;
    XRAM[5911] = 8'b0;
    XRAM[5912] = 8'b0;
    XRAM[5913] = 8'b0;
    XRAM[5914] = 8'b0;
    XRAM[5915] = 8'b0;
    XRAM[5916] = 8'b0;
    XRAM[5917] = 8'b0;
    XRAM[5918] = 8'b0;
    XRAM[5919] = 8'b0;
    XRAM[5920] = 8'b0;
    XRAM[5921] = 8'b0;
    XRAM[5922] = 8'b0;
    XRAM[5923] = 8'b0;
    XRAM[5924] = 8'b0;
    XRAM[5925] = 8'b0;
    XRAM[5926] = 8'b0;
    XRAM[5927] = 8'b0;
    XRAM[5928] = 8'b0;
    XRAM[5929] = 8'b0;
    XRAM[5930] = 8'b0;
    XRAM[5931] = 8'b0;
    XRAM[5932] = 8'b0;
    XRAM[5933] = 8'b0;
    XRAM[5934] = 8'b0;
    XRAM[5935] = 8'b0;
    XRAM[5936] = 8'b0;
    XRAM[5937] = 8'b0;
    XRAM[5938] = 8'b0;
    XRAM[5939] = 8'b0;
    XRAM[5940] = 8'b0;
    XRAM[5941] = 8'b0;
    XRAM[5942] = 8'b0;
    XRAM[5943] = 8'b0;
    XRAM[5944] = 8'b0;
    XRAM[5945] = 8'b0;
    XRAM[5946] = 8'b0;
    XRAM[5947] = 8'b0;
    XRAM[5948] = 8'b0;
    XRAM[5949] = 8'b0;
    XRAM[5950] = 8'b0;
    XRAM[5951] = 8'b0;
    XRAM[5952] = 8'b0;
    XRAM[5953] = 8'b0;
    XRAM[5954] = 8'b0;
    XRAM[5955] = 8'b0;
    XRAM[5956] = 8'b0;
    XRAM[5957] = 8'b0;
    XRAM[5958] = 8'b0;
    XRAM[5959] = 8'b0;
    XRAM[5960] = 8'b0;
    XRAM[5961] = 8'b0;
    XRAM[5962] = 8'b0;
    XRAM[5963] = 8'b0;
    XRAM[5964] = 8'b0;
    XRAM[5965] = 8'b0;
    XRAM[5966] = 8'b0;
    XRAM[5967] = 8'b0;
    XRAM[5968] = 8'b0;
    XRAM[5969] = 8'b0;
    XRAM[5970] = 8'b0;
    XRAM[5971] = 8'b0;
    XRAM[5972] = 8'b0;
    XRAM[5973] = 8'b0;
    XRAM[5974] = 8'b0;
    XRAM[5975] = 8'b0;
    XRAM[5976] = 8'b0;
    XRAM[5977] = 8'b0;
    XRAM[5978] = 8'b0;
    XRAM[5979] = 8'b0;
    XRAM[5980] = 8'b0;
    XRAM[5981] = 8'b0;
    XRAM[5982] = 8'b0;
    XRAM[5983] = 8'b0;
    XRAM[5984] = 8'b0;
    XRAM[5985] = 8'b0;
    XRAM[5986] = 8'b0;
    XRAM[5987] = 8'b0;
    XRAM[5988] = 8'b0;
    XRAM[5989] = 8'b0;
    XRAM[5990] = 8'b0;
    XRAM[5991] = 8'b0;
    XRAM[5992] = 8'b0;
    XRAM[5993] = 8'b0;
    XRAM[5994] = 8'b0;
    XRAM[5995] = 8'b0;
    XRAM[5996] = 8'b0;
    XRAM[5997] = 8'b0;
    XRAM[5998] = 8'b0;
    XRAM[5999] = 8'b0;
    XRAM[6000] = 8'b0;
    XRAM[6001] = 8'b0;
    XRAM[6002] = 8'b0;
    XRAM[6003] = 8'b0;
    XRAM[6004] = 8'b0;
    XRAM[6005] = 8'b0;
    XRAM[6006] = 8'b0;
    XRAM[6007] = 8'b0;
    XRAM[6008] = 8'b0;
    XRAM[6009] = 8'b0;
    XRAM[6010] = 8'b0;
    XRAM[6011] = 8'b0;
    XRAM[6012] = 8'b0;
    XRAM[6013] = 8'b0;
    XRAM[6014] = 8'b0;
    XRAM[6015] = 8'b0;
    XRAM[6016] = 8'b0;
    XRAM[6017] = 8'b0;
    XRAM[6018] = 8'b0;
    XRAM[6019] = 8'b0;
    XRAM[6020] = 8'b0;
    XRAM[6021] = 8'b0;
    XRAM[6022] = 8'b0;
    XRAM[6023] = 8'b0;
    XRAM[6024] = 8'b0;
    XRAM[6025] = 8'b0;
    XRAM[6026] = 8'b0;
    XRAM[6027] = 8'b0;
    XRAM[6028] = 8'b0;
    XRAM[6029] = 8'b0;
    XRAM[6030] = 8'b0;
    XRAM[6031] = 8'b0;
    XRAM[6032] = 8'b0;
    XRAM[6033] = 8'b0;
    XRAM[6034] = 8'b0;
    XRAM[6035] = 8'b0;
    XRAM[6036] = 8'b0;
    XRAM[6037] = 8'b0;
    XRAM[6038] = 8'b0;
    XRAM[6039] = 8'b0;
    XRAM[6040] = 8'b0;
    XRAM[6041] = 8'b0;
    XRAM[6042] = 8'b0;
    XRAM[6043] = 8'b0;
    XRAM[6044] = 8'b0;
    XRAM[6045] = 8'b0;
    XRAM[6046] = 8'b0;
    XRAM[6047] = 8'b0;
    XRAM[6048] = 8'b0;
    XRAM[6049] = 8'b0;
    XRAM[6050] = 8'b0;
    XRAM[6051] = 8'b0;
    XRAM[6052] = 8'b0;
    XRAM[6053] = 8'b0;
    XRAM[6054] = 8'b0;
    XRAM[6055] = 8'b0;
    XRAM[6056] = 8'b0;
    XRAM[6057] = 8'b0;
    XRAM[6058] = 8'b0;
    XRAM[6059] = 8'b0;
    XRAM[6060] = 8'b0;
    XRAM[6061] = 8'b0;
    XRAM[6062] = 8'b0;
    XRAM[6063] = 8'b0;
    XRAM[6064] = 8'b0;
    XRAM[6065] = 8'b0;
    XRAM[6066] = 8'b0;
    XRAM[6067] = 8'b0;
    XRAM[6068] = 8'b0;
    XRAM[6069] = 8'b0;
    XRAM[6070] = 8'b0;
    XRAM[6071] = 8'b0;
    XRAM[6072] = 8'b0;
    XRAM[6073] = 8'b0;
    XRAM[6074] = 8'b0;
    XRAM[6075] = 8'b0;
    XRAM[6076] = 8'b0;
    XRAM[6077] = 8'b0;
    XRAM[6078] = 8'b0;
    XRAM[6079] = 8'b0;
    XRAM[6080] = 8'b0;
    XRAM[6081] = 8'b0;
    XRAM[6082] = 8'b0;
    XRAM[6083] = 8'b0;
    XRAM[6084] = 8'b0;
    XRAM[6085] = 8'b0;
    XRAM[6086] = 8'b0;
    XRAM[6087] = 8'b0;
    XRAM[6088] = 8'b0;
    XRAM[6089] = 8'b0;
    XRAM[6090] = 8'b0;
    XRAM[6091] = 8'b0;
    XRAM[6092] = 8'b0;
    XRAM[6093] = 8'b0;
    XRAM[6094] = 8'b0;
    XRAM[6095] = 8'b0;
    XRAM[6096] = 8'b0;
    XRAM[6097] = 8'b0;
    XRAM[6098] = 8'b0;
    XRAM[6099] = 8'b0;
    XRAM[6100] = 8'b0;
    XRAM[6101] = 8'b0;
    XRAM[6102] = 8'b0;
    XRAM[6103] = 8'b0;
    XRAM[6104] = 8'b0;
    XRAM[6105] = 8'b0;
    XRAM[6106] = 8'b0;
    XRAM[6107] = 8'b0;
    XRAM[6108] = 8'b0;
    XRAM[6109] = 8'b0;
    XRAM[6110] = 8'b0;
    XRAM[6111] = 8'b0;
    XRAM[6112] = 8'b0;
    XRAM[6113] = 8'b0;
    XRAM[6114] = 8'b0;
    XRAM[6115] = 8'b0;
    XRAM[6116] = 8'b0;
    XRAM[6117] = 8'b0;
    XRAM[6118] = 8'b0;
    XRAM[6119] = 8'b0;
    XRAM[6120] = 8'b0;
    XRAM[6121] = 8'b0;
    XRAM[6122] = 8'b0;
    XRAM[6123] = 8'b0;
    XRAM[6124] = 8'b0;
    XRAM[6125] = 8'b0;
    XRAM[6126] = 8'b0;
    XRAM[6127] = 8'b0;
    XRAM[6128] = 8'b0;
    XRAM[6129] = 8'b0;
    XRAM[6130] = 8'b0;
    XRAM[6131] = 8'b0;
    XRAM[6132] = 8'b0;
    XRAM[6133] = 8'b0;
    XRAM[6134] = 8'b0;
    XRAM[6135] = 8'b0;
    XRAM[6136] = 8'b0;
    XRAM[6137] = 8'b0;
    XRAM[6138] = 8'b0;
    XRAM[6139] = 8'b0;
    XRAM[6140] = 8'b0;
    XRAM[6141] = 8'b0;
    XRAM[6142] = 8'b0;
    XRAM[6143] = 8'b0;
    XRAM[6144] = 8'b0;
    XRAM[6145] = 8'b0;
    XRAM[6146] = 8'b0;
    XRAM[6147] = 8'b0;
    XRAM[6148] = 8'b0;
    XRAM[6149] = 8'b0;
    XRAM[6150] = 8'b0;
    XRAM[6151] = 8'b0;
    XRAM[6152] = 8'b0;
    XRAM[6153] = 8'b0;
    XRAM[6154] = 8'b0;
    XRAM[6155] = 8'b0;
    XRAM[6156] = 8'b0;
    XRAM[6157] = 8'b0;
    XRAM[6158] = 8'b0;
    XRAM[6159] = 8'b0;
    XRAM[6160] = 8'b0;
    XRAM[6161] = 8'b0;
    XRAM[6162] = 8'b0;
    XRAM[6163] = 8'b0;
    XRAM[6164] = 8'b0;
    XRAM[6165] = 8'b0;
    XRAM[6166] = 8'b0;
    XRAM[6167] = 8'b0;
    XRAM[6168] = 8'b0;
    XRAM[6169] = 8'b0;
    XRAM[6170] = 8'b0;
    XRAM[6171] = 8'b0;
    XRAM[6172] = 8'b0;
    XRAM[6173] = 8'b0;
    XRAM[6174] = 8'b0;
    XRAM[6175] = 8'b0;
    XRAM[6176] = 8'b0;
    XRAM[6177] = 8'b0;
    XRAM[6178] = 8'b0;
    XRAM[6179] = 8'b0;
    XRAM[6180] = 8'b0;
    XRAM[6181] = 8'b0;
    XRAM[6182] = 8'b0;
    XRAM[6183] = 8'b0;
    XRAM[6184] = 8'b0;
    XRAM[6185] = 8'b0;
    XRAM[6186] = 8'b0;
    XRAM[6187] = 8'b0;
    XRAM[6188] = 8'b0;
    XRAM[6189] = 8'b0;
    XRAM[6190] = 8'b0;
    XRAM[6191] = 8'b0;
    XRAM[6192] = 8'b0;
    XRAM[6193] = 8'b0;
    XRAM[6194] = 8'b0;
    XRAM[6195] = 8'b0;
    XRAM[6196] = 8'b0;
    XRAM[6197] = 8'b0;
    XRAM[6198] = 8'b0;
    XRAM[6199] = 8'b0;
    XRAM[6200] = 8'b0;
    XRAM[6201] = 8'b0;
    XRAM[6202] = 8'b0;
    XRAM[6203] = 8'b0;
    XRAM[6204] = 8'b0;
    XRAM[6205] = 8'b0;
    XRAM[6206] = 8'b0;
    XRAM[6207] = 8'b0;
    XRAM[6208] = 8'b0;
    XRAM[6209] = 8'b0;
    XRAM[6210] = 8'b0;
    XRAM[6211] = 8'b0;
    XRAM[6212] = 8'b0;
    XRAM[6213] = 8'b0;
    XRAM[6214] = 8'b0;
    XRAM[6215] = 8'b0;
    XRAM[6216] = 8'b0;
    XRAM[6217] = 8'b0;
    XRAM[6218] = 8'b0;
    XRAM[6219] = 8'b0;
    XRAM[6220] = 8'b0;
    XRAM[6221] = 8'b0;
    XRAM[6222] = 8'b0;
    XRAM[6223] = 8'b0;
    XRAM[6224] = 8'b0;
    XRAM[6225] = 8'b0;
    XRAM[6226] = 8'b0;
    XRAM[6227] = 8'b0;
    XRAM[6228] = 8'b0;
    XRAM[6229] = 8'b0;
    XRAM[6230] = 8'b0;
    XRAM[6231] = 8'b0;
    XRAM[6232] = 8'b0;
    XRAM[6233] = 8'b0;
    XRAM[6234] = 8'b0;
    XRAM[6235] = 8'b0;
    XRAM[6236] = 8'b0;
    XRAM[6237] = 8'b0;
    XRAM[6238] = 8'b0;
    XRAM[6239] = 8'b0;
    XRAM[6240] = 8'b0;
    XRAM[6241] = 8'b0;
    XRAM[6242] = 8'b0;
    XRAM[6243] = 8'b0;
    XRAM[6244] = 8'b0;
    XRAM[6245] = 8'b0;
    XRAM[6246] = 8'b0;
    XRAM[6247] = 8'b0;
    XRAM[6248] = 8'b0;
    XRAM[6249] = 8'b0;
    XRAM[6250] = 8'b0;
    XRAM[6251] = 8'b0;
    XRAM[6252] = 8'b0;
    XRAM[6253] = 8'b0;
    XRAM[6254] = 8'b0;
    XRAM[6255] = 8'b0;
    XRAM[6256] = 8'b0;
    XRAM[6257] = 8'b0;
    XRAM[6258] = 8'b0;
    XRAM[6259] = 8'b0;
    XRAM[6260] = 8'b0;
    XRAM[6261] = 8'b0;
    XRAM[6262] = 8'b0;
    XRAM[6263] = 8'b0;
    XRAM[6264] = 8'b0;
    XRAM[6265] = 8'b0;
    XRAM[6266] = 8'b0;
    XRAM[6267] = 8'b0;
    XRAM[6268] = 8'b0;
    XRAM[6269] = 8'b0;
    XRAM[6270] = 8'b0;
    XRAM[6271] = 8'b0;
    XRAM[6272] = 8'b0;
    XRAM[6273] = 8'b0;
    XRAM[6274] = 8'b0;
    XRAM[6275] = 8'b0;
    XRAM[6276] = 8'b0;
    XRAM[6277] = 8'b0;
    XRAM[6278] = 8'b0;
    XRAM[6279] = 8'b0;
    XRAM[6280] = 8'b0;
    XRAM[6281] = 8'b0;
    XRAM[6282] = 8'b0;
    XRAM[6283] = 8'b0;
    XRAM[6284] = 8'b0;
    XRAM[6285] = 8'b0;
    XRAM[6286] = 8'b0;
    XRAM[6287] = 8'b0;
    XRAM[6288] = 8'b0;
    XRAM[6289] = 8'b0;
    XRAM[6290] = 8'b0;
    XRAM[6291] = 8'b0;
    XRAM[6292] = 8'b0;
    XRAM[6293] = 8'b0;
    XRAM[6294] = 8'b0;
    XRAM[6295] = 8'b0;
    XRAM[6296] = 8'b0;
    XRAM[6297] = 8'b0;
    XRAM[6298] = 8'b0;
    XRAM[6299] = 8'b0;
    XRAM[6300] = 8'b0;
    XRAM[6301] = 8'b0;
    XRAM[6302] = 8'b0;
    XRAM[6303] = 8'b0;
    XRAM[6304] = 8'b0;
    XRAM[6305] = 8'b0;
    XRAM[6306] = 8'b0;
    XRAM[6307] = 8'b0;
    XRAM[6308] = 8'b0;
    XRAM[6309] = 8'b0;
    XRAM[6310] = 8'b0;
    XRAM[6311] = 8'b0;
    XRAM[6312] = 8'b0;
    XRAM[6313] = 8'b0;
    XRAM[6314] = 8'b0;
    XRAM[6315] = 8'b0;
    XRAM[6316] = 8'b0;
    XRAM[6317] = 8'b0;
    XRAM[6318] = 8'b0;
    XRAM[6319] = 8'b0;
    XRAM[6320] = 8'b0;
    XRAM[6321] = 8'b0;
    XRAM[6322] = 8'b0;
    XRAM[6323] = 8'b0;
    XRAM[6324] = 8'b0;
    XRAM[6325] = 8'b0;
    XRAM[6326] = 8'b0;
    XRAM[6327] = 8'b0;
    XRAM[6328] = 8'b0;
    XRAM[6329] = 8'b0;
    XRAM[6330] = 8'b0;
    XRAM[6331] = 8'b0;
    XRAM[6332] = 8'b0;
    XRAM[6333] = 8'b0;
    XRAM[6334] = 8'b0;
    XRAM[6335] = 8'b0;
    XRAM[6336] = 8'b0;
    XRAM[6337] = 8'b0;
    XRAM[6338] = 8'b0;
    XRAM[6339] = 8'b0;
    XRAM[6340] = 8'b0;
    XRAM[6341] = 8'b0;
    XRAM[6342] = 8'b0;
    XRAM[6343] = 8'b0;
    XRAM[6344] = 8'b0;
    XRAM[6345] = 8'b0;
    XRAM[6346] = 8'b0;
    XRAM[6347] = 8'b0;
    XRAM[6348] = 8'b0;
    XRAM[6349] = 8'b0;
    XRAM[6350] = 8'b0;
    XRAM[6351] = 8'b0;
    XRAM[6352] = 8'b0;
    XRAM[6353] = 8'b0;
    XRAM[6354] = 8'b0;
    XRAM[6355] = 8'b0;
    XRAM[6356] = 8'b0;
    XRAM[6357] = 8'b0;
    XRAM[6358] = 8'b0;
    XRAM[6359] = 8'b0;
    XRAM[6360] = 8'b0;
    XRAM[6361] = 8'b0;
    XRAM[6362] = 8'b0;
    XRAM[6363] = 8'b0;
    XRAM[6364] = 8'b0;
    XRAM[6365] = 8'b0;
    XRAM[6366] = 8'b0;
    XRAM[6367] = 8'b0;
    XRAM[6368] = 8'b0;
    XRAM[6369] = 8'b0;
    XRAM[6370] = 8'b0;
    XRAM[6371] = 8'b0;
    XRAM[6372] = 8'b0;
    XRAM[6373] = 8'b0;
    XRAM[6374] = 8'b0;
    XRAM[6375] = 8'b0;
    XRAM[6376] = 8'b0;
    XRAM[6377] = 8'b0;
    XRAM[6378] = 8'b0;
    XRAM[6379] = 8'b0;
    XRAM[6380] = 8'b0;
    XRAM[6381] = 8'b0;
    XRAM[6382] = 8'b0;
    XRAM[6383] = 8'b0;
    XRAM[6384] = 8'b0;
    XRAM[6385] = 8'b0;
    XRAM[6386] = 8'b0;
    XRAM[6387] = 8'b0;
    XRAM[6388] = 8'b0;
    XRAM[6389] = 8'b0;
    XRAM[6390] = 8'b0;
    XRAM[6391] = 8'b0;
    XRAM[6392] = 8'b0;
    XRAM[6393] = 8'b0;
    XRAM[6394] = 8'b0;
    XRAM[6395] = 8'b0;
    XRAM[6396] = 8'b0;
    XRAM[6397] = 8'b0;
    XRAM[6398] = 8'b0;
    XRAM[6399] = 8'b0;
    XRAM[6400] = 8'b0;
    XRAM[6401] = 8'b0;
    XRAM[6402] = 8'b0;
    XRAM[6403] = 8'b0;
    XRAM[6404] = 8'b0;
    XRAM[6405] = 8'b0;
    XRAM[6406] = 8'b0;
    XRAM[6407] = 8'b0;
    XRAM[6408] = 8'b0;
    XRAM[6409] = 8'b0;
    XRAM[6410] = 8'b0;
    XRAM[6411] = 8'b0;
    XRAM[6412] = 8'b0;
    XRAM[6413] = 8'b0;
    XRAM[6414] = 8'b0;
    XRAM[6415] = 8'b0;
    XRAM[6416] = 8'b0;
    XRAM[6417] = 8'b0;
    XRAM[6418] = 8'b0;
    XRAM[6419] = 8'b0;
    XRAM[6420] = 8'b0;
    XRAM[6421] = 8'b0;
    XRAM[6422] = 8'b0;
    XRAM[6423] = 8'b0;
    XRAM[6424] = 8'b0;
    XRAM[6425] = 8'b0;
    XRAM[6426] = 8'b0;
    XRAM[6427] = 8'b0;
    XRAM[6428] = 8'b0;
    XRAM[6429] = 8'b0;
    XRAM[6430] = 8'b0;
    XRAM[6431] = 8'b0;
    XRAM[6432] = 8'b0;
    XRAM[6433] = 8'b0;
    XRAM[6434] = 8'b0;
    XRAM[6435] = 8'b0;
    XRAM[6436] = 8'b0;
    XRAM[6437] = 8'b0;
    XRAM[6438] = 8'b0;
    XRAM[6439] = 8'b0;
    XRAM[6440] = 8'b0;
    XRAM[6441] = 8'b0;
    XRAM[6442] = 8'b0;
    XRAM[6443] = 8'b0;
    XRAM[6444] = 8'b0;
    XRAM[6445] = 8'b0;
    XRAM[6446] = 8'b0;
    XRAM[6447] = 8'b0;
    XRAM[6448] = 8'b0;
    XRAM[6449] = 8'b0;
    XRAM[6450] = 8'b0;
    XRAM[6451] = 8'b0;
    XRAM[6452] = 8'b0;
    XRAM[6453] = 8'b0;
    XRAM[6454] = 8'b0;
    XRAM[6455] = 8'b0;
    XRAM[6456] = 8'b0;
    XRAM[6457] = 8'b0;
    XRAM[6458] = 8'b0;
    XRAM[6459] = 8'b0;
    XRAM[6460] = 8'b0;
    XRAM[6461] = 8'b0;
    XRAM[6462] = 8'b0;
    XRAM[6463] = 8'b0;
    XRAM[6464] = 8'b0;
    XRAM[6465] = 8'b0;
    XRAM[6466] = 8'b0;
    XRAM[6467] = 8'b0;
    XRAM[6468] = 8'b0;
    XRAM[6469] = 8'b0;
    XRAM[6470] = 8'b0;
    XRAM[6471] = 8'b0;
    XRAM[6472] = 8'b0;
    XRAM[6473] = 8'b0;
    XRAM[6474] = 8'b0;
    XRAM[6475] = 8'b0;
    XRAM[6476] = 8'b0;
    XRAM[6477] = 8'b0;
    XRAM[6478] = 8'b0;
    XRAM[6479] = 8'b0;
    XRAM[6480] = 8'b0;
    XRAM[6481] = 8'b0;
    XRAM[6482] = 8'b0;
    XRAM[6483] = 8'b0;
    XRAM[6484] = 8'b0;
    XRAM[6485] = 8'b0;
    XRAM[6486] = 8'b0;
    XRAM[6487] = 8'b0;
    XRAM[6488] = 8'b0;
    XRAM[6489] = 8'b0;
    XRAM[6490] = 8'b0;
    XRAM[6491] = 8'b0;
    XRAM[6492] = 8'b0;
    XRAM[6493] = 8'b0;
    XRAM[6494] = 8'b0;
    XRAM[6495] = 8'b0;
    XRAM[6496] = 8'b0;
    XRAM[6497] = 8'b0;
    XRAM[6498] = 8'b0;
    XRAM[6499] = 8'b0;
    XRAM[6500] = 8'b0;
    XRAM[6501] = 8'b0;
    XRAM[6502] = 8'b0;
    XRAM[6503] = 8'b0;
    XRAM[6504] = 8'b0;
    XRAM[6505] = 8'b0;
    XRAM[6506] = 8'b0;
    XRAM[6507] = 8'b0;
    XRAM[6508] = 8'b0;
    XRAM[6509] = 8'b0;
    XRAM[6510] = 8'b0;
    XRAM[6511] = 8'b0;
    XRAM[6512] = 8'b0;
    XRAM[6513] = 8'b0;
    XRAM[6514] = 8'b0;
    XRAM[6515] = 8'b0;
    XRAM[6516] = 8'b0;
    XRAM[6517] = 8'b0;
    XRAM[6518] = 8'b0;
    XRAM[6519] = 8'b0;
    XRAM[6520] = 8'b0;
    XRAM[6521] = 8'b0;
    XRAM[6522] = 8'b0;
    XRAM[6523] = 8'b0;
    XRAM[6524] = 8'b0;
    XRAM[6525] = 8'b0;
    XRAM[6526] = 8'b0;
    XRAM[6527] = 8'b0;
    XRAM[6528] = 8'b0;
    XRAM[6529] = 8'b0;
    XRAM[6530] = 8'b0;
    XRAM[6531] = 8'b0;
    XRAM[6532] = 8'b0;
    XRAM[6533] = 8'b0;
    XRAM[6534] = 8'b0;
    XRAM[6535] = 8'b0;
    XRAM[6536] = 8'b0;
    XRAM[6537] = 8'b0;
    XRAM[6538] = 8'b0;
    XRAM[6539] = 8'b0;
    XRAM[6540] = 8'b0;
    XRAM[6541] = 8'b0;
    XRAM[6542] = 8'b0;
    XRAM[6543] = 8'b0;
    XRAM[6544] = 8'b0;
    XRAM[6545] = 8'b0;
    XRAM[6546] = 8'b0;
    XRAM[6547] = 8'b0;
    XRAM[6548] = 8'b0;
    XRAM[6549] = 8'b0;
    XRAM[6550] = 8'b0;
    XRAM[6551] = 8'b0;
    XRAM[6552] = 8'b0;
    XRAM[6553] = 8'b0;
    XRAM[6554] = 8'b0;
    XRAM[6555] = 8'b0;
    XRAM[6556] = 8'b0;
    XRAM[6557] = 8'b0;
    XRAM[6558] = 8'b0;
    XRAM[6559] = 8'b0;
    XRAM[6560] = 8'b0;
    XRAM[6561] = 8'b0;
    XRAM[6562] = 8'b0;
    XRAM[6563] = 8'b0;
    XRAM[6564] = 8'b0;
    XRAM[6565] = 8'b0;
    XRAM[6566] = 8'b0;
    XRAM[6567] = 8'b0;
    XRAM[6568] = 8'b0;
    XRAM[6569] = 8'b0;
    XRAM[6570] = 8'b0;
    XRAM[6571] = 8'b0;
    XRAM[6572] = 8'b0;
    XRAM[6573] = 8'b0;
    XRAM[6574] = 8'b0;
    XRAM[6575] = 8'b0;
    XRAM[6576] = 8'b0;
    XRAM[6577] = 8'b0;
    XRAM[6578] = 8'b0;
    XRAM[6579] = 8'b0;
    XRAM[6580] = 8'b0;
    XRAM[6581] = 8'b0;
    XRAM[6582] = 8'b0;
    XRAM[6583] = 8'b0;
    XRAM[6584] = 8'b0;
    XRAM[6585] = 8'b0;
    XRAM[6586] = 8'b0;
    XRAM[6587] = 8'b0;
    XRAM[6588] = 8'b0;
    XRAM[6589] = 8'b0;
    XRAM[6590] = 8'b0;
    XRAM[6591] = 8'b0;
    XRAM[6592] = 8'b0;
    XRAM[6593] = 8'b0;
    XRAM[6594] = 8'b0;
    XRAM[6595] = 8'b0;
    XRAM[6596] = 8'b0;
    XRAM[6597] = 8'b0;
    XRAM[6598] = 8'b0;
    XRAM[6599] = 8'b0;
    XRAM[6600] = 8'b0;
    XRAM[6601] = 8'b0;
    XRAM[6602] = 8'b0;
    XRAM[6603] = 8'b0;
    XRAM[6604] = 8'b0;
    XRAM[6605] = 8'b0;
    XRAM[6606] = 8'b0;
    XRAM[6607] = 8'b0;
    XRAM[6608] = 8'b0;
    XRAM[6609] = 8'b0;
    XRAM[6610] = 8'b0;
    XRAM[6611] = 8'b0;
    XRAM[6612] = 8'b0;
    XRAM[6613] = 8'b0;
    XRAM[6614] = 8'b0;
    XRAM[6615] = 8'b0;
    XRAM[6616] = 8'b0;
    XRAM[6617] = 8'b0;
    XRAM[6618] = 8'b0;
    XRAM[6619] = 8'b0;
    XRAM[6620] = 8'b0;
    XRAM[6621] = 8'b0;
    XRAM[6622] = 8'b0;
    XRAM[6623] = 8'b0;
    XRAM[6624] = 8'b0;
    XRAM[6625] = 8'b0;
    XRAM[6626] = 8'b0;
    XRAM[6627] = 8'b0;
    XRAM[6628] = 8'b0;
    XRAM[6629] = 8'b0;
    XRAM[6630] = 8'b0;
    XRAM[6631] = 8'b0;
    XRAM[6632] = 8'b0;
    XRAM[6633] = 8'b0;
    XRAM[6634] = 8'b0;
    XRAM[6635] = 8'b0;
    XRAM[6636] = 8'b0;
    XRAM[6637] = 8'b0;
    XRAM[6638] = 8'b0;
    XRAM[6639] = 8'b0;
    XRAM[6640] = 8'b0;
    XRAM[6641] = 8'b0;
    XRAM[6642] = 8'b0;
    XRAM[6643] = 8'b0;
    XRAM[6644] = 8'b0;
    XRAM[6645] = 8'b0;
    XRAM[6646] = 8'b0;
    XRAM[6647] = 8'b0;
    XRAM[6648] = 8'b0;
    XRAM[6649] = 8'b0;
    XRAM[6650] = 8'b0;
    XRAM[6651] = 8'b0;
    XRAM[6652] = 8'b0;
    XRAM[6653] = 8'b0;
    XRAM[6654] = 8'b0;
    XRAM[6655] = 8'b0;
    XRAM[6656] = 8'b0;
    XRAM[6657] = 8'b0;
    XRAM[6658] = 8'b0;
    XRAM[6659] = 8'b0;
    XRAM[6660] = 8'b0;
    XRAM[6661] = 8'b0;
    XRAM[6662] = 8'b0;
    XRAM[6663] = 8'b0;
    XRAM[6664] = 8'b0;
    XRAM[6665] = 8'b0;
    XRAM[6666] = 8'b0;
    XRAM[6667] = 8'b0;
    XRAM[6668] = 8'b0;
    XRAM[6669] = 8'b0;
    XRAM[6670] = 8'b0;
    XRAM[6671] = 8'b0;
    XRAM[6672] = 8'b0;
    XRAM[6673] = 8'b0;
    XRAM[6674] = 8'b0;
    XRAM[6675] = 8'b0;
    XRAM[6676] = 8'b0;
    XRAM[6677] = 8'b0;
    XRAM[6678] = 8'b0;
    XRAM[6679] = 8'b0;
    XRAM[6680] = 8'b0;
    XRAM[6681] = 8'b0;
    XRAM[6682] = 8'b0;
    XRAM[6683] = 8'b0;
    XRAM[6684] = 8'b0;
    XRAM[6685] = 8'b0;
    XRAM[6686] = 8'b0;
    XRAM[6687] = 8'b0;
    XRAM[6688] = 8'b0;
    XRAM[6689] = 8'b0;
    XRAM[6690] = 8'b0;
    XRAM[6691] = 8'b0;
    XRAM[6692] = 8'b0;
    XRAM[6693] = 8'b0;
    XRAM[6694] = 8'b0;
    XRAM[6695] = 8'b0;
    XRAM[6696] = 8'b0;
    XRAM[6697] = 8'b0;
    XRAM[6698] = 8'b0;
    XRAM[6699] = 8'b0;
    XRAM[6700] = 8'b0;
    XRAM[6701] = 8'b0;
    XRAM[6702] = 8'b0;
    XRAM[6703] = 8'b0;
    XRAM[6704] = 8'b0;
    XRAM[6705] = 8'b0;
    XRAM[6706] = 8'b0;
    XRAM[6707] = 8'b0;
    XRAM[6708] = 8'b0;
    XRAM[6709] = 8'b0;
    XRAM[6710] = 8'b0;
    XRAM[6711] = 8'b0;
    XRAM[6712] = 8'b0;
    XRAM[6713] = 8'b0;
    XRAM[6714] = 8'b0;
    XRAM[6715] = 8'b0;
    XRAM[6716] = 8'b0;
    XRAM[6717] = 8'b0;
    XRAM[6718] = 8'b0;
    XRAM[6719] = 8'b0;
    XRAM[6720] = 8'b0;
    XRAM[6721] = 8'b0;
    XRAM[6722] = 8'b0;
    XRAM[6723] = 8'b0;
    XRAM[6724] = 8'b0;
    XRAM[6725] = 8'b0;
    XRAM[6726] = 8'b0;
    XRAM[6727] = 8'b0;
    XRAM[6728] = 8'b0;
    XRAM[6729] = 8'b0;
    XRAM[6730] = 8'b0;
    XRAM[6731] = 8'b0;
    XRAM[6732] = 8'b0;
    XRAM[6733] = 8'b0;
    XRAM[6734] = 8'b0;
    XRAM[6735] = 8'b0;
    XRAM[6736] = 8'b0;
    XRAM[6737] = 8'b0;
    XRAM[6738] = 8'b0;
    XRAM[6739] = 8'b0;
    XRAM[6740] = 8'b0;
    XRAM[6741] = 8'b0;
    XRAM[6742] = 8'b0;
    XRAM[6743] = 8'b0;
    XRAM[6744] = 8'b0;
    XRAM[6745] = 8'b0;
    XRAM[6746] = 8'b0;
    XRAM[6747] = 8'b0;
    XRAM[6748] = 8'b0;
    XRAM[6749] = 8'b0;
    XRAM[6750] = 8'b0;
    XRAM[6751] = 8'b0;
    XRAM[6752] = 8'b0;
    XRAM[6753] = 8'b0;
    XRAM[6754] = 8'b0;
    XRAM[6755] = 8'b0;
    XRAM[6756] = 8'b0;
    XRAM[6757] = 8'b0;
    XRAM[6758] = 8'b0;
    XRAM[6759] = 8'b0;
    XRAM[6760] = 8'b0;
    XRAM[6761] = 8'b0;
    XRAM[6762] = 8'b0;
    XRAM[6763] = 8'b0;
    XRAM[6764] = 8'b0;
    XRAM[6765] = 8'b0;
    XRAM[6766] = 8'b0;
    XRAM[6767] = 8'b0;
    XRAM[6768] = 8'b0;
    XRAM[6769] = 8'b0;
    XRAM[6770] = 8'b0;
    XRAM[6771] = 8'b0;
    XRAM[6772] = 8'b0;
    XRAM[6773] = 8'b0;
    XRAM[6774] = 8'b0;
    XRAM[6775] = 8'b0;
    XRAM[6776] = 8'b0;
    XRAM[6777] = 8'b0;
    XRAM[6778] = 8'b0;
    XRAM[6779] = 8'b0;
    XRAM[6780] = 8'b0;
    XRAM[6781] = 8'b0;
    XRAM[6782] = 8'b0;
    XRAM[6783] = 8'b0;
    XRAM[6784] = 8'b0;
    XRAM[6785] = 8'b0;
    XRAM[6786] = 8'b0;
    XRAM[6787] = 8'b0;
    XRAM[6788] = 8'b0;
    XRAM[6789] = 8'b0;
    XRAM[6790] = 8'b0;
    XRAM[6791] = 8'b0;
    XRAM[6792] = 8'b0;
    XRAM[6793] = 8'b0;
    XRAM[6794] = 8'b0;
    XRAM[6795] = 8'b0;
    XRAM[6796] = 8'b0;
    XRAM[6797] = 8'b0;
    XRAM[6798] = 8'b0;
    XRAM[6799] = 8'b0;
    XRAM[6800] = 8'b0;
    XRAM[6801] = 8'b0;
    XRAM[6802] = 8'b0;
    XRAM[6803] = 8'b0;
    XRAM[6804] = 8'b0;
    XRAM[6805] = 8'b0;
    XRAM[6806] = 8'b0;
    XRAM[6807] = 8'b0;
    XRAM[6808] = 8'b0;
    XRAM[6809] = 8'b0;
    XRAM[6810] = 8'b0;
    XRAM[6811] = 8'b0;
    XRAM[6812] = 8'b0;
    XRAM[6813] = 8'b0;
    XRAM[6814] = 8'b0;
    XRAM[6815] = 8'b0;
    XRAM[6816] = 8'b0;
    XRAM[6817] = 8'b0;
    XRAM[6818] = 8'b0;
    XRAM[6819] = 8'b0;
    XRAM[6820] = 8'b0;
    XRAM[6821] = 8'b0;
    XRAM[6822] = 8'b0;
    XRAM[6823] = 8'b0;
    XRAM[6824] = 8'b0;
    XRAM[6825] = 8'b0;
    XRAM[6826] = 8'b0;
    XRAM[6827] = 8'b0;
    XRAM[6828] = 8'b0;
    XRAM[6829] = 8'b0;
    XRAM[6830] = 8'b0;
    XRAM[6831] = 8'b0;
    XRAM[6832] = 8'b0;
    XRAM[6833] = 8'b0;
    XRAM[6834] = 8'b0;
    XRAM[6835] = 8'b0;
    XRAM[6836] = 8'b0;
    XRAM[6837] = 8'b0;
    XRAM[6838] = 8'b0;
    XRAM[6839] = 8'b0;
    XRAM[6840] = 8'b0;
    XRAM[6841] = 8'b0;
    XRAM[6842] = 8'b0;
    XRAM[6843] = 8'b0;
    XRAM[6844] = 8'b0;
    XRAM[6845] = 8'b0;
    XRAM[6846] = 8'b0;
    XRAM[6847] = 8'b0;
    XRAM[6848] = 8'b0;
    XRAM[6849] = 8'b0;
    XRAM[6850] = 8'b0;
    XRAM[6851] = 8'b0;
    XRAM[6852] = 8'b0;
    XRAM[6853] = 8'b0;
    XRAM[6854] = 8'b0;
    XRAM[6855] = 8'b0;
    XRAM[6856] = 8'b0;
    XRAM[6857] = 8'b0;
    XRAM[6858] = 8'b0;
    XRAM[6859] = 8'b0;
    XRAM[6860] = 8'b0;
    XRAM[6861] = 8'b0;
    XRAM[6862] = 8'b0;
    XRAM[6863] = 8'b0;
    XRAM[6864] = 8'b0;
    XRAM[6865] = 8'b0;
    XRAM[6866] = 8'b0;
    XRAM[6867] = 8'b0;
    XRAM[6868] = 8'b0;
    XRAM[6869] = 8'b0;
    XRAM[6870] = 8'b0;
    XRAM[6871] = 8'b0;
    XRAM[6872] = 8'b0;
    XRAM[6873] = 8'b0;
    XRAM[6874] = 8'b0;
    XRAM[6875] = 8'b0;
    XRAM[6876] = 8'b0;
    XRAM[6877] = 8'b0;
    XRAM[6878] = 8'b0;
    XRAM[6879] = 8'b0;
    XRAM[6880] = 8'b0;
    XRAM[6881] = 8'b0;
    XRAM[6882] = 8'b0;
    XRAM[6883] = 8'b0;
    XRAM[6884] = 8'b0;
    XRAM[6885] = 8'b0;
    XRAM[6886] = 8'b0;
    XRAM[6887] = 8'b0;
    XRAM[6888] = 8'b0;
    XRAM[6889] = 8'b0;
    XRAM[6890] = 8'b0;
    XRAM[6891] = 8'b0;
    XRAM[6892] = 8'b0;
    XRAM[6893] = 8'b0;
    XRAM[6894] = 8'b0;
    XRAM[6895] = 8'b0;
    XRAM[6896] = 8'b0;
    XRAM[6897] = 8'b0;
    XRAM[6898] = 8'b0;
    XRAM[6899] = 8'b0;
    XRAM[6900] = 8'b0;
    XRAM[6901] = 8'b0;
    XRAM[6902] = 8'b0;
    XRAM[6903] = 8'b0;
    XRAM[6904] = 8'b0;
    XRAM[6905] = 8'b0;
    XRAM[6906] = 8'b0;
    XRAM[6907] = 8'b0;
    XRAM[6908] = 8'b0;
    XRAM[6909] = 8'b0;
    XRAM[6910] = 8'b0;
    XRAM[6911] = 8'b0;
    XRAM[6912] = 8'b0;
    XRAM[6913] = 8'b0;
    XRAM[6914] = 8'b0;
    XRAM[6915] = 8'b0;
    XRAM[6916] = 8'b0;
    XRAM[6917] = 8'b0;
    XRAM[6918] = 8'b0;
    XRAM[6919] = 8'b0;
    XRAM[6920] = 8'b0;
    XRAM[6921] = 8'b0;
    XRAM[6922] = 8'b0;
    XRAM[6923] = 8'b0;
    XRAM[6924] = 8'b0;
    XRAM[6925] = 8'b0;
    XRAM[6926] = 8'b0;
    XRAM[6927] = 8'b0;
    XRAM[6928] = 8'b0;
    XRAM[6929] = 8'b0;
    XRAM[6930] = 8'b0;
    XRAM[6931] = 8'b0;
    XRAM[6932] = 8'b0;
    XRAM[6933] = 8'b0;
    XRAM[6934] = 8'b0;
    XRAM[6935] = 8'b0;
    XRAM[6936] = 8'b0;
    XRAM[6937] = 8'b0;
    XRAM[6938] = 8'b0;
    XRAM[6939] = 8'b0;
    XRAM[6940] = 8'b0;
    XRAM[6941] = 8'b0;
    XRAM[6942] = 8'b0;
    XRAM[6943] = 8'b0;
    XRAM[6944] = 8'b0;
    XRAM[6945] = 8'b0;
    XRAM[6946] = 8'b0;
    XRAM[6947] = 8'b0;
    XRAM[6948] = 8'b0;
    XRAM[6949] = 8'b0;
    XRAM[6950] = 8'b0;
    XRAM[6951] = 8'b0;
    XRAM[6952] = 8'b0;
    XRAM[6953] = 8'b0;
    XRAM[6954] = 8'b0;
    XRAM[6955] = 8'b0;
    XRAM[6956] = 8'b0;
    XRAM[6957] = 8'b0;
    XRAM[6958] = 8'b0;
    XRAM[6959] = 8'b0;
    XRAM[6960] = 8'b0;
    XRAM[6961] = 8'b0;
    XRAM[6962] = 8'b0;
    XRAM[6963] = 8'b0;
    XRAM[6964] = 8'b0;
    XRAM[6965] = 8'b0;
    XRAM[6966] = 8'b0;
    XRAM[6967] = 8'b0;
    XRAM[6968] = 8'b0;
    XRAM[6969] = 8'b0;
    XRAM[6970] = 8'b0;
    XRAM[6971] = 8'b0;
    XRAM[6972] = 8'b0;
    XRAM[6973] = 8'b0;
    XRAM[6974] = 8'b0;
    XRAM[6975] = 8'b0;
    XRAM[6976] = 8'b0;
    XRAM[6977] = 8'b0;
    XRAM[6978] = 8'b0;
    XRAM[6979] = 8'b0;
    XRAM[6980] = 8'b0;
    XRAM[6981] = 8'b0;
    XRAM[6982] = 8'b0;
    XRAM[6983] = 8'b0;
    XRAM[6984] = 8'b0;
    XRAM[6985] = 8'b0;
    XRAM[6986] = 8'b0;
    XRAM[6987] = 8'b0;
    XRAM[6988] = 8'b0;
    XRAM[6989] = 8'b0;
    XRAM[6990] = 8'b0;
    XRAM[6991] = 8'b0;
    XRAM[6992] = 8'b0;
    XRAM[6993] = 8'b0;
    XRAM[6994] = 8'b0;
    XRAM[6995] = 8'b0;
    XRAM[6996] = 8'b0;
    XRAM[6997] = 8'b0;
    XRAM[6998] = 8'b0;
    XRAM[6999] = 8'b0;
    XRAM[7000] = 8'b0;
    XRAM[7001] = 8'b0;
    XRAM[7002] = 8'b0;
    XRAM[7003] = 8'b0;
    XRAM[7004] = 8'b0;
    XRAM[7005] = 8'b0;
    XRAM[7006] = 8'b0;
    XRAM[7007] = 8'b0;
    XRAM[7008] = 8'b0;
    XRAM[7009] = 8'b0;
    XRAM[7010] = 8'b0;
    XRAM[7011] = 8'b0;
    XRAM[7012] = 8'b0;
    XRAM[7013] = 8'b0;
    XRAM[7014] = 8'b0;
    XRAM[7015] = 8'b0;
    XRAM[7016] = 8'b0;
    XRAM[7017] = 8'b0;
    XRAM[7018] = 8'b0;
    XRAM[7019] = 8'b0;
    XRAM[7020] = 8'b0;
    XRAM[7021] = 8'b0;
    XRAM[7022] = 8'b0;
    XRAM[7023] = 8'b0;
    XRAM[7024] = 8'b0;
    XRAM[7025] = 8'b0;
    XRAM[7026] = 8'b0;
    XRAM[7027] = 8'b0;
    XRAM[7028] = 8'b0;
    XRAM[7029] = 8'b0;
    XRAM[7030] = 8'b0;
    XRAM[7031] = 8'b0;
    XRAM[7032] = 8'b0;
    XRAM[7033] = 8'b0;
    XRAM[7034] = 8'b0;
    XRAM[7035] = 8'b0;
    XRAM[7036] = 8'b0;
    XRAM[7037] = 8'b0;
    XRAM[7038] = 8'b0;
    XRAM[7039] = 8'b0;
    XRAM[7040] = 8'b0;
    XRAM[7041] = 8'b0;
    XRAM[7042] = 8'b0;
    XRAM[7043] = 8'b0;
    XRAM[7044] = 8'b0;
    XRAM[7045] = 8'b0;
    XRAM[7046] = 8'b0;
    XRAM[7047] = 8'b0;
    XRAM[7048] = 8'b0;
    XRAM[7049] = 8'b0;
    XRAM[7050] = 8'b0;
    XRAM[7051] = 8'b0;
    XRAM[7052] = 8'b0;
    XRAM[7053] = 8'b0;
    XRAM[7054] = 8'b0;
    XRAM[7055] = 8'b0;
    XRAM[7056] = 8'b0;
    XRAM[7057] = 8'b0;
    XRAM[7058] = 8'b0;
    XRAM[7059] = 8'b0;
    XRAM[7060] = 8'b0;
    XRAM[7061] = 8'b0;
    XRAM[7062] = 8'b0;
    XRAM[7063] = 8'b0;
    XRAM[7064] = 8'b0;
    XRAM[7065] = 8'b0;
    XRAM[7066] = 8'b0;
    XRAM[7067] = 8'b0;
    XRAM[7068] = 8'b0;
    XRAM[7069] = 8'b0;
    XRAM[7070] = 8'b0;
    XRAM[7071] = 8'b0;
    XRAM[7072] = 8'b0;
    XRAM[7073] = 8'b0;
    XRAM[7074] = 8'b0;
    XRAM[7075] = 8'b0;
    XRAM[7076] = 8'b0;
    XRAM[7077] = 8'b0;
    XRAM[7078] = 8'b0;
    XRAM[7079] = 8'b0;
    XRAM[7080] = 8'b0;
    XRAM[7081] = 8'b0;
    XRAM[7082] = 8'b0;
    XRAM[7083] = 8'b0;
    XRAM[7084] = 8'b0;
    XRAM[7085] = 8'b0;
    XRAM[7086] = 8'b0;
    XRAM[7087] = 8'b0;
    XRAM[7088] = 8'b0;
    XRAM[7089] = 8'b0;
    XRAM[7090] = 8'b0;
    XRAM[7091] = 8'b0;
    XRAM[7092] = 8'b0;
    XRAM[7093] = 8'b0;
    XRAM[7094] = 8'b0;
    XRAM[7095] = 8'b0;
    XRAM[7096] = 8'b0;
    XRAM[7097] = 8'b0;
    XRAM[7098] = 8'b0;
    XRAM[7099] = 8'b0;
    XRAM[7100] = 8'b0;
    XRAM[7101] = 8'b0;
    XRAM[7102] = 8'b0;
    XRAM[7103] = 8'b0;
    XRAM[7104] = 8'b0;
    XRAM[7105] = 8'b0;
    XRAM[7106] = 8'b0;
    XRAM[7107] = 8'b0;
    XRAM[7108] = 8'b0;
    XRAM[7109] = 8'b0;
    XRAM[7110] = 8'b0;
    XRAM[7111] = 8'b0;
    XRAM[7112] = 8'b0;
    XRAM[7113] = 8'b0;
    XRAM[7114] = 8'b0;
    XRAM[7115] = 8'b0;
    XRAM[7116] = 8'b0;
    XRAM[7117] = 8'b0;
    XRAM[7118] = 8'b0;
    XRAM[7119] = 8'b0;
    XRAM[7120] = 8'b0;
    XRAM[7121] = 8'b0;
    XRAM[7122] = 8'b0;
    XRAM[7123] = 8'b0;
    XRAM[7124] = 8'b0;
    XRAM[7125] = 8'b0;
    XRAM[7126] = 8'b0;
    XRAM[7127] = 8'b0;
    XRAM[7128] = 8'b0;
    XRAM[7129] = 8'b0;
    XRAM[7130] = 8'b0;
    XRAM[7131] = 8'b0;
    XRAM[7132] = 8'b0;
    XRAM[7133] = 8'b0;
    XRAM[7134] = 8'b0;
    XRAM[7135] = 8'b0;
    XRAM[7136] = 8'b0;
    XRAM[7137] = 8'b0;
    XRAM[7138] = 8'b0;
    XRAM[7139] = 8'b0;
    XRAM[7140] = 8'b0;
    XRAM[7141] = 8'b0;
    XRAM[7142] = 8'b0;
    XRAM[7143] = 8'b0;
    XRAM[7144] = 8'b0;
    XRAM[7145] = 8'b0;
    XRAM[7146] = 8'b0;
    XRAM[7147] = 8'b0;
    XRAM[7148] = 8'b0;
    XRAM[7149] = 8'b0;
    XRAM[7150] = 8'b0;
    XRAM[7151] = 8'b0;
    XRAM[7152] = 8'b0;
    XRAM[7153] = 8'b0;
    XRAM[7154] = 8'b0;
    XRAM[7155] = 8'b0;
    XRAM[7156] = 8'b0;
    XRAM[7157] = 8'b0;
    XRAM[7158] = 8'b0;
    XRAM[7159] = 8'b0;
    XRAM[7160] = 8'b0;
    XRAM[7161] = 8'b0;
    XRAM[7162] = 8'b0;
    XRAM[7163] = 8'b0;
    XRAM[7164] = 8'b0;
    XRAM[7165] = 8'b0;
    XRAM[7166] = 8'b0;
    XRAM[7167] = 8'b0;
    XRAM[7168] = 8'b0;
    XRAM[7169] = 8'b0;
    XRAM[7170] = 8'b0;
    XRAM[7171] = 8'b0;
    XRAM[7172] = 8'b0;
    XRAM[7173] = 8'b0;
    XRAM[7174] = 8'b0;
    XRAM[7175] = 8'b0;
    XRAM[7176] = 8'b0;
    XRAM[7177] = 8'b0;
    XRAM[7178] = 8'b0;
    XRAM[7179] = 8'b0;
    XRAM[7180] = 8'b0;
    XRAM[7181] = 8'b0;
    XRAM[7182] = 8'b0;
    XRAM[7183] = 8'b0;
    XRAM[7184] = 8'b0;
    XRAM[7185] = 8'b0;
    XRAM[7186] = 8'b0;
    XRAM[7187] = 8'b0;
    XRAM[7188] = 8'b0;
    XRAM[7189] = 8'b0;
    XRAM[7190] = 8'b0;
    XRAM[7191] = 8'b0;
    XRAM[7192] = 8'b0;
    XRAM[7193] = 8'b0;
    XRAM[7194] = 8'b0;
    XRAM[7195] = 8'b0;
    XRAM[7196] = 8'b0;
    XRAM[7197] = 8'b0;
    XRAM[7198] = 8'b0;
    XRAM[7199] = 8'b0;
    XRAM[7200] = 8'b0;
    XRAM[7201] = 8'b0;
    XRAM[7202] = 8'b0;
    XRAM[7203] = 8'b0;
    XRAM[7204] = 8'b0;
    XRAM[7205] = 8'b0;
    XRAM[7206] = 8'b0;
    XRAM[7207] = 8'b0;
    XRAM[7208] = 8'b0;
    XRAM[7209] = 8'b0;
    XRAM[7210] = 8'b0;
    XRAM[7211] = 8'b0;
    XRAM[7212] = 8'b0;
    XRAM[7213] = 8'b0;
    XRAM[7214] = 8'b0;
    XRAM[7215] = 8'b0;
    XRAM[7216] = 8'b0;
    XRAM[7217] = 8'b0;
    XRAM[7218] = 8'b0;
    XRAM[7219] = 8'b0;
    XRAM[7220] = 8'b0;
    XRAM[7221] = 8'b0;
    XRAM[7222] = 8'b0;
    XRAM[7223] = 8'b0;
    XRAM[7224] = 8'b0;
    XRAM[7225] = 8'b0;
    XRAM[7226] = 8'b0;
    XRAM[7227] = 8'b0;
    XRAM[7228] = 8'b0;
    XRAM[7229] = 8'b0;
    XRAM[7230] = 8'b0;
    XRAM[7231] = 8'b0;
    XRAM[7232] = 8'b0;
    XRAM[7233] = 8'b0;
    XRAM[7234] = 8'b0;
    XRAM[7235] = 8'b0;
    XRAM[7236] = 8'b0;
    XRAM[7237] = 8'b0;
    XRAM[7238] = 8'b0;
    XRAM[7239] = 8'b0;
    XRAM[7240] = 8'b0;
    XRAM[7241] = 8'b0;
    XRAM[7242] = 8'b0;
    XRAM[7243] = 8'b0;
    XRAM[7244] = 8'b0;
    XRAM[7245] = 8'b0;
    XRAM[7246] = 8'b0;
    XRAM[7247] = 8'b0;
    XRAM[7248] = 8'b0;
    XRAM[7249] = 8'b0;
    XRAM[7250] = 8'b0;
    XRAM[7251] = 8'b0;
    XRAM[7252] = 8'b0;
    XRAM[7253] = 8'b0;
    XRAM[7254] = 8'b0;
    XRAM[7255] = 8'b0;
    XRAM[7256] = 8'b0;
    XRAM[7257] = 8'b0;
    XRAM[7258] = 8'b0;
    XRAM[7259] = 8'b0;
    XRAM[7260] = 8'b0;
    XRAM[7261] = 8'b0;
    XRAM[7262] = 8'b0;
    XRAM[7263] = 8'b0;
    XRAM[7264] = 8'b0;
    XRAM[7265] = 8'b0;
    XRAM[7266] = 8'b0;
    XRAM[7267] = 8'b0;
    XRAM[7268] = 8'b0;
    XRAM[7269] = 8'b0;
    XRAM[7270] = 8'b0;
    XRAM[7271] = 8'b0;
    XRAM[7272] = 8'b0;
    XRAM[7273] = 8'b0;
    XRAM[7274] = 8'b0;
    XRAM[7275] = 8'b0;
    XRAM[7276] = 8'b0;
    XRAM[7277] = 8'b0;
    XRAM[7278] = 8'b0;
    XRAM[7279] = 8'b0;
    XRAM[7280] = 8'b0;
    XRAM[7281] = 8'b0;
    XRAM[7282] = 8'b0;
    XRAM[7283] = 8'b0;
    XRAM[7284] = 8'b0;
    XRAM[7285] = 8'b0;
    XRAM[7286] = 8'b0;
    XRAM[7287] = 8'b0;
    XRAM[7288] = 8'b0;
    XRAM[7289] = 8'b0;
    XRAM[7290] = 8'b0;
    XRAM[7291] = 8'b0;
    XRAM[7292] = 8'b0;
    XRAM[7293] = 8'b0;
    XRAM[7294] = 8'b0;
    XRAM[7295] = 8'b0;
    XRAM[7296] = 8'b0;
    XRAM[7297] = 8'b0;
    XRAM[7298] = 8'b0;
    XRAM[7299] = 8'b0;
    XRAM[7300] = 8'b0;
    XRAM[7301] = 8'b0;
    XRAM[7302] = 8'b0;
    XRAM[7303] = 8'b0;
    XRAM[7304] = 8'b0;
    XRAM[7305] = 8'b0;
    XRAM[7306] = 8'b0;
    XRAM[7307] = 8'b0;
    XRAM[7308] = 8'b0;
    XRAM[7309] = 8'b0;
    XRAM[7310] = 8'b0;
    XRAM[7311] = 8'b0;
    XRAM[7312] = 8'b0;
    XRAM[7313] = 8'b0;
    XRAM[7314] = 8'b0;
    XRAM[7315] = 8'b0;
    XRAM[7316] = 8'b0;
    XRAM[7317] = 8'b0;
    XRAM[7318] = 8'b0;
    XRAM[7319] = 8'b0;
    XRAM[7320] = 8'b0;
    XRAM[7321] = 8'b0;
    XRAM[7322] = 8'b0;
    XRAM[7323] = 8'b0;
    XRAM[7324] = 8'b0;
    XRAM[7325] = 8'b0;
    XRAM[7326] = 8'b0;
    XRAM[7327] = 8'b0;
    XRAM[7328] = 8'b0;
    XRAM[7329] = 8'b0;
    XRAM[7330] = 8'b0;
    XRAM[7331] = 8'b0;
    XRAM[7332] = 8'b0;
    XRAM[7333] = 8'b0;
    XRAM[7334] = 8'b0;
    XRAM[7335] = 8'b0;
    XRAM[7336] = 8'b0;
    XRAM[7337] = 8'b0;
    XRAM[7338] = 8'b0;
    XRAM[7339] = 8'b0;
    XRAM[7340] = 8'b0;
    XRAM[7341] = 8'b0;
    XRAM[7342] = 8'b0;
    XRAM[7343] = 8'b0;
    XRAM[7344] = 8'b0;
    XRAM[7345] = 8'b0;
    XRAM[7346] = 8'b0;
    XRAM[7347] = 8'b0;
    XRAM[7348] = 8'b0;
    XRAM[7349] = 8'b0;
    XRAM[7350] = 8'b0;
    XRAM[7351] = 8'b0;
    XRAM[7352] = 8'b0;
    XRAM[7353] = 8'b0;
    XRAM[7354] = 8'b0;
    XRAM[7355] = 8'b0;
    XRAM[7356] = 8'b0;
    XRAM[7357] = 8'b0;
    XRAM[7358] = 8'b0;
    XRAM[7359] = 8'b0;
    XRAM[7360] = 8'b0;
    XRAM[7361] = 8'b0;
    XRAM[7362] = 8'b0;
    XRAM[7363] = 8'b0;
    XRAM[7364] = 8'b0;
    XRAM[7365] = 8'b0;
    XRAM[7366] = 8'b0;
    XRAM[7367] = 8'b0;
    XRAM[7368] = 8'b0;
    XRAM[7369] = 8'b0;
    XRAM[7370] = 8'b0;
    XRAM[7371] = 8'b0;
    XRAM[7372] = 8'b0;
    XRAM[7373] = 8'b0;
    XRAM[7374] = 8'b0;
    XRAM[7375] = 8'b0;
    XRAM[7376] = 8'b0;
    XRAM[7377] = 8'b0;
    XRAM[7378] = 8'b0;
    XRAM[7379] = 8'b0;
    XRAM[7380] = 8'b0;
    XRAM[7381] = 8'b0;
    XRAM[7382] = 8'b0;
    XRAM[7383] = 8'b0;
    XRAM[7384] = 8'b0;
    XRAM[7385] = 8'b0;
    XRAM[7386] = 8'b0;
    XRAM[7387] = 8'b0;
    XRAM[7388] = 8'b0;
    XRAM[7389] = 8'b0;
    XRAM[7390] = 8'b0;
    XRAM[7391] = 8'b0;
    XRAM[7392] = 8'b0;
    XRAM[7393] = 8'b0;
    XRAM[7394] = 8'b0;
    XRAM[7395] = 8'b0;
    XRAM[7396] = 8'b0;
    XRAM[7397] = 8'b0;
    XRAM[7398] = 8'b0;
    XRAM[7399] = 8'b0;
    XRAM[7400] = 8'b0;
    XRAM[7401] = 8'b0;
    XRAM[7402] = 8'b0;
    XRAM[7403] = 8'b0;
    XRAM[7404] = 8'b0;
    XRAM[7405] = 8'b0;
    XRAM[7406] = 8'b0;
    XRAM[7407] = 8'b0;
    XRAM[7408] = 8'b0;
    XRAM[7409] = 8'b0;
    XRAM[7410] = 8'b0;
    XRAM[7411] = 8'b0;
    XRAM[7412] = 8'b0;
    XRAM[7413] = 8'b0;
    XRAM[7414] = 8'b0;
    XRAM[7415] = 8'b0;
    XRAM[7416] = 8'b0;
    XRAM[7417] = 8'b0;
    XRAM[7418] = 8'b0;
    XRAM[7419] = 8'b0;
    XRAM[7420] = 8'b0;
    XRAM[7421] = 8'b0;
    XRAM[7422] = 8'b0;
    XRAM[7423] = 8'b0;
    XRAM[7424] = 8'b0;
    XRAM[7425] = 8'b0;
    XRAM[7426] = 8'b0;
    XRAM[7427] = 8'b0;
    XRAM[7428] = 8'b0;
    XRAM[7429] = 8'b0;
    XRAM[7430] = 8'b0;
    XRAM[7431] = 8'b0;
    XRAM[7432] = 8'b0;
    XRAM[7433] = 8'b0;
    XRAM[7434] = 8'b0;
    XRAM[7435] = 8'b0;
    XRAM[7436] = 8'b0;
    XRAM[7437] = 8'b0;
    XRAM[7438] = 8'b0;
    XRAM[7439] = 8'b0;
    XRAM[7440] = 8'b0;
    XRAM[7441] = 8'b0;
    XRAM[7442] = 8'b0;
    XRAM[7443] = 8'b0;
    XRAM[7444] = 8'b0;
    XRAM[7445] = 8'b0;
    XRAM[7446] = 8'b0;
    XRAM[7447] = 8'b0;
    XRAM[7448] = 8'b0;
    XRAM[7449] = 8'b0;
    XRAM[7450] = 8'b0;
    XRAM[7451] = 8'b0;
    XRAM[7452] = 8'b0;
    XRAM[7453] = 8'b0;
    XRAM[7454] = 8'b0;
    XRAM[7455] = 8'b0;
    XRAM[7456] = 8'b0;
    XRAM[7457] = 8'b0;
    XRAM[7458] = 8'b0;
    XRAM[7459] = 8'b0;
    XRAM[7460] = 8'b0;
    XRAM[7461] = 8'b0;
    XRAM[7462] = 8'b0;
    XRAM[7463] = 8'b0;
    XRAM[7464] = 8'b0;
    XRAM[7465] = 8'b0;
    XRAM[7466] = 8'b0;
    XRAM[7467] = 8'b0;
    XRAM[7468] = 8'b0;
    XRAM[7469] = 8'b0;
    XRAM[7470] = 8'b0;
    XRAM[7471] = 8'b0;
    XRAM[7472] = 8'b0;
    XRAM[7473] = 8'b0;
    XRAM[7474] = 8'b0;
    XRAM[7475] = 8'b0;
    XRAM[7476] = 8'b0;
    XRAM[7477] = 8'b0;
    XRAM[7478] = 8'b0;
    XRAM[7479] = 8'b0;
    XRAM[7480] = 8'b0;
    XRAM[7481] = 8'b0;
    XRAM[7482] = 8'b0;
    XRAM[7483] = 8'b0;
    XRAM[7484] = 8'b0;
    XRAM[7485] = 8'b0;
    XRAM[7486] = 8'b0;
    XRAM[7487] = 8'b0;
    XRAM[7488] = 8'b0;
    XRAM[7489] = 8'b0;
    XRAM[7490] = 8'b0;
    XRAM[7491] = 8'b0;
    XRAM[7492] = 8'b0;
    XRAM[7493] = 8'b0;
    XRAM[7494] = 8'b0;
    XRAM[7495] = 8'b0;
    XRAM[7496] = 8'b0;
    XRAM[7497] = 8'b0;
    XRAM[7498] = 8'b0;
    XRAM[7499] = 8'b0;
    XRAM[7500] = 8'b0;
    XRAM[7501] = 8'b0;
    XRAM[7502] = 8'b0;
    XRAM[7503] = 8'b0;
    XRAM[7504] = 8'b0;
    XRAM[7505] = 8'b0;
    XRAM[7506] = 8'b0;
    XRAM[7507] = 8'b0;
    XRAM[7508] = 8'b0;
    XRAM[7509] = 8'b0;
    XRAM[7510] = 8'b0;
    XRAM[7511] = 8'b0;
    XRAM[7512] = 8'b0;
    XRAM[7513] = 8'b0;
    XRAM[7514] = 8'b0;
    XRAM[7515] = 8'b0;
    XRAM[7516] = 8'b0;
    XRAM[7517] = 8'b0;
    XRAM[7518] = 8'b0;
    XRAM[7519] = 8'b0;
    XRAM[7520] = 8'b0;
    XRAM[7521] = 8'b0;
    XRAM[7522] = 8'b0;
    XRAM[7523] = 8'b0;
    XRAM[7524] = 8'b0;
    XRAM[7525] = 8'b0;
    XRAM[7526] = 8'b0;
    XRAM[7527] = 8'b0;
    XRAM[7528] = 8'b0;
    XRAM[7529] = 8'b0;
    XRAM[7530] = 8'b0;
    XRAM[7531] = 8'b0;
    XRAM[7532] = 8'b0;
    XRAM[7533] = 8'b0;
    XRAM[7534] = 8'b0;
    XRAM[7535] = 8'b0;
    XRAM[7536] = 8'b0;
    XRAM[7537] = 8'b0;
    XRAM[7538] = 8'b0;
    XRAM[7539] = 8'b0;
    XRAM[7540] = 8'b0;
    XRAM[7541] = 8'b0;
    XRAM[7542] = 8'b0;
    XRAM[7543] = 8'b0;
    XRAM[7544] = 8'b0;
    XRAM[7545] = 8'b0;
    XRAM[7546] = 8'b0;
    XRAM[7547] = 8'b0;
    XRAM[7548] = 8'b0;
    XRAM[7549] = 8'b0;
    XRAM[7550] = 8'b0;
    XRAM[7551] = 8'b0;
    XRAM[7552] = 8'b0;
    XRAM[7553] = 8'b0;
    XRAM[7554] = 8'b0;
    XRAM[7555] = 8'b0;
    XRAM[7556] = 8'b0;
    XRAM[7557] = 8'b0;
    XRAM[7558] = 8'b0;
    XRAM[7559] = 8'b0;
    XRAM[7560] = 8'b0;
    XRAM[7561] = 8'b0;
    XRAM[7562] = 8'b0;
    XRAM[7563] = 8'b0;
    XRAM[7564] = 8'b0;
    XRAM[7565] = 8'b0;
    XRAM[7566] = 8'b0;
    XRAM[7567] = 8'b0;
    XRAM[7568] = 8'b0;
    XRAM[7569] = 8'b0;
    XRAM[7570] = 8'b0;
    XRAM[7571] = 8'b0;
    XRAM[7572] = 8'b0;
    XRAM[7573] = 8'b0;
    XRAM[7574] = 8'b0;
    XRAM[7575] = 8'b0;
    XRAM[7576] = 8'b0;
    XRAM[7577] = 8'b0;
    XRAM[7578] = 8'b0;
    XRAM[7579] = 8'b0;
    XRAM[7580] = 8'b0;
    XRAM[7581] = 8'b0;
    XRAM[7582] = 8'b0;
    XRAM[7583] = 8'b0;
    XRAM[7584] = 8'b0;
    XRAM[7585] = 8'b0;
    XRAM[7586] = 8'b0;
    XRAM[7587] = 8'b0;
    XRAM[7588] = 8'b0;
    XRAM[7589] = 8'b0;
    XRAM[7590] = 8'b0;
    XRAM[7591] = 8'b0;
    XRAM[7592] = 8'b0;
    XRAM[7593] = 8'b0;
    XRAM[7594] = 8'b0;
    XRAM[7595] = 8'b0;
    XRAM[7596] = 8'b0;
    XRAM[7597] = 8'b0;
    XRAM[7598] = 8'b0;
    XRAM[7599] = 8'b0;
    XRAM[7600] = 8'b0;
    XRAM[7601] = 8'b0;
    XRAM[7602] = 8'b0;
    XRAM[7603] = 8'b0;
    XRAM[7604] = 8'b0;
    XRAM[7605] = 8'b0;
    XRAM[7606] = 8'b0;
    XRAM[7607] = 8'b0;
    XRAM[7608] = 8'b0;
    XRAM[7609] = 8'b0;
    XRAM[7610] = 8'b0;
    XRAM[7611] = 8'b0;
    XRAM[7612] = 8'b0;
    XRAM[7613] = 8'b0;
    XRAM[7614] = 8'b0;
    XRAM[7615] = 8'b0;
    XRAM[7616] = 8'b0;
    XRAM[7617] = 8'b0;
    XRAM[7618] = 8'b0;
    XRAM[7619] = 8'b0;
    XRAM[7620] = 8'b0;
    XRAM[7621] = 8'b0;
    XRAM[7622] = 8'b0;
    XRAM[7623] = 8'b0;
    XRAM[7624] = 8'b0;
    XRAM[7625] = 8'b0;
    XRAM[7626] = 8'b0;
    XRAM[7627] = 8'b0;
    XRAM[7628] = 8'b0;
    XRAM[7629] = 8'b0;
    XRAM[7630] = 8'b0;
    XRAM[7631] = 8'b0;
    XRAM[7632] = 8'b0;
    XRAM[7633] = 8'b0;
    XRAM[7634] = 8'b0;
    XRAM[7635] = 8'b0;
    XRAM[7636] = 8'b0;
    XRAM[7637] = 8'b0;
    XRAM[7638] = 8'b0;
    XRAM[7639] = 8'b0;
    XRAM[7640] = 8'b0;
    XRAM[7641] = 8'b0;
    XRAM[7642] = 8'b0;
    XRAM[7643] = 8'b0;
    XRAM[7644] = 8'b0;
    XRAM[7645] = 8'b0;
    XRAM[7646] = 8'b0;
    XRAM[7647] = 8'b0;
    XRAM[7648] = 8'b0;
    XRAM[7649] = 8'b0;
    XRAM[7650] = 8'b0;
    XRAM[7651] = 8'b0;
    XRAM[7652] = 8'b0;
    XRAM[7653] = 8'b0;
    XRAM[7654] = 8'b0;
    XRAM[7655] = 8'b0;
    XRAM[7656] = 8'b0;
    XRAM[7657] = 8'b0;
    XRAM[7658] = 8'b0;
    XRAM[7659] = 8'b0;
    XRAM[7660] = 8'b0;
    XRAM[7661] = 8'b0;
    XRAM[7662] = 8'b0;
    XRAM[7663] = 8'b0;
    XRAM[7664] = 8'b0;
    XRAM[7665] = 8'b0;
    XRAM[7666] = 8'b0;
    XRAM[7667] = 8'b0;
    XRAM[7668] = 8'b0;
    XRAM[7669] = 8'b0;
    XRAM[7670] = 8'b0;
    XRAM[7671] = 8'b0;
    XRAM[7672] = 8'b0;
    XRAM[7673] = 8'b0;
    XRAM[7674] = 8'b0;
    XRAM[7675] = 8'b0;
    XRAM[7676] = 8'b0;
    XRAM[7677] = 8'b0;
    XRAM[7678] = 8'b0;
    XRAM[7679] = 8'b0;
    XRAM[7680] = 8'b0;
    XRAM[7681] = 8'b0;
    XRAM[7682] = 8'b0;
    XRAM[7683] = 8'b0;
    XRAM[7684] = 8'b0;
    XRAM[7685] = 8'b0;
    XRAM[7686] = 8'b0;
    XRAM[7687] = 8'b0;
    XRAM[7688] = 8'b0;
    XRAM[7689] = 8'b0;
    XRAM[7690] = 8'b0;
    XRAM[7691] = 8'b0;
    XRAM[7692] = 8'b0;
    XRAM[7693] = 8'b0;
    XRAM[7694] = 8'b0;
    XRAM[7695] = 8'b0;
    XRAM[7696] = 8'b0;
    XRAM[7697] = 8'b0;
    XRAM[7698] = 8'b0;
    XRAM[7699] = 8'b0;
    XRAM[7700] = 8'b0;
    XRAM[7701] = 8'b0;
    XRAM[7702] = 8'b0;
    XRAM[7703] = 8'b0;
    XRAM[7704] = 8'b0;
    XRAM[7705] = 8'b0;
    XRAM[7706] = 8'b0;
    XRAM[7707] = 8'b0;
    XRAM[7708] = 8'b0;
    XRAM[7709] = 8'b0;
    XRAM[7710] = 8'b0;
    XRAM[7711] = 8'b0;
    XRAM[7712] = 8'b0;
    XRAM[7713] = 8'b0;
    XRAM[7714] = 8'b0;
    XRAM[7715] = 8'b0;
    XRAM[7716] = 8'b0;
    XRAM[7717] = 8'b0;
    XRAM[7718] = 8'b0;
    XRAM[7719] = 8'b0;
    XRAM[7720] = 8'b0;
    XRAM[7721] = 8'b0;
    XRAM[7722] = 8'b0;
    XRAM[7723] = 8'b0;
    XRAM[7724] = 8'b0;
    XRAM[7725] = 8'b0;
    XRAM[7726] = 8'b0;
    XRAM[7727] = 8'b0;
    XRAM[7728] = 8'b0;
    XRAM[7729] = 8'b0;
    XRAM[7730] = 8'b0;
    XRAM[7731] = 8'b0;
    XRAM[7732] = 8'b0;
    XRAM[7733] = 8'b0;
    XRAM[7734] = 8'b0;
    XRAM[7735] = 8'b0;
    XRAM[7736] = 8'b0;
    XRAM[7737] = 8'b0;
    XRAM[7738] = 8'b0;
    XRAM[7739] = 8'b0;
    XRAM[7740] = 8'b0;
    XRAM[7741] = 8'b0;
    XRAM[7742] = 8'b0;
    XRAM[7743] = 8'b0;
    XRAM[7744] = 8'b0;
    XRAM[7745] = 8'b0;
    XRAM[7746] = 8'b0;
    XRAM[7747] = 8'b0;
    XRAM[7748] = 8'b0;
    XRAM[7749] = 8'b0;
    XRAM[7750] = 8'b0;
    XRAM[7751] = 8'b0;
    XRAM[7752] = 8'b0;
    XRAM[7753] = 8'b0;
    XRAM[7754] = 8'b0;
    XRAM[7755] = 8'b0;
    XRAM[7756] = 8'b0;
    XRAM[7757] = 8'b0;
    XRAM[7758] = 8'b0;
    XRAM[7759] = 8'b0;
    XRAM[7760] = 8'b0;
    XRAM[7761] = 8'b0;
    XRAM[7762] = 8'b0;
    XRAM[7763] = 8'b0;
    XRAM[7764] = 8'b0;
    XRAM[7765] = 8'b0;
    XRAM[7766] = 8'b0;
    XRAM[7767] = 8'b0;
    XRAM[7768] = 8'b0;
    XRAM[7769] = 8'b0;
    XRAM[7770] = 8'b0;
    XRAM[7771] = 8'b0;
    XRAM[7772] = 8'b0;
    XRAM[7773] = 8'b0;
    XRAM[7774] = 8'b0;
    XRAM[7775] = 8'b0;
    XRAM[7776] = 8'b0;
    XRAM[7777] = 8'b0;
    XRAM[7778] = 8'b0;
    XRAM[7779] = 8'b0;
    XRAM[7780] = 8'b0;
    XRAM[7781] = 8'b0;
    XRAM[7782] = 8'b0;
    XRAM[7783] = 8'b0;
    XRAM[7784] = 8'b0;
    XRAM[7785] = 8'b0;
    XRAM[7786] = 8'b0;
    XRAM[7787] = 8'b0;
    XRAM[7788] = 8'b0;
    XRAM[7789] = 8'b0;
    XRAM[7790] = 8'b0;
    XRAM[7791] = 8'b0;
    XRAM[7792] = 8'b0;
    XRAM[7793] = 8'b0;
    XRAM[7794] = 8'b0;
    XRAM[7795] = 8'b0;
    XRAM[7796] = 8'b0;
    XRAM[7797] = 8'b0;
    XRAM[7798] = 8'b0;
    XRAM[7799] = 8'b0;
    XRAM[7800] = 8'b0;
    XRAM[7801] = 8'b0;
    XRAM[7802] = 8'b0;
    XRAM[7803] = 8'b0;
    XRAM[7804] = 8'b0;
    XRAM[7805] = 8'b0;
    XRAM[7806] = 8'b0;
    XRAM[7807] = 8'b0;
    XRAM[7808] = 8'b0;
    XRAM[7809] = 8'b0;
    XRAM[7810] = 8'b0;
    XRAM[7811] = 8'b0;
    XRAM[7812] = 8'b0;
    XRAM[7813] = 8'b0;
    XRAM[7814] = 8'b0;
    XRAM[7815] = 8'b0;
    XRAM[7816] = 8'b0;
    XRAM[7817] = 8'b0;
    XRAM[7818] = 8'b0;
    XRAM[7819] = 8'b0;
    XRAM[7820] = 8'b0;
    XRAM[7821] = 8'b0;
    XRAM[7822] = 8'b0;
    XRAM[7823] = 8'b0;
    XRAM[7824] = 8'b0;
    XRAM[7825] = 8'b0;
    XRAM[7826] = 8'b0;
    XRAM[7827] = 8'b0;
    XRAM[7828] = 8'b0;
    XRAM[7829] = 8'b0;
    XRAM[7830] = 8'b0;
    XRAM[7831] = 8'b0;
    XRAM[7832] = 8'b0;
    XRAM[7833] = 8'b0;
    XRAM[7834] = 8'b0;
    XRAM[7835] = 8'b0;
    XRAM[7836] = 8'b0;
    XRAM[7837] = 8'b0;
    XRAM[7838] = 8'b0;
    XRAM[7839] = 8'b0;
    XRAM[7840] = 8'b0;
    XRAM[7841] = 8'b0;
    XRAM[7842] = 8'b0;
    XRAM[7843] = 8'b0;
    XRAM[7844] = 8'b0;
    XRAM[7845] = 8'b0;
    XRAM[7846] = 8'b0;
    XRAM[7847] = 8'b0;
    XRAM[7848] = 8'b0;
    XRAM[7849] = 8'b0;
    XRAM[7850] = 8'b0;
    XRAM[7851] = 8'b0;
    XRAM[7852] = 8'b0;
    XRAM[7853] = 8'b0;
    XRAM[7854] = 8'b0;
    XRAM[7855] = 8'b0;
    XRAM[7856] = 8'b0;
    XRAM[7857] = 8'b0;
    XRAM[7858] = 8'b0;
    XRAM[7859] = 8'b0;
    XRAM[7860] = 8'b0;
    XRAM[7861] = 8'b0;
    XRAM[7862] = 8'b0;
    XRAM[7863] = 8'b0;
    XRAM[7864] = 8'b0;
    XRAM[7865] = 8'b0;
    XRAM[7866] = 8'b0;
    XRAM[7867] = 8'b0;
    XRAM[7868] = 8'b0;
    XRAM[7869] = 8'b0;
    XRAM[7870] = 8'b0;
    XRAM[7871] = 8'b0;
    XRAM[7872] = 8'b0;
    XRAM[7873] = 8'b0;
    XRAM[7874] = 8'b0;
    XRAM[7875] = 8'b0;
    XRAM[7876] = 8'b0;
    XRAM[7877] = 8'b0;
    XRAM[7878] = 8'b0;
    XRAM[7879] = 8'b0;
    XRAM[7880] = 8'b0;
    XRAM[7881] = 8'b0;
    XRAM[7882] = 8'b0;
    XRAM[7883] = 8'b0;
    XRAM[7884] = 8'b0;
    XRAM[7885] = 8'b0;
    XRAM[7886] = 8'b0;
    XRAM[7887] = 8'b0;
    XRAM[7888] = 8'b0;
    XRAM[7889] = 8'b0;
    XRAM[7890] = 8'b0;
    XRAM[7891] = 8'b0;
    XRAM[7892] = 8'b0;
    XRAM[7893] = 8'b0;
    XRAM[7894] = 8'b0;
    XRAM[7895] = 8'b0;
    XRAM[7896] = 8'b0;
    XRAM[7897] = 8'b0;
    XRAM[7898] = 8'b0;
    XRAM[7899] = 8'b0;
    XRAM[7900] = 8'b0;
    XRAM[7901] = 8'b0;
    XRAM[7902] = 8'b0;
    XRAM[7903] = 8'b0;
    XRAM[7904] = 8'b0;
    XRAM[7905] = 8'b0;
    XRAM[7906] = 8'b0;
    XRAM[7907] = 8'b0;
    XRAM[7908] = 8'b0;
    XRAM[7909] = 8'b0;
    XRAM[7910] = 8'b0;
    XRAM[7911] = 8'b0;
    XRAM[7912] = 8'b0;
    XRAM[7913] = 8'b0;
    XRAM[7914] = 8'b0;
    XRAM[7915] = 8'b0;
    XRAM[7916] = 8'b0;
    XRAM[7917] = 8'b0;
    XRAM[7918] = 8'b0;
    XRAM[7919] = 8'b0;
    XRAM[7920] = 8'b0;
    XRAM[7921] = 8'b0;
    XRAM[7922] = 8'b0;
    XRAM[7923] = 8'b0;
    XRAM[7924] = 8'b0;
    XRAM[7925] = 8'b0;
    XRAM[7926] = 8'b0;
    XRAM[7927] = 8'b0;
    XRAM[7928] = 8'b0;
    XRAM[7929] = 8'b0;
    XRAM[7930] = 8'b0;
    XRAM[7931] = 8'b0;
    XRAM[7932] = 8'b0;
    XRAM[7933] = 8'b0;
    XRAM[7934] = 8'b0;
    XRAM[7935] = 8'b0;
    XRAM[7936] = 8'b0;
    XRAM[7937] = 8'b0;
    XRAM[7938] = 8'b0;
    XRAM[7939] = 8'b0;
    XRAM[7940] = 8'b0;
    XRAM[7941] = 8'b0;
    XRAM[7942] = 8'b0;
    XRAM[7943] = 8'b0;
    XRAM[7944] = 8'b0;
    XRAM[7945] = 8'b0;
    XRAM[7946] = 8'b0;
    XRAM[7947] = 8'b0;
    XRAM[7948] = 8'b0;
    XRAM[7949] = 8'b0;
    XRAM[7950] = 8'b0;
    XRAM[7951] = 8'b0;
    XRAM[7952] = 8'b0;
    XRAM[7953] = 8'b0;
    XRAM[7954] = 8'b0;
    XRAM[7955] = 8'b0;
    XRAM[7956] = 8'b0;
    XRAM[7957] = 8'b0;
    XRAM[7958] = 8'b0;
    XRAM[7959] = 8'b0;
    XRAM[7960] = 8'b0;
    XRAM[7961] = 8'b0;
    XRAM[7962] = 8'b0;
    XRAM[7963] = 8'b0;
    XRAM[7964] = 8'b0;
    XRAM[7965] = 8'b0;
    XRAM[7966] = 8'b0;
    XRAM[7967] = 8'b0;
    XRAM[7968] = 8'b0;
    XRAM[7969] = 8'b0;
    XRAM[7970] = 8'b0;
    XRAM[7971] = 8'b0;
    XRAM[7972] = 8'b0;
    XRAM[7973] = 8'b0;
    XRAM[7974] = 8'b0;
    XRAM[7975] = 8'b0;
    XRAM[7976] = 8'b0;
    XRAM[7977] = 8'b0;
    XRAM[7978] = 8'b0;
    XRAM[7979] = 8'b0;
    XRAM[7980] = 8'b0;
    XRAM[7981] = 8'b0;
    XRAM[7982] = 8'b0;
    XRAM[7983] = 8'b0;
    XRAM[7984] = 8'b0;
    XRAM[7985] = 8'b0;
    XRAM[7986] = 8'b0;
    XRAM[7987] = 8'b0;
    XRAM[7988] = 8'b0;
    XRAM[7989] = 8'b0;
    XRAM[7990] = 8'b0;
    XRAM[7991] = 8'b0;
    XRAM[7992] = 8'b0;
    XRAM[7993] = 8'b0;
    XRAM[7994] = 8'b0;
    XRAM[7995] = 8'b0;
    XRAM[7996] = 8'b0;
    XRAM[7997] = 8'b0;
    XRAM[7998] = 8'b0;
    XRAM[7999] = 8'b0;
    XRAM[8000] = 8'b0;
    XRAM[8001] = 8'b0;
    XRAM[8002] = 8'b0;
    XRAM[8003] = 8'b0;
    XRAM[8004] = 8'b0;
    XRAM[8005] = 8'b0;
    XRAM[8006] = 8'b0;
    XRAM[8007] = 8'b0;
    XRAM[8008] = 8'b0;
    XRAM[8009] = 8'b0;
    XRAM[8010] = 8'b0;
    XRAM[8011] = 8'b0;
    XRAM[8012] = 8'b0;
    XRAM[8013] = 8'b0;
    XRAM[8014] = 8'b0;
    XRAM[8015] = 8'b0;
    XRAM[8016] = 8'b0;
    XRAM[8017] = 8'b0;
    XRAM[8018] = 8'b0;
    XRAM[8019] = 8'b0;
    XRAM[8020] = 8'b0;
    XRAM[8021] = 8'b0;
    XRAM[8022] = 8'b0;
    XRAM[8023] = 8'b0;
    XRAM[8024] = 8'b0;
    XRAM[8025] = 8'b0;
    XRAM[8026] = 8'b0;
    XRAM[8027] = 8'b0;
    XRAM[8028] = 8'b0;
    XRAM[8029] = 8'b0;
    XRAM[8030] = 8'b0;
    XRAM[8031] = 8'b0;
    XRAM[8032] = 8'b0;
    XRAM[8033] = 8'b0;
    XRAM[8034] = 8'b0;
    XRAM[8035] = 8'b0;
    XRAM[8036] = 8'b0;
    XRAM[8037] = 8'b0;
    XRAM[8038] = 8'b0;
    XRAM[8039] = 8'b0;
    XRAM[8040] = 8'b0;
    XRAM[8041] = 8'b0;
    XRAM[8042] = 8'b0;
    XRAM[8043] = 8'b0;
    XRAM[8044] = 8'b0;
    XRAM[8045] = 8'b0;
    XRAM[8046] = 8'b0;
    XRAM[8047] = 8'b0;
    XRAM[8048] = 8'b0;
    XRAM[8049] = 8'b0;
    XRAM[8050] = 8'b0;
    XRAM[8051] = 8'b0;
    XRAM[8052] = 8'b0;
    XRAM[8053] = 8'b0;
    XRAM[8054] = 8'b0;
    XRAM[8055] = 8'b0;
    XRAM[8056] = 8'b0;
    XRAM[8057] = 8'b0;
    XRAM[8058] = 8'b0;
    XRAM[8059] = 8'b0;
    XRAM[8060] = 8'b0;
    XRAM[8061] = 8'b0;
    XRAM[8062] = 8'b0;
    XRAM[8063] = 8'b0;
    XRAM[8064] = 8'b0;
    XRAM[8065] = 8'b0;
    XRAM[8066] = 8'b0;
    XRAM[8067] = 8'b0;
    XRAM[8068] = 8'b0;
    XRAM[8069] = 8'b0;
    XRAM[8070] = 8'b0;
    XRAM[8071] = 8'b0;
    XRAM[8072] = 8'b0;
    XRAM[8073] = 8'b0;
    XRAM[8074] = 8'b0;
    XRAM[8075] = 8'b0;
    XRAM[8076] = 8'b0;
    XRAM[8077] = 8'b0;
    XRAM[8078] = 8'b0;
    XRAM[8079] = 8'b0;
    XRAM[8080] = 8'b0;
    XRAM[8081] = 8'b0;
    XRAM[8082] = 8'b0;
    XRAM[8083] = 8'b0;
    XRAM[8084] = 8'b0;
    XRAM[8085] = 8'b0;
    XRAM[8086] = 8'b0;
    XRAM[8087] = 8'b0;
    XRAM[8088] = 8'b0;
    XRAM[8089] = 8'b0;
    XRAM[8090] = 8'b0;
    XRAM[8091] = 8'b0;
    XRAM[8092] = 8'b0;
    XRAM[8093] = 8'b0;
    XRAM[8094] = 8'b0;
    XRAM[8095] = 8'b0;
    XRAM[8096] = 8'b0;
    XRAM[8097] = 8'b0;
    XRAM[8098] = 8'b0;
    XRAM[8099] = 8'b0;
    XRAM[8100] = 8'b0;
    XRAM[8101] = 8'b0;
    XRAM[8102] = 8'b0;
    XRAM[8103] = 8'b0;
    XRAM[8104] = 8'b0;
    XRAM[8105] = 8'b0;
    XRAM[8106] = 8'b0;
    XRAM[8107] = 8'b0;
    XRAM[8108] = 8'b0;
    XRAM[8109] = 8'b0;
    XRAM[8110] = 8'b0;
    XRAM[8111] = 8'b0;
    XRAM[8112] = 8'b0;
    XRAM[8113] = 8'b0;
    XRAM[8114] = 8'b0;
    XRAM[8115] = 8'b0;
    XRAM[8116] = 8'b0;
    XRAM[8117] = 8'b0;
    XRAM[8118] = 8'b0;
    XRAM[8119] = 8'b0;
    XRAM[8120] = 8'b0;
    XRAM[8121] = 8'b0;
    XRAM[8122] = 8'b0;
    XRAM[8123] = 8'b0;
    XRAM[8124] = 8'b0;
    XRAM[8125] = 8'b0;
    XRAM[8126] = 8'b0;
    XRAM[8127] = 8'b0;
    XRAM[8128] = 8'b0;
    XRAM[8129] = 8'b0;
    XRAM[8130] = 8'b0;
    XRAM[8131] = 8'b0;
    XRAM[8132] = 8'b0;
    XRAM[8133] = 8'b0;
    XRAM[8134] = 8'b0;
    XRAM[8135] = 8'b0;
    XRAM[8136] = 8'b0;
    XRAM[8137] = 8'b0;
    XRAM[8138] = 8'b0;
    XRAM[8139] = 8'b0;
    XRAM[8140] = 8'b0;
    XRAM[8141] = 8'b0;
    XRAM[8142] = 8'b0;
    XRAM[8143] = 8'b0;
    XRAM[8144] = 8'b0;
    XRAM[8145] = 8'b0;
    XRAM[8146] = 8'b0;
    XRAM[8147] = 8'b0;
    XRAM[8148] = 8'b0;
    XRAM[8149] = 8'b0;
    XRAM[8150] = 8'b0;
    XRAM[8151] = 8'b0;
    XRAM[8152] = 8'b0;
    XRAM[8153] = 8'b0;
    XRAM[8154] = 8'b0;
    XRAM[8155] = 8'b0;
    XRAM[8156] = 8'b0;
    XRAM[8157] = 8'b0;
    XRAM[8158] = 8'b0;
    XRAM[8159] = 8'b0;
    XRAM[8160] = 8'b0;
    XRAM[8161] = 8'b0;
    XRAM[8162] = 8'b0;
    XRAM[8163] = 8'b0;
    XRAM[8164] = 8'b0;
    XRAM[8165] = 8'b0;
    XRAM[8166] = 8'b0;
    XRAM[8167] = 8'b0;
    XRAM[8168] = 8'b0;
    XRAM[8169] = 8'b0;
    XRAM[8170] = 8'b0;
    XRAM[8171] = 8'b0;
    XRAM[8172] = 8'b0;
    XRAM[8173] = 8'b0;
    XRAM[8174] = 8'b0;
    XRAM[8175] = 8'b0;
    XRAM[8176] = 8'b0;
    XRAM[8177] = 8'b0;
    XRAM[8178] = 8'b0;
    XRAM[8179] = 8'b0;
    XRAM[8180] = 8'b0;
    XRAM[8181] = 8'b0;
    XRAM[8182] = 8'b0;
    XRAM[8183] = 8'b0;
    XRAM[8184] = 8'b0;
    XRAM[8185] = 8'b0;
    XRAM[8186] = 8'b0;
    XRAM[8187] = 8'b0;
    XRAM[8188] = 8'b0;
    XRAM[8189] = 8'b0;
    XRAM[8190] = 8'b0;
    XRAM[8191] = 8'b0;
    XRAM[8192] = 8'b0;
    XRAM[8193] = 8'b0;
    XRAM[8194] = 8'b0;
    XRAM[8195] = 8'b0;
    XRAM[8196] = 8'b0;
    XRAM[8197] = 8'b0;
    XRAM[8198] = 8'b0;
    XRAM[8199] = 8'b0;
    XRAM[8200] = 8'b0;
    XRAM[8201] = 8'b0;
    XRAM[8202] = 8'b0;
    XRAM[8203] = 8'b0;
    XRAM[8204] = 8'b0;
    XRAM[8205] = 8'b0;
    XRAM[8206] = 8'b0;
    XRAM[8207] = 8'b0;
    XRAM[8208] = 8'b0;
    XRAM[8209] = 8'b0;
    XRAM[8210] = 8'b0;
    XRAM[8211] = 8'b0;
    XRAM[8212] = 8'b0;
    XRAM[8213] = 8'b0;
    XRAM[8214] = 8'b0;
    XRAM[8215] = 8'b0;
    XRAM[8216] = 8'b0;
    XRAM[8217] = 8'b0;
    XRAM[8218] = 8'b0;
    XRAM[8219] = 8'b0;
    XRAM[8220] = 8'b0;
    XRAM[8221] = 8'b0;
    XRAM[8222] = 8'b0;
    XRAM[8223] = 8'b0;
    XRAM[8224] = 8'b0;
    XRAM[8225] = 8'b0;
    XRAM[8226] = 8'b0;
    XRAM[8227] = 8'b0;
    XRAM[8228] = 8'b0;
    XRAM[8229] = 8'b0;
    XRAM[8230] = 8'b0;
    XRAM[8231] = 8'b0;
    XRAM[8232] = 8'b0;
    XRAM[8233] = 8'b0;
    XRAM[8234] = 8'b0;
    XRAM[8235] = 8'b0;
    XRAM[8236] = 8'b0;
    XRAM[8237] = 8'b0;
    XRAM[8238] = 8'b0;
    XRAM[8239] = 8'b0;
    XRAM[8240] = 8'b0;
    XRAM[8241] = 8'b0;
    XRAM[8242] = 8'b0;
    XRAM[8243] = 8'b0;
    XRAM[8244] = 8'b0;
    XRAM[8245] = 8'b0;
    XRAM[8246] = 8'b0;
    XRAM[8247] = 8'b0;
    XRAM[8248] = 8'b0;
    XRAM[8249] = 8'b0;
    XRAM[8250] = 8'b0;
    XRAM[8251] = 8'b0;
    XRAM[8252] = 8'b0;
    XRAM[8253] = 8'b0;
    XRAM[8254] = 8'b0;
    XRAM[8255] = 8'b0;
    XRAM[8256] = 8'b0;
    XRAM[8257] = 8'b0;
    XRAM[8258] = 8'b0;
    XRAM[8259] = 8'b0;
    XRAM[8260] = 8'b0;
    XRAM[8261] = 8'b0;
    XRAM[8262] = 8'b0;
    XRAM[8263] = 8'b0;
    XRAM[8264] = 8'b0;
    XRAM[8265] = 8'b0;
    XRAM[8266] = 8'b0;
    XRAM[8267] = 8'b0;
    XRAM[8268] = 8'b0;
    XRAM[8269] = 8'b0;
    XRAM[8270] = 8'b0;
    XRAM[8271] = 8'b0;
    XRAM[8272] = 8'b0;
    XRAM[8273] = 8'b0;
    XRAM[8274] = 8'b0;
    XRAM[8275] = 8'b0;
    XRAM[8276] = 8'b0;
    XRAM[8277] = 8'b0;
    XRAM[8278] = 8'b0;
    XRAM[8279] = 8'b0;
    XRAM[8280] = 8'b0;
    XRAM[8281] = 8'b0;
    XRAM[8282] = 8'b0;
    XRAM[8283] = 8'b0;
    XRAM[8284] = 8'b0;
    XRAM[8285] = 8'b0;
    XRAM[8286] = 8'b0;
    XRAM[8287] = 8'b0;
    XRAM[8288] = 8'b0;
    XRAM[8289] = 8'b0;
    XRAM[8290] = 8'b0;
    XRAM[8291] = 8'b0;
    XRAM[8292] = 8'b0;
    XRAM[8293] = 8'b0;
    XRAM[8294] = 8'b0;
    XRAM[8295] = 8'b0;
    XRAM[8296] = 8'b0;
    XRAM[8297] = 8'b0;
    XRAM[8298] = 8'b0;
    XRAM[8299] = 8'b0;
    XRAM[8300] = 8'b0;
    XRAM[8301] = 8'b0;
    XRAM[8302] = 8'b0;
    XRAM[8303] = 8'b0;
    XRAM[8304] = 8'b0;
    XRAM[8305] = 8'b0;
    XRAM[8306] = 8'b0;
    XRAM[8307] = 8'b0;
    XRAM[8308] = 8'b0;
    XRAM[8309] = 8'b0;
    XRAM[8310] = 8'b0;
    XRAM[8311] = 8'b0;
    XRAM[8312] = 8'b0;
    XRAM[8313] = 8'b0;
    XRAM[8314] = 8'b0;
    XRAM[8315] = 8'b0;
    XRAM[8316] = 8'b0;
    XRAM[8317] = 8'b0;
    XRAM[8318] = 8'b0;
    XRAM[8319] = 8'b0;
    XRAM[8320] = 8'b0;
    XRAM[8321] = 8'b0;
    XRAM[8322] = 8'b0;
    XRAM[8323] = 8'b0;
    XRAM[8324] = 8'b0;
    XRAM[8325] = 8'b0;
    XRAM[8326] = 8'b0;
    XRAM[8327] = 8'b0;
    XRAM[8328] = 8'b0;
    XRAM[8329] = 8'b0;
    XRAM[8330] = 8'b0;
    XRAM[8331] = 8'b0;
    XRAM[8332] = 8'b0;
    XRAM[8333] = 8'b0;
    XRAM[8334] = 8'b0;
    XRAM[8335] = 8'b0;
    XRAM[8336] = 8'b0;
    XRAM[8337] = 8'b0;
    XRAM[8338] = 8'b0;
    XRAM[8339] = 8'b0;
    XRAM[8340] = 8'b0;
    XRAM[8341] = 8'b0;
    XRAM[8342] = 8'b0;
    XRAM[8343] = 8'b0;
    XRAM[8344] = 8'b0;
    XRAM[8345] = 8'b0;
    XRAM[8346] = 8'b0;
    XRAM[8347] = 8'b0;
    XRAM[8348] = 8'b0;
    XRAM[8349] = 8'b0;
    XRAM[8350] = 8'b0;
    XRAM[8351] = 8'b0;
    XRAM[8352] = 8'b0;
    XRAM[8353] = 8'b0;
    XRAM[8354] = 8'b0;
    XRAM[8355] = 8'b0;
    XRAM[8356] = 8'b0;
    XRAM[8357] = 8'b0;
    XRAM[8358] = 8'b0;
    XRAM[8359] = 8'b0;
    XRAM[8360] = 8'b0;
    XRAM[8361] = 8'b0;
    XRAM[8362] = 8'b0;
    XRAM[8363] = 8'b0;
    XRAM[8364] = 8'b0;
    XRAM[8365] = 8'b0;
    XRAM[8366] = 8'b0;
    XRAM[8367] = 8'b0;
    XRAM[8368] = 8'b0;
    XRAM[8369] = 8'b0;
    XRAM[8370] = 8'b0;
    XRAM[8371] = 8'b0;
    XRAM[8372] = 8'b0;
    XRAM[8373] = 8'b0;
    XRAM[8374] = 8'b0;
    XRAM[8375] = 8'b0;
    XRAM[8376] = 8'b0;
    XRAM[8377] = 8'b0;
    XRAM[8378] = 8'b0;
    XRAM[8379] = 8'b0;
    XRAM[8380] = 8'b0;
    XRAM[8381] = 8'b0;
    XRAM[8382] = 8'b0;
    XRAM[8383] = 8'b0;
    XRAM[8384] = 8'b0;
    XRAM[8385] = 8'b0;
    XRAM[8386] = 8'b0;
    XRAM[8387] = 8'b0;
    XRAM[8388] = 8'b0;
    XRAM[8389] = 8'b0;
    XRAM[8390] = 8'b0;
    XRAM[8391] = 8'b0;
    XRAM[8392] = 8'b0;
    XRAM[8393] = 8'b0;
    XRAM[8394] = 8'b0;
    XRAM[8395] = 8'b0;
    XRAM[8396] = 8'b0;
    XRAM[8397] = 8'b0;
    XRAM[8398] = 8'b0;
    XRAM[8399] = 8'b0;
    XRAM[8400] = 8'b0;
    XRAM[8401] = 8'b0;
    XRAM[8402] = 8'b0;
    XRAM[8403] = 8'b0;
    XRAM[8404] = 8'b0;
    XRAM[8405] = 8'b0;
    XRAM[8406] = 8'b0;
    XRAM[8407] = 8'b0;
    XRAM[8408] = 8'b0;
    XRAM[8409] = 8'b0;
    XRAM[8410] = 8'b0;
    XRAM[8411] = 8'b0;
    XRAM[8412] = 8'b0;
    XRAM[8413] = 8'b0;
    XRAM[8414] = 8'b0;
    XRAM[8415] = 8'b0;
    XRAM[8416] = 8'b0;
    XRAM[8417] = 8'b0;
    XRAM[8418] = 8'b0;
    XRAM[8419] = 8'b0;
    XRAM[8420] = 8'b0;
    XRAM[8421] = 8'b0;
    XRAM[8422] = 8'b0;
    XRAM[8423] = 8'b0;
    XRAM[8424] = 8'b0;
    XRAM[8425] = 8'b0;
    XRAM[8426] = 8'b0;
    XRAM[8427] = 8'b0;
    XRAM[8428] = 8'b0;
    XRAM[8429] = 8'b0;
    XRAM[8430] = 8'b0;
    XRAM[8431] = 8'b0;
    XRAM[8432] = 8'b0;
    XRAM[8433] = 8'b0;
    XRAM[8434] = 8'b0;
    XRAM[8435] = 8'b0;
    XRAM[8436] = 8'b0;
    XRAM[8437] = 8'b0;
    XRAM[8438] = 8'b0;
    XRAM[8439] = 8'b0;
    XRAM[8440] = 8'b0;
    XRAM[8441] = 8'b0;
    XRAM[8442] = 8'b0;
    XRAM[8443] = 8'b0;
    XRAM[8444] = 8'b0;
    XRAM[8445] = 8'b0;
    XRAM[8446] = 8'b0;
    XRAM[8447] = 8'b0;
    XRAM[8448] = 8'b0;
    XRAM[8449] = 8'b0;
    XRAM[8450] = 8'b0;
    XRAM[8451] = 8'b0;
    XRAM[8452] = 8'b0;
    XRAM[8453] = 8'b0;
    XRAM[8454] = 8'b0;
    XRAM[8455] = 8'b0;
    XRAM[8456] = 8'b0;
    XRAM[8457] = 8'b0;
    XRAM[8458] = 8'b0;
    XRAM[8459] = 8'b0;
    XRAM[8460] = 8'b0;
    XRAM[8461] = 8'b0;
    XRAM[8462] = 8'b0;
    XRAM[8463] = 8'b0;
    XRAM[8464] = 8'b0;
    XRAM[8465] = 8'b0;
    XRAM[8466] = 8'b0;
    XRAM[8467] = 8'b0;
    XRAM[8468] = 8'b0;
    XRAM[8469] = 8'b0;
    XRAM[8470] = 8'b0;
    XRAM[8471] = 8'b0;
    XRAM[8472] = 8'b0;
    XRAM[8473] = 8'b0;
    XRAM[8474] = 8'b0;
    XRAM[8475] = 8'b0;
    XRAM[8476] = 8'b0;
    XRAM[8477] = 8'b0;
    XRAM[8478] = 8'b0;
    XRAM[8479] = 8'b0;
    XRAM[8480] = 8'b0;
    XRAM[8481] = 8'b0;
    XRAM[8482] = 8'b0;
    XRAM[8483] = 8'b0;
    XRAM[8484] = 8'b0;
    XRAM[8485] = 8'b0;
    XRAM[8486] = 8'b0;
    XRAM[8487] = 8'b0;
    XRAM[8488] = 8'b0;
    XRAM[8489] = 8'b0;
    XRAM[8490] = 8'b0;
    XRAM[8491] = 8'b0;
    XRAM[8492] = 8'b0;
    XRAM[8493] = 8'b0;
    XRAM[8494] = 8'b0;
    XRAM[8495] = 8'b0;
    XRAM[8496] = 8'b0;
    XRAM[8497] = 8'b0;
    XRAM[8498] = 8'b0;
    XRAM[8499] = 8'b0;
    XRAM[8500] = 8'b0;
    XRAM[8501] = 8'b0;
    XRAM[8502] = 8'b0;
    XRAM[8503] = 8'b0;
    XRAM[8504] = 8'b0;
    XRAM[8505] = 8'b0;
    XRAM[8506] = 8'b0;
    XRAM[8507] = 8'b0;
    XRAM[8508] = 8'b0;
    XRAM[8509] = 8'b0;
    XRAM[8510] = 8'b0;
    XRAM[8511] = 8'b0;
    XRAM[8512] = 8'b0;
    XRAM[8513] = 8'b0;
    XRAM[8514] = 8'b0;
    XRAM[8515] = 8'b0;
    XRAM[8516] = 8'b0;
    XRAM[8517] = 8'b0;
    XRAM[8518] = 8'b0;
    XRAM[8519] = 8'b0;
    XRAM[8520] = 8'b0;
    XRAM[8521] = 8'b0;
    XRAM[8522] = 8'b0;
    XRAM[8523] = 8'b0;
    XRAM[8524] = 8'b0;
    XRAM[8525] = 8'b0;
    XRAM[8526] = 8'b0;
    XRAM[8527] = 8'b0;
    XRAM[8528] = 8'b0;
    XRAM[8529] = 8'b0;
    XRAM[8530] = 8'b0;
    XRAM[8531] = 8'b0;
    XRAM[8532] = 8'b0;
    XRAM[8533] = 8'b0;
    XRAM[8534] = 8'b0;
    XRAM[8535] = 8'b0;
    XRAM[8536] = 8'b0;
    XRAM[8537] = 8'b0;
    XRAM[8538] = 8'b0;
    XRAM[8539] = 8'b0;
    XRAM[8540] = 8'b0;
    XRAM[8541] = 8'b0;
    XRAM[8542] = 8'b0;
    XRAM[8543] = 8'b0;
    XRAM[8544] = 8'b0;
    XRAM[8545] = 8'b0;
    XRAM[8546] = 8'b0;
    XRAM[8547] = 8'b0;
    XRAM[8548] = 8'b0;
    XRAM[8549] = 8'b0;
    XRAM[8550] = 8'b0;
    XRAM[8551] = 8'b0;
    XRAM[8552] = 8'b0;
    XRAM[8553] = 8'b0;
    XRAM[8554] = 8'b0;
    XRAM[8555] = 8'b0;
    XRAM[8556] = 8'b0;
    XRAM[8557] = 8'b0;
    XRAM[8558] = 8'b0;
    XRAM[8559] = 8'b0;
    XRAM[8560] = 8'b0;
    XRAM[8561] = 8'b0;
    XRAM[8562] = 8'b0;
    XRAM[8563] = 8'b0;
    XRAM[8564] = 8'b0;
    XRAM[8565] = 8'b0;
    XRAM[8566] = 8'b0;
    XRAM[8567] = 8'b0;
    XRAM[8568] = 8'b0;
    XRAM[8569] = 8'b0;
    XRAM[8570] = 8'b0;
    XRAM[8571] = 8'b0;
    XRAM[8572] = 8'b0;
    XRAM[8573] = 8'b0;
    XRAM[8574] = 8'b0;
    XRAM[8575] = 8'b0;
    XRAM[8576] = 8'b0;
    XRAM[8577] = 8'b0;
    XRAM[8578] = 8'b0;
    XRAM[8579] = 8'b0;
    XRAM[8580] = 8'b0;
    XRAM[8581] = 8'b0;
    XRAM[8582] = 8'b0;
    XRAM[8583] = 8'b0;
    XRAM[8584] = 8'b0;
    XRAM[8585] = 8'b0;
    XRAM[8586] = 8'b0;
    XRAM[8587] = 8'b0;
    XRAM[8588] = 8'b0;
    XRAM[8589] = 8'b0;
    XRAM[8590] = 8'b0;
    XRAM[8591] = 8'b0;
    XRAM[8592] = 8'b0;
    XRAM[8593] = 8'b0;
    XRAM[8594] = 8'b0;
    XRAM[8595] = 8'b0;
    XRAM[8596] = 8'b0;
    XRAM[8597] = 8'b0;
    XRAM[8598] = 8'b0;
    XRAM[8599] = 8'b0;
    XRAM[8600] = 8'b0;
    XRAM[8601] = 8'b0;
    XRAM[8602] = 8'b0;
    XRAM[8603] = 8'b0;
    XRAM[8604] = 8'b0;
    XRAM[8605] = 8'b0;
    XRAM[8606] = 8'b0;
    XRAM[8607] = 8'b0;
    XRAM[8608] = 8'b0;
    XRAM[8609] = 8'b0;
    XRAM[8610] = 8'b0;
    XRAM[8611] = 8'b0;
    XRAM[8612] = 8'b0;
    XRAM[8613] = 8'b0;
    XRAM[8614] = 8'b0;
    XRAM[8615] = 8'b0;
    XRAM[8616] = 8'b0;
    XRAM[8617] = 8'b0;
    XRAM[8618] = 8'b0;
    XRAM[8619] = 8'b0;
    XRAM[8620] = 8'b0;
    XRAM[8621] = 8'b0;
    XRAM[8622] = 8'b0;
    XRAM[8623] = 8'b0;
    XRAM[8624] = 8'b0;
    XRAM[8625] = 8'b0;
    XRAM[8626] = 8'b0;
    XRAM[8627] = 8'b0;
    XRAM[8628] = 8'b0;
    XRAM[8629] = 8'b0;
    XRAM[8630] = 8'b0;
    XRAM[8631] = 8'b0;
    XRAM[8632] = 8'b0;
    XRAM[8633] = 8'b0;
    XRAM[8634] = 8'b0;
    XRAM[8635] = 8'b0;
    XRAM[8636] = 8'b0;
    XRAM[8637] = 8'b0;
    XRAM[8638] = 8'b0;
    XRAM[8639] = 8'b0;
    XRAM[8640] = 8'b0;
    XRAM[8641] = 8'b0;
    XRAM[8642] = 8'b0;
    XRAM[8643] = 8'b0;
    XRAM[8644] = 8'b0;
    XRAM[8645] = 8'b0;
    XRAM[8646] = 8'b0;
    XRAM[8647] = 8'b0;
    XRAM[8648] = 8'b0;
    XRAM[8649] = 8'b0;
    XRAM[8650] = 8'b0;
    XRAM[8651] = 8'b0;
    XRAM[8652] = 8'b0;
    XRAM[8653] = 8'b0;
    XRAM[8654] = 8'b0;
    XRAM[8655] = 8'b0;
    XRAM[8656] = 8'b0;
    XRAM[8657] = 8'b0;
    XRAM[8658] = 8'b0;
    XRAM[8659] = 8'b0;
    XRAM[8660] = 8'b0;
    XRAM[8661] = 8'b0;
    XRAM[8662] = 8'b0;
    XRAM[8663] = 8'b0;
    XRAM[8664] = 8'b0;
    XRAM[8665] = 8'b0;
    XRAM[8666] = 8'b0;
    XRAM[8667] = 8'b0;
    XRAM[8668] = 8'b0;
    XRAM[8669] = 8'b0;
    XRAM[8670] = 8'b0;
    XRAM[8671] = 8'b0;
    XRAM[8672] = 8'b0;
    XRAM[8673] = 8'b0;
    XRAM[8674] = 8'b0;
    XRAM[8675] = 8'b0;
    XRAM[8676] = 8'b0;
    XRAM[8677] = 8'b0;
    XRAM[8678] = 8'b0;
    XRAM[8679] = 8'b0;
    XRAM[8680] = 8'b0;
    XRAM[8681] = 8'b0;
    XRAM[8682] = 8'b0;
    XRAM[8683] = 8'b0;
    XRAM[8684] = 8'b0;
    XRAM[8685] = 8'b0;
    XRAM[8686] = 8'b0;
    XRAM[8687] = 8'b0;
    XRAM[8688] = 8'b0;
    XRAM[8689] = 8'b0;
    XRAM[8690] = 8'b0;
    XRAM[8691] = 8'b0;
    XRAM[8692] = 8'b0;
    XRAM[8693] = 8'b0;
    XRAM[8694] = 8'b0;
    XRAM[8695] = 8'b0;
    XRAM[8696] = 8'b0;
    XRAM[8697] = 8'b0;
    XRAM[8698] = 8'b0;
    XRAM[8699] = 8'b0;
    XRAM[8700] = 8'b0;
    XRAM[8701] = 8'b0;
    XRAM[8702] = 8'b0;
    XRAM[8703] = 8'b0;
    XRAM[8704] = 8'b0;
    XRAM[8705] = 8'b0;
    XRAM[8706] = 8'b0;
    XRAM[8707] = 8'b0;
    XRAM[8708] = 8'b0;
    XRAM[8709] = 8'b0;
    XRAM[8710] = 8'b0;
    XRAM[8711] = 8'b0;
    XRAM[8712] = 8'b0;
    XRAM[8713] = 8'b0;
    XRAM[8714] = 8'b0;
    XRAM[8715] = 8'b0;
    XRAM[8716] = 8'b0;
    XRAM[8717] = 8'b0;
    XRAM[8718] = 8'b0;
    XRAM[8719] = 8'b0;
    XRAM[8720] = 8'b0;
    XRAM[8721] = 8'b0;
    XRAM[8722] = 8'b0;
    XRAM[8723] = 8'b0;
    XRAM[8724] = 8'b0;
    XRAM[8725] = 8'b0;
    XRAM[8726] = 8'b0;
    XRAM[8727] = 8'b0;
    XRAM[8728] = 8'b0;
    XRAM[8729] = 8'b0;
    XRAM[8730] = 8'b0;
    XRAM[8731] = 8'b0;
    XRAM[8732] = 8'b0;
    XRAM[8733] = 8'b0;
    XRAM[8734] = 8'b0;
    XRAM[8735] = 8'b0;
    XRAM[8736] = 8'b0;
    XRAM[8737] = 8'b0;
    XRAM[8738] = 8'b0;
    XRAM[8739] = 8'b0;
    XRAM[8740] = 8'b0;
    XRAM[8741] = 8'b0;
    XRAM[8742] = 8'b0;
    XRAM[8743] = 8'b0;
    XRAM[8744] = 8'b0;
    XRAM[8745] = 8'b0;
    XRAM[8746] = 8'b0;
    XRAM[8747] = 8'b0;
    XRAM[8748] = 8'b0;
    XRAM[8749] = 8'b0;
    XRAM[8750] = 8'b0;
    XRAM[8751] = 8'b0;
    XRAM[8752] = 8'b0;
    XRAM[8753] = 8'b0;
    XRAM[8754] = 8'b0;
    XRAM[8755] = 8'b0;
    XRAM[8756] = 8'b0;
    XRAM[8757] = 8'b0;
    XRAM[8758] = 8'b0;
    XRAM[8759] = 8'b0;
    XRAM[8760] = 8'b0;
    XRAM[8761] = 8'b0;
    XRAM[8762] = 8'b0;
    XRAM[8763] = 8'b0;
    XRAM[8764] = 8'b0;
    XRAM[8765] = 8'b0;
    XRAM[8766] = 8'b0;
    XRAM[8767] = 8'b0;
    XRAM[8768] = 8'b0;
    XRAM[8769] = 8'b0;
    XRAM[8770] = 8'b0;
    XRAM[8771] = 8'b0;
    XRAM[8772] = 8'b0;
    XRAM[8773] = 8'b0;
    XRAM[8774] = 8'b0;
    XRAM[8775] = 8'b0;
    XRAM[8776] = 8'b0;
    XRAM[8777] = 8'b0;
    XRAM[8778] = 8'b0;
    XRAM[8779] = 8'b0;
    XRAM[8780] = 8'b0;
    XRAM[8781] = 8'b0;
    XRAM[8782] = 8'b0;
    XRAM[8783] = 8'b0;
    XRAM[8784] = 8'b0;
    XRAM[8785] = 8'b0;
    XRAM[8786] = 8'b0;
    XRAM[8787] = 8'b0;
    XRAM[8788] = 8'b0;
    XRAM[8789] = 8'b0;
    XRAM[8790] = 8'b0;
    XRAM[8791] = 8'b0;
    XRAM[8792] = 8'b0;
    XRAM[8793] = 8'b0;
    XRAM[8794] = 8'b0;
    XRAM[8795] = 8'b0;
    XRAM[8796] = 8'b0;
    XRAM[8797] = 8'b0;
    XRAM[8798] = 8'b0;
    XRAM[8799] = 8'b0;
    XRAM[8800] = 8'b0;
    XRAM[8801] = 8'b0;
    XRAM[8802] = 8'b0;
    XRAM[8803] = 8'b0;
    XRAM[8804] = 8'b0;
    XRAM[8805] = 8'b0;
    XRAM[8806] = 8'b0;
    XRAM[8807] = 8'b0;
    XRAM[8808] = 8'b0;
    XRAM[8809] = 8'b0;
    XRAM[8810] = 8'b0;
    XRAM[8811] = 8'b0;
    XRAM[8812] = 8'b0;
    XRAM[8813] = 8'b0;
    XRAM[8814] = 8'b0;
    XRAM[8815] = 8'b0;
    XRAM[8816] = 8'b0;
    XRAM[8817] = 8'b0;
    XRAM[8818] = 8'b0;
    XRAM[8819] = 8'b0;
    XRAM[8820] = 8'b0;
    XRAM[8821] = 8'b0;
    XRAM[8822] = 8'b0;
    XRAM[8823] = 8'b0;
    XRAM[8824] = 8'b0;
    XRAM[8825] = 8'b0;
    XRAM[8826] = 8'b0;
    XRAM[8827] = 8'b0;
    XRAM[8828] = 8'b0;
    XRAM[8829] = 8'b0;
    XRAM[8830] = 8'b0;
    XRAM[8831] = 8'b0;
    XRAM[8832] = 8'b0;
    XRAM[8833] = 8'b0;
    XRAM[8834] = 8'b0;
    XRAM[8835] = 8'b0;
    XRAM[8836] = 8'b0;
    XRAM[8837] = 8'b0;
    XRAM[8838] = 8'b0;
    XRAM[8839] = 8'b0;
    XRAM[8840] = 8'b0;
    XRAM[8841] = 8'b0;
    XRAM[8842] = 8'b0;
    XRAM[8843] = 8'b0;
    XRAM[8844] = 8'b0;
    XRAM[8845] = 8'b0;
    XRAM[8846] = 8'b0;
    XRAM[8847] = 8'b0;
    XRAM[8848] = 8'b0;
    XRAM[8849] = 8'b0;
    XRAM[8850] = 8'b0;
    XRAM[8851] = 8'b0;
    XRAM[8852] = 8'b0;
    XRAM[8853] = 8'b0;
    XRAM[8854] = 8'b0;
    XRAM[8855] = 8'b0;
    XRAM[8856] = 8'b0;
    XRAM[8857] = 8'b0;
    XRAM[8858] = 8'b0;
    XRAM[8859] = 8'b0;
    XRAM[8860] = 8'b0;
    XRAM[8861] = 8'b0;
    XRAM[8862] = 8'b0;
    XRAM[8863] = 8'b0;
    XRAM[8864] = 8'b0;
    XRAM[8865] = 8'b0;
    XRAM[8866] = 8'b0;
    XRAM[8867] = 8'b0;
    XRAM[8868] = 8'b0;
    XRAM[8869] = 8'b0;
    XRAM[8870] = 8'b0;
    XRAM[8871] = 8'b0;
    XRAM[8872] = 8'b0;
    XRAM[8873] = 8'b0;
    XRAM[8874] = 8'b0;
    XRAM[8875] = 8'b0;
    XRAM[8876] = 8'b0;
    XRAM[8877] = 8'b0;
    XRAM[8878] = 8'b0;
    XRAM[8879] = 8'b0;
    XRAM[8880] = 8'b0;
    XRAM[8881] = 8'b0;
    XRAM[8882] = 8'b0;
    XRAM[8883] = 8'b0;
    XRAM[8884] = 8'b0;
    XRAM[8885] = 8'b0;
    XRAM[8886] = 8'b0;
    XRAM[8887] = 8'b0;
    XRAM[8888] = 8'b0;
    XRAM[8889] = 8'b0;
    XRAM[8890] = 8'b0;
    XRAM[8891] = 8'b0;
    XRAM[8892] = 8'b0;
    XRAM[8893] = 8'b0;
    XRAM[8894] = 8'b0;
    XRAM[8895] = 8'b0;
    XRAM[8896] = 8'b0;
    XRAM[8897] = 8'b0;
    XRAM[8898] = 8'b0;
    XRAM[8899] = 8'b0;
    XRAM[8900] = 8'b0;
    XRAM[8901] = 8'b0;
    XRAM[8902] = 8'b0;
    XRAM[8903] = 8'b0;
    XRAM[8904] = 8'b0;
    XRAM[8905] = 8'b0;
    XRAM[8906] = 8'b0;
    XRAM[8907] = 8'b0;
    XRAM[8908] = 8'b0;
    XRAM[8909] = 8'b0;
    XRAM[8910] = 8'b0;
    XRAM[8911] = 8'b0;
    XRAM[8912] = 8'b0;
    XRAM[8913] = 8'b0;
    XRAM[8914] = 8'b0;
    XRAM[8915] = 8'b0;
    XRAM[8916] = 8'b0;
    XRAM[8917] = 8'b0;
    XRAM[8918] = 8'b0;
    XRAM[8919] = 8'b0;
    XRAM[8920] = 8'b0;
    XRAM[8921] = 8'b0;
    XRAM[8922] = 8'b0;
    XRAM[8923] = 8'b0;
    XRAM[8924] = 8'b0;
    XRAM[8925] = 8'b0;
    XRAM[8926] = 8'b0;
    XRAM[8927] = 8'b0;
    XRAM[8928] = 8'b0;
    XRAM[8929] = 8'b0;
    XRAM[8930] = 8'b0;
    XRAM[8931] = 8'b0;
    XRAM[8932] = 8'b0;
    XRAM[8933] = 8'b0;
    XRAM[8934] = 8'b0;
    XRAM[8935] = 8'b0;
    XRAM[8936] = 8'b0;
    XRAM[8937] = 8'b0;
    XRAM[8938] = 8'b0;
    XRAM[8939] = 8'b0;
    XRAM[8940] = 8'b0;
    XRAM[8941] = 8'b0;
    XRAM[8942] = 8'b0;
    XRAM[8943] = 8'b0;
    XRAM[8944] = 8'b0;
    XRAM[8945] = 8'b0;
    XRAM[8946] = 8'b0;
    XRAM[8947] = 8'b0;
    XRAM[8948] = 8'b0;
    XRAM[8949] = 8'b0;
    XRAM[8950] = 8'b0;
    XRAM[8951] = 8'b0;
    XRAM[8952] = 8'b0;
    XRAM[8953] = 8'b0;
    XRAM[8954] = 8'b0;
    XRAM[8955] = 8'b0;
    XRAM[8956] = 8'b0;
    XRAM[8957] = 8'b0;
    XRAM[8958] = 8'b0;
    XRAM[8959] = 8'b0;
    XRAM[8960] = 8'b0;
    XRAM[8961] = 8'b0;
    XRAM[8962] = 8'b0;
    XRAM[8963] = 8'b0;
    XRAM[8964] = 8'b0;
    XRAM[8965] = 8'b0;
    XRAM[8966] = 8'b0;
    XRAM[8967] = 8'b0;
    XRAM[8968] = 8'b0;
    XRAM[8969] = 8'b0;
    XRAM[8970] = 8'b0;
    XRAM[8971] = 8'b0;
    XRAM[8972] = 8'b0;
    XRAM[8973] = 8'b0;
    XRAM[8974] = 8'b0;
    XRAM[8975] = 8'b0;
    XRAM[8976] = 8'b0;
    XRAM[8977] = 8'b0;
    XRAM[8978] = 8'b0;
    XRAM[8979] = 8'b0;
    XRAM[8980] = 8'b0;
    XRAM[8981] = 8'b0;
    XRAM[8982] = 8'b0;
    XRAM[8983] = 8'b0;
    XRAM[8984] = 8'b0;
    XRAM[8985] = 8'b0;
    XRAM[8986] = 8'b0;
    XRAM[8987] = 8'b0;
    XRAM[8988] = 8'b0;
    XRAM[8989] = 8'b0;
    XRAM[8990] = 8'b0;
    XRAM[8991] = 8'b0;
    XRAM[8992] = 8'b0;
    XRAM[8993] = 8'b0;
    XRAM[8994] = 8'b0;
    XRAM[8995] = 8'b0;
    XRAM[8996] = 8'b0;
    XRAM[8997] = 8'b0;
    XRAM[8998] = 8'b0;
    XRAM[8999] = 8'b0;
    XRAM[9000] = 8'b0;
    XRAM[9001] = 8'b0;
    XRAM[9002] = 8'b0;
    XRAM[9003] = 8'b0;
    XRAM[9004] = 8'b0;
    XRAM[9005] = 8'b0;
    XRAM[9006] = 8'b0;
    XRAM[9007] = 8'b0;
    XRAM[9008] = 8'b0;
    XRAM[9009] = 8'b0;
    XRAM[9010] = 8'b0;
    XRAM[9011] = 8'b0;
    XRAM[9012] = 8'b0;
    XRAM[9013] = 8'b0;
    XRAM[9014] = 8'b0;
    XRAM[9015] = 8'b0;
    XRAM[9016] = 8'b0;
    XRAM[9017] = 8'b0;
    XRAM[9018] = 8'b0;
    XRAM[9019] = 8'b0;
    XRAM[9020] = 8'b0;
    XRAM[9021] = 8'b0;
    XRAM[9022] = 8'b0;
    XRAM[9023] = 8'b0;
    XRAM[9024] = 8'b0;
    XRAM[9025] = 8'b0;
    XRAM[9026] = 8'b0;
    XRAM[9027] = 8'b0;
    XRAM[9028] = 8'b0;
    XRAM[9029] = 8'b0;
    XRAM[9030] = 8'b0;
    XRAM[9031] = 8'b0;
    XRAM[9032] = 8'b0;
    XRAM[9033] = 8'b0;
    XRAM[9034] = 8'b0;
    XRAM[9035] = 8'b0;
    XRAM[9036] = 8'b0;
    XRAM[9037] = 8'b0;
    XRAM[9038] = 8'b0;
    XRAM[9039] = 8'b0;
    XRAM[9040] = 8'b0;
    XRAM[9041] = 8'b0;
    XRAM[9042] = 8'b0;
    XRAM[9043] = 8'b0;
    XRAM[9044] = 8'b0;
    XRAM[9045] = 8'b0;
    XRAM[9046] = 8'b0;
    XRAM[9047] = 8'b0;
    XRAM[9048] = 8'b0;
    XRAM[9049] = 8'b0;
    XRAM[9050] = 8'b0;
    XRAM[9051] = 8'b0;
    XRAM[9052] = 8'b0;
    XRAM[9053] = 8'b0;
    XRAM[9054] = 8'b0;
    XRAM[9055] = 8'b0;
    XRAM[9056] = 8'b0;
    XRAM[9057] = 8'b0;
    XRAM[9058] = 8'b0;
    XRAM[9059] = 8'b0;
    XRAM[9060] = 8'b0;
    XRAM[9061] = 8'b0;
    XRAM[9062] = 8'b0;
    XRAM[9063] = 8'b0;
    XRAM[9064] = 8'b0;
    XRAM[9065] = 8'b0;
    XRAM[9066] = 8'b0;
    XRAM[9067] = 8'b0;
    XRAM[9068] = 8'b0;
    XRAM[9069] = 8'b0;
    XRAM[9070] = 8'b0;
    XRAM[9071] = 8'b0;
    XRAM[9072] = 8'b0;
    XRAM[9073] = 8'b0;
    XRAM[9074] = 8'b0;
    XRAM[9075] = 8'b0;
    XRAM[9076] = 8'b0;
    XRAM[9077] = 8'b0;
    XRAM[9078] = 8'b0;
    XRAM[9079] = 8'b0;
    XRAM[9080] = 8'b0;
    XRAM[9081] = 8'b0;
    XRAM[9082] = 8'b0;
    XRAM[9083] = 8'b0;
    XRAM[9084] = 8'b0;
    XRAM[9085] = 8'b0;
    XRAM[9086] = 8'b0;
    XRAM[9087] = 8'b0;
    XRAM[9088] = 8'b0;
    XRAM[9089] = 8'b0;
    XRAM[9090] = 8'b0;
    XRAM[9091] = 8'b0;
    XRAM[9092] = 8'b0;
    XRAM[9093] = 8'b0;
    XRAM[9094] = 8'b0;
    XRAM[9095] = 8'b0;
    XRAM[9096] = 8'b0;
    XRAM[9097] = 8'b0;
    XRAM[9098] = 8'b0;
    XRAM[9099] = 8'b0;
    XRAM[9100] = 8'b0;
    XRAM[9101] = 8'b0;
    XRAM[9102] = 8'b0;
    XRAM[9103] = 8'b0;
    XRAM[9104] = 8'b0;
    XRAM[9105] = 8'b0;
    XRAM[9106] = 8'b0;
    XRAM[9107] = 8'b0;
    XRAM[9108] = 8'b0;
    XRAM[9109] = 8'b0;
    XRAM[9110] = 8'b0;
    XRAM[9111] = 8'b0;
    XRAM[9112] = 8'b0;
    XRAM[9113] = 8'b0;
    XRAM[9114] = 8'b0;
    XRAM[9115] = 8'b0;
    XRAM[9116] = 8'b0;
    XRAM[9117] = 8'b0;
    XRAM[9118] = 8'b0;
    XRAM[9119] = 8'b0;
    XRAM[9120] = 8'b0;
    XRAM[9121] = 8'b0;
    XRAM[9122] = 8'b0;
    XRAM[9123] = 8'b0;
    XRAM[9124] = 8'b0;
    XRAM[9125] = 8'b0;
    XRAM[9126] = 8'b0;
    XRAM[9127] = 8'b0;
    XRAM[9128] = 8'b0;
    XRAM[9129] = 8'b0;
    XRAM[9130] = 8'b0;
    XRAM[9131] = 8'b0;
    XRAM[9132] = 8'b0;
    XRAM[9133] = 8'b0;
    XRAM[9134] = 8'b0;
    XRAM[9135] = 8'b0;
    XRAM[9136] = 8'b0;
    XRAM[9137] = 8'b0;
    XRAM[9138] = 8'b0;
    XRAM[9139] = 8'b0;
    XRAM[9140] = 8'b0;
    XRAM[9141] = 8'b0;
    XRAM[9142] = 8'b0;
    XRAM[9143] = 8'b0;
    XRAM[9144] = 8'b0;
    XRAM[9145] = 8'b0;
    XRAM[9146] = 8'b0;
    XRAM[9147] = 8'b0;
    XRAM[9148] = 8'b0;
    XRAM[9149] = 8'b0;
    XRAM[9150] = 8'b0;
    XRAM[9151] = 8'b0;
    XRAM[9152] = 8'b0;
    XRAM[9153] = 8'b0;
    XRAM[9154] = 8'b0;
    XRAM[9155] = 8'b0;
    XRAM[9156] = 8'b0;
    XRAM[9157] = 8'b0;
    XRAM[9158] = 8'b0;
    XRAM[9159] = 8'b0;
    XRAM[9160] = 8'b0;
    XRAM[9161] = 8'b0;
    XRAM[9162] = 8'b0;
    XRAM[9163] = 8'b0;
    XRAM[9164] = 8'b0;
    XRAM[9165] = 8'b0;
    XRAM[9166] = 8'b0;
    XRAM[9167] = 8'b0;
    XRAM[9168] = 8'b0;
    XRAM[9169] = 8'b0;
    XRAM[9170] = 8'b0;
    XRAM[9171] = 8'b0;
    XRAM[9172] = 8'b0;
    XRAM[9173] = 8'b0;
    XRAM[9174] = 8'b0;
    XRAM[9175] = 8'b0;
    XRAM[9176] = 8'b0;
    XRAM[9177] = 8'b0;
    XRAM[9178] = 8'b0;
    XRAM[9179] = 8'b0;
    XRAM[9180] = 8'b0;
    XRAM[9181] = 8'b0;
    XRAM[9182] = 8'b0;
    XRAM[9183] = 8'b0;
    XRAM[9184] = 8'b0;
    XRAM[9185] = 8'b0;
    XRAM[9186] = 8'b0;
    XRAM[9187] = 8'b0;
    XRAM[9188] = 8'b0;
    XRAM[9189] = 8'b0;
    XRAM[9190] = 8'b0;
    XRAM[9191] = 8'b0;
    XRAM[9192] = 8'b0;
    XRAM[9193] = 8'b0;
    XRAM[9194] = 8'b0;
    XRAM[9195] = 8'b0;
    XRAM[9196] = 8'b0;
    XRAM[9197] = 8'b0;
    XRAM[9198] = 8'b0;
    XRAM[9199] = 8'b0;
    XRAM[9200] = 8'b0;
    XRAM[9201] = 8'b0;
    XRAM[9202] = 8'b0;
    XRAM[9203] = 8'b0;
    XRAM[9204] = 8'b0;
    XRAM[9205] = 8'b0;
    XRAM[9206] = 8'b0;
    XRAM[9207] = 8'b0;
    XRAM[9208] = 8'b0;
    XRAM[9209] = 8'b0;
    XRAM[9210] = 8'b0;
    XRAM[9211] = 8'b0;
    XRAM[9212] = 8'b0;
    XRAM[9213] = 8'b0;
    XRAM[9214] = 8'b0;
    XRAM[9215] = 8'b0;
    XRAM[9216] = 8'b0;
    XRAM[9217] = 8'b0;
    XRAM[9218] = 8'b0;
    XRAM[9219] = 8'b0;
    XRAM[9220] = 8'b0;
    XRAM[9221] = 8'b0;
    XRAM[9222] = 8'b0;
    XRAM[9223] = 8'b0;
    XRAM[9224] = 8'b0;
    XRAM[9225] = 8'b0;
    XRAM[9226] = 8'b0;
    XRAM[9227] = 8'b0;
    XRAM[9228] = 8'b0;
    XRAM[9229] = 8'b0;
    XRAM[9230] = 8'b0;
    XRAM[9231] = 8'b0;
    XRAM[9232] = 8'b0;
    XRAM[9233] = 8'b0;
    XRAM[9234] = 8'b0;
    XRAM[9235] = 8'b0;
    XRAM[9236] = 8'b0;
    XRAM[9237] = 8'b0;
    XRAM[9238] = 8'b0;
    XRAM[9239] = 8'b0;
    XRAM[9240] = 8'b0;
    XRAM[9241] = 8'b0;
    XRAM[9242] = 8'b0;
    XRAM[9243] = 8'b0;
    XRAM[9244] = 8'b0;
    XRAM[9245] = 8'b0;
    XRAM[9246] = 8'b0;
    XRAM[9247] = 8'b0;
    XRAM[9248] = 8'b0;
    XRAM[9249] = 8'b0;
    XRAM[9250] = 8'b0;
    XRAM[9251] = 8'b0;
    XRAM[9252] = 8'b0;
    XRAM[9253] = 8'b0;
    XRAM[9254] = 8'b0;
    XRAM[9255] = 8'b0;
    XRAM[9256] = 8'b0;
    XRAM[9257] = 8'b0;
    XRAM[9258] = 8'b0;
    XRAM[9259] = 8'b0;
    XRAM[9260] = 8'b0;
    XRAM[9261] = 8'b0;
    XRAM[9262] = 8'b0;
    XRAM[9263] = 8'b0;
    XRAM[9264] = 8'b0;
    XRAM[9265] = 8'b0;
    XRAM[9266] = 8'b0;
    XRAM[9267] = 8'b0;
    XRAM[9268] = 8'b0;
    XRAM[9269] = 8'b0;
    XRAM[9270] = 8'b0;
    XRAM[9271] = 8'b0;
    XRAM[9272] = 8'b0;
    XRAM[9273] = 8'b0;
    XRAM[9274] = 8'b0;
    XRAM[9275] = 8'b0;
    XRAM[9276] = 8'b0;
    XRAM[9277] = 8'b0;
    XRAM[9278] = 8'b0;
    XRAM[9279] = 8'b0;
    XRAM[9280] = 8'b0;
    XRAM[9281] = 8'b0;
    XRAM[9282] = 8'b0;
    XRAM[9283] = 8'b0;
    XRAM[9284] = 8'b0;
    XRAM[9285] = 8'b0;
    XRAM[9286] = 8'b0;
    XRAM[9287] = 8'b0;
    XRAM[9288] = 8'b0;
    XRAM[9289] = 8'b0;
    XRAM[9290] = 8'b0;
    XRAM[9291] = 8'b0;
    XRAM[9292] = 8'b0;
    XRAM[9293] = 8'b0;
    XRAM[9294] = 8'b0;
    XRAM[9295] = 8'b0;
    XRAM[9296] = 8'b0;
    XRAM[9297] = 8'b0;
    XRAM[9298] = 8'b0;
    XRAM[9299] = 8'b0;
    XRAM[9300] = 8'b0;
    XRAM[9301] = 8'b0;
    XRAM[9302] = 8'b0;
    XRAM[9303] = 8'b0;
    XRAM[9304] = 8'b0;
    XRAM[9305] = 8'b0;
    XRAM[9306] = 8'b0;
    XRAM[9307] = 8'b0;
    XRAM[9308] = 8'b0;
    XRAM[9309] = 8'b0;
    XRAM[9310] = 8'b0;
    XRAM[9311] = 8'b0;
    XRAM[9312] = 8'b0;
    XRAM[9313] = 8'b0;
    XRAM[9314] = 8'b0;
    XRAM[9315] = 8'b0;
    XRAM[9316] = 8'b0;
    XRAM[9317] = 8'b0;
    XRAM[9318] = 8'b0;
    XRAM[9319] = 8'b0;
    XRAM[9320] = 8'b0;
    XRAM[9321] = 8'b0;
    XRAM[9322] = 8'b0;
    XRAM[9323] = 8'b0;
    XRAM[9324] = 8'b0;
    XRAM[9325] = 8'b0;
    XRAM[9326] = 8'b0;
    XRAM[9327] = 8'b0;
    XRAM[9328] = 8'b0;
    XRAM[9329] = 8'b0;
    XRAM[9330] = 8'b0;
    XRAM[9331] = 8'b0;
    XRAM[9332] = 8'b0;
    XRAM[9333] = 8'b0;
    XRAM[9334] = 8'b0;
    XRAM[9335] = 8'b0;
    XRAM[9336] = 8'b0;
    XRAM[9337] = 8'b0;
    XRAM[9338] = 8'b0;
    XRAM[9339] = 8'b0;
    XRAM[9340] = 8'b0;
    XRAM[9341] = 8'b0;
    XRAM[9342] = 8'b0;
    XRAM[9343] = 8'b0;
    XRAM[9344] = 8'b0;
    XRAM[9345] = 8'b0;
    XRAM[9346] = 8'b0;
    XRAM[9347] = 8'b0;
    XRAM[9348] = 8'b0;
    XRAM[9349] = 8'b0;
    XRAM[9350] = 8'b0;
    XRAM[9351] = 8'b0;
    XRAM[9352] = 8'b0;
    XRAM[9353] = 8'b0;
    XRAM[9354] = 8'b0;
    XRAM[9355] = 8'b0;
    XRAM[9356] = 8'b0;
    XRAM[9357] = 8'b0;
    XRAM[9358] = 8'b0;
    XRAM[9359] = 8'b0;
    XRAM[9360] = 8'b0;
    XRAM[9361] = 8'b0;
    XRAM[9362] = 8'b0;
    XRAM[9363] = 8'b0;
    XRAM[9364] = 8'b0;
    XRAM[9365] = 8'b0;
    XRAM[9366] = 8'b0;
    XRAM[9367] = 8'b0;
    XRAM[9368] = 8'b0;
    XRAM[9369] = 8'b0;
    XRAM[9370] = 8'b0;
    XRAM[9371] = 8'b0;
    XRAM[9372] = 8'b0;
    XRAM[9373] = 8'b0;
    XRAM[9374] = 8'b0;
    XRAM[9375] = 8'b0;
    XRAM[9376] = 8'b0;
    XRAM[9377] = 8'b0;
    XRAM[9378] = 8'b0;
    XRAM[9379] = 8'b0;
    XRAM[9380] = 8'b0;
    XRAM[9381] = 8'b0;
    XRAM[9382] = 8'b0;
    XRAM[9383] = 8'b0;
    XRAM[9384] = 8'b0;
    XRAM[9385] = 8'b0;
    XRAM[9386] = 8'b0;
    XRAM[9387] = 8'b0;
    XRAM[9388] = 8'b0;
    XRAM[9389] = 8'b0;
    XRAM[9390] = 8'b0;
    XRAM[9391] = 8'b0;
    XRAM[9392] = 8'b0;
    XRAM[9393] = 8'b0;
    XRAM[9394] = 8'b0;
    XRAM[9395] = 8'b0;
    XRAM[9396] = 8'b0;
    XRAM[9397] = 8'b0;
    XRAM[9398] = 8'b0;
    XRAM[9399] = 8'b0;
    XRAM[9400] = 8'b0;
    XRAM[9401] = 8'b0;
    XRAM[9402] = 8'b0;
    XRAM[9403] = 8'b0;
    XRAM[9404] = 8'b0;
    XRAM[9405] = 8'b0;
    XRAM[9406] = 8'b0;
    XRAM[9407] = 8'b0;
    XRAM[9408] = 8'b0;
    XRAM[9409] = 8'b0;
    XRAM[9410] = 8'b0;
    XRAM[9411] = 8'b0;
    XRAM[9412] = 8'b0;
    XRAM[9413] = 8'b0;
    XRAM[9414] = 8'b0;
    XRAM[9415] = 8'b0;
    XRAM[9416] = 8'b0;
    XRAM[9417] = 8'b0;
    XRAM[9418] = 8'b0;
    XRAM[9419] = 8'b0;
    XRAM[9420] = 8'b0;
    XRAM[9421] = 8'b0;
    XRAM[9422] = 8'b0;
    XRAM[9423] = 8'b0;
    XRAM[9424] = 8'b0;
    XRAM[9425] = 8'b0;
    XRAM[9426] = 8'b0;
    XRAM[9427] = 8'b0;
    XRAM[9428] = 8'b0;
    XRAM[9429] = 8'b0;
    XRAM[9430] = 8'b0;
    XRAM[9431] = 8'b0;
    XRAM[9432] = 8'b0;
    XRAM[9433] = 8'b0;
    XRAM[9434] = 8'b0;
    XRAM[9435] = 8'b0;
    XRAM[9436] = 8'b0;
    XRAM[9437] = 8'b0;
    XRAM[9438] = 8'b0;
    XRAM[9439] = 8'b0;
    XRAM[9440] = 8'b0;
    XRAM[9441] = 8'b0;
    XRAM[9442] = 8'b0;
    XRAM[9443] = 8'b0;
    XRAM[9444] = 8'b0;
    XRAM[9445] = 8'b0;
    XRAM[9446] = 8'b0;
    XRAM[9447] = 8'b0;
    XRAM[9448] = 8'b0;
    XRAM[9449] = 8'b0;
    XRAM[9450] = 8'b0;
    XRAM[9451] = 8'b0;
    XRAM[9452] = 8'b0;
    XRAM[9453] = 8'b0;
    XRAM[9454] = 8'b0;
    XRAM[9455] = 8'b0;
    XRAM[9456] = 8'b0;
    XRAM[9457] = 8'b0;
    XRAM[9458] = 8'b0;
    XRAM[9459] = 8'b0;
    XRAM[9460] = 8'b0;
    XRAM[9461] = 8'b0;
    XRAM[9462] = 8'b0;
    XRAM[9463] = 8'b0;
    XRAM[9464] = 8'b0;
    XRAM[9465] = 8'b0;
    XRAM[9466] = 8'b0;
    XRAM[9467] = 8'b0;
    XRAM[9468] = 8'b0;
    XRAM[9469] = 8'b0;
    XRAM[9470] = 8'b0;
    XRAM[9471] = 8'b0;
    XRAM[9472] = 8'b0;
    XRAM[9473] = 8'b0;
    XRAM[9474] = 8'b0;
    XRAM[9475] = 8'b0;
    XRAM[9476] = 8'b0;
    XRAM[9477] = 8'b0;
    XRAM[9478] = 8'b0;
    XRAM[9479] = 8'b0;
    XRAM[9480] = 8'b0;
    XRAM[9481] = 8'b0;
    XRAM[9482] = 8'b0;
    XRAM[9483] = 8'b0;
    XRAM[9484] = 8'b0;
    XRAM[9485] = 8'b0;
    XRAM[9486] = 8'b0;
    XRAM[9487] = 8'b0;
    XRAM[9488] = 8'b0;
    XRAM[9489] = 8'b0;
    XRAM[9490] = 8'b0;
    XRAM[9491] = 8'b0;
    XRAM[9492] = 8'b0;
    XRAM[9493] = 8'b0;
    XRAM[9494] = 8'b0;
    XRAM[9495] = 8'b0;
    XRAM[9496] = 8'b0;
    XRAM[9497] = 8'b0;
    XRAM[9498] = 8'b0;
    XRAM[9499] = 8'b0;
    XRAM[9500] = 8'b0;
    XRAM[9501] = 8'b0;
    XRAM[9502] = 8'b0;
    XRAM[9503] = 8'b0;
    XRAM[9504] = 8'b0;
    XRAM[9505] = 8'b0;
    XRAM[9506] = 8'b0;
    XRAM[9507] = 8'b0;
    XRAM[9508] = 8'b0;
    XRAM[9509] = 8'b0;
    XRAM[9510] = 8'b0;
    XRAM[9511] = 8'b0;
    XRAM[9512] = 8'b0;
    XRAM[9513] = 8'b0;
    XRAM[9514] = 8'b0;
    XRAM[9515] = 8'b0;
    XRAM[9516] = 8'b0;
    XRAM[9517] = 8'b0;
    XRAM[9518] = 8'b0;
    XRAM[9519] = 8'b0;
    XRAM[9520] = 8'b0;
    XRAM[9521] = 8'b0;
    XRAM[9522] = 8'b0;
    XRAM[9523] = 8'b0;
    XRAM[9524] = 8'b0;
    XRAM[9525] = 8'b0;
    XRAM[9526] = 8'b0;
    XRAM[9527] = 8'b0;
    XRAM[9528] = 8'b0;
    XRAM[9529] = 8'b0;
    XRAM[9530] = 8'b0;
    XRAM[9531] = 8'b0;
    XRAM[9532] = 8'b0;
    XRAM[9533] = 8'b0;
    XRAM[9534] = 8'b0;
    XRAM[9535] = 8'b0;
    XRAM[9536] = 8'b0;
    XRAM[9537] = 8'b0;
    XRAM[9538] = 8'b0;
    XRAM[9539] = 8'b0;
    XRAM[9540] = 8'b0;
    XRAM[9541] = 8'b0;
    XRAM[9542] = 8'b0;
    XRAM[9543] = 8'b0;
    XRAM[9544] = 8'b0;
    XRAM[9545] = 8'b0;
    XRAM[9546] = 8'b0;
    XRAM[9547] = 8'b0;
    XRAM[9548] = 8'b0;
    XRAM[9549] = 8'b0;
    XRAM[9550] = 8'b0;
    XRAM[9551] = 8'b0;
    XRAM[9552] = 8'b0;
    XRAM[9553] = 8'b0;
    XRAM[9554] = 8'b0;
    XRAM[9555] = 8'b0;
    XRAM[9556] = 8'b0;
    XRAM[9557] = 8'b0;
    XRAM[9558] = 8'b0;
    XRAM[9559] = 8'b0;
    XRAM[9560] = 8'b0;
    XRAM[9561] = 8'b0;
    XRAM[9562] = 8'b0;
    XRAM[9563] = 8'b0;
    XRAM[9564] = 8'b0;
    XRAM[9565] = 8'b0;
    XRAM[9566] = 8'b0;
    XRAM[9567] = 8'b0;
    XRAM[9568] = 8'b0;
    XRAM[9569] = 8'b0;
    XRAM[9570] = 8'b0;
    XRAM[9571] = 8'b0;
    XRAM[9572] = 8'b0;
    XRAM[9573] = 8'b0;
    XRAM[9574] = 8'b0;
    XRAM[9575] = 8'b0;
    XRAM[9576] = 8'b0;
    XRAM[9577] = 8'b0;
    XRAM[9578] = 8'b0;
    XRAM[9579] = 8'b0;
    XRAM[9580] = 8'b0;
    XRAM[9581] = 8'b0;
    XRAM[9582] = 8'b0;
    XRAM[9583] = 8'b0;
    XRAM[9584] = 8'b0;
    XRAM[9585] = 8'b0;
    XRAM[9586] = 8'b0;
    XRAM[9587] = 8'b0;
    XRAM[9588] = 8'b0;
    XRAM[9589] = 8'b0;
    XRAM[9590] = 8'b0;
    XRAM[9591] = 8'b0;
    XRAM[9592] = 8'b0;
    XRAM[9593] = 8'b0;
    XRAM[9594] = 8'b0;
    XRAM[9595] = 8'b0;
    XRAM[9596] = 8'b0;
    XRAM[9597] = 8'b0;
    XRAM[9598] = 8'b0;
    XRAM[9599] = 8'b0;
    XRAM[9600] = 8'b0;
    XRAM[9601] = 8'b0;
    XRAM[9602] = 8'b0;
    XRAM[9603] = 8'b0;
    XRAM[9604] = 8'b0;
    XRAM[9605] = 8'b0;
    XRAM[9606] = 8'b0;
    XRAM[9607] = 8'b0;
    XRAM[9608] = 8'b0;
    XRAM[9609] = 8'b0;
    XRAM[9610] = 8'b0;
    XRAM[9611] = 8'b0;
    XRAM[9612] = 8'b0;
    XRAM[9613] = 8'b0;
    XRAM[9614] = 8'b0;
    XRAM[9615] = 8'b0;
    XRAM[9616] = 8'b0;
    XRAM[9617] = 8'b0;
    XRAM[9618] = 8'b0;
    XRAM[9619] = 8'b0;
    XRAM[9620] = 8'b0;
    XRAM[9621] = 8'b0;
    XRAM[9622] = 8'b0;
    XRAM[9623] = 8'b0;
    XRAM[9624] = 8'b0;
    XRAM[9625] = 8'b0;
    XRAM[9626] = 8'b0;
    XRAM[9627] = 8'b0;
    XRAM[9628] = 8'b0;
    XRAM[9629] = 8'b0;
    XRAM[9630] = 8'b0;
    XRAM[9631] = 8'b0;
    XRAM[9632] = 8'b0;
    XRAM[9633] = 8'b0;
    XRAM[9634] = 8'b0;
    XRAM[9635] = 8'b0;
    XRAM[9636] = 8'b0;
    XRAM[9637] = 8'b0;
    XRAM[9638] = 8'b0;
    XRAM[9639] = 8'b0;
    XRAM[9640] = 8'b0;
    XRAM[9641] = 8'b0;
    XRAM[9642] = 8'b0;
    XRAM[9643] = 8'b0;
    XRAM[9644] = 8'b0;
    XRAM[9645] = 8'b0;
    XRAM[9646] = 8'b0;
    XRAM[9647] = 8'b0;
    XRAM[9648] = 8'b0;
    XRAM[9649] = 8'b0;
    XRAM[9650] = 8'b0;
    XRAM[9651] = 8'b0;
    XRAM[9652] = 8'b0;
    XRAM[9653] = 8'b0;
    XRAM[9654] = 8'b0;
    XRAM[9655] = 8'b0;
    XRAM[9656] = 8'b0;
    XRAM[9657] = 8'b0;
    XRAM[9658] = 8'b0;
    XRAM[9659] = 8'b0;
    XRAM[9660] = 8'b0;
    XRAM[9661] = 8'b0;
    XRAM[9662] = 8'b0;
    XRAM[9663] = 8'b0;
    XRAM[9664] = 8'b0;
    XRAM[9665] = 8'b0;
    XRAM[9666] = 8'b0;
    XRAM[9667] = 8'b0;
    XRAM[9668] = 8'b0;
    XRAM[9669] = 8'b0;
    XRAM[9670] = 8'b0;
    XRAM[9671] = 8'b0;
    XRAM[9672] = 8'b0;
    XRAM[9673] = 8'b0;
    XRAM[9674] = 8'b0;
    XRAM[9675] = 8'b0;
    XRAM[9676] = 8'b0;
    XRAM[9677] = 8'b0;
    XRAM[9678] = 8'b0;
    XRAM[9679] = 8'b0;
    XRAM[9680] = 8'b0;
    XRAM[9681] = 8'b0;
    XRAM[9682] = 8'b0;
    XRAM[9683] = 8'b0;
    XRAM[9684] = 8'b0;
    XRAM[9685] = 8'b0;
    XRAM[9686] = 8'b0;
    XRAM[9687] = 8'b0;
    XRAM[9688] = 8'b0;
    XRAM[9689] = 8'b0;
    XRAM[9690] = 8'b0;
    XRAM[9691] = 8'b0;
    XRAM[9692] = 8'b0;
    XRAM[9693] = 8'b0;
    XRAM[9694] = 8'b0;
    XRAM[9695] = 8'b0;
    XRAM[9696] = 8'b0;
    XRAM[9697] = 8'b0;
    XRAM[9698] = 8'b0;
    XRAM[9699] = 8'b0;
    XRAM[9700] = 8'b0;
    XRAM[9701] = 8'b0;
    XRAM[9702] = 8'b0;
    XRAM[9703] = 8'b0;
    XRAM[9704] = 8'b0;
    XRAM[9705] = 8'b0;
    XRAM[9706] = 8'b0;
    XRAM[9707] = 8'b0;
    XRAM[9708] = 8'b0;
    XRAM[9709] = 8'b0;
    XRAM[9710] = 8'b0;
    XRAM[9711] = 8'b0;
    XRAM[9712] = 8'b0;
    XRAM[9713] = 8'b0;
    XRAM[9714] = 8'b0;
    XRAM[9715] = 8'b0;
    XRAM[9716] = 8'b0;
    XRAM[9717] = 8'b0;
    XRAM[9718] = 8'b0;
    XRAM[9719] = 8'b0;
    XRAM[9720] = 8'b0;
    XRAM[9721] = 8'b0;
    XRAM[9722] = 8'b0;
    XRAM[9723] = 8'b0;
    XRAM[9724] = 8'b0;
    XRAM[9725] = 8'b0;
    XRAM[9726] = 8'b0;
    XRAM[9727] = 8'b0;
    XRAM[9728] = 8'b0;
    XRAM[9729] = 8'b0;
    XRAM[9730] = 8'b0;
    XRAM[9731] = 8'b0;
    XRAM[9732] = 8'b0;
    XRAM[9733] = 8'b0;
    XRAM[9734] = 8'b0;
    XRAM[9735] = 8'b0;
    XRAM[9736] = 8'b0;
    XRAM[9737] = 8'b0;
    XRAM[9738] = 8'b0;
    XRAM[9739] = 8'b0;
    XRAM[9740] = 8'b0;
    XRAM[9741] = 8'b0;
    XRAM[9742] = 8'b0;
    XRAM[9743] = 8'b0;
    XRAM[9744] = 8'b0;
    XRAM[9745] = 8'b0;
    XRAM[9746] = 8'b0;
    XRAM[9747] = 8'b0;
    XRAM[9748] = 8'b0;
    XRAM[9749] = 8'b0;
    XRAM[9750] = 8'b0;
    XRAM[9751] = 8'b0;
    XRAM[9752] = 8'b0;
    XRAM[9753] = 8'b0;
    XRAM[9754] = 8'b0;
    XRAM[9755] = 8'b0;
    XRAM[9756] = 8'b0;
    XRAM[9757] = 8'b0;
    XRAM[9758] = 8'b0;
    XRAM[9759] = 8'b0;
    XRAM[9760] = 8'b0;
    XRAM[9761] = 8'b0;
    XRAM[9762] = 8'b0;
    XRAM[9763] = 8'b0;
    XRAM[9764] = 8'b0;
    XRAM[9765] = 8'b0;
    XRAM[9766] = 8'b0;
    XRAM[9767] = 8'b0;
    XRAM[9768] = 8'b0;
    XRAM[9769] = 8'b0;
    XRAM[9770] = 8'b0;
    XRAM[9771] = 8'b0;
    XRAM[9772] = 8'b0;
    XRAM[9773] = 8'b0;
    XRAM[9774] = 8'b0;
    XRAM[9775] = 8'b0;
    XRAM[9776] = 8'b0;
    XRAM[9777] = 8'b0;
    XRAM[9778] = 8'b0;
    XRAM[9779] = 8'b0;
    XRAM[9780] = 8'b0;
    XRAM[9781] = 8'b0;
    XRAM[9782] = 8'b0;
    XRAM[9783] = 8'b0;
    XRAM[9784] = 8'b0;
    XRAM[9785] = 8'b0;
    XRAM[9786] = 8'b0;
    XRAM[9787] = 8'b0;
    XRAM[9788] = 8'b0;
    XRAM[9789] = 8'b0;
    XRAM[9790] = 8'b0;
    XRAM[9791] = 8'b0;
    XRAM[9792] = 8'b0;
    XRAM[9793] = 8'b0;
    XRAM[9794] = 8'b0;
    XRAM[9795] = 8'b0;
    XRAM[9796] = 8'b0;
    XRAM[9797] = 8'b0;
    XRAM[9798] = 8'b0;
    XRAM[9799] = 8'b0;
    XRAM[9800] = 8'b0;
    XRAM[9801] = 8'b0;
    XRAM[9802] = 8'b0;
    XRAM[9803] = 8'b0;
    XRAM[9804] = 8'b0;
    XRAM[9805] = 8'b0;
    XRAM[9806] = 8'b0;
    XRAM[9807] = 8'b0;
    XRAM[9808] = 8'b0;
    XRAM[9809] = 8'b0;
    XRAM[9810] = 8'b0;
    XRAM[9811] = 8'b0;
    XRAM[9812] = 8'b0;
    XRAM[9813] = 8'b0;
    XRAM[9814] = 8'b0;
    XRAM[9815] = 8'b0;
    XRAM[9816] = 8'b0;
    XRAM[9817] = 8'b0;
    XRAM[9818] = 8'b0;
    XRAM[9819] = 8'b0;
    XRAM[9820] = 8'b0;
    XRAM[9821] = 8'b0;
    XRAM[9822] = 8'b0;
    XRAM[9823] = 8'b0;
    XRAM[9824] = 8'b0;
    XRAM[9825] = 8'b0;
    XRAM[9826] = 8'b0;
    XRAM[9827] = 8'b0;
    XRAM[9828] = 8'b0;
    XRAM[9829] = 8'b0;
    XRAM[9830] = 8'b0;
    XRAM[9831] = 8'b0;
    XRAM[9832] = 8'b0;
    XRAM[9833] = 8'b0;
    XRAM[9834] = 8'b0;
    XRAM[9835] = 8'b0;
    XRAM[9836] = 8'b0;
    XRAM[9837] = 8'b0;
    XRAM[9838] = 8'b0;
    XRAM[9839] = 8'b0;
    XRAM[9840] = 8'b0;
    XRAM[9841] = 8'b0;
    XRAM[9842] = 8'b0;
    XRAM[9843] = 8'b0;
    XRAM[9844] = 8'b0;
    XRAM[9845] = 8'b0;
    XRAM[9846] = 8'b0;
    XRAM[9847] = 8'b0;
    XRAM[9848] = 8'b0;
    XRAM[9849] = 8'b0;
    XRAM[9850] = 8'b0;
    XRAM[9851] = 8'b0;
    XRAM[9852] = 8'b0;
    XRAM[9853] = 8'b0;
    XRAM[9854] = 8'b0;
    XRAM[9855] = 8'b0;
    XRAM[9856] = 8'b0;
    XRAM[9857] = 8'b0;
    XRAM[9858] = 8'b0;
    XRAM[9859] = 8'b0;
    XRAM[9860] = 8'b0;
    XRAM[9861] = 8'b0;
    XRAM[9862] = 8'b0;
    XRAM[9863] = 8'b0;
    XRAM[9864] = 8'b0;
    XRAM[9865] = 8'b0;
    XRAM[9866] = 8'b0;
    XRAM[9867] = 8'b0;
    XRAM[9868] = 8'b0;
    XRAM[9869] = 8'b0;
    XRAM[9870] = 8'b0;
    XRAM[9871] = 8'b0;
    XRAM[9872] = 8'b0;
    XRAM[9873] = 8'b0;
    XRAM[9874] = 8'b0;
    XRAM[9875] = 8'b0;
    XRAM[9876] = 8'b0;
    XRAM[9877] = 8'b0;
    XRAM[9878] = 8'b0;
    XRAM[9879] = 8'b0;
    XRAM[9880] = 8'b0;
    XRAM[9881] = 8'b0;
    XRAM[9882] = 8'b0;
    XRAM[9883] = 8'b0;
    XRAM[9884] = 8'b0;
    XRAM[9885] = 8'b0;
    XRAM[9886] = 8'b0;
    XRAM[9887] = 8'b0;
    XRAM[9888] = 8'b0;
    XRAM[9889] = 8'b0;
    XRAM[9890] = 8'b0;
    XRAM[9891] = 8'b0;
    XRAM[9892] = 8'b0;
    XRAM[9893] = 8'b0;
    XRAM[9894] = 8'b0;
    XRAM[9895] = 8'b0;
    XRAM[9896] = 8'b0;
    XRAM[9897] = 8'b0;
    XRAM[9898] = 8'b0;
    XRAM[9899] = 8'b0;
    XRAM[9900] = 8'b0;
    XRAM[9901] = 8'b0;
    XRAM[9902] = 8'b0;
    XRAM[9903] = 8'b0;
    XRAM[9904] = 8'b0;
    XRAM[9905] = 8'b0;
    XRAM[9906] = 8'b0;
    XRAM[9907] = 8'b0;
    XRAM[9908] = 8'b0;
    XRAM[9909] = 8'b0;
    XRAM[9910] = 8'b0;
    XRAM[9911] = 8'b0;
    XRAM[9912] = 8'b0;
    XRAM[9913] = 8'b0;
    XRAM[9914] = 8'b0;
    XRAM[9915] = 8'b0;
    XRAM[9916] = 8'b0;
    XRAM[9917] = 8'b0;
    XRAM[9918] = 8'b0;
    XRAM[9919] = 8'b0;
    XRAM[9920] = 8'b0;
    XRAM[9921] = 8'b0;
    XRAM[9922] = 8'b0;
    XRAM[9923] = 8'b0;
    XRAM[9924] = 8'b0;
    XRAM[9925] = 8'b0;
    XRAM[9926] = 8'b0;
    XRAM[9927] = 8'b0;
    XRAM[9928] = 8'b0;
    XRAM[9929] = 8'b0;
    XRAM[9930] = 8'b0;
    XRAM[9931] = 8'b0;
    XRAM[9932] = 8'b0;
    XRAM[9933] = 8'b0;
    XRAM[9934] = 8'b0;
    XRAM[9935] = 8'b0;
    XRAM[9936] = 8'b0;
    XRAM[9937] = 8'b0;
    XRAM[9938] = 8'b0;
    XRAM[9939] = 8'b0;
    XRAM[9940] = 8'b0;
    XRAM[9941] = 8'b0;
    XRAM[9942] = 8'b0;
    XRAM[9943] = 8'b0;
    XRAM[9944] = 8'b0;
    XRAM[9945] = 8'b0;
    XRAM[9946] = 8'b0;
    XRAM[9947] = 8'b0;
    XRAM[9948] = 8'b0;
    XRAM[9949] = 8'b0;
    XRAM[9950] = 8'b0;
    XRAM[9951] = 8'b0;
    XRAM[9952] = 8'b0;
    XRAM[9953] = 8'b0;
    XRAM[9954] = 8'b0;
    XRAM[9955] = 8'b0;
    XRAM[9956] = 8'b0;
    XRAM[9957] = 8'b0;
    XRAM[9958] = 8'b0;
    XRAM[9959] = 8'b0;
    XRAM[9960] = 8'b0;
    XRAM[9961] = 8'b0;
    XRAM[9962] = 8'b0;
    XRAM[9963] = 8'b0;
    XRAM[9964] = 8'b0;
    XRAM[9965] = 8'b0;
    XRAM[9966] = 8'b0;
    XRAM[9967] = 8'b0;
    XRAM[9968] = 8'b0;
    XRAM[9969] = 8'b0;
    XRAM[9970] = 8'b0;
    XRAM[9971] = 8'b0;
    XRAM[9972] = 8'b0;
    XRAM[9973] = 8'b0;
    XRAM[9974] = 8'b0;
    XRAM[9975] = 8'b0;
    XRAM[9976] = 8'b0;
    XRAM[9977] = 8'b0;
    XRAM[9978] = 8'b0;
    XRAM[9979] = 8'b0;
    XRAM[9980] = 8'b0;
    XRAM[9981] = 8'b0;
    XRAM[9982] = 8'b0;
    XRAM[9983] = 8'b0;
    XRAM[9984] = 8'b0;
    XRAM[9985] = 8'b0;
    XRAM[9986] = 8'b0;
    XRAM[9987] = 8'b0;
    XRAM[9988] = 8'b0;
    XRAM[9989] = 8'b0;
    XRAM[9990] = 8'b0;
    XRAM[9991] = 8'b0;
    XRAM[9992] = 8'b0;
    XRAM[9993] = 8'b0;
    XRAM[9994] = 8'b0;
    XRAM[9995] = 8'b0;
    XRAM[9996] = 8'b0;
    XRAM[9997] = 8'b0;
    XRAM[9998] = 8'b0;
    XRAM[9999] = 8'b0;
    XRAM[10000] = 8'b0;
    XRAM[10001] = 8'b0;
    XRAM[10002] = 8'b0;
    XRAM[10003] = 8'b0;
    XRAM[10004] = 8'b0;
    XRAM[10005] = 8'b0;
    XRAM[10006] = 8'b0;
    XRAM[10007] = 8'b0;
    XRAM[10008] = 8'b0;
    XRAM[10009] = 8'b0;
    XRAM[10010] = 8'b0;
    XRAM[10011] = 8'b0;
    XRAM[10012] = 8'b0;
    XRAM[10013] = 8'b0;
    XRAM[10014] = 8'b0;
    XRAM[10015] = 8'b0;
    XRAM[10016] = 8'b0;
    XRAM[10017] = 8'b0;
    XRAM[10018] = 8'b0;
    XRAM[10019] = 8'b0;
    XRAM[10020] = 8'b0;
    XRAM[10021] = 8'b0;
    XRAM[10022] = 8'b0;
    XRAM[10023] = 8'b0;
    XRAM[10024] = 8'b0;
    XRAM[10025] = 8'b0;
    XRAM[10026] = 8'b0;
    XRAM[10027] = 8'b0;
    XRAM[10028] = 8'b0;
    XRAM[10029] = 8'b0;
    XRAM[10030] = 8'b0;
    XRAM[10031] = 8'b0;
    XRAM[10032] = 8'b0;
    XRAM[10033] = 8'b0;
    XRAM[10034] = 8'b0;
    XRAM[10035] = 8'b0;
    XRAM[10036] = 8'b0;
    XRAM[10037] = 8'b0;
    XRAM[10038] = 8'b0;
    XRAM[10039] = 8'b0;
    XRAM[10040] = 8'b0;
    XRAM[10041] = 8'b0;
    XRAM[10042] = 8'b0;
    XRAM[10043] = 8'b0;
    XRAM[10044] = 8'b0;
    XRAM[10045] = 8'b0;
    XRAM[10046] = 8'b0;
    XRAM[10047] = 8'b0;
    XRAM[10048] = 8'b0;
    XRAM[10049] = 8'b0;
    XRAM[10050] = 8'b0;
    XRAM[10051] = 8'b0;
    XRAM[10052] = 8'b0;
    XRAM[10053] = 8'b0;
    XRAM[10054] = 8'b0;
    XRAM[10055] = 8'b0;
    XRAM[10056] = 8'b0;
    XRAM[10057] = 8'b0;
    XRAM[10058] = 8'b0;
    XRAM[10059] = 8'b0;
    XRAM[10060] = 8'b0;
    XRAM[10061] = 8'b0;
    XRAM[10062] = 8'b0;
    XRAM[10063] = 8'b0;
    XRAM[10064] = 8'b0;
    XRAM[10065] = 8'b0;
    XRAM[10066] = 8'b0;
    XRAM[10067] = 8'b0;
    XRAM[10068] = 8'b0;
    XRAM[10069] = 8'b0;
    XRAM[10070] = 8'b0;
    XRAM[10071] = 8'b0;
    XRAM[10072] = 8'b0;
    XRAM[10073] = 8'b0;
    XRAM[10074] = 8'b0;
    XRAM[10075] = 8'b0;
    XRAM[10076] = 8'b0;
    XRAM[10077] = 8'b0;
    XRAM[10078] = 8'b0;
    XRAM[10079] = 8'b0;
    XRAM[10080] = 8'b0;
    XRAM[10081] = 8'b0;
    XRAM[10082] = 8'b0;
    XRAM[10083] = 8'b0;
    XRAM[10084] = 8'b0;
    XRAM[10085] = 8'b0;
    XRAM[10086] = 8'b0;
    XRAM[10087] = 8'b0;
    XRAM[10088] = 8'b0;
    XRAM[10089] = 8'b0;
    XRAM[10090] = 8'b0;
    XRAM[10091] = 8'b0;
    XRAM[10092] = 8'b0;
    XRAM[10093] = 8'b0;
    XRAM[10094] = 8'b0;
    XRAM[10095] = 8'b0;
    XRAM[10096] = 8'b0;
    XRAM[10097] = 8'b0;
    XRAM[10098] = 8'b0;
    XRAM[10099] = 8'b0;
    XRAM[10100] = 8'b0;
    XRAM[10101] = 8'b0;
    XRAM[10102] = 8'b0;
    XRAM[10103] = 8'b0;
    XRAM[10104] = 8'b0;
    XRAM[10105] = 8'b0;
    XRAM[10106] = 8'b0;
    XRAM[10107] = 8'b0;
    XRAM[10108] = 8'b0;
    XRAM[10109] = 8'b0;
    XRAM[10110] = 8'b0;
    XRAM[10111] = 8'b0;
    XRAM[10112] = 8'b0;
    XRAM[10113] = 8'b0;
    XRAM[10114] = 8'b0;
    XRAM[10115] = 8'b0;
    XRAM[10116] = 8'b0;
    XRAM[10117] = 8'b0;
    XRAM[10118] = 8'b0;
    XRAM[10119] = 8'b0;
    XRAM[10120] = 8'b0;
    XRAM[10121] = 8'b0;
    XRAM[10122] = 8'b0;
    XRAM[10123] = 8'b0;
    XRAM[10124] = 8'b0;
    XRAM[10125] = 8'b0;
    XRAM[10126] = 8'b0;
    XRAM[10127] = 8'b0;
    XRAM[10128] = 8'b0;
    XRAM[10129] = 8'b0;
    XRAM[10130] = 8'b0;
    XRAM[10131] = 8'b0;
    XRAM[10132] = 8'b0;
    XRAM[10133] = 8'b0;
    XRAM[10134] = 8'b0;
    XRAM[10135] = 8'b0;
    XRAM[10136] = 8'b0;
    XRAM[10137] = 8'b0;
    XRAM[10138] = 8'b0;
    XRAM[10139] = 8'b0;
    XRAM[10140] = 8'b0;
    XRAM[10141] = 8'b0;
    XRAM[10142] = 8'b0;
    XRAM[10143] = 8'b0;
    XRAM[10144] = 8'b0;
    XRAM[10145] = 8'b0;
    XRAM[10146] = 8'b0;
    XRAM[10147] = 8'b0;
    XRAM[10148] = 8'b0;
    XRAM[10149] = 8'b0;
    XRAM[10150] = 8'b0;
    XRAM[10151] = 8'b0;
    XRAM[10152] = 8'b0;
    XRAM[10153] = 8'b0;
    XRAM[10154] = 8'b0;
    XRAM[10155] = 8'b0;
    XRAM[10156] = 8'b0;
    XRAM[10157] = 8'b0;
    XRAM[10158] = 8'b0;
    XRAM[10159] = 8'b0;
    XRAM[10160] = 8'b0;
    XRAM[10161] = 8'b0;
    XRAM[10162] = 8'b0;
    XRAM[10163] = 8'b0;
    XRAM[10164] = 8'b0;
    XRAM[10165] = 8'b0;
    XRAM[10166] = 8'b0;
    XRAM[10167] = 8'b0;
    XRAM[10168] = 8'b0;
    XRAM[10169] = 8'b0;
    XRAM[10170] = 8'b0;
    XRAM[10171] = 8'b0;
    XRAM[10172] = 8'b0;
    XRAM[10173] = 8'b0;
    XRAM[10174] = 8'b0;
    XRAM[10175] = 8'b0;
    XRAM[10176] = 8'b0;
    XRAM[10177] = 8'b0;
    XRAM[10178] = 8'b0;
    XRAM[10179] = 8'b0;
    XRAM[10180] = 8'b0;
    XRAM[10181] = 8'b0;
    XRAM[10182] = 8'b0;
    XRAM[10183] = 8'b0;
    XRAM[10184] = 8'b0;
    XRAM[10185] = 8'b0;
    XRAM[10186] = 8'b0;
    XRAM[10187] = 8'b0;
    XRAM[10188] = 8'b0;
    XRAM[10189] = 8'b0;
    XRAM[10190] = 8'b0;
    XRAM[10191] = 8'b0;
    XRAM[10192] = 8'b0;
    XRAM[10193] = 8'b0;
    XRAM[10194] = 8'b0;
    XRAM[10195] = 8'b0;
    XRAM[10196] = 8'b0;
    XRAM[10197] = 8'b0;
    XRAM[10198] = 8'b0;
    XRAM[10199] = 8'b0;
    XRAM[10200] = 8'b0;
    XRAM[10201] = 8'b0;
    XRAM[10202] = 8'b0;
    XRAM[10203] = 8'b0;
    XRAM[10204] = 8'b0;
    XRAM[10205] = 8'b0;
    XRAM[10206] = 8'b0;
    XRAM[10207] = 8'b0;
    XRAM[10208] = 8'b0;
    XRAM[10209] = 8'b0;
    XRAM[10210] = 8'b0;
    XRAM[10211] = 8'b0;
    XRAM[10212] = 8'b0;
    XRAM[10213] = 8'b0;
    XRAM[10214] = 8'b0;
    XRAM[10215] = 8'b0;
    XRAM[10216] = 8'b0;
    XRAM[10217] = 8'b0;
    XRAM[10218] = 8'b0;
    XRAM[10219] = 8'b0;
    XRAM[10220] = 8'b0;
    XRAM[10221] = 8'b0;
    XRAM[10222] = 8'b0;
    XRAM[10223] = 8'b0;
    XRAM[10224] = 8'b0;
    XRAM[10225] = 8'b0;
    XRAM[10226] = 8'b0;
    XRAM[10227] = 8'b0;
    XRAM[10228] = 8'b0;
    XRAM[10229] = 8'b0;
    XRAM[10230] = 8'b0;
    XRAM[10231] = 8'b0;
    XRAM[10232] = 8'b0;
    XRAM[10233] = 8'b0;
    XRAM[10234] = 8'b0;
    XRAM[10235] = 8'b0;
    XRAM[10236] = 8'b0;
    XRAM[10237] = 8'b0;
    XRAM[10238] = 8'b0;
    XRAM[10239] = 8'b0;
    XRAM[10240] = 8'b0;
    XRAM[10241] = 8'b0;
    XRAM[10242] = 8'b0;
    XRAM[10243] = 8'b0;
    XRAM[10244] = 8'b0;
    XRAM[10245] = 8'b0;
    XRAM[10246] = 8'b0;
    XRAM[10247] = 8'b0;
    XRAM[10248] = 8'b0;
    XRAM[10249] = 8'b0;
    XRAM[10250] = 8'b0;
    XRAM[10251] = 8'b0;
    XRAM[10252] = 8'b0;
    XRAM[10253] = 8'b0;
    XRAM[10254] = 8'b0;
    XRAM[10255] = 8'b0;
    XRAM[10256] = 8'b0;
    XRAM[10257] = 8'b0;
    XRAM[10258] = 8'b0;
    XRAM[10259] = 8'b0;
    XRAM[10260] = 8'b0;
    XRAM[10261] = 8'b0;
    XRAM[10262] = 8'b0;
    XRAM[10263] = 8'b0;
    XRAM[10264] = 8'b0;
    XRAM[10265] = 8'b0;
    XRAM[10266] = 8'b0;
    XRAM[10267] = 8'b0;
    XRAM[10268] = 8'b0;
    XRAM[10269] = 8'b0;
    XRAM[10270] = 8'b0;
    XRAM[10271] = 8'b0;
    XRAM[10272] = 8'b0;
    XRAM[10273] = 8'b0;
    XRAM[10274] = 8'b0;
    XRAM[10275] = 8'b0;
    XRAM[10276] = 8'b0;
    XRAM[10277] = 8'b0;
    XRAM[10278] = 8'b0;
    XRAM[10279] = 8'b0;
    XRAM[10280] = 8'b0;
    XRAM[10281] = 8'b0;
    XRAM[10282] = 8'b0;
    XRAM[10283] = 8'b0;
    XRAM[10284] = 8'b0;
    XRAM[10285] = 8'b0;
    XRAM[10286] = 8'b0;
    XRAM[10287] = 8'b0;
    XRAM[10288] = 8'b0;
    XRAM[10289] = 8'b0;
    XRAM[10290] = 8'b0;
    XRAM[10291] = 8'b0;
    XRAM[10292] = 8'b0;
    XRAM[10293] = 8'b0;
    XRAM[10294] = 8'b0;
    XRAM[10295] = 8'b0;
    XRAM[10296] = 8'b0;
    XRAM[10297] = 8'b0;
    XRAM[10298] = 8'b0;
    XRAM[10299] = 8'b0;
    XRAM[10300] = 8'b0;
    XRAM[10301] = 8'b0;
    XRAM[10302] = 8'b0;
    XRAM[10303] = 8'b0;
    XRAM[10304] = 8'b0;
    XRAM[10305] = 8'b0;
    XRAM[10306] = 8'b0;
    XRAM[10307] = 8'b0;
    XRAM[10308] = 8'b0;
    XRAM[10309] = 8'b0;
    XRAM[10310] = 8'b0;
    XRAM[10311] = 8'b0;
    XRAM[10312] = 8'b0;
    XRAM[10313] = 8'b0;
    XRAM[10314] = 8'b0;
    XRAM[10315] = 8'b0;
    XRAM[10316] = 8'b0;
    XRAM[10317] = 8'b0;
    XRAM[10318] = 8'b0;
    XRAM[10319] = 8'b0;
    XRAM[10320] = 8'b0;
    XRAM[10321] = 8'b0;
    XRAM[10322] = 8'b0;
    XRAM[10323] = 8'b0;
    XRAM[10324] = 8'b0;
    XRAM[10325] = 8'b0;
    XRAM[10326] = 8'b0;
    XRAM[10327] = 8'b0;
    XRAM[10328] = 8'b0;
    XRAM[10329] = 8'b0;
    XRAM[10330] = 8'b0;
    XRAM[10331] = 8'b0;
    XRAM[10332] = 8'b0;
    XRAM[10333] = 8'b0;
    XRAM[10334] = 8'b0;
    XRAM[10335] = 8'b0;
    XRAM[10336] = 8'b0;
    XRAM[10337] = 8'b0;
    XRAM[10338] = 8'b0;
    XRAM[10339] = 8'b0;
    XRAM[10340] = 8'b0;
    XRAM[10341] = 8'b0;
    XRAM[10342] = 8'b0;
    XRAM[10343] = 8'b0;
    XRAM[10344] = 8'b0;
    XRAM[10345] = 8'b0;
    XRAM[10346] = 8'b0;
    XRAM[10347] = 8'b0;
    XRAM[10348] = 8'b0;
    XRAM[10349] = 8'b0;
    XRAM[10350] = 8'b0;
    XRAM[10351] = 8'b0;
    XRAM[10352] = 8'b0;
    XRAM[10353] = 8'b0;
    XRAM[10354] = 8'b0;
    XRAM[10355] = 8'b0;
    XRAM[10356] = 8'b0;
    XRAM[10357] = 8'b0;
    XRAM[10358] = 8'b0;
    XRAM[10359] = 8'b0;
    XRAM[10360] = 8'b0;
    XRAM[10361] = 8'b0;
    XRAM[10362] = 8'b0;
    XRAM[10363] = 8'b0;
    XRAM[10364] = 8'b0;
    XRAM[10365] = 8'b0;
    XRAM[10366] = 8'b0;
    XRAM[10367] = 8'b0;
    XRAM[10368] = 8'b0;
    XRAM[10369] = 8'b0;
    XRAM[10370] = 8'b0;
    XRAM[10371] = 8'b0;
    XRAM[10372] = 8'b0;
    XRAM[10373] = 8'b0;
    XRAM[10374] = 8'b0;
    XRAM[10375] = 8'b0;
    XRAM[10376] = 8'b0;
    XRAM[10377] = 8'b0;
    XRAM[10378] = 8'b0;
    XRAM[10379] = 8'b0;
    XRAM[10380] = 8'b0;
    XRAM[10381] = 8'b0;
    XRAM[10382] = 8'b0;
    XRAM[10383] = 8'b0;
    XRAM[10384] = 8'b0;
    XRAM[10385] = 8'b0;
    XRAM[10386] = 8'b0;
    XRAM[10387] = 8'b0;
    XRAM[10388] = 8'b0;
    XRAM[10389] = 8'b0;
    XRAM[10390] = 8'b0;
    XRAM[10391] = 8'b0;
    XRAM[10392] = 8'b0;
    XRAM[10393] = 8'b0;
    XRAM[10394] = 8'b0;
    XRAM[10395] = 8'b0;
    XRAM[10396] = 8'b0;
    XRAM[10397] = 8'b0;
    XRAM[10398] = 8'b0;
    XRAM[10399] = 8'b0;
    XRAM[10400] = 8'b0;
    XRAM[10401] = 8'b0;
    XRAM[10402] = 8'b0;
    XRAM[10403] = 8'b0;
    XRAM[10404] = 8'b0;
    XRAM[10405] = 8'b0;
    XRAM[10406] = 8'b0;
    XRAM[10407] = 8'b0;
    XRAM[10408] = 8'b0;
    XRAM[10409] = 8'b0;
    XRAM[10410] = 8'b0;
    XRAM[10411] = 8'b0;
    XRAM[10412] = 8'b0;
    XRAM[10413] = 8'b0;
    XRAM[10414] = 8'b0;
    XRAM[10415] = 8'b0;
    XRAM[10416] = 8'b0;
    XRAM[10417] = 8'b0;
    XRAM[10418] = 8'b0;
    XRAM[10419] = 8'b0;
    XRAM[10420] = 8'b0;
    XRAM[10421] = 8'b0;
    XRAM[10422] = 8'b0;
    XRAM[10423] = 8'b0;
    XRAM[10424] = 8'b0;
    XRAM[10425] = 8'b0;
    XRAM[10426] = 8'b0;
    XRAM[10427] = 8'b0;
    XRAM[10428] = 8'b0;
    XRAM[10429] = 8'b0;
    XRAM[10430] = 8'b0;
    XRAM[10431] = 8'b0;
    XRAM[10432] = 8'b0;
    XRAM[10433] = 8'b0;
    XRAM[10434] = 8'b0;
    XRAM[10435] = 8'b0;
    XRAM[10436] = 8'b0;
    XRAM[10437] = 8'b0;
    XRAM[10438] = 8'b0;
    XRAM[10439] = 8'b0;
    XRAM[10440] = 8'b0;
    XRAM[10441] = 8'b0;
    XRAM[10442] = 8'b0;
    XRAM[10443] = 8'b0;
    XRAM[10444] = 8'b0;
    XRAM[10445] = 8'b0;
    XRAM[10446] = 8'b0;
    XRAM[10447] = 8'b0;
    XRAM[10448] = 8'b0;
    XRAM[10449] = 8'b0;
    XRAM[10450] = 8'b0;
    XRAM[10451] = 8'b0;
    XRAM[10452] = 8'b0;
    XRAM[10453] = 8'b0;
    XRAM[10454] = 8'b0;
    XRAM[10455] = 8'b0;
    XRAM[10456] = 8'b0;
    XRAM[10457] = 8'b0;
    XRAM[10458] = 8'b0;
    XRAM[10459] = 8'b0;
    XRAM[10460] = 8'b0;
    XRAM[10461] = 8'b0;
    XRAM[10462] = 8'b0;
    XRAM[10463] = 8'b0;
    XRAM[10464] = 8'b0;
    XRAM[10465] = 8'b0;
    XRAM[10466] = 8'b0;
    XRAM[10467] = 8'b0;
    XRAM[10468] = 8'b0;
    XRAM[10469] = 8'b0;
    XRAM[10470] = 8'b0;
    XRAM[10471] = 8'b0;
    XRAM[10472] = 8'b0;
    XRAM[10473] = 8'b0;
    XRAM[10474] = 8'b0;
    XRAM[10475] = 8'b0;
    XRAM[10476] = 8'b0;
    XRAM[10477] = 8'b0;
    XRAM[10478] = 8'b0;
    XRAM[10479] = 8'b0;
    XRAM[10480] = 8'b0;
    XRAM[10481] = 8'b0;
    XRAM[10482] = 8'b0;
    XRAM[10483] = 8'b0;
    XRAM[10484] = 8'b0;
    XRAM[10485] = 8'b0;
    XRAM[10486] = 8'b0;
    XRAM[10487] = 8'b0;
    XRAM[10488] = 8'b0;
    XRAM[10489] = 8'b0;
    XRAM[10490] = 8'b0;
    XRAM[10491] = 8'b0;
    XRAM[10492] = 8'b0;
    XRAM[10493] = 8'b0;
    XRAM[10494] = 8'b0;
    XRAM[10495] = 8'b0;
    XRAM[10496] = 8'b0;
    XRAM[10497] = 8'b0;
    XRAM[10498] = 8'b0;
    XRAM[10499] = 8'b0;
    XRAM[10500] = 8'b0;
    XRAM[10501] = 8'b0;
    XRAM[10502] = 8'b0;
    XRAM[10503] = 8'b0;
    XRAM[10504] = 8'b0;
    XRAM[10505] = 8'b0;
    XRAM[10506] = 8'b0;
    XRAM[10507] = 8'b0;
    XRAM[10508] = 8'b0;
    XRAM[10509] = 8'b0;
    XRAM[10510] = 8'b0;
    XRAM[10511] = 8'b0;
    XRAM[10512] = 8'b0;
    XRAM[10513] = 8'b0;
    XRAM[10514] = 8'b0;
    XRAM[10515] = 8'b0;
    XRAM[10516] = 8'b0;
    XRAM[10517] = 8'b0;
    XRAM[10518] = 8'b0;
    XRAM[10519] = 8'b0;
    XRAM[10520] = 8'b0;
    XRAM[10521] = 8'b0;
    XRAM[10522] = 8'b0;
    XRAM[10523] = 8'b0;
    XRAM[10524] = 8'b0;
    XRAM[10525] = 8'b0;
    XRAM[10526] = 8'b0;
    XRAM[10527] = 8'b0;
    XRAM[10528] = 8'b0;
    XRAM[10529] = 8'b0;
    XRAM[10530] = 8'b0;
    XRAM[10531] = 8'b0;
    XRAM[10532] = 8'b0;
    XRAM[10533] = 8'b0;
    XRAM[10534] = 8'b0;
    XRAM[10535] = 8'b0;
    XRAM[10536] = 8'b0;
    XRAM[10537] = 8'b0;
    XRAM[10538] = 8'b0;
    XRAM[10539] = 8'b0;
    XRAM[10540] = 8'b0;
    XRAM[10541] = 8'b0;
    XRAM[10542] = 8'b0;
    XRAM[10543] = 8'b0;
    XRAM[10544] = 8'b0;
    XRAM[10545] = 8'b0;
    XRAM[10546] = 8'b0;
    XRAM[10547] = 8'b0;
    XRAM[10548] = 8'b0;
    XRAM[10549] = 8'b0;
    XRAM[10550] = 8'b0;
    XRAM[10551] = 8'b0;
    XRAM[10552] = 8'b0;
    XRAM[10553] = 8'b0;
    XRAM[10554] = 8'b0;
    XRAM[10555] = 8'b0;
    XRAM[10556] = 8'b0;
    XRAM[10557] = 8'b0;
    XRAM[10558] = 8'b0;
    XRAM[10559] = 8'b0;
    XRAM[10560] = 8'b0;
    XRAM[10561] = 8'b0;
    XRAM[10562] = 8'b0;
    XRAM[10563] = 8'b0;
    XRAM[10564] = 8'b0;
    XRAM[10565] = 8'b0;
    XRAM[10566] = 8'b0;
    XRAM[10567] = 8'b0;
    XRAM[10568] = 8'b0;
    XRAM[10569] = 8'b0;
    XRAM[10570] = 8'b0;
    XRAM[10571] = 8'b0;
    XRAM[10572] = 8'b0;
    XRAM[10573] = 8'b0;
    XRAM[10574] = 8'b0;
    XRAM[10575] = 8'b0;
    XRAM[10576] = 8'b0;
    XRAM[10577] = 8'b0;
    XRAM[10578] = 8'b0;
    XRAM[10579] = 8'b0;
    XRAM[10580] = 8'b0;
    XRAM[10581] = 8'b0;
    XRAM[10582] = 8'b0;
    XRAM[10583] = 8'b0;
    XRAM[10584] = 8'b0;
    XRAM[10585] = 8'b0;
    XRAM[10586] = 8'b0;
    XRAM[10587] = 8'b0;
    XRAM[10588] = 8'b0;
    XRAM[10589] = 8'b0;
    XRAM[10590] = 8'b0;
    XRAM[10591] = 8'b0;
    XRAM[10592] = 8'b0;
    XRAM[10593] = 8'b0;
    XRAM[10594] = 8'b0;
    XRAM[10595] = 8'b0;
    XRAM[10596] = 8'b0;
    XRAM[10597] = 8'b0;
    XRAM[10598] = 8'b0;
    XRAM[10599] = 8'b0;
    XRAM[10600] = 8'b0;
    XRAM[10601] = 8'b0;
    XRAM[10602] = 8'b0;
    XRAM[10603] = 8'b0;
    XRAM[10604] = 8'b0;
    XRAM[10605] = 8'b0;
    XRAM[10606] = 8'b0;
    XRAM[10607] = 8'b0;
    XRAM[10608] = 8'b0;
    XRAM[10609] = 8'b0;
    XRAM[10610] = 8'b0;
    XRAM[10611] = 8'b0;
    XRAM[10612] = 8'b0;
    XRAM[10613] = 8'b0;
    XRAM[10614] = 8'b0;
    XRAM[10615] = 8'b0;
    XRAM[10616] = 8'b0;
    XRAM[10617] = 8'b0;
    XRAM[10618] = 8'b0;
    XRAM[10619] = 8'b0;
    XRAM[10620] = 8'b0;
    XRAM[10621] = 8'b0;
    XRAM[10622] = 8'b0;
    XRAM[10623] = 8'b0;
    XRAM[10624] = 8'b0;
    XRAM[10625] = 8'b0;
    XRAM[10626] = 8'b0;
    XRAM[10627] = 8'b0;
    XRAM[10628] = 8'b0;
    XRAM[10629] = 8'b0;
    XRAM[10630] = 8'b0;
    XRAM[10631] = 8'b0;
    XRAM[10632] = 8'b0;
    XRAM[10633] = 8'b0;
    XRAM[10634] = 8'b0;
    XRAM[10635] = 8'b0;
    XRAM[10636] = 8'b0;
    XRAM[10637] = 8'b0;
    XRAM[10638] = 8'b0;
    XRAM[10639] = 8'b0;
    XRAM[10640] = 8'b0;
    XRAM[10641] = 8'b0;
    XRAM[10642] = 8'b0;
    XRAM[10643] = 8'b0;
    XRAM[10644] = 8'b0;
    XRAM[10645] = 8'b0;
    XRAM[10646] = 8'b0;
    XRAM[10647] = 8'b0;
    XRAM[10648] = 8'b0;
    XRAM[10649] = 8'b0;
    XRAM[10650] = 8'b0;
    XRAM[10651] = 8'b0;
    XRAM[10652] = 8'b0;
    XRAM[10653] = 8'b0;
    XRAM[10654] = 8'b0;
    XRAM[10655] = 8'b0;
    XRAM[10656] = 8'b0;
    XRAM[10657] = 8'b0;
    XRAM[10658] = 8'b0;
    XRAM[10659] = 8'b0;
    XRAM[10660] = 8'b0;
    XRAM[10661] = 8'b0;
    XRAM[10662] = 8'b0;
    XRAM[10663] = 8'b0;
    XRAM[10664] = 8'b0;
    XRAM[10665] = 8'b0;
    XRAM[10666] = 8'b0;
    XRAM[10667] = 8'b0;
    XRAM[10668] = 8'b0;
    XRAM[10669] = 8'b0;
    XRAM[10670] = 8'b0;
    XRAM[10671] = 8'b0;
    XRAM[10672] = 8'b0;
    XRAM[10673] = 8'b0;
    XRAM[10674] = 8'b0;
    XRAM[10675] = 8'b0;
    XRAM[10676] = 8'b0;
    XRAM[10677] = 8'b0;
    XRAM[10678] = 8'b0;
    XRAM[10679] = 8'b0;
    XRAM[10680] = 8'b0;
    XRAM[10681] = 8'b0;
    XRAM[10682] = 8'b0;
    XRAM[10683] = 8'b0;
    XRAM[10684] = 8'b0;
    XRAM[10685] = 8'b0;
    XRAM[10686] = 8'b0;
    XRAM[10687] = 8'b0;
    XRAM[10688] = 8'b0;
    XRAM[10689] = 8'b0;
    XRAM[10690] = 8'b0;
    XRAM[10691] = 8'b0;
    XRAM[10692] = 8'b0;
    XRAM[10693] = 8'b0;
    XRAM[10694] = 8'b0;
    XRAM[10695] = 8'b0;
    XRAM[10696] = 8'b0;
    XRAM[10697] = 8'b0;
    XRAM[10698] = 8'b0;
    XRAM[10699] = 8'b0;
    XRAM[10700] = 8'b0;
    XRAM[10701] = 8'b0;
    XRAM[10702] = 8'b0;
    XRAM[10703] = 8'b0;
    XRAM[10704] = 8'b0;
    XRAM[10705] = 8'b0;
    XRAM[10706] = 8'b0;
    XRAM[10707] = 8'b0;
    XRAM[10708] = 8'b0;
    XRAM[10709] = 8'b0;
    XRAM[10710] = 8'b0;
    XRAM[10711] = 8'b0;
    XRAM[10712] = 8'b0;
    XRAM[10713] = 8'b0;
    XRAM[10714] = 8'b0;
    XRAM[10715] = 8'b0;
    XRAM[10716] = 8'b0;
    XRAM[10717] = 8'b0;
    XRAM[10718] = 8'b0;
    XRAM[10719] = 8'b0;
    XRAM[10720] = 8'b0;
    XRAM[10721] = 8'b0;
    XRAM[10722] = 8'b0;
    XRAM[10723] = 8'b0;
    XRAM[10724] = 8'b0;
    XRAM[10725] = 8'b0;
    XRAM[10726] = 8'b0;
    XRAM[10727] = 8'b0;
    XRAM[10728] = 8'b0;
    XRAM[10729] = 8'b0;
    XRAM[10730] = 8'b0;
    XRAM[10731] = 8'b0;
    XRAM[10732] = 8'b0;
    XRAM[10733] = 8'b0;
    XRAM[10734] = 8'b0;
    XRAM[10735] = 8'b0;
    XRAM[10736] = 8'b0;
    XRAM[10737] = 8'b0;
    XRAM[10738] = 8'b0;
    XRAM[10739] = 8'b0;
    XRAM[10740] = 8'b0;
    XRAM[10741] = 8'b0;
    XRAM[10742] = 8'b0;
    XRAM[10743] = 8'b0;
    XRAM[10744] = 8'b0;
    XRAM[10745] = 8'b0;
    XRAM[10746] = 8'b0;
    XRAM[10747] = 8'b0;
    XRAM[10748] = 8'b0;
    XRAM[10749] = 8'b0;
    XRAM[10750] = 8'b0;
    XRAM[10751] = 8'b0;
    XRAM[10752] = 8'b0;
    XRAM[10753] = 8'b0;
    XRAM[10754] = 8'b0;
    XRAM[10755] = 8'b0;
    XRAM[10756] = 8'b0;
    XRAM[10757] = 8'b0;
    XRAM[10758] = 8'b0;
    XRAM[10759] = 8'b0;
    XRAM[10760] = 8'b0;
    XRAM[10761] = 8'b0;
    XRAM[10762] = 8'b0;
    XRAM[10763] = 8'b0;
    XRAM[10764] = 8'b0;
    XRAM[10765] = 8'b0;
    XRAM[10766] = 8'b0;
    XRAM[10767] = 8'b0;
    XRAM[10768] = 8'b0;
    XRAM[10769] = 8'b0;
    XRAM[10770] = 8'b0;
    XRAM[10771] = 8'b0;
    XRAM[10772] = 8'b0;
    XRAM[10773] = 8'b0;
    XRAM[10774] = 8'b0;
    XRAM[10775] = 8'b0;
    XRAM[10776] = 8'b0;
    XRAM[10777] = 8'b0;
    XRAM[10778] = 8'b0;
    XRAM[10779] = 8'b0;
    XRAM[10780] = 8'b0;
    XRAM[10781] = 8'b0;
    XRAM[10782] = 8'b0;
    XRAM[10783] = 8'b0;
    XRAM[10784] = 8'b0;
    XRAM[10785] = 8'b0;
    XRAM[10786] = 8'b0;
    XRAM[10787] = 8'b0;
    XRAM[10788] = 8'b0;
    XRAM[10789] = 8'b0;
    XRAM[10790] = 8'b0;
    XRAM[10791] = 8'b0;
    XRAM[10792] = 8'b0;
    XRAM[10793] = 8'b0;
    XRAM[10794] = 8'b0;
    XRAM[10795] = 8'b0;
    XRAM[10796] = 8'b0;
    XRAM[10797] = 8'b0;
    XRAM[10798] = 8'b0;
    XRAM[10799] = 8'b0;
    XRAM[10800] = 8'b0;
    XRAM[10801] = 8'b0;
    XRAM[10802] = 8'b0;
    XRAM[10803] = 8'b0;
    XRAM[10804] = 8'b0;
    XRAM[10805] = 8'b0;
    XRAM[10806] = 8'b0;
    XRAM[10807] = 8'b0;
    XRAM[10808] = 8'b0;
    XRAM[10809] = 8'b0;
    XRAM[10810] = 8'b0;
    XRAM[10811] = 8'b0;
    XRAM[10812] = 8'b0;
    XRAM[10813] = 8'b0;
    XRAM[10814] = 8'b0;
    XRAM[10815] = 8'b0;
    XRAM[10816] = 8'b0;
    XRAM[10817] = 8'b0;
    XRAM[10818] = 8'b0;
    XRAM[10819] = 8'b0;
    XRAM[10820] = 8'b0;
    XRAM[10821] = 8'b0;
    XRAM[10822] = 8'b0;
    XRAM[10823] = 8'b0;
    XRAM[10824] = 8'b0;
    XRAM[10825] = 8'b0;
    XRAM[10826] = 8'b0;
    XRAM[10827] = 8'b0;
    XRAM[10828] = 8'b0;
    XRAM[10829] = 8'b0;
    XRAM[10830] = 8'b0;
    XRAM[10831] = 8'b0;
    XRAM[10832] = 8'b0;
    XRAM[10833] = 8'b0;
    XRAM[10834] = 8'b0;
    XRAM[10835] = 8'b0;
    XRAM[10836] = 8'b0;
    XRAM[10837] = 8'b0;
    XRAM[10838] = 8'b0;
    XRAM[10839] = 8'b0;
    XRAM[10840] = 8'b0;
    XRAM[10841] = 8'b0;
    XRAM[10842] = 8'b0;
    XRAM[10843] = 8'b0;
    XRAM[10844] = 8'b0;
    XRAM[10845] = 8'b0;
    XRAM[10846] = 8'b0;
    XRAM[10847] = 8'b0;
    XRAM[10848] = 8'b0;
    XRAM[10849] = 8'b0;
    XRAM[10850] = 8'b0;
    XRAM[10851] = 8'b0;
    XRAM[10852] = 8'b0;
    XRAM[10853] = 8'b0;
    XRAM[10854] = 8'b0;
    XRAM[10855] = 8'b0;
    XRAM[10856] = 8'b0;
    XRAM[10857] = 8'b0;
    XRAM[10858] = 8'b0;
    XRAM[10859] = 8'b0;
    XRAM[10860] = 8'b0;
    XRAM[10861] = 8'b0;
    XRAM[10862] = 8'b0;
    XRAM[10863] = 8'b0;
    XRAM[10864] = 8'b0;
    XRAM[10865] = 8'b0;
    XRAM[10866] = 8'b0;
    XRAM[10867] = 8'b0;
    XRAM[10868] = 8'b0;
    XRAM[10869] = 8'b0;
    XRAM[10870] = 8'b0;
    XRAM[10871] = 8'b0;
    XRAM[10872] = 8'b0;
    XRAM[10873] = 8'b0;
    XRAM[10874] = 8'b0;
    XRAM[10875] = 8'b0;
    XRAM[10876] = 8'b0;
    XRAM[10877] = 8'b0;
    XRAM[10878] = 8'b0;
    XRAM[10879] = 8'b0;
    XRAM[10880] = 8'b0;
    XRAM[10881] = 8'b0;
    XRAM[10882] = 8'b0;
    XRAM[10883] = 8'b0;
    XRAM[10884] = 8'b0;
    XRAM[10885] = 8'b0;
    XRAM[10886] = 8'b0;
    XRAM[10887] = 8'b0;
    XRAM[10888] = 8'b0;
    XRAM[10889] = 8'b0;
    XRAM[10890] = 8'b0;
    XRAM[10891] = 8'b0;
    XRAM[10892] = 8'b0;
    XRAM[10893] = 8'b0;
    XRAM[10894] = 8'b0;
    XRAM[10895] = 8'b0;
    XRAM[10896] = 8'b0;
    XRAM[10897] = 8'b0;
    XRAM[10898] = 8'b0;
    XRAM[10899] = 8'b0;
    XRAM[10900] = 8'b0;
    XRAM[10901] = 8'b0;
    XRAM[10902] = 8'b0;
    XRAM[10903] = 8'b0;
    XRAM[10904] = 8'b0;
    XRAM[10905] = 8'b0;
    XRAM[10906] = 8'b0;
    XRAM[10907] = 8'b0;
    XRAM[10908] = 8'b0;
    XRAM[10909] = 8'b0;
    XRAM[10910] = 8'b0;
    XRAM[10911] = 8'b0;
    XRAM[10912] = 8'b0;
    XRAM[10913] = 8'b0;
    XRAM[10914] = 8'b0;
    XRAM[10915] = 8'b0;
    XRAM[10916] = 8'b0;
    XRAM[10917] = 8'b0;
    XRAM[10918] = 8'b0;
    XRAM[10919] = 8'b0;
    XRAM[10920] = 8'b0;
    XRAM[10921] = 8'b0;
    XRAM[10922] = 8'b0;
    XRAM[10923] = 8'b0;
    XRAM[10924] = 8'b0;
    XRAM[10925] = 8'b0;
    XRAM[10926] = 8'b0;
    XRAM[10927] = 8'b0;
    XRAM[10928] = 8'b0;
    XRAM[10929] = 8'b0;
    XRAM[10930] = 8'b0;
    XRAM[10931] = 8'b0;
    XRAM[10932] = 8'b0;
    XRAM[10933] = 8'b0;
    XRAM[10934] = 8'b0;
    XRAM[10935] = 8'b0;
    XRAM[10936] = 8'b0;
    XRAM[10937] = 8'b0;
    XRAM[10938] = 8'b0;
    XRAM[10939] = 8'b0;
    XRAM[10940] = 8'b0;
    XRAM[10941] = 8'b0;
    XRAM[10942] = 8'b0;
    XRAM[10943] = 8'b0;
    XRAM[10944] = 8'b0;
    XRAM[10945] = 8'b0;
    XRAM[10946] = 8'b0;
    XRAM[10947] = 8'b0;
    XRAM[10948] = 8'b0;
    XRAM[10949] = 8'b0;
    XRAM[10950] = 8'b0;
    XRAM[10951] = 8'b0;
    XRAM[10952] = 8'b0;
    XRAM[10953] = 8'b0;
    XRAM[10954] = 8'b0;
    XRAM[10955] = 8'b0;
    XRAM[10956] = 8'b0;
    XRAM[10957] = 8'b0;
    XRAM[10958] = 8'b0;
    XRAM[10959] = 8'b0;
    XRAM[10960] = 8'b0;
    XRAM[10961] = 8'b0;
    XRAM[10962] = 8'b0;
    XRAM[10963] = 8'b0;
    XRAM[10964] = 8'b0;
    XRAM[10965] = 8'b0;
    XRAM[10966] = 8'b0;
    XRAM[10967] = 8'b0;
    XRAM[10968] = 8'b0;
    XRAM[10969] = 8'b0;
    XRAM[10970] = 8'b0;
    XRAM[10971] = 8'b0;
    XRAM[10972] = 8'b0;
    XRAM[10973] = 8'b0;
    XRAM[10974] = 8'b0;
    XRAM[10975] = 8'b0;
    XRAM[10976] = 8'b0;
    XRAM[10977] = 8'b0;
    XRAM[10978] = 8'b0;
    XRAM[10979] = 8'b0;
    XRAM[10980] = 8'b0;
    XRAM[10981] = 8'b0;
    XRAM[10982] = 8'b0;
    XRAM[10983] = 8'b0;
    XRAM[10984] = 8'b0;
    XRAM[10985] = 8'b0;
    XRAM[10986] = 8'b0;
    XRAM[10987] = 8'b0;
    XRAM[10988] = 8'b0;
    XRAM[10989] = 8'b0;
    XRAM[10990] = 8'b0;
    XRAM[10991] = 8'b0;
    XRAM[10992] = 8'b0;
    XRAM[10993] = 8'b0;
    XRAM[10994] = 8'b0;
    XRAM[10995] = 8'b0;
    XRAM[10996] = 8'b0;
    XRAM[10997] = 8'b0;
    XRAM[10998] = 8'b0;
    XRAM[10999] = 8'b0;
    XRAM[11000] = 8'b0;
    XRAM[11001] = 8'b0;
    XRAM[11002] = 8'b0;
    XRAM[11003] = 8'b0;
    XRAM[11004] = 8'b0;
    XRAM[11005] = 8'b0;
    XRAM[11006] = 8'b0;
    XRAM[11007] = 8'b0;
    XRAM[11008] = 8'b0;
    XRAM[11009] = 8'b0;
    XRAM[11010] = 8'b0;
    XRAM[11011] = 8'b0;
    XRAM[11012] = 8'b0;
    XRAM[11013] = 8'b0;
    XRAM[11014] = 8'b0;
    XRAM[11015] = 8'b0;
    XRAM[11016] = 8'b0;
    XRAM[11017] = 8'b0;
    XRAM[11018] = 8'b0;
    XRAM[11019] = 8'b0;
    XRAM[11020] = 8'b0;
    XRAM[11021] = 8'b0;
    XRAM[11022] = 8'b0;
    XRAM[11023] = 8'b0;
    XRAM[11024] = 8'b0;
    XRAM[11025] = 8'b0;
    XRAM[11026] = 8'b0;
    XRAM[11027] = 8'b0;
    XRAM[11028] = 8'b0;
    XRAM[11029] = 8'b0;
    XRAM[11030] = 8'b0;
    XRAM[11031] = 8'b0;
    XRAM[11032] = 8'b0;
    XRAM[11033] = 8'b0;
    XRAM[11034] = 8'b0;
    XRAM[11035] = 8'b0;
    XRAM[11036] = 8'b0;
    XRAM[11037] = 8'b0;
    XRAM[11038] = 8'b0;
    XRAM[11039] = 8'b0;
    XRAM[11040] = 8'b0;
    XRAM[11041] = 8'b0;
    XRAM[11042] = 8'b0;
    XRAM[11043] = 8'b0;
    XRAM[11044] = 8'b0;
    XRAM[11045] = 8'b0;
    XRAM[11046] = 8'b0;
    XRAM[11047] = 8'b0;
    XRAM[11048] = 8'b0;
    XRAM[11049] = 8'b0;
    XRAM[11050] = 8'b0;
    XRAM[11051] = 8'b0;
    XRAM[11052] = 8'b0;
    XRAM[11053] = 8'b0;
    XRAM[11054] = 8'b0;
    XRAM[11055] = 8'b0;
    XRAM[11056] = 8'b0;
    XRAM[11057] = 8'b0;
    XRAM[11058] = 8'b0;
    XRAM[11059] = 8'b0;
    XRAM[11060] = 8'b0;
    XRAM[11061] = 8'b0;
    XRAM[11062] = 8'b0;
    XRAM[11063] = 8'b0;
    XRAM[11064] = 8'b0;
    XRAM[11065] = 8'b0;
    XRAM[11066] = 8'b0;
    XRAM[11067] = 8'b0;
    XRAM[11068] = 8'b0;
    XRAM[11069] = 8'b0;
    XRAM[11070] = 8'b0;
    XRAM[11071] = 8'b0;
    XRAM[11072] = 8'b0;
    XRAM[11073] = 8'b0;
    XRAM[11074] = 8'b0;
    XRAM[11075] = 8'b0;
    XRAM[11076] = 8'b0;
    XRAM[11077] = 8'b0;
    XRAM[11078] = 8'b0;
    XRAM[11079] = 8'b0;
    XRAM[11080] = 8'b0;
    XRAM[11081] = 8'b0;
    XRAM[11082] = 8'b0;
    XRAM[11083] = 8'b0;
    XRAM[11084] = 8'b0;
    XRAM[11085] = 8'b0;
    XRAM[11086] = 8'b0;
    XRAM[11087] = 8'b0;
    XRAM[11088] = 8'b0;
    XRAM[11089] = 8'b0;
    XRAM[11090] = 8'b0;
    XRAM[11091] = 8'b0;
    XRAM[11092] = 8'b0;
    XRAM[11093] = 8'b0;
    XRAM[11094] = 8'b0;
    XRAM[11095] = 8'b0;
    XRAM[11096] = 8'b0;
    XRAM[11097] = 8'b0;
    XRAM[11098] = 8'b0;
    XRAM[11099] = 8'b0;
    XRAM[11100] = 8'b0;
    XRAM[11101] = 8'b0;
    XRAM[11102] = 8'b0;
    XRAM[11103] = 8'b0;
    XRAM[11104] = 8'b0;
    XRAM[11105] = 8'b0;
    XRAM[11106] = 8'b0;
    XRAM[11107] = 8'b0;
    XRAM[11108] = 8'b0;
    XRAM[11109] = 8'b0;
    XRAM[11110] = 8'b0;
    XRAM[11111] = 8'b0;
    XRAM[11112] = 8'b0;
    XRAM[11113] = 8'b0;
    XRAM[11114] = 8'b0;
    XRAM[11115] = 8'b0;
    XRAM[11116] = 8'b0;
    XRAM[11117] = 8'b0;
    XRAM[11118] = 8'b0;
    XRAM[11119] = 8'b0;
    XRAM[11120] = 8'b0;
    XRAM[11121] = 8'b0;
    XRAM[11122] = 8'b0;
    XRAM[11123] = 8'b0;
    XRAM[11124] = 8'b0;
    XRAM[11125] = 8'b0;
    XRAM[11126] = 8'b0;
    XRAM[11127] = 8'b0;
    XRAM[11128] = 8'b0;
    XRAM[11129] = 8'b0;
    XRAM[11130] = 8'b0;
    XRAM[11131] = 8'b0;
    XRAM[11132] = 8'b0;
    XRAM[11133] = 8'b0;
    XRAM[11134] = 8'b0;
    XRAM[11135] = 8'b0;
    XRAM[11136] = 8'b0;
    XRAM[11137] = 8'b0;
    XRAM[11138] = 8'b0;
    XRAM[11139] = 8'b0;
    XRAM[11140] = 8'b0;
    XRAM[11141] = 8'b0;
    XRAM[11142] = 8'b0;
    XRAM[11143] = 8'b0;
    XRAM[11144] = 8'b0;
    XRAM[11145] = 8'b0;
    XRAM[11146] = 8'b0;
    XRAM[11147] = 8'b0;
    XRAM[11148] = 8'b0;
    XRAM[11149] = 8'b0;
    XRAM[11150] = 8'b0;
    XRAM[11151] = 8'b0;
    XRAM[11152] = 8'b0;
    XRAM[11153] = 8'b0;
    XRAM[11154] = 8'b0;
    XRAM[11155] = 8'b0;
    XRAM[11156] = 8'b0;
    XRAM[11157] = 8'b0;
    XRAM[11158] = 8'b0;
    XRAM[11159] = 8'b0;
    XRAM[11160] = 8'b0;
    XRAM[11161] = 8'b0;
    XRAM[11162] = 8'b0;
    XRAM[11163] = 8'b0;
    XRAM[11164] = 8'b0;
    XRAM[11165] = 8'b0;
    XRAM[11166] = 8'b0;
    XRAM[11167] = 8'b0;
    XRAM[11168] = 8'b0;
    XRAM[11169] = 8'b0;
    XRAM[11170] = 8'b0;
    XRAM[11171] = 8'b0;
    XRAM[11172] = 8'b0;
    XRAM[11173] = 8'b0;
    XRAM[11174] = 8'b0;
    XRAM[11175] = 8'b0;
    XRAM[11176] = 8'b0;
    XRAM[11177] = 8'b0;
    XRAM[11178] = 8'b0;
    XRAM[11179] = 8'b0;
    XRAM[11180] = 8'b0;
    XRAM[11181] = 8'b0;
    XRAM[11182] = 8'b0;
    XRAM[11183] = 8'b0;
    XRAM[11184] = 8'b0;
    XRAM[11185] = 8'b0;
    XRAM[11186] = 8'b0;
    XRAM[11187] = 8'b0;
    XRAM[11188] = 8'b0;
    XRAM[11189] = 8'b0;
    XRAM[11190] = 8'b0;
    XRAM[11191] = 8'b0;
    XRAM[11192] = 8'b0;
    XRAM[11193] = 8'b0;
    XRAM[11194] = 8'b0;
    XRAM[11195] = 8'b0;
    XRAM[11196] = 8'b0;
    XRAM[11197] = 8'b0;
    XRAM[11198] = 8'b0;
    XRAM[11199] = 8'b0;
    XRAM[11200] = 8'b0;
    XRAM[11201] = 8'b0;
    XRAM[11202] = 8'b0;
    XRAM[11203] = 8'b0;
    XRAM[11204] = 8'b0;
    XRAM[11205] = 8'b0;
    XRAM[11206] = 8'b0;
    XRAM[11207] = 8'b0;
    XRAM[11208] = 8'b0;
    XRAM[11209] = 8'b0;
    XRAM[11210] = 8'b0;
    XRAM[11211] = 8'b0;
    XRAM[11212] = 8'b0;
    XRAM[11213] = 8'b0;
    XRAM[11214] = 8'b0;
    XRAM[11215] = 8'b0;
    XRAM[11216] = 8'b0;
    XRAM[11217] = 8'b0;
    XRAM[11218] = 8'b0;
    XRAM[11219] = 8'b0;
    XRAM[11220] = 8'b0;
    XRAM[11221] = 8'b0;
    XRAM[11222] = 8'b0;
    XRAM[11223] = 8'b0;
    XRAM[11224] = 8'b0;
    XRAM[11225] = 8'b0;
    XRAM[11226] = 8'b0;
    XRAM[11227] = 8'b0;
    XRAM[11228] = 8'b0;
    XRAM[11229] = 8'b0;
    XRAM[11230] = 8'b0;
    XRAM[11231] = 8'b0;
    XRAM[11232] = 8'b0;
    XRAM[11233] = 8'b0;
    XRAM[11234] = 8'b0;
    XRAM[11235] = 8'b0;
    XRAM[11236] = 8'b0;
    XRAM[11237] = 8'b0;
    XRAM[11238] = 8'b0;
    XRAM[11239] = 8'b0;
    XRAM[11240] = 8'b0;
    XRAM[11241] = 8'b0;
    XRAM[11242] = 8'b0;
    XRAM[11243] = 8'b0;
    XRAM[11244] = 8'b0;
    XRAM[11245] = 8'b0;
    XRAM[11246] = 8'b0;
    XRAM[11247] = 8'b0;
    XRAM[11248] = 8'b0;
    XRAM[11249] = 8'b0;
    XRAM[11250] = 8'b0;
    XRAM[11251] = 8'b0;
    XRAM[11252] = 8'b0;
    XRAM[11253] = 8'b0;
    XRAM[11254] = 8'b0;
    XRAM[11255] = 8'b0;
    XRAM[11256] = 8'b0;
    XRAM[11257] = 8'b0;
    XRAM[11258] = 8'b0;
    XRAM[11259] = 8'b0;
    XRAM[11260] = 8'b0;
    XRAM[11261] = 8'b0;
    XRAM[11262] = 8'b0;
    XRAM[11263] = 8'b0;
    XRAM[11264] = 8'b0;
    XRAM[11265] = 8'b0;
    XRAM[11266] = 8'b0;
    XRAM[11267] = 8'b0;
    XRAM[11268] = 8'b0;
    XRAM[11269] = 8'b0;
    XRAM[11270] = 8'b0;
    XRAM[11271] = 8'b0;
    XRAM[11272] = 8'b0;
    XRAM[11273] = 8'b0;
    XRAM[11274] = 8'b0;
    XRAM[11275] = 8'b0;
    XRAM[11276] = 8'b0;
    XRAM[11277] = 8'b0;
    XRAM[11278] = 8'b0;
    XRAM[11279] = 8'b0;
    XRAM[11280] = 8'b0;
    XRAM[11281] = 8'b0;
    XRAM[11282] = 8'b0;
    XRAM[11283] = 8'b0;
    XRAM[11284] = 8'b0;
    XRAM[11285] = 8'b0;
    XRAM[11286] = 8'b0;
    XRAM[11287] = 8'b0;
    XRAM[11288] = 8'b0;
    XRAM[11289] = 8'b0;
    XRAM[11290] = 8'b0;
    XRAM[11291] = 8'b0;
    XRAM[11292] = 8'b0;
    XRAM[11293] = 8'b0;
    XRAM[11294] = 8'b0;
    XRAM[11295] = 8'b0;
    XRAM[11296] = 8'b0;
    XRAM[11297] = 8'b0;
    XRAM[11298] = 8'b0;
    XRAM[11299] = 8'b0;
    XRAM[11300] = 8'b0;
    XRAM[11301] = 8'b0;
    XRAM[11302] = 8'b0;
    XRAM[11303] = 8'b0;
    XRAM[11304] = 8'b0;
    XRAM[11305] = 8'b0;
    XRAM[11306] = 8'b0;
    XRAM[11307] = 8'b0;
    XRAM[11308] = 8'b0;
    XRAM[11309] = 8'b0;
    XRAM[11310] = 8'b0;
    XRAM[11311] = 8'b0;
    XRAM[11312] = 8'b0;
    XRAM[11313] = 8'b0;
    XRAM[11314] = 8'b0;
    XRAM[11315] = 8'b0;
    XRAM[11316] = 8'b0;
    XRAM[11317] = 8'b0;
    XRAM[11318] = 8'b0;
    XRAM[11319] = 8'b0;
    XRAM[11320] = 8'b0;
    XRAM[11321] = 8'b0;
    XRAM[11322] = 8'b0;
    XRAM[11323] = 8'b0;
    XRAM[11324] = 8'b0;
    XRAM[11325] = 8'b0;
    XRAM[11326] = 8'b0;
    XRAM[11327] = 8'b0;
    XRAM[11328] = 8'b0;
    XRAM[11329] = 8'b0;
    XRAM[11330] = 8'b0;
    XRAM[11331] = 8'b0;
    XRAM[11332] = 8'b0;
    XRAM[11333] = 8'b0;
    XRAM[11334] = 8'b0;
    XRAM[11335] = 8'b0;
    XRAM[11336] = 8'b0;
    XRAM[11337] = 8'b0;
    XRAM[11338] = 8'b0;
    XRAM[11339] = 8'b0;
    XRAM[11340] = 8'b0;
    XRAM[11341] = 8'b0;
    XRAM[11342] = 8'b0;
    XRAM[11343] = 8'b0;
    XRAM[11344] = 8'b0;
    XRAM[11345] = 8'b0;
    XRAM[11346] = 8'b0;
    XRAM[11347] = 8'b0;
    XRAM[11348] = 8'b0;
    XRAM[11349] = 8'b0;
    XRAM[11350] = 8'b0;
    XRAM[11351] = 8'b0;
    XRAM[11352] = 8'b0;
    XRAM[11353] = 8'b0;
    XRAM[11354] = 8'b0;
    XRAM[11355] = 8'b0;
    XRAM[11356] = 8'b0;
    XRAM[11357] = 8'b0;
    XRAM[11358] = 8'b0;
    XRAM[11359] = 8'b0;
    XRAM[11360] = 8'b0;
    XRAM[11361] = 8'b0;
    XRAM[11362] = 8'b0;
    XRAM[11363] = 8'b0;
    XRAM[11364] = 8'b0;
    XRAM[11365] = 8'b0;
    XRAM[11366] = 8'b0;
    XRAM[11367] = 8'b0;
    XRAM[11368] = 8'b0;
    XRAM[11369] = 8'b0;
    XRAM[11370] = 8'b0;
    XRAM[11371] = 8'b0;
    XRAM[11372] = 8'b0;
    XRAM[11373] = 8'b0;
    XRAM[11374] = 8'b0;
    XRAM[11375] = 8'b0;
    XRAM[11376] = 8'b0;
    XRAM[11377] = 8'b0;
    XRAM[11378] = 8'b0;
    XRAM[11379] = 8'b0;
    XRAM[11380] = 8'b0;
    XRAM[11381] = 8'b0;
    XRAM[11382] = 8'b0;
    XRAM[11383] = 8'b0;
    XRAM[11384] = 8'b0;
    XRAM[11385] = 8'b0;
    XRAM[11386] = 8'b0;
    XRAM[11387] = 8'b0;
    XRAM[11388] = 8'b0;
    XRAM[11389] = 8'b0;
    XRAM[11390] = 8'b0;
    XRAM[11391] = 8'b0;
    XRAM[11392] = 8'b0;
    XRAM[11393] = 8'b0;
    XRAM[11394] = 8'b0;
    XRAM[11395] = 8'b0;
    XRAM[11396] = 8'b0;
    XRAM[11397] = 8'b0;
    XRAM[11398] = 8'b0;
    XRAM[11399] = 8'b0;
    XRAM[11400] = 8'b0;
    XRAM[11401] = 8'b0;
    XRAM[11402] = 8'b0;
    XRAM[11403] = 8'b0;
    XRAM[11404] = 8'b0;
    XRAM[11405] = 8'b0;
    XRAM[11406] = 8'b0;
    XRAM[11407] = 8'b0;
    XRAM[11408] = 8'b0;
    XRAM[11409] = 8'b0;
    XRAM[11410] = 8'b0;
    XRAM[11411] = 8'b0;
    XRAM[11412] = 8'b0;
    XRAM[11413] = 8'b0;
    XRAM[11414] = 8'b0;
    XRAM[11415] = 8'b0;
    XRAM[11416] = 8'b0;
    XRAM[11417] = 8'b0;
    XRAM[11418] = 8'b0;
    XRAM[11419] = 8'b0;
    XRAM[11420] = 8'b0;
    XRAM[11421] = 8'b0;
    XRAM[11422] = 8'b0;
    XRAM[11423] = 8'b0;
    XRAM[11424] = 8'b0;
    XRAM[11425] = 8'b0;
    XRAM[11426] = 8'b0;
    XRAM[11427] = 8'b0;
    XRAM[11428] = 8'b0;
    XRAM[11429] = 8'b0;
    XRAM[11430] = 8'b0;
    XRAM[11431] = 8'b0;
    XRAM[11432] = 8'b0;
    XRAM[11433] = 8'b0;
    XRAM[11434] = 8'b0;
    XRAM[11435] = 8'b0;
    XRAM[11436] = 8'b0;
    XRAM[11437] = 8'b0;
    XRAM[11438] = 8'b0;
    XRAM[11439] = 8'b0;
    XRAM[11440] = 8'b0;
    XRAM[11441] = 8'b0;
    XRAM[11442] = 8'b0;
    XRAM[11443] = 8'b0;
    XRAM[11444] = 8'b0;
    XRAM[11445] = 8'b0;
    XRAM[11446] = 8'b0;
    XRAM[11447] = 8'b0;
    XRAM[11448] = 8'b0;
    XRAM[11449] = 8'b0;
    XRAM[11450] = 8'b0;
    XRAM[11451] = 8'b0;
    XRAM[11452] = 8'b0;
    XRAM[11453] = 8'b0;
    XRAM[11454] = 8'b0;
    XRAM[11455] = 8'b0;
    XRAM[11456] = 8'b0;
    XRAM[11457] = 8'b0;
    XRAM[11458] = 8'b0;
    XRAM[11459] = 8'b0;
    XRAM[11460] = 8'b0;
    XRAM[11461] = 8'b0;
    XRAM[11462] = 8'b0;
    XRAM[11463] = 8'b0;
    XRAM[11464] = 8'b0;
    XRAM[11465] = 8'b0;
    XRAM[11466] = 8'b0;
    XRAM[11467] = 8'b0;
    XRAM[11468] = 8'b0;
    XRAM[11469] = 8'b0;
    XRAM[11470] = 8'b0;
    XRAM[11471] = 8'b0;
    XRAM[11472] = 8'b0;
    XRAM[11473] = 8'b0;
    XRAM[11474] = 8'b0;
    XRAM[11475] = 8'b0;
    XRAM[11476] = 8'b0;
    XRAM[11477] = 8'b0;
    XRAM[11478] = 8'b0;
    XRAM[11479] = 8'b0;
    XRAM[11480] = 8'b0;
    XRAM[11481] = 8'b0;
    XRAM[11482] = 8'b0;
    XRAM[11483] = 8'b0;
    XRAM[11484] = 8'b0;
    XRAM[11485] = 8'b0;
    XRAM[11486] = 8'b0;
    XRAM[11487] = 8'b0;
    XRAM[11488] = 8'b0;
    XRAM[11489] = 8'b0;
    XRAM[11490] = 8'b0;
    XRAM[11491] = 8'b0;
    XRAM[11492] = 8'b0;
    XRAM[11493] = 8'b0;
    XRAM[11494] = 8'b0;
    XRAM[11495] = 8'b0;
    XRAM[11496] = 8'b0;
    XRAM[11497] = 8'b0;
    XRAM[11498] = 8'b0;
    XRAM[11499] = 8'b0;
    XRAM[11500] = 8'b0;
    XRAM[11501] = 8'b0;
    XRAM[11502] = 8'b0;
    XRAM[11503] = 8'b0;
    XRAM[11504] = 8'b0;
    XRAM[11505] = 8'b0;
    XRAM[11506] = 8'b0;
    XRAM[11507] = 8'b0;
    XRAM[11508] = 8'b0;
    XRAM[11509] = 8'b0;
    XRAM[11510] = 8'b0;
    XRAM[11511] = 8'b0;
    XRAM[11512] = 8'b0;
    XRAM[11513] = 8'b0;
    XRAM[11514] = 8'b0;
    XRAM[11515] = 8'b0;
    XRAM[11516] = 8'b0;
    XRAM[11517] = 8'b0;
    XRAM[11518] = 8'b0;
    XRAM[11519] = 8'b0;
    XRAM[11520] = 8'b0;
    XRAM[11521] = 8'b0;
    XRAM[11522] = 8'b0;
    XRAM[11523] = 8'b0;
    XRAM[11524] = 8'b0;
    XRAM[11525] = 8'b0;
    XRAM[11526] = 8'b0;
    XRAM[11527] = 8'b0;
    XRAM[11528] = 8'b0;
    XRAM[11529] = 8'b0;
    XRAM[11530] = 8'b0;
    XRAM[11531] = 8'b0;
    XRAM[11532] = 8'b0;
    XRAM[11533] = 8'b0;
    XRAM[11534] = 8'b0;
    XRAM[11535] = 8'b0;
    XRAM[11536] = 8'b0;
    XRAM[11537] = 8'b0;
    XRAM[11538] = 8'b0;
    XRAM[11539] = 8'b0;
    XRAM[11540] = 8'b0;
    XRAM[11541] = 8'b0;
    XRAM[11542] = 8'b0;
    XRAM[11543] = 8'b0;
    XRAM[11544] = 8'b0;
    XRAM[11545] = 8'b0;
    XRAM[11546] = 8'b0;
    XRAM[11547] = 8'b0;
    XRAM[11548] = 8'b0;
    XRAM[11549] = 8'b0;
    XRAM[11550] = 8'b0;
    XRAM[11551] = 8'b0;
    XRAM[11552] = 8'b0;
    XRAM[11553] = 8'b0;
    XRAM[11554] = 8'b0;
    XRAM[11555] = 8'b0;
    XRAM[11556] = 8'b0;
    XRAM[11557] = 8'b0;
    XRAM[11558] = 8'b0;
    XRAM[11559] = 8'b0;
    XRAM[11560] = 8'b0;
    XRAM[11561] = 8'b0;
    XRAM[11562] = 8'b0;
    XRAM[11563] = 8'b0;
    XRAM[11564] = 8'b0;
    XRAM[11565] = 8'b0;
    XRAM[11566] = 8'b0;
    XRAM[11567] = 8'b0;
    XRAM[11568] = 8'b0;
    XRAM[11569] = 8'b0;
    XRAM[11570] = 8'b0;
    XRAM[11571] = 8'b0;
    XRAM[11572] = 8'b0;
    XRAM[11573] = 8'b0;
    XRAM[11574] = 8'b0;
    XRAM[11575] = 8'b0;
    XRAM[11576] = 8'b0;
    XRAM[11577] = 8'b0;
    XRAM[11578] = 8'b0;
    XRAM[11579] = 8'b0;
    XRAM[11580] = 8'b0;
    XRAM[11581] = 8'b0;
    XRAM[11582] = 8'b0;
    XRAM[11583] = 8'b0;
    XRAM[11584] = 8'b0;
    XRAM[11585] = 8'b0;
    XRAM[11586] = 8'b0;
    XRAM[11587] = 8'b0;
    XRAM[11588] = 8'b0;
    XRAM[11589] = 8'b0;
    XRAM[11590] = 8'b0;
    XRAM[11591] = 8'b0;
    XRAM[11592] = 8'b0;
    XRAM[11593] = 8'b0;
    XRAM[11594] = 8'b0;
    XRAM[11595] = 8'b0;
    XRAM[11596] = 8'b0;
    XRAM[11597] = 8'b0;
    XRAM[11598] = 8'b0;
    XRAM[11599] = 8'b0;
    XRAM[11600] = 8'b0;
    XRAM[11601] = 8'b0;
    XRAM[11602] = 8'b0;
    XRAM[11603] = 8'b0;
    XRAM[11604] = 8'b0;
    XRAM[11605] = 8'b0;
    XRAM[11606] = 8'b0;
    XRAM[11607] = 8'b0;
    XRAM[11608] = 8'b0;
    XRAM[11609] = 8'b0;
    XRAM[11610] = 8'b0;
    XRAM[11611] = 8'b0;
    XRAM[11612] = 8'b0;
    XRAM[11613] = 8'b0;
    XRAM[11614] = 8'b0;
    XRAM[11615] = 8'b0;
    XRAM[11616] = 8'b0;
    XRAM[11617] = 8'b0;
    XRAM[11618] = 8'b0;
    XRAM[11619] = 8'b0;
    XRAM[11620] = 8'b0;
    XRAM[11621] = 8'b0;
    XRAM[11622] = 8'b0;
    XRAM[11623] = 8'b0;
    XRAM[11624] = 8'b0;
    XRAM[11625] = 8'b0;
    XRAM[11626] = 8'b0;
    XRAM[11627] = 8'b0;
    XRAM[11628] = 8'b0;
    XRAM[11629] = 8'b0;
    XRAM[11630] = 8'b0;
    XRAM[11631] = 8'b0;
    XRAM[11632] = 8'b0;
    XRAM[11633] = 8'b0;
    XRAM[11634] = 8'b0;
    XRAM[11635] = 8'b0;
    XRAM[11636] = 8'b0;
    XRAM[11637] = 8'b0;
    XRAM[11638] = 8'b0;
    XRAM[11639] = 8'b0;
    XRAM[11640] = 8'b0;
    XRAM[11641] = 8'b0;
    XRAM[11642] = 8'b0;
    XRAM[11643] = 8'b0;
    XRAM[11644] = 8'b0;
    XRAM[11645] = 8'b0;
    XRAM[11646] = 8'b0;
    XRAM[11647] = 8'b0;
    XRAM[11648] = 8'b0;
    XRAM[11649] = 8'b0;
    XRAM[11650] = 8'b0;
    XRAM[11651] = 8'b0;
    XRAM[11652] = 8'b0;
    XRAM[11653] = 8'b0;
    XRAM[11654] = 8'b0;
    XRAM[11655] = 8'b0;
    XRAM[11656] = 8'b0;
    XRAM[11657] = 8'b0;
    XRAM[11658] = 8'b0;
    XRAM[11659] = 8'b0;
    XRAM[11660] = 8'b0;
    XRAM[11661] = 8'b0;
    XRAM[11662] = 8'b0;
    XRAM[11663] = 8'b0;
    XRAM[11664] = 8'b0;
    XRAM[11665] = 8'b0;
    XRAM[11666] = 8'b0;
    XRAM[11667] = 8'b0;
    XRAM[11668] = 8'b0;
    XRAM[11669] = 8'b0;
    XRAM[11670] = 8'b0;
    XRAM[11671] = 8'b0;
    XRAM[11672] = 8'b0;
    XRAM[11673] = 8'b0;
    XRAM[11674] = 8'b0;
    XRAM[11675] = 8'b0;
    XRAM[11676] = 8'b0;
    XRAM[11677] = 8'b0;
    XRAM[11678] = 8'b0;
    XRAM[11679] = 8'b0;
    XRAM[11680] = 8'b0;
    XRAM[11681] = 8'b0;
    XRAM[11682] = 8'b0;
    XRAM[11683] = 8'b0;
    XRAM[11684] = 8'b0;
    XRAM[11685] = 8'b0;
    XRAM[11686] = 8'b0;
    XRAM[11687] = 8'b0;
    XRAM[11688] = 8'b0;
    XRAM[11689] = 8'b0;
    XRAM[11690] = 8'b0;
    XRAM[11691] = 8'b0;
    XRAM[11692] = 8'b0;
    XRAM[11693] = 8'b0;
    XRAM[11694] = 8'b0;
    XRAM[11695] = 8'b0;
    XRAM[11696] = 8'b0;
    XRAM[11697] = 8'b0;
    XRAM[11698] = 8'b0;
    XRAM[11699] = 8'b0;
    XRAM[11700] = 8'b0;
    XRAM[11701] = 8'b0;
    XRAM[11702] = 8'b0;
    XRAM[11703] = 8'b0;
    XRAM[11704] = 8'b0;
    XRAM[11705] = 8'b0;
    XRAM[11706] = 8'b0;
    XRAM[11707] = 8'b0;
    XRAM[11708] = 8'b0;
    XRAM[11709] = 8'b0;
    XRAM[11710] = 8'b0;
    XRAM[11711] = 8'b0;
    XRAM[11712] = 8'b0;
    XRAM[11713] = 8'b0;
    XRAM[11714] = 8'b0;
    XRAM[11715] = 8'b0;
    XRAM[11716] = 8'b0;
    XRAM[11717] = 8'b0;
    XRAM[11718] = 8'b0;
    XRAM[11719] = 8'b0;
    XRAM[11720] = 8'b0;
    XRAM[11721] = 8'b0;
    XRAM[11722] = 8'b0;
    XRAM[11723] = 8'b0;
    XRAM[11724] = 8'b0;
    XRAM[11725] = 8'b0;
    XRAM[11726] = 8'b0;
    XRAM[11727] = 8'b0;
    XRAM[11728] = 8'b0;
    XRAM[11729] = 8'b0;
    XRAM[11730] = 8'b0;
    XRAM[11731] = 8'b0;
    XRAM[11732] = 8'b0;
    XRAM[11733] = 8'b0;
    XRAM[11734] = 8'b0;
    XRAM[11735] = 8'b0;
    XRAM[11736] = 8'b0;
    XRAM[11737] = 8'b0;
    XRAM[11738] = 8'b0;
    XRAM[11739] = 8'b0;
    XRAM[11740] = 8'b0;
    XRAM[11741] = 8'b0;
    XRAM[11742] = 8'b0;
    XRAM[11743] = 8'b0;
    XRAM[11744] = 8'b0;
    XRAM[11745] = 8'b0;
    XRAM[11746] = 8'b0;
    XRAM[11747] = 8'b0;
    XRAM[11748] = 8'b0;
    XRAM[11749] = 8'b0;
    XRAM[11750] = 8'b0;
    XRAM[11751] = 8'b0;
    XRAM[11752] = 8'b0;
    XRAM[11753] = 8'b0;
    XRAM[11754] = 8'b0;
    XRAM[11755] = 8'b0;
    XRAM[11756] = 8'b0;
    XRAM[11757] = 8'b0;
    XRAM[11758] = 8'b0;
    XRAM[11759] = 8'b0;
    XRAM[11760] = 8'b0;
    XRAM[11761] = 8'b0;
    XRAM[11762] = 8'b0;
    XRAM[11763] = 8'b0;
    XRAM[11764] = 8'b0;
    XRAM[11765] = 8'b0;
    XRAM[11766] = 8'b0;
    XRAM[11767] = 8'b0;
    XRAM[11768] = 8'b0;
    XRAM[11769] = 8'b0;
    XRAM[11770] = 8'b0;
    XRAM[11771] = 8'b0;
    XRAM[11772] = 8'b0;
    XRAM[11773] = 8'b0;
    XRAM[11774] = 8'b0;
    XRAM[11775] = 8'b0;
    XRAM[11776] = 8'b0;
    XRAM[11777] = 8'b0;
    XRAM[11778] = 8'b0;
    XRAM[11779] = 8'b0;
    XRAM[11780] = 8'b0;
    XRAM[11781] = 8'b0;
    XRAM[11782] = 8'b0;
    XRAM[11783] = 8'b0;
    XRAM[11784] = 8'b0;
    XRAM[11785] = 8'b0;
    XRAM[11786] = 8'b0;
    XRAM[11787] = 8'b0;
    XRAM[11788] = 8'b0;
    XRAM[11789] = 8'b0;
    XRAM[11790] = 8'b0;
    XRAM[11791] = 8'b0;
    XRAM[11792] = 8'b0;
    XRAM[11793] = 8'b0;
    XRAM[11794] = 8'b0;
    XRAM[11795] = 8'b0;
    XRAM[11796] = 8'b0;
    XRAM[11797] = 8'b0;
    XRAM[11798] = 8'b0;
    XRAM[11799] = 8'b0;
    XRAM[11800] = 8'b0;
    XRAM[11801] = 8'b0;
    XRAM[11802] = 8'b0;
    XRAM[11803] = 8'b0;
    XRAM[11804] = 8'b0;
    XRAM[11805] = 8'b0;
    XRAM[11806] = 8'b0;
    XRAM[11807] = 8'b0;
    XRAM[11808] = 8'b0;
    XRAM[11809] = 8'b0;
    XRAM[11810] = 8'b0;
    XRAM[11811] = 8'b0;
    XRAM[11812] = 8'b0;
    XRAM[11813] = 8'b0;
    XRAM[11814] = 8'b0;
    XRAM[11815] = 8'b0;
    XRAM[11816] = 8'b0;
    XRAM[11817] = 8'b0;
    XRAM[11818] = 8'b0;
    XRAM[11819] = 8'b0;
    XRAM[11820] = 8'b0;
    XRAM[11821] = 8'b0;
    XRAM[11822] = 8'b0;
    XRAM[11823] = 8'b0;
    XRAM[11824] = 8'b0;
    XRAM[11825] = 8'b0;
    XRAM[11826] = 8'b0;
    XRAM[11827] = 8'b0;
    XRAM[11828] = 8'b0;
    XRAM[11829] = 8'b0;
    XRAM[11830] = 8'b0;
    XRAM[11831] = 8'b0;
    XRAM[11832] = 8'b0;
    XRAM[11833] = 8'b0;
    XRAM[11834] = 8'b0;
    XRAM[11835] = 8'b0;
    XRAM[11836] = 8'b0;
    XRAM[11837] = 8'b0;
    XRAM[11838] = 8'b0;
    XRAM[11839] = 8'b0;
    XRAM[11840] = 8'b0;
    XRAM[11841] = 8'b0;
    XRAM[11842] = 8'b0;
    XRAM[11843] = 8'b0;
    XRAM[11844] = 8'b0;
    XRAM[11845] = 8'b0;
    XRAM[11846] = 8'b0;
    XRAM[11847] = 8'b0;
    XRAM[11848] = 8'b0;
    XRAM[11849] = 8'b0;
    XRAM[11850] = 8'b0;
    XRAM[11851] = 8'b0;
    XRAM[11852] = 8'b0;
    XRAM[11853] = 8'b0;
    XRAM[11854] = 8'b0;
    XRAM[11855] = 8'b0;
    XRAM[11856] = 8'b0;
    XRAM[11857] = 8'b0;
    XRAM[11858] = 8'b0;
    XRAM[11859] = 8'b0;
    XRAM[11860] = 8'b0;
    XRAM[11861] = 8'b0;
    XRAM[11862] = 8'b0;
    XRAM[11863] = 8'b0;
    XRAM[11864] = 8'b0;
    XRAM[11865] = 8'b0;
    XRAM[11866] = 8'b0;
    XRAM[11867] = 8'b0;
    XRAM[11868] = 8'b0;
    XRAM[11869] = 8'b0;
    XRAM[11870] = 8'b0;
    XRAM[11871] = 8'b0;
    XRAM[11872] = 8'b0;
    XRAM[11873] = 8'b0;
    XRAM[11874] = 8'b0;
    XRAM[11875] = 8'b0;
    XRAM[11876] = 8'b0;
    XRAM[11877] = 8'b0;
    XRAM[11878] = 8'b0;
    XRAM[11879] = 8'b0;
    XRAM[11880] = 8'b0;
    XRAM[11881] = 8'b0;
    XRAM[11882] = 8'b0;
    XRAM[11883] = 8'b0;
    XRAM[11884] = 8'b0;
    XRAM[11885] = 8'b0;
    XRAM[11886] = 8'b0;
    XRAM[11887] = 8'b0;
    XRAM[11888] = 8'b0;
    XRAM[11889] = 8'b0;
    XRAM[11890] = 8'b0;
    XRAM[11891] = 8'b0;
    XRAM[11892] = 8'b0;
    XRAM[11893] = 8'b0;
    XRAM[11894] = 8'b0;
    XRAM[11895] = 8'b0;
    XRAM[11896] = 8'b0;
    XRAM[11897] = 8'b0;
    XRAM[11898] = 8'b0;
    XRAM[11899] = 8'b0;
    XRAM[11900] = 8'b0;
    XRAM[11901] = 8'b0;
    XRAM[11902] = 8'b0;
    XRAM[11903] = 8'b0;
    XRAM[11904] = 8'b0;
    XRAM[11905] = 8'b0;
    XRAM[11906] = 8'b0;
    XRAM[11907] = 8'b0;
    XRAM[11908] = 8'b0;
    XRAM[11909] = 8'b0;
    XRAM[11910] = 8'b0;
    XRAM[11911] = 8'b0;
    XRAM[11912] = 8'b0;
    XRAM[11913] = 8'b0;
    XRAM[11914] = 8'b0;
    XRAM[11915] = 8'b0;
    XRAM[11916] = 8'b0;
    XRAM[11917] = 8'b0;
    XRAM[11918] = 8'b0;
    XRAM[11919] = 8'b0;
    XRAM[11920] = 8'b0;
    XRAM[11921] = 8'b0;
    XRAM[11922] = 8'b0;
    XRAM[11923] = 8'b0;
    XRAM[11924] = 8'b0;
    XRAM[11925] = 8'b0;
    XRAM[11926] = 8'b0;
    XRAM[11927] = 8'b0;
    XRAM[11928] = 8'b0;
    XRAM[11929] = 8'b0;
    XRAM[11930] = 8'b0;
    XRAM[11931] = 8'b0;
    XRAM[11932] = 8'b0;
    XRAM[11933] = 8'b0;
    XRAM[11934] = 8'b0;
    XRAM[11935] = 8'b0;
    XRAM[11936] = 8'b0;
    XRAM[11937] = 8'b0;
    XRAM[11938] = 8'b0;
    XRAM[11939] = 8'b0;
    XRAM[11940] = 8'b0;
    XRAM[11941] = 8'b0;
    XRAM[11942] = 8'b0;
    XRAM[11943] = 8'b0;
    XRAM[11944] = 8'b0;
    XRAM[11945] = 8'b0;
    XRAM[11946] = 8'b0;
    XRAM[11947] = 8'b0;
    XRAM[11948] = 8'b0;
    XRAM[11949] = 8'b0;
    XRAM[11950] = 8'b0;
    XRAM[11951] = 8'b0;
    XRAM[11952] = 8'b0;
    XRAM[11953] = 8'b0;
    XRAM[11954] = 8'b0;
    XRAM[11955] = 8'b0;
    XRAM[11956] = 8'b0;
    XRAM[11957] = 8'b0;
    XRAM[11958] = 8'b0;
    XRAM[11959] = 8'b0;
    XRAM[11960] = 8'b0;
    XRAM[11961] = 8'b0;
    XRAM[11962] = 8'b0;
    XRAM[11963] = 8'b0;
    XRAM[11964] = 8'b0;
    XRAM[11965] = 8'b0;
    XRAM[11966] = 8'b0;
    XRAM[11967] = 8'b0;
    XRAM[11968] = 8'b0;
    XRAM[11969] = 8'b0;
    XRAM[11970] = 8'b0;
    XRAM[11971] = 8'b0;
    XRAM[11972] = 8'b0;
    XRAM[11973] = 8'b0;
    XRAM[11974] = 8'b0;
    XRAM[11975] = 8'b0;
    XRAM[11976] = 8'b0;
    XRAM[11977] = 8'b0;
    XRAM[11978] = 8'b0;
    XRAM[11979] = 8'b0;
    XRAM[11980] = 8'b0;
    XRAM[11981] = 8'b0;
    XRAM[11982] = 8'b0;
    XRAM[11983] = 8'b0;
    XRAM[11984] = 8'b0;
    XRAM[11985] = 8'b0;
    XRAM[11986] = 8'b0;
    XRAM[11987] = 8'b0;
    XRAM[11988] = 8'b0;
    XRAM[11989] = 8'b0;
    XRAM[11990] = 8'b0;
    XRAM[11991] = 8'b0;
    XRAM[11992] = 8'b0;
    XRAM[11993] = 8'b0;
    XRAM[11994] = 8'b0;
    XRAM[11995] = 8'b0;
    XRAM[11996] = 8'b0;
    XRAM[11997] = 8'b0;
    XRAM[11998] = 8'b0;
    XRAM[11999] = 8'b0;
    XRAM[12000] = 8'b0;
    XRAM[12001] = 8'b0;
    XRAM[12002] = 8'b0;
    XRAM[12003] = 8'b0;
    XRAM[12004] = 8'b0;
    XRAM[12005] = 8'b0;
    XRAM[12006] = 8'b0;
    XRAM[12007] = 8'b0;
    XRAM[12008] = 8'b0;
    XRAM[12009] = 8'b0;
    XRAM[12010] = 8'b0;
    XRAM[12011] = 8'b0;
    XRAM[12012] = 8'b0;
    XRAM[12013] = 8'b0;
    XRAM[12014] = 8'b0;
    XRAM[12015] = 8'b0;
    XRAM[12016] = 8'b0;
    XRAM[12017] = 8'b0;
    XRAM[12018] = 8'b0;
    XRAM[12019] = 8'b0;
    XRAM[12020] = 8'b0;
    XRAM[12021] = 8'b0;
    XRAM[12022] = 8'b0;
    XRAM[12023] = 8'b0;
    XRAM[12024] = 8'b0;
    XRAM[12025] = 8'b0;
    XRAM[12026] = 8'b0;
    XRAM[12027] = 8'b0;
    XRAM[12028] = 8'b0;
    XRAM[12029] = 8'b0;
    XRAM[12030] = 8'b0;
    XRAM[12031] = 8'b0;
    XRAM[12032] = 8'b0;
    XRAM[12033] = 8'b0;
    XRAM[12034] = 8'b0;
    XRAM[12035] = 8'b0;
    XRAM[12036] = 8'b0;
    XRAM[12037] = 8'b0;
    XRAM[12038] = 8'b0;
    XRAM[12039] = 8'b0;
    XRAM[12040] = 8'b0;
    XRAM[12041] = 8'b0;
    XRAM[12042] = 8'b0;
    XRAM[12043] = 8'b0;
    XRAM[12044] = 8'b0;
    XRAM[12045] = 8'b0;
    XRAM[12046] = 8'b0;
    XRAM[12047] = 8'b0;
    XRAM[12048] = 8'b0;
    XRAM[12049] = 8'b0;
    XRAM[12050] = 8'b0;
    XRAM[12051] = 8'b0;
    XRAM[12052] = 8'b0;
    XRAM[12053] = 8'b0;
    XRAM[12054] = 8'b0;
    XRAM[12055] = 8'b0;
    XRAM[12056] = 8'b0;
    XRAM[12057] = 8'b0;
    XRAM[12058] = 8'b0;
    XRAM[12059] = 8'b0;
    XRAM[12060] = 8'b0;
    XRAM[12061] = 8'b0;
    XRAM[12062] = 8'b0;
    XRAM[12063] = 8'b0;
    XRAM[12064] = 8'b0;
    XRAM[12065] = 8'b0;
    XRAM[12066] = 8'b0;
    XRAM[12067] = 8'b0;
    XRAM[12068] = 8'b0;
    XRAM[12069] = 8'b0;
    XRAM[12070] = 8'b0;
    XRAM[12071] = 8'b0;
    XRAM[12072] = 8'b0;
    XRAM[12073] = 8'b0;
    XRAM[12074] = 8'b0;
    XRAM[12075] = 8'b0;
    XRAM[12076] = 8'b0;
    XRAM[12077] = 8'b0;
    XRAM[12078] = 8'b0;
    XRAM[12079] = 8'b0;
    XRAM[12080] = 8'b0;
    XRAM[12081] = 8'b0;
    XRAM[12082] = 8'b0;
    XRAM[12083] = 8'b0;
    XRAM[12084] = 8'b0;
    XRAM[12085] = 8'b0;
    XRAM[12086] = 8'b0;
    XRAM[12087] = 8'b0;
    XRAM[12088] = 8'b0;
    XRAM[12089] = 8'b0;
    XRAM[12090] = 8'b0;
    XRAM[12091] = 8'b0;
    XRAM[12092] = 8'b0;
    XRAM[12093] = 8'b0;
    XRAM[12094] = 8'b0;
    XRAM[12095] = 8'b0;
    XRAM[12096] = 8'b0;
    XRAM[12097] = 8'b0;
    XRAM[12098] = 8'b0;
    XRAM[12099] = 8'b0;
    XRAM[12100] = 8'b0;
    XRAM[12101] = 8'b0;
    XRAM[12102] = 8'b0;
    XRAM[12103] = 8'b0;
    XRAM[12104] = 8'b0;
    XRAM[12105] = 8'b0;
    XRAM[12106] = 8'b0;
    XRAM[12107] = 8'b0;
    XRAM[12108] = 8'b0;
    XRAM[12109] = 8'b0;
    XRAM[12110] = 8'b0;
    XRAM[12111] = 8'b0;
    XRAM[12112] = 8'b0;
    XRAM[12113] = 8'b0;
    XRAM[12114] = 8'b0;
    XRAM[12115] = 8'b0;
    XRAM[12116] = 8'b0;
    XRAM[12117] = 8'b0;
    XRAM[12118] = 8'b0;
    XRAM[12119] = 8'b0;
    XRAM[12120] = 8'b0;
    XRAM[12121] = 8'b0;
    XRAM[12122] = 8'b0;
    XRAM[12123] = 8'b0;
    XRAM[12124] = 8'b0;
    XRAM[12125] = 8'b0;
    XRAM[12126] = 8'b0;
    XRAM[12127] = 8'b0;
    XRAM[12128] = 8'b0;
    XRAM[12129] = 8'b0;
    XRAM[12130] = 8'b0;
    XRAM[12131] = 8'b0;
    XRAM[12132] = 8'b0;
    XRAM[12133] = 8'b0;
    XRAM[12134] = 8'b0;
    XRAM[12135] = 8'b0;
    XRAM[12136] = 8'b0;
    XRAM[12137] = 8'b0;
    XRAM[12138] = 8'b0;
    XRAM[12139] = 8'b0;
    XRAM[12140] = 8'b0;
    XRAM[12141] = 8'b0;
    XRAM[12142] = 8'b0;
    XRAM[12143] = 8'b0;
    XRAM[12144] = 8'b0;
    XRAM[12145] = 8'b0;
    XRAM[12146] = 8'b0;
    XRAM[12147] = 8'b0;
    XRAM[12148] = 8'b0;
    XRAM[12149] = 8'b0;
    XRAM[12150] = 8'b0;
    XRAM[12151] = 8'b0;
    XRAM[12152] = 8'b0;
    XRAM[12153] = 8'b0;
    XRAM[12154] = 8'b0;
    XRAM[12155] = 8'b0;
    XRAM[12156] = 8'b0;
    XRAM[12157] = 8'b0;
    XRAM[12158] = 8'b0;
    XRAM[12159] = 8'b0;
    XRAM[12160] = 8'b0;
    XRAM[12161] = 8'b0;
    XRAM[12162] = 8'b0;
    XRAM[12163] = 8'b0;
    XRAM[12164] = 8'b0;
    XRAM[12165] = 8'b0;
    XRAM[12166] = 8'b0;
    XRAM[12167] = 8'b0;
    XRAM[12168] = 8'b0;
    XRAM[12169] = 8'b0;
    XRAM[12170] = 8'b0;
    XRAM[12171] = 8'b0;
    XRAM[12172] = 8'b0;
    XRAM[12173] = 8'b0;
    XRAM[12174] = 8'b0;
    XRAM[12175] = 8'b0;
    XRAM[12176] = 8'b0;
    XRAM[12177] = 8'b0;
    XRAM[12178] = 8'b0;
    XRAM[12179] = 8'b0;
    XRAM[12180] = 8'b0;
    XRAM[12181] = 8'b0;
    XRAM[12182] = 8'b0;
    XRAM[12183] = 8'b0;
    XRAM[12184] = 8'b0;
    XRAM[12185] = 8'b0;
    XRAM[12186] = 8'b0;
    XRAM[12187] = 8'b0;
    XRAM[12188] = 8'b0;
    XRAM[12189] = 8'b0;
    XRAM[12190] = 8'b0;
    XRAM[12191] = 8'b0;
    XRAM[12192] = 8'b0;
    XRAM[12193] = 8'b0;
    XRAM[12194] = 8'b0;
    XRAM[12195] = 8'b0;
    XRAM[12196] = 8'b0;
    XRAM[12197] = 8'b0;
    XRAM[12198] = 8'b0;
    XRAM[12199] = 8'b0;
    XRAM[12200] = 8'b0;
    XRAM[12201] = 8'b0;
    XRAM[12202] = 8'b0;
    XRAM[12203] = 8'b0;
    XRAM[12204] = 8'b0;
    XRAM[12205] = 8'b0;
    XRAM[12206] = 8'b0;
    XRAM[12207] = 8'b0;
    XRAM[12208] = 8'b0;
    XRAM[12209] = 8'b0;
    XRAM[12210] = 8'b0;
    XRAM[12211] = 8'b0;
    XRAM[12212] = 8'b0;
    XRAM[12213] = 8'b0;
    XRAM[12214] = 8'b0;
    XRAM[12215] = 8'b0;
    XRAM[12216] = 8'b0;
    XRAM[12217] = 8'b0;
    XRAM[12218] = 8'b0;
    XRAM[12219] = 8'b0;
    XRAM[12220] = 8'b0;
    XRAM[12221] = 8'b0;
    XRAM[12222] = 8'b0;
    XRAM[12223] = 8'b0;
    XRAM[12224] = 8'b0;
    XRAM[12225] = 8'b0;
    XRAM[12226] = 8'b0;
    XRAM[12227] = 8'b0;
    XRAM[12228] = 8'b0;
    XRAM[12229] = 8'b0;
    XRAM[12230] = 8'b0;
    XRAM[12231] = 8'b0;
    XRAM[12232] = 8'b0;
    XRAM[12233] = 8'b0;
    XRAM[12234] = 8'b0;
    XRAM[12235] = 8'b0;
    XRAM[12236] = 8'b0;
    XRAM[12237] = 8'b0;
    XRAM[12238] = 8'b0;
    XRAM[12239] = 8'b0;
    XRAM[12240] = 8'b0;
    XRAM[12241] = 8'b0;
    XRAM[12242] = 8'b0;
    XRAM[12243] = 8'b0;
    XRAM[12244] = 8'b0;
    XRAM[12245] = 8'b0;
    XRAM[12246] = 8'b0;
    XRAM[12247] = 8'b0;
    XRAM[12248] = 8'b0;
    XRAM[12249] = 8'b0;
    XRAM[12250] = 8'b0;
    XRAM[12251] = 8'b0;
    XRAM[12252] = 8'b0;
    XRAM[12253] = 8'b0;
    XRAM[12254] = 8'b0;
    XRAM[12255] = 8'b0;
    XRAM[12256] = 8'b0;
    XRAM[12257] = 8'b0;
    XRAM[12258] = 8'b0;
    XRAM[12259] = 8'b0;
    XRAM[12260] = 8'b0;
    XRAM[12261] = 8'b0;
    XRAM[12262] = 8'b0;
    XRAM[12263] = 8'b0;
    XRAM[12264] = 8'b0;
    XRAM[12265] = 8'b0;
    XRAM[12266] = 8'b0;
    XRAM[12267] = 8'b0;
    XRAM[12268] = 8'b0;
    XRAM[12269] = 8'b0;
    XRAM[12270] = 8'b0;
    XRAM[12271] = 8'b0;
    XRAM[12272] = 8'b0;
    XRAM[12273] = 8'b0;
    XRAM[12274] = 8'b0;
    XRAM[12275] = 8'b0;
    XRAM[12276] = 8'b0;
    XRAM[12277] = 8'b0;
    XRAM[12278] = 8'b0;
    XRAM[12279] = 8'b0;
    XRAM[12280] = 8'b0;
    XRAM[12281] = 8'b0;
    XRAM[12282] = 8'b0;
    XRAM[12283] = 8'b0;
    XRAM[12284] = 8'b0;
    XRAM[12285] = 8'b0;
    XRAM[12286] = 8'b0;
    XRAM[12287] = 8'b0;
    XRAM[12288] = 8'b0;
    XRAM[12289] = 8'b0;
    XRAM[12290] = 8'b0;
    XRAM[12291] = 8'b0;
    XRAM[12292] = 8'b0;
    XRAM[12293] = 8'b0;
    XRAM[12294] = 8'b0;
    XRAM[12295] = 8'b0;
    XRAM[12296] = 8'b0;
    XRAM[12297] = 8'b0;
    XRAM[12298] = 8'b0;
    XRAM[12299] = 8'b0;
    XRAM[12300] = 8'b0;
    XRAM[12301] = 8'b0;
    XRAM[12302] = 8'b0;
    XRAM[12303] = 8'b0;
    XRAM[12304] = 8'b0;
    XRAM[12305] = 8'b0;
    XRAM[12306] = 8'b0;
    XRAM[12307] = 8'b0;
    XRAM[12308] = 8'b0;
    XRAM[12309] = 8'b0;
    XRAM[12310] = 8'b0;
    XRAM[12311] = 8'b0;
    XRAM[12312] = 8'b0;
    XRAM[12313] = 8'b0;
    XRAM[12314] = 8'b0;
    XRAM[12315] = 8'b0;
    XRAM[12316] = 8'b0;
    XRAM[12317] = 8'b0;
    XRAM[12318] = 8'b0;
    XRAM[12319] = 8'b0;
    XRAM[12320] = 8'b0;
    XRAM[12321] = 8'b0;
    XRAM[12322] = 8'b0;
    XRAM[12323] = 8'b0;
    XRAM[12324] = 8'b0;
    XRAM[12325] = 8'b0;
    XRAM[12326] = 8'b0;
    XRAM[12327] = 8'b0;
    XRAM[12328] = 8'b0;
    XRAM[12329] = 8'b0;
    XRAM[12330] = 8'b0;
    XRAM[12331] = 8'b0;
    XRAM[12332] = 8'b0;
    XRAM[12333] = 8'b0;
    XRAM[12334] = 8'b0;
    XRAM[12335] = 8'b0;
    XRAM[12336] = 8'b0;
    XRAM[12337] = 8'b0;
    XRAM[12338] = 8'b0;
    XRAM[12339] = 8'b0;
    XRAM[12340] = 8'b0;
    XRAM[12341] = 8'b0;
    XRAM[12342] = 8'b0;
    XRAM[12343] = 8'b0;
    XRAM[12344] = 8'b0;
    XRAM[12345] = 8'b0;
    XRAM[12346] = 8'b0;
    XRAM[12347] = 8'b0;
    XRAM[12348] = 8'b0;
    XRAM[12349] = 8'b0;
    XRAM[12350] = 8'b0;
    XRAM[12351] = 8'b0;
    XRAM[12352] = 8'b0;
    XRAM[12353] = 8'b0;
    XRAM[12354] = 8'b0;
    XRAM[12355] = 8'b0;
    XRAM[12356] = 8'b0;
    XRAM[12357] = 8'b0;
    XRAM[12358] = 8'b0;
    XRAM[12359] = 8'b0;
    XRAM[12360] = 8'b0;
    XRAM[12361] = 8'b0;
    XRAM[12362] = 8'b0;
    XRAM[12363] = 8'b0;
    XRAM[12364] = 8'b0;
    XRAM[12365] = 8'b0;
    XRAM[12366] = 8'b0;
    XRAM[12367] = 8'b0;
    XRAM[12368] = 8'b0;
    XRAM[12369] = 8'b0;
    XRAM[12370] = 8'b0;
    XRAM[12371] = 8'b0;
    XRAM[12372] = 8'b0;
    XRAM[12373] = 8'b0;
    XRAM[12374] = 8'b0;
    XRAM[12375] = 8'b0;
    XRAM[12376] = 8'b0;
    XRAM[12377] = 8'b0;
    XRAM[12378] = 8'b0;
    XRAM[12379] = 8'b0;
    XRAM[12380] = 8'b0;
    XRAM[12381] = 8'b0;
    XRAM[12382] = 8'b0;
    XRAM[12383] = 8'b0;
    XRAM[12384] = 8'b0;
    XRAM[12385] = 8'b0;
    XRAM[12386] = 8'b0;
    XRAM[12387] = 8'b0;
    XRAM[12388] = 8'b0;
    XRAM[12389] = 8'b0;
    XRAM[12390] = 8'b0;
    XRAM[12391] = 8'b0;
    XRAM[12392] = 8'b0;
    XRAM[12393] = 8'b0;
    XRAM[12394] = 8'b0;
    XRAM[12395] = 8'b0;
    XRAM[12396] = 8'b0;
    XRAM[12397] = 8'b0;
    XRAM[12398] = 8'b0;
    XRAM[12399] = 8'b0;
    XRAM[12400] = 8'b0;
    XRAM[12401] = 8'b0;
    XRAM[12402] = 8'b0;
    XRAM[12403] = 8'b0;
    XRAM[12404] = 8'b0;
    XRAM[12405] = 8'b0;
    XRAM[12406] = 8'b0;
    XRAM[12407] = 8'b0;
    XRAM[12408] = 8'b0;
    XRAM[12409] = 8'b0;
    XRAM[12410] = 8'b0;
    XRAM[12411] = 8'b0;
    XRAM[12412] = 8'b0;
    XRAM[12413] = 8'b0;
    XRAM[12414] = 8'b0;
    XRAM[12415] = 8'b0;
    XRAM[12416] = 8'b0;
    XRAM[12417] = 8'b0;
    XRAM[12418] = 8'b0;
    XRAM[12419] = 8'b0;
    XRAM[12420] = 8'b0;
    XRAM[12421] = 8'b0;
    XRAM[12422] = 8'b0;
    XRAM[12423] = 8'b0;
    XRAM[12424] = 8'b0;
    XRAM[12425] = 8'b0;
    XRAM[12426] = 8'b0;
    XRAM[12427] = 8'b0;
    XRAM[12428] = 8'b0;
    XRAM[12429] = 8'b0;
    XRAM[12430] = 8'b0;
    XRAM[12431] = 8'b0;
    XRAM[12432] = 8'b0;
    XRAM[12433] = 8'b0;
    XRAM[12434] = 8'b0;
    XRAM[12435] = 8'b0;
    XRAM[12436] = 8'b0;
    XRAM[12437] = 8'b0;
    XRAM[12438] = 8'b0;
    XRAM[12439] = 8'b0;
    XRAM[12440] = 8'b0;
    XRAM[12441] = 8'b0;
    XRAM[12442] = 8'b0;
    XRAM[12443] = 8'b0;
    XRAM[12444] = 8'b0;
    XRAM[12445] = 8'b0;
    XRAM[12446] = 8'b0;
    XRAM[12447] = 8'b0;
    XRAM[12448] = 8'b0;
    XRAM[12449] = 8'b0;
    XRAM[12450] = 8'b0;
    XRAM[12451] = 8'b0;
    XRAM[12452] = 8'b0;
    XRAM[12453] = 8'b0;
    XRAM[12454] = 8'b0;
    XRAM[12455] = 8'b0;
    XRAM[12456] = 8'b0;
    XRAM[12457] = 8'b0;
    XRAM[12458] = 8'b0;
    XRAM[12459] = 8'b0;
    XRAM[12460] = 8'b0;
    XRAM[12461] = 8'b0;
    XRAM[12462] = 8'b0;
    XRAM[12463] = 8'b0;
    XRAM[12464] = 8'b0;
    XRAM[12465] = 8'b0;
    XRAM[12466] = 8'b0;
    XRAM[12467] = 8'b0;
    XRAM[12468] = 8'b0;
    XRAM[12469] = 8'b0;
    XRAM[12470] = 8'b0;
    XRAM[12471] = 8'b0;
    XRAM[12472] = 8'b0;
    XRAM[12473] = 8'b0;
    XRAM[12474] = 8'b0;
    XRAM[12475] = 8'b0;
    XRAM[12476] = 8'b0;
    XRAM[12477] = 8'b0;
    XRAM[12478] = 8'b0;
    XRAM[12479] = 8'b0;
    XRAM[12480] = 8'b0;
    XRAM[12481] = 8'b0;
    XRAM[12482] = 8'b0;
    XRAM[12483] = 8'b0;
    XRAM[12484] = 8'b0;
    XRAM[12485] = 8'b0;
    XRAM[12486] = 8'b0;
    XRAM[12487] = 8'b0;
    XRAM[12488] = 8'b0;
    XRAM[12489] = 8'b0;
    XRAM[12490] = 8'b0;
    XRAM[12491] = 8'b0;
    XRAM[12492] = 8'b0;
    XRAM[12493] = 8'b0;
    XRAM[12494] = 8'b0;
    XRAM[12495] = 8'b0;
    XRAM[12496] = 8'b0;
    XRAM[12497] = 8'b0;
    XRAM[12498] = 8'b0;
    XRAM[12499] = 8'b0;
    XRAM[12500] = 8'b0;
    XRAM[12501] = 8'b0;
    XRAM[12502] = 8'b0;
    XRAM[12503] = 8'b0;
    XRAM[12504] = 8'b0;
    XRAM[12505] = 8'b0;
    XRAM[12506] = 8'b0;
    XRAM[12507] = 8'b0;
    XRAM[12508] = 8'b0;
    XRAM[12509] = 8'b0;
    XRAM[12510] = 8'b0;
    XRAM[12511] = 8'b0;
    XRAM[12512] = 8'b0;
    XRAM[12513] = 8'b0;
    XRAM[12514] = 8'b0;
    XRAM[12515] = 8'b0;
    XRAM[12516] = 8'b0;
    XRAM[12517] = 8'b0;
    XRAM[12518] = 8'b0;
    XRAM[12519] = 8'b0;
    XRAM[12520] = 8'b0;
    XRAM[12521] = 8'b0;
    XRAM[12522] = 8'b0;
    XRAM[12523] = 8'b0;
    XRAM[12524] = 8'b0;
    XRAM[12525] = 8'b0;
    XRAM[12526] = 8'b0;
    XRAM[12527] = 8'b0;
    XRAM[12528] = 8'b0;
    XRAM[12529] = 8'b0;
    XRAM[12530] = 8'b0;
    XRAM[12531] = 8'b0;
    XRAM[12532] = 8'b0;
    XRAM[12533] = 8'b0;
    XRAM[12534] = 8'b0;
    XRAM[12535] = 8'b0;
    XRAM[12536] = 8'b0;
    XRAM[12537] = 8'b0;
    XRAM[12538] = 8'b0;
    XRAM[12539] = 8'b0;
    XRAM[12540] = 8'b0;
    XRAM[12541] = 8'b0;
    XRAM[12542] = 8'b0;
    XRAM[12543] = 8'b0;
    XRAM[12544] = 8'b0;
    XRAM[12545] = 8'b0;
    XRAM[12546] = 8'b0;
    XRAM[12547] = 8'b0;
    XRAM[12548] = 8'b0;
    XRAM[12549] = 8'b0;
    XRAM[12550] = 8'b0;
    XRAM[12551] = 8'b0;
    XRAM[12552] = 8'b0;
    XRAM[12553] = 8'b0;
    XRAM[12554] = 8'b0;
    XRAM[12555] = 8'b0;
    XRAM[12556] = 8'b0;
    XRAM[12557] = 8'b0;
    XRAM[12558] = 8'b0;
    XRAM[12559] = 8'b0;
    XRAM[12560] = 8'b0;
    XRAM[12561] = 8'b0;
    XRAM[12562] = 8'b0;
    XRAM[12563] = 8'b0;
    XRAM[12564] = 8'b0;
    XRAM[12565] = 8'b0;
    XRAM[12566] = 8'b0;
    XRAM[12567] = 8'b0;
    XRAM[12568] = 8'b0;
    XRAM[12569] = 8'b0;
    XRAM[12570] = 8'b0;
    XRAM[12571] = 8'b0;
    XRAM[12572] = 8'b0;
    XRAM[12573] = 8'b0;
    XRAM[12574] = 8'b0;
    XRAM[12575] = 8'b0;
    XRAM[12576] = 8'b0;
    XRAM[12577] = 8'b0;
    XRAM[12578] = 8'b0;
    XRAM[12579] = 8'b0;
    XRAM[12580] = 8'b0;
    XRAM[12581] = 8'b0;
    XRAM[12582] = 8'b0;
    XRAM[12583] = 8'b0;
    XRAM[12584] = 8'b0;
    XRAM[12585] = 8'b0;
    XRAM[12586] = 8'b0;
    XRAM[12587] = 8'b0;
    XRAM[12588] = 8'b0;
    XRAM[12589] = 8'b0;
    XRAM[12590] = 8'b0;
    XRAM[12591] = 8'b0;
    XRAM[12592] = 8'b0;
    XRAM[12593] = 8'b0;
    XRAM[12594] = 8'b0;
    XRAM[12595] = 8'b0;
    XRAM[12596] = 8'b0;
    XRAM[12597] = 8'b0;
    XRAM[12598] = 8'b0;
    XRAM[12599] = 8'b0;
    XRAM[12600] = 8'b0;
    XRAM[12601] = 8'b0;
    XRAM[12602] = 8'b0;
    XRAM[12603] = 8'b0;
    XRAM[12604] = 8'b0;
    XRAM[12605] = 8'b0;
    XRAM[12606] = 8'b0;
    XRAM[12607] = 8'b0;
    XRAM[12608] = 8'b0;
    XRAM[12609] = 8'b0;
    XRAM[12610] = 8'b0;
    XRAM[12611] = 8'b0;
    XRAM[12612] = 8'b0;
    XRAM[12613] = 8'b0;
    XRAM[12614] = 8'b0;
    XRAM[12615] = 8'b0;
    XRAM[12616] = 8'b0;
    XRAM[12617] = 8'b0;
    XRAM[12618] = 8'b0;
    XRAM[12619] = 8'b0;
    XRAM[12620] = 8'b0;
    XRAM[12621] = 8'b0;
    XRAM[12622] = 8'b0;
    XRAM[12623] = 8'b0;
    XRAM[12624] = 8'b0;
    XRAM[12625] = 8'b0;
    XRAM[12626] = 8'b0;
    XRAM[12627] = 8'b0;
    XRAM[12628] = 8'b0;
    XRAM[12629] = 8'b0;
    XRAM[12630] = 8'b0;
    XRAM[12631] = 8'b0;
    XRAM[12632] = 8'b0;
    XRAM[12633] = 8'b0;
    XRAM[12634] = 8'b0;
    XRAM[12635] = 8'b0;
    XRAM[12636] = 8'b0;
    XRAM[12637] = 8'b0;
    XRAM[12638] = 8'b0;
    XRAM[12639] = 8'b0;
    XRAM[12640] = 8'b0;
    XRAM[12641] = 8'b0;
    XRAM[12642] = 8'b0;
    XRAM[12643] = 8'b0;
    XRAM[12644] = 8'b0;
    XRAM[12645] = 8'b0;
    XRAM[12646] = 8'b0;
    XRAM[12647] = 8'b0;
    XRAM[12648] = 8'b0;
    XRAM[12649] = 8'b0;
    XRAM[12650] = 8'b0;
    XRAM[12651] = 8'b0;
    XRAM[12652] = 8'b0;
    XRAM[12653] = 8'b0;
    XRAM[12654] = 8'b0;
    XRAM[12655] = 8'b0;
    XRAM[12656] = 8'b0;
    XRAM[12657] = 8'b0;
    XRAM[12658] = 8'b0;
    XRAM[12659] = 8'b0;
    XRAM[12660] = 8'b0;
    XRAM[12661] = 8'b0;
    XRAM[12662] = 8'b0;
    XRAM[12663] = 8'b0;
    XRAM[12664] = 8'b0;
    XRAM[12665] = 8'b0;
    XRAM[12666] = 8'b0;
    XRAM[12667] = 8'b0;
    XRAM[12668] = 8'b0;
    XRAM[12669] = 8'b0;
    XRAM[12670] = 8'b0;
    XRAM[12671] = 8'b0;
    XRAM[12672] = 8'b0;
    XRAM[12673] = 8'b0;
    XRAM[12674] = 8'b0;
    XRAM[12675] = 8'b0;
    XRAM[12676] = 8'b0;
    XRAM[12677] = 8'b0;
    XRAM[12678] = 8'b0;
    XRAM[12679] = 8'b0;
    XRAM[12680] = 8'b0;
    XRAM[12681] = 8'b0;
    XRAM[12682] = 8'b0;
    XRAM[12683] = 8'b0;
    XRAM[12684] = 8'b0;
    XRAM[12685] = 8'b0;
    XRAM[12686] = 8'b0;
    XRAM[12687] = 8'b0;
    XRAM[12688] = 8'b0;
    XRAM[12689] = 8'b0;
    XRAM[12690] = 8'b0;
    XRAM[12691] = 8'b0;
    XRAM[12692] = 8'b0;
    XRAM[12693] = 8'b0;
    XRAM[12694] = 8'b0;
    XRAM[12695] = 8'b0;
    XRAM[12696] = 8'b0;
    XRAM[12697] = 8'b0;
    XRAM[12698] = 8'b0;
    XRAM[12699] = 8'b0;
    XRAM[12700] = 8'b0;
    XRAM[12701] = 8'b0;
    XRAM[12702] = 8'b0;
    XRAM[12703] = 8'b0;
    XRAM[12704] = 8'b0;
    XRAM[12705] = 8'b0;
    XRAM[12706] = 8'b0;
    XRAM[12707] = 8'b0;
    XRAM[12708] = 8'b0;
    XRAM[12709] = 8'b0;
    XRAM[12710] = 8'b0;
    XRAM[12711] = 8'b0;
    XRAM[12712] = 8'b0;
    XRAM[12713] = 8'b0;
    XRAM[12714] = 8'b0;
    XRAM[12715] = 8'b0;
    XRAM[12716] = 8'b0;
    XRAM[12717] = 8'b0;
    XRAM[12718] = 8'b0;
    XRAM[12719] = 8'b0;
    XRAM[12720] = 8'b0;
    XRAM[12721] = 8'b0;
    XRAM[12722] = 8'b0;
    XRAM[12723] = 8'b0;
    XRAM[12724] = 8'b0;
    XRAM[12725] = 8'b0;
    XRAM[12726] = 8'b0;
    XRAM[12727] = 8'b0;
    XRAM[12728] = 8'b0;
    XRAM[12729] = 8'b0;
    XRAM[12730] = 8'b0;
    XRAM[12731] = 8'b0;
    XRAM[12732] = 8'b0;
    XRAM[12733] = 8'b0;
    XRAM[12734] = 8'b0;
    XRAM[12735] = 8'b0;
    XRAM[12736] = 8'b0;
    XRAM[12737] = 8'b0;
    XRAM[12738] = 8'b0;
    XRAM[12739] = 8'b0;
    XRAM[12740] = 8'b0;
    XRAM[12741] = 8'b0;
    XRAM[12742] = 8'b0;
    XRAM[12743] = 8'b0;
    XRAM[12744] = 8'b0;
    XRAM[12745] = 8'b0;
    XRAM[12746] = 8'b0;
    XRAM[12747] = 8'b0;
    XRAM[12748] = 8'b0;
    XRAM[12749] = 8'b0;
    XRAM[12750] = 8'b0;
    XRAM[12751] = 8'b0;
    XRAM[12752] = 8'b0;
    XRAM[12753] = 8'b0;
    XRAM[12754] = 8'b0;
    XRAM[12755] = 8'b0;
    XRAM[12756] = 8'b0;
    XRAM[12757] = 8'b0;
    XRAM[12758] = 8'b0;
    XRAM[12759] = 8'b0;
    XRAM[12760] = 8'b0;
    XRAM[12761] = 8'b0;
    XRAM[12762] = 8'b0;
    XRAM[12763] = 8'b0;
    XRAM[12764] = 8'b0;
    XRAM[12765] = 8'b0;
    XRAM[12766] = 8'b0;
    XRAM[12767] = 8'b0;
    XRAM[12768] = 8'b0;
    XRAM[12769] = 8'b0;
    XRAM[12770] = 8'b0;
    XRAM[12771] = 8'b0;
    XRAM[12772] = 8'b0;
    XRAM[12773] = 8'b0;
    XRAM[12774] = 8'b0;
    XRAM[12775] = 8'b0;
    XRAM[12776] = 8'b0;
    XRAM[12777] = 8'b0;
    XRAM[12778] = 8'b0;
    XRAM[12779] = 8'b0;
    XRAM[12780] = 8'b0;
    XRAM[12781] = 8'b0;
    XRAM[12782] = 8'b0;
    XRAM[12783] = 8'b0;
    XRAM[12784] = 8'b0;
    XRAM[12785] = 8'b0;
    XRAM[12786] = 8'b0;
    XRAM[12787] = 8'b0;
    XRAM[12788] = 8'b0;
    XRAM[12789] = 8'b0;
    XRAM[12790] = 8'b0;
    XRAM[12791] = 8'b0;
    XRAM[12792] = 8'b0;
    XRAM[12793] = 8'b0;
    XRAM[12794] = 8'b0;
    XRAM[12795] = 8'b0;
    XRAM[12796] = 8'b0;
    XRAM[12797] = 8'b0;
    XRAM[12798] = 8'b0;
    XRAM[12799] = 8'b0;
    XRAM[12800] = 8'b0;
    XRAM[12801] = 8'b0;
    XRAM[12802] = 8'b0;
    XRAM[12803] = 8'b0;
    XRAM[12804] = 8'b0;
    XRAM[12805] = 8'b0;
    XRAM[12806] = 8'b0;
    XRAM[12807] = 8'b0;
    XRAM[12808] = 8'b0;
    XRAM[12809] = 8'b0;
    XRAM[12810] = 8'b0;
    XRAM[12811] = 8'b0;
    XRAM[12812] = 8'b0;
    XRAM[12813] = 8'b0;
    XRAM[12814] = 8'b0;
    XRAM[12815] = 8'b0;
    XRAM[12816] = 8'b0;
    XRAM[12817] = 8'b0;
    XRAM[12818] = 8'b0;
    XRAM[12819] = 8'b0;
    XRAM[12820] = 8'b0;
    XRAM[12821] = 8'b0;
    XRAM[12822] = 8'b0;
    XRAM[12823] = 8'b0;
    XRAM[12824] = 8'b0;
    XRAM[12825] = 8'b0;
    XRAM[12826] = 8'b0;
    XRAM[12827] = 8'b0;
    XRAM[12828] = 8'b0;
    XRAM[12829] = 8'b0;
    XRAM[12830] = 8'b0;
    XRAM[12831] = 8'b0;
    XRAM[12832] = 8'b0;
    XRAM[12833] = 8'b0;
    XRAM[12834] = 8'b0;
    XRAM[12835] = 8'b0;
    XRAM[12836] = 8'b0;
    XRAM[12837] = 8'b0;
    XRAM[12838] = 8'b0;
    XRAM[12839] = 8'b0;
    XRAM[12840] = 8'b0;
    XRAM[12841] = 8'b0;
    XRAM[12842] = 8'b0;
    XRAM[12843] = 8'b0;
    XRAM[12844] = 8'b0;
    XRAM[12845] = 8'b0;
    XRAM[12846] = 8'b0;
    XRAM[12847] = 8'b0;
    XRAM[12848] = 8'b0;
    XRAM[12849] = 8'b0;
    XRAM[12850] = 8'b0;
    XRAM[12851] = 8'b0;
    XRAM[12852] = 8'b0;
    XRAM[12853] = 8'b0;
    XRAM[12854] = 8'b0;
    XRAM[12855] = 8'b0;
    XRAM[12856] = 8'b0;
    XRAM[12857] = 8'b0;
    XRAM[12858] = 8'b0;
    XRAM[12859] = 8'b0;
    XRAM[12860] = 8'b0;
    XRAM[12861] = 8'b0;
    XRAM[12862] = 8'b0;
    XRAM[12863] = 8'b0;
    XRAM[12864] = 8'b0;
    XRAM[12865] = 8'b0;
    XRAM[12866] = 8'b0;
    XRAM[12867] = 8'b0;
    XRAM[12868] = 8'b0;
    XRAM[12869] = 8'b0;
    XRAM[12870] = 8'b0;
    XRAM[12871] = 8'b0;
    XRAM[12872] = 8'b0;
    XRAM[12873] = 8'b0;
    XRAM[12874] = 8'b0;
    XRAM[12875] = 8'b0;
    XRAM[12876] = 8'b0;
    XRAM[12877] = 8'b0;
    XRAM[12878] = 8'b0;
    XRAM[12879] = 8'b0;
    XRAM[12880] = 8'b0;
    XRAM[12881] = 8'b0;
    XRAM[12882] = 8'b0;
    XRAM[12883] = 8'b0;
    XRAM[12884] = 8'b0;
    XRAM[12885] = 8'b0;
    XRAM[12886] = 8'b0;
    XRAM[12887] = 8'b0;
    XRAM[12888] = 8'b0;
    XRAM[12889] = 8'b0;
    XRAM[12890] = 8'b0;
    XRAM[12891] = 8'b0;
    XRAM[12892] = 8'b0;
    XRAM[12893] = 8'b0;
    XRAM[12894] = 8'b0;
    XRAM[12895] = 8'b0;
    XRAM[12896] = 8'b0;
    XRAM[12897] = 8'b0;
    XRAM[12898] = 8'b0;
    XRAM[12899] = 8'b0;
    XRAM[12900] = 8'b0;
    XRAM[12901] = 8'b0;
    XRAM[12902] = 8'b0;
    XRAM[12903] = 8'b0;
    XRAM[12904] = 8'b0;
    XRAM[12905] = 8'b0;
    XRAM[12906] = 8'b0;
    XRAM[12907] = 8'b0;
    XRAM[12908] = 8'b0;
    XRAM[12909] = 8'b0;
    XRAM[12910] = 8'b0;
    XRAM[12911] = 8'b0;
    XRAM[12912] = 8'b0;
    XRAM[12913] = 8'b0;
    XRAM[12914] = 8'b0;
    XRAM[12915] = 8'b0;
    XRAM[12916] = 8'b0;
    XRAM[12917] = 8'b0;
    XRAM[12918] = 8'b0;
    XRAM[12919] = 8'b0;
    XRAM[12920] = 8'b0;
    XRAM[12921] = 8'b0;
    XRAM[12922] = 8'b0;
    XRAM[12923] = 8'b0;
    XRAM[12924] = 8'b0;
    XRAM[12925] = 8'b0;
    XRAM[12926] = 8'b0;
    XRAM[12927] = 8'b0;
    XRAM[12928] = 8'b0;
    XRAM[12929] = 8'b0;
    XRAM[12930] = 8'b0;
    XRAM[12931] = 8'b0;
    XRAM[12932] = 8'b0;
    XRAM[12933] = 8'b0;
    XRAM[12934] = 8'b0;
    XRAM[12935] = 8'b0;
    XRAM[12936] = 8'b0;
    XRAM[12937] = 8'b0;
    XRAM[12938] = 8'b0;
    XRAM[12939] = 8'b0;
    XRAM[12940] = 8'b0;
    XRAM[12941] = 8'b0;
    XRAM[12942] = 8'b0;
    XRAM[12943] = 8'b0;
    XRAM[12944] = 8'b0;
    XRAM[12945] = 8'b0;
    XRAM[12946] = 8'b0;
    XRAM[12947] = 8'b0;
    XRAM[12948] = 8'b0;
    XRAM[12949] = 8'b0;
    XRAM[12950] = 8'b0;
    XRAM[12951] = 8'b0;
    XRAM[12952] = 8'b0;
    XRAM[12953] = 8'b0;
    XRAM[12954] = 8'b0;
    XRAM[12955] = 8'b0;
    XRAM[12956] = 8'b0;
    XRAM[12957] = 8'b0;
    XRAM[12958] = 8'b0;
    XRAM[12959] = 8'b0;
    XRAM[12960] = 8'b0;
    XRAM[12961] = 8'b0;
    XRAM[12962] = 8'b0;
    XRAM[12963] = 8'b0;
    XRAM[12964] = 8'b0;
    XRAM[12965] = 8'b0;
    XRAM[12966] = 8'b0;
    XRAM[12967] = 8'b0;
    XRAM[12968] = 8'b0;
    XRAM[12969] = 8'b0;
    XRAM[12970] = 8'b0;
    XRAM[12971] = 8'b0;
    XRAM[12972] = 8'b0;
    XRAM[12973] = 8'b0;
    XRAM[12974] = 8'b0;
    XRAM[12975] = 8'b0;
    XRAM[12976] = 8'b0;
    XRAM[12977] = 8'b0;
    XRAM[12978] = 8'b0;
    XRAM[12979] = 8'b0;
    XRAM[12980] = 8'b0;
    XRAM[12981] = 8'b0;
    XRAM[12982] = 8'b0;
    XRAM[12983] = 8'b0;
    XRAM[12984] = 8'b0;
    XRAM[12985] = 8'b0;
    XRAM[12986] = 8'b0;
    XRAM[12987] = 8'b0;
    XRAM[12988] = 8'b0;
    XRAM[12989] = 8'b0;
    XRAM[12990] = 8'b0;
    XRAM[12991] = 8'b0;
    XRAM[12992] = 8'b0;
    XRAM[12993] = 8'b0;
    XRAM[12994] = 8'b0;
    XRAM[12995] = 8'b0;
    XRAM[12996] = 8'b0;
    XRAM[12997] = 8'b0;
    XRAM[12998] = 8'b0;
    XRAM[12999] = 8'b0;
    XRAM[13000] = 8'b0;
    XRAM[13001] = 8'b0;
    XRAM[13002] = 8'b0;
    XRAM[13003] = 8'b0;
    XRAM[13004] = 8'b0;
    XRAM[13005] = 8'b0;
    XRAM[13006] = 8'b0;
    XRAM[13007] = 8'b0;
    XRAM[13008] = 8'b0;
    XRAM[13009] = 8'b0;
    XRAM[13010] = 8'b0;
    XRAM[13011] = 8'b0;
    XRAM[13012] = 8'b0;
    XRAM[13013] = 8'b0;
    XRAM[13014] = 8'b0;
    XRAM[13015] = 8'b0;
    XRAM[13016] = 8'b0;
    XRAM[13017] = 8'b0;
    XRAM[13018] = 8'b0;
    XRAM[13019] = 8'b0;
    XRAM[13020] = 8'b0;
    XRAM[13021] = 8'b0;
    XRAM[13022] = 8'b0;
    XRAM[13023] = 8'b0;
    XRAM[13024] = 8'b0;
    XRAM[13025] = 8'b0;
    XRAM[13026] = 8'b0;
    XRAM[13027] = 8'b0;
    XRAM[13028] = 8'b0;
    XRAM[13029] = 8'b0;
    XRAM[13030] = 8'b0;
    XRAM[13031] = 8'b0;
    XRAM[13032] = 8'b0;
    XRAM[13033] = 8'b0;
    XRAM[13034] = 8'b0;
    XRAM[13035] = 8'b0;
    XRAM[13036] = 8'b0;
    XRAM[13037] = 8'b0;
    XRAM[13038] = 8'b0;
    XRAM[13039] = 8'b0;
    XRAM[13040] = 8'b0;
    XRAM[13041] = 8'b0;
    XRAM[13042] = 8'b0;
    XRAM[13043] = 8'b0;
    XRAM[13044] = 8'b0;
    XRAM[13045] = 8'b0;
    XRAM[13046] = 8'b0;
    XRAM[13047] = 8'b0;
    XRAM[13048] = 8'b0;
    XRAM[13049] = 8'b0;
    XRAM[13050] = 8'b0;
    XRAM[13051] = 8'b0;
    XRAM[13052] = 8'b0;
    XRAM[13053] = 8'b0;
    XRAM[13054] = 8'b0;
    XRAM[13055] = 8'b0;
    XRAM[13056] = 8'b0;
    XRAM[13057] = 8'b0;
    XRAM[13058] = 8'b0;
    XRAM[13059] = 8'b0;
    XRAM[13060] = 8'b0;
    XRAM[13061] = 8'b0;
    XRAM[13062] = 8'b0;
    XRAM[13063] = 8'b0;
    XRAM[13064] = 8'b0;
    XRAM[13065] = 8'b0;
    XRAM[13066] = 8'b0;
    XRAM[13067] = 8'b0;
    XRAM[13068] = 8'b0;
    XRAM[13069] = 8'b0;
    XRAM[13070] = 8'b0;
    XRAM[13071] = 8'b0;
    XRAM[13072] = 8'b0;
    XRAM[13073] = 8'b0;
    XRAM[13074] = 8'b0;
    XRAM[13075] = 8'b0;
    XRAM[13076] = 8'b0;
    XRAM[13077] = 8'b0;
    XRAM[13078] = 8'b0;
    XRAM[13079] = 8'b0;
    XRAM[13080] = 8'b0;
    XRAM[13081] = 8'b0;
    XRAM[13082] = 8'b0;
    XRAM[13083] = 8'b0;
    XRAM[13084] = 8'b0;
    XRAM[13085] = 8'b0;
    XRAM[13086] = 8'b0;
    XRAM[13087] = 8'b0;
    XRAM[13088] = 8'b0;
    XRAM[13089] = 8'b0;
    XRAM[13090] = 8'b0;
    XRAM[13091] = 8'b0;
    XRAM[13092] = 8'b0;
    XRAM[13093] = 8'b0;
    XRAM[13094] = 8'b0;
    XRAM[13095] = 8'b0;
    XRAM[13096] = 8'b0;
    XRAM[13097] = 8'b0;
    XRAM[13098] = 8'b0;
    XRAM[13099] = 8'b0;
    XRAM[13100] = 8'b0;
    XRAM[13101] = 8'b0;
    XRAM[13102] = 8'b0;
    XRAM[13103] = 8'b0;
    XRAM[13104] = 8'b0;
    XRAM[13105] = 8'b0;
    XRAM[13106] = 8'b0;
    XRAM[13107] = 8'b0;
    XRAM[13108] = 8'b0;
    XRAM[13109] = 8'b0;
    XRAM[13110] = 8'b0;
    XRAM[13111] = 8'b0;
    XRAM[13112] = 8'b0;
    XRAM[13113] = 8'b0;
    XRAM[13114] = 8'b0;
    XRAM[13115] = 8'b0;
    XRAM[13116] = 8'b0;
    XRAM[13117] = 8'b0;
    XRAM[13118] = 8'b0;
    XRAM[13119] = 8'b0;
    XRAM[13120] = 8'b0;
    XRAM[13121] = 8'b0;
    XRAM[13122] = 8'b0;
    XRAM[13123] = 8'b0;
    XRAM[13124] = 8'b0;
    XRAM[13125] = 8'b0;
    XRAM[13126] = 8'b0;
    XRAM[13127] = 8'b0;
    XRAM[13128] = 8'b0;
    XRAM[13129] = 8'b0;
    XRAM[13130] = 8'b0;
    XRAM[13131] = 8'b0;
    XRAM[13132] = 8'b0;
    XRAM[13133] = 8'b0;
    XRAM[13134] = 8'b0;
    XRAM[13135] = 8'b0;
    XRAM[13136] = 8'b0;
    XRAM[13137] = 8'b0;
    XRAM[13138] = 8'b0;
    XRAM[13139] = 8'b0;
    XRAM[13140] = 8'b0;
    XRAM[13141] = 8'b0;
    XRAM[13142] = 8'b0;
    XRAM[13143] = 8'b0;
    XRAM[13144] = 8'b0;
    XRAM[13145] = 8'b0;
    XRAM[13146] = 8'b0;
    XRAM[13147] = 8'b0;
    XRAM[13148] = 8'b0;
    XRAM[13149] = 8'b0;
    XRAM[13150] = 8'b0;
    XRAM[13151] = 8'b0;
    XRAM[13152] = 8'b0;
    XRAM[13153] = 8'b0;
    XRAM[13154] = 8'b0;
    XRAM[13155] = 8'b0;
    XRAM[13156] = 8'b0;
    XRAM[13157] = 8'b0;
    XRAM[13158] = 8'b0;
    XRAM[13159] = 8'b0;
    XRAM[13160] = 8'b0;
    XRAM[13161] = 8'b0;
    XRAM[13162] = 8'b0;
    XRAM[13163] = 8'b0;
    XRAM[13164] = 8'b0;
    XRAM[13165] = 8'b0;
    XRAM[13166] = 8'b0;
    XRAM[13167] = 8'b0;
    XRAM[13168] = 8'b0;
    XRAM[13169] = 8'b0;
    XRAM[13170] = 8'b0;
    XRAM[13171] = 8'b0;
    XRAM[13172] = 8'b0;
    XRAM[13173] = 8'b0;
    XRAM[13174] = 8'b0;
    XRAM[13175] = 8'b0;
    XRAM[13176] = 8'b0;
    XRAM[13177] = 8'b0;
    XRAM[13178] = 8'b0;
    XRAM[13179] = 8'b0;
    XRAM[13180] = 8'b0;
    XRAM[13181] = 8'b0;
    XRAM[13182] = 8'b0;
    XRAM[13183] = 8'b0;
    XRAM[13184] = 8'b0;
    XRAM[13185] = 8'b0;
    XRAM[13186] = 8'b0;
    XRAM[13187] = 8'b0;
    XRAM[13188] = 8'b0;
    XRAM[13189] = 8'b0;
    XRAM[13190] = 8'b0;
    XRAM[13191] = 8'b0;
    XRAM[13192] = 8'b0;
    XRAM[13193] = 8'b0;
    XRAM[13194] = 8'b0;
    XRAM[13195] = 8'b0;
    XRAM[13196] = 8'b0;
    XRAM[13197] = 8'b0;
    XRAM[13198] = 8'b0;
    XRAM[13199] = 8'b0;
    XRAM[13200] = 8'b0;
    XRAM[13201] = 8'b0;
    XRAM[13202] = 8'b0;
    XRAM[13203] = 8'b0;
    XRAM[13204] = 8'b0;
    XRAM[13205] = 8'b0;
    XRAM[13206] = 8'b0;
    XRAM[13207] = 8'b0;
    XRAM[13208] = 8'b0;
    XRAM[13209] = 8'b0;
    XRAM[13210] = 8'b0;
    XRAM[13211] = 8'b0;
    XRAM[13212] = 8'b0;
    XRAM[13213] = 8'b0;
    XRAM[13214] = 8'b0;
    XRAM[13215] = 8'b0;
    XRAM[13216] = 8'b0;
    XRAM[13217] = 8'b0;
    XRAM[13218] = 8'b0;
    XRAM[13219] = 8'b0;
    XRAM[13220] = 8'b0;
    XRAM[13221] = 8'b0;
    XRAM[13222] = 8'b0;
    XRAM[13223] = 8'b0;
    XRAM[13224] = 8'b0;
    XRAM[13225] = 8'b0;
    XRAM[13226] = 8'b0;
    XRAM[13227] = 8'b0;
    XRAM[13228] = 8'b0;
    XRAM[13229] = 8'b0;
    XRAM[13230] = 8'b0;
    XRAM[13231] = 8'b0;
    XRAM[13232] = 8'b0;
    XRAM[13233] = 8'b0;
    XRAM[13234] = 8'b0;
    XRAM[13235] = 8'b0;
    XRAM[13236] = 8'b0;
    XRAM[13237] = 8'b0;
    XRAM[13238] = 8'b0;
    XRAM[13239] = 8'b0;
    XRAM[13240] = 8'b0;
    XRAM[13241] = 8'b0;
    XRAM[13242] = 8'b0;
    XRAM[13243] = 8'b0;
    XRAM[13244] = 8'b0;
    XRAM[13245] = 8'b0;
    XRAM[13246] = 8'b0;
    XRAM[13247] = 8'b0;
    XRAM[13248] = 8'b0;
    XRAM[13249] = 8'b0;
    XRAM[13250] = 8'b0;
    XRAM[13251] = 8'b0;
    XRAM[13252] = 8'b0;
    XRAM[13253] = 8'b0;
    XRAM[13254] = 8'b0;
    XRAM[13255] = 8'b0;
    XRAM[13256] = 8'b0;
    XRAM[13257] = 8'b0;
    XRAM[13258] = 8'b0;
    XRAM[13259] = 8'b0;
    XRAM[13260] = 8'b0;
    XRAM[13261] = 8'b0;
    XRAM[13262] = 8'b0;
    XRAM[13263] = 8'b0;
    XRAM[13264] = 8'b0;
    XRAM[13265] = 8'b0;
    XRAM[13266] = 8'b0;
    XRAM[13267] = 8'b0;
    XRAM[13268] = 8'b0;
    XRAM[13269] = 8'b0;
    XRAM[13270] = 8'b0;
    XRAM[13271] = 8'b0;
    XRAM[13272] = 8'b0;
    XRAM[13273] = 8'b0;
    XRAM[13274] = 8'b0;
    XRAM[13275] = 8'b0;
    XRAM[13276] = 8'b0;
    XRAM[13277] = 8'b0;
    XRAM[13278] = 8'b0;
    XRAM[13279] = 8'b0;
    XRAM[13280] = 8'b0;
    XRAM[13281] = 8'b0;
    XRAM[13282] = 8'b0;
    XRAM[13283] = 8'b0;
    XRAM[13284] = 8'b0;
    XRAM[13285] = 8'b0;
    XRAM[13286] = 8'b0;
    XRAM[13287] = 8'b0;
    XRAM[13288] = 8'b0;
    XRAM[13289] = 8'b0;
    XRAM[13290] = 8'b0;
    XRAM[13291] = 8'b0;
    XRAM[13292] = 8'b0;
    XRAM[13293] = 8'b0;
    XRAM[13294] = 8'b0;
    XRAM[13295] = 8'b0;
    XRAM[13296] = 8'b0;
    XRAM[13297] = 8'b0;
    XRAM[13298] = 8'b0;
    XRAM[13299] = 8'b0;
    XRAM[13300] = 8'b0;
    XRAM[13301] = 8'b0;
    XRAM[13302] = 8'b0;
    XRAM[13303] = 8'b0;
    XRAM[13304] = 8'b0;
    XRAM[13305] = 8'b0;
    XRAM[13306] = 8'b0;
    XRAM[13307] = 8'b0;
    XRAM[13308] = 8'b0;
    XRAM[13309] = 8'b0;
    XRAM[13310] = 8'b0;
    XRAM[13311] = 8'b0;
    XRAM[13312] = 8'b0;
    XRAM[13313] = 8'b0;
    XRAM[13314] = 8'b0;
    XRAM[13315] = 8'b0;
    XRAM[13316] = 8'b0;
    XRAM[13317] = 8'b0;
    XRAM[13318] = 8'b0;
    XRAM[13319] = 8'b0;
    XRAM[13320] = 8'b0;
    XRAM[13321] = 8'b0;
    XRAM[13322] = 8'b0;
    XRAM[13323] = 8'b0;
    XRAM[13324] = 8'b0;
    XRAM[13325] = 8'b0;
    XRAM[13326] = 8'b0;
    XRAM[13327] = 8'b0;
    XRAM[13328] = 8'b0;
    XRAM[13329] = 8'b0;
    XRAM[13330] = 8'b0;
    XRAM[13331] = 8'b0;
    XRAM[13332] = 8'b0;
    XRAM[13333] = 8'b0;
    XRAM[13334] = 8'b0;
    XRAM[13335] = 8'b0;
    XRAM[13336] = 8'b0;
    XRAM[13337] = 8'b0;
    XRAM[13338] = 8'b0;
    XRAM[13339] = 8'b0;
    XRAM[13340] = 8'b0;
    XRAM[13341] = 8'b0;
    XRAM[13342] = 8'b0;
    XRAM[13343] = 8'b0;
    XRAM[13344] = 8'b0;
    XRAM[13345] = 8'b0;
    XRAM[13346] = 8'b0;
    XRAM[13347] = 8'b0;
    XRAM[13348] = 8'b0;
    XRAM[13349] = 8'b0;
    XRAM[13350] = 8'b0;
    XRAM[13351] = 8'b0;
    XRAM[13352] = 8'b0;
    XRAM[13353] = 8'b0;
    XRAM[13354] = 8'b0;
    XRAM[13355] = 8'b0;
    XRAM[13356] = 8'b0;
    XRAM[13357] = 8'b0;
    XRAM[13358] = 8'b0;
    XRAM[13359] = 8'b0;
    XRAM[13360] = 8'b0;
    XRAM[13361] = 8'b0;
    XRAM[13362] = 8'b0;
    XRAM[13363] = 8'b0;
    XRAM[13364] = 8'b0;
    XRAM[13365] = 8'b0;
    XRAM[13366] = 8'b0;
    XRAM[13367] = 8'b0;
    XRAM[13368] = 8'b0;
    XRAM[13369] = 8'b0;
    XRAM[13370] = 8'b0;
    XRAM[13371] = 8'b0;
    XRAM[13372] = 8'b0;
    XRAM[13373] = 8'b0;
    XRAM[13374] = 8'b0;
    XRAM[13375] = 8'b0;
    XRAM[13376] = 8'b0;
    XRAM[13377] = 8'b0;
    XRAM[13378] = 8'b0;
    XRAM[13379] = 8'b0;
    XRAM[13380] = 8'b0;
    XRAM[13381] = 8'b0;
    XRAM[13382] = 8'b0;
    XRAM[13383] = 8'b0;
    XRAM[13384] = 8'b0;
    XRAM[13385] = 8'b0;
    XRAM[13386] = 8'b0;
    XRAM[13387] = 8'b0;
    XRAM[13388] = 8'b0;
    XRAM[13389] = 8'b0;
    XRAM[13390] = 8'b0;
    XRAM[13391] = 8'b0;
    XRAM[13392] = 8'b0;
    XRAM[13393] = 8'b0;
    XRAM[13394] = 8'b0;
    XRAM[13395] = 8'b0;
    XRAM[13396] = 8'b0;
    XRAM[13397] = 8'b0;
    XRAM[13398] = 8'b0;
    XRAM[13399] = 8'b0;
    XRAM[13400] = 8'b0;
    XRAM[13401] = 8'b0;
    XRAM[13402] = 8'b0;
    XRAM[13403] = 8'b0;
    XRAM[13404] = 8'b0;
    XRAM[13405] = 8'b0;
    XRAM[13406] = 8'b0;
    XRAM[13407] = 8'b0;
    XRAM[13408] = 8'b0;
    XRAM[13409] = 8'b0;
    XRAM[13410] = 8'b0;
    XRAM[13411] = 8'b0;
    XRAM[13412] = 8'b0;
    XRAM[13413] = 8'b0;
    XRAM[13414] = 8'b0;
    XRAM[13415] = 8'b0;
    XRAM[13416] = 8'b0;
    XRAM[13417] = 8'b0;
    XRAM[13418] = 8'b0;
    XRAM[13419] = 8'b0;
    XRAM[13420] = 8'b0;
    XRAM[13421] = 8'b0;
    XRAM[13422] = 8'b0;
    XRAM[13423] = 8'b0;
    XRAM[13424] = 8'b0;
    XRAM[13425] = 8'b0;
    XRAM[13426] = 8'b0;
    XRAM[13427] = 8'b0;
    XRAM[13428] = 8'b0;
    XRAM[13429] = 8'b0;
    XRAM[13430] = 8'b0;
    XRAM[13431] = 8'b0;
    XRAM[13432] = 8'b0;
    XRAM[13433] = 8'b0;
    XRAM[13434] = 8'b0;
    XRAM[13435] = 8'b0;
    XRAM[13436] = 8'b0;
    XRAM[13437] = 8'b0;
    XRAM[13438] = 8'b0;
    XRAM[13439] = 8'b0;
    XRAM[13440] = 8'b0;
    XRAM[13441] = 8'b0;
    XRAM[13442] = 8'b0;
    XRAM[13443] = 8'b0;
    XRAM[13444] = 8'b0;
    XRAM[13445] = 8'b0;
    XRAM[13446] = 8'b0;
    XRAM[13447] = 8'b0;
    XRAM[13448] = 8'b0;
    XRAM[13449] = 8'b0;
    XRAM[13450] = 8'b0;
    XRAM[13451] = 8'b0;
    XRAM[13452] = 8'b0;
    XRAM[13453] = 8'b0;
    XRAM[13454] = 8'b0;
    XRAM[13455] = 8'b0;
    XRAM[13456] = 8'b0;
    XRAM[13457] = 8'b0;
    XRAM[13458] = 8'b0;
    XRAM[13459] = 8'b0;
    XRAM[13460] = 8'b0;
    XRAM[13461] = 8'b0;
    XRAM[13462] = 8'b0;
    XRAM[13463] = 8'b0;
    XRAM[13464] = 8'b0;
    XRAM[13465] = 8'b0;
    XRAM[13466] = 8'b0;
    XRAM[13467] = 8'b0;
    XRAM[13468] = 8'b0;
    XRAM[13469] = 8'b0;
    XRAM[13470] = 8'b0;
    XRAM[13471] = 8'b0;
    XRAM[13472] = 8'b0;
    XRAM[13473] = 8'b0;
    XRAM[13474] = 8'b0;
    XRAM[13475] = 8'b0;
    XRAM[13476] = 8'b0;
    XRAM[13477] = 8'b0;
    XRAM[13478] = 8'b0;
    XRAM[13479] = 8'b0;
    XRAM[13480] = 8'b0;
    XRAM[13481] = 8'b0;
    XRAM[13482] = 8'b0;
    XRAM[13483] = 8'b0;
    XRAM[13484] = 8'b0;
    XRAM[13485] = 8'b0;
    XRAM[13486] = 8'b0;
    XRAM[13487] = 8'b0;
    XRAM[13488] = 8'b0;
    XRAM[13489] = 8'b0;
    XRAM[13490] = 8'b0;
    XRAM[13491] = 8'b0;
    XRAM[13492] = 8'b0;
    XRAM[13493] = 8'b0;
    XRAM[13494] = 8'b0;
    XRAM[13495] = 8'b0;
    XRAM[13496] = 8'b0;
    XRAM[13497] = 8'b0;
    XRAM[13498] = 8'b0;
    XRAM[13499] = 8'b0;
    XRAM[13500] = 8'b0;
    XRAM[13501] = 8'b0;
    XRAM[13502] = 8'b0;
    XRAM[13503] = 8'b0;
    XRAM[13504] = 8'b0;
    XRAM[13505] = 8'b0;
    XRAM[13506] = 8'b0;
    XRAM[13507] = 8'b0;
    XRAM[13508] = 8'b0;
    XRAM[13509] = 8'b0;
    XRAM[13510] = 8'b0;
    XRAM[13511] = 8'b0;
    XRAM[13512] = 8'b0;
    XRAM[13513] = 8'b0;
    XRAM[13514] = 8'b0;
    XRAM[13515] = 8'b0;
    XRAM[13516] = 8'b0;
    XRAM[13517] = 8'b0;
    XRAM[13518] = 8'b0;
    XRAM[13519] = 8'b0;
    XRAM[13520] = 8'b0;
    XRAM[13521] = 8'b0;
    XRAM[13522] = 8'b0;
    XRAM[13523] = 8'b0;
    XRAM[13524] = 8'b0;
    XRAM[13525] = 8'b0;
    XRAM[13526] = 8'b0;
    XRAM[13527] = 8'b0;
    XRAM[13528] = 8'b0;
    XRAM[13529] = 8'b0;
    XRAM[13530] = 8'b0;
    XRAM[13531] = 8'b0;
    XRAM[13532] = 8'b0;
    XRAM[13533] = 8'b0;
    XRAM[13534] = 8'b0;
    XRAM[13535] = 8'b0;
    XRAM[13536] = 8'b0;
    XRAM[13537] = 8'b0;
    XRAM[13538] = 8'b0;
    XRAM[13539] = 8'b0;
    XRAM[13540] = 8'b0;
    XRAM[13541] = 8'b0;
    XRAM[13542] = 8'b0;
    XRAM[13543] = 8'b0;
    XRAM[13544] = 8'b0;
    XRAM[13545] = 8'b0;
    XRAM[13546] = 8'b0;
    XRAM[13547] = 8'b0;
    XRAM[13548] = 8'b0;
    XRAM[13549] = 8'b0;
    XRAM[13550] = 8'b0;
    XRAM[13551] = 8'b0;
    XRAM[13552] = 8'b0;
    XRAM[13553] = 8'b0;
    XRAM[13554] = 8'b0;
    XRAM[13555] = 8'b0;
    XRAM[13556] = 8'b0;
    XRAM[13557] = 8'b0;
    XRAM[13558] = 8'b0;
    XRAM[13559] = 8'b0;
    XRAM[13560] = 8'b0;
    XRAM[13561] = 8'b0;
    XRAM[13562] = 8'b0;
    XRAM[13563] = 8'b0;
    XRAM[13564] = 8'b0;
    XRAM[13565] = 8'b0;
    XRAM[13566] = 8'b0;
    XRAM[13567] = 8'b0;
    XRAM[13568] = 8'b0;
    XRAM[13569] = 8'b0;
    XRAM[13570] = 8'b0;
    XRAM[13571] = 8'b0;
    XRAM[13572] = 8'b0;
    XRAM[13573] = 8'b0;
    XRAM[13574] = 8'b0;
    XRAM[13575] = 8'b0;
    XRAM[13576] = 8'b0;
    XRAM[13577] = 8'b0;
    XRAM[13578] = 8'b0;
    XRAM[13579] = 8'b0;
    XRAM[13580] = 8'b0;
    XRAM[13581] = 8'b0;
    XRAM[13582] = 8'b0;
    XRAM[13583] = 8'b0;
    XRAM[13584] = 8'b0;
    XRAM[13585] = 8'b0;
    XRAM[13586] = 8'b0;
    XRAM[13587] = 8'b0;
    XRAM[13588] = 8'b0;
    XRAM[13589] = 8'b0;
    XRAM[13590] = 8'b0;
    XRAM[13591] = 8'b0;
    XRAM[13592] = 8'b0;
    XRAM[13593] = 8'b0;
    XRAM[13594] = 8'b0;
    XRAM[13595] = 8'b0;
    XRAM[13596] = 8'b0;
    XRAM[13597] = 8'b0;
    XRAM[13598] = 8'b0;
    XRAM[13599] = 8'b0;
    XRAM[13600] = 8'b0;
    XRAM[13601] = 8'b0;
    XRAM[13602] = 8'b0;
    XRAM[13603] = 8'b0;
    XRAM[13604] = 8'b0;
    XRAM[13605] = 8'b0;
    XRAM[13606] = 8'b0;
    XRAM[13607] = 8'b0;
    XRAM[13608] = 8'b0;
    XRAM[13609] = 8'b0;
    XRAM[13610] = 8'b0;
    XRAM[13611] = 8'b0;
    XRAM[13612] = 8'b0;
    XRAM[13613] = 8'b0;
    XRAM[13614] = 8'b0;
    XRAM[13615] = 8'b0;
    XRAM[13616] = 8'b0;
    XRAM[13617] = 8'b0;
    XRAM[13618] = 8'b0;
    XRAM[13619] = 8'b0;
    XRAM[13620] = 8'b0;
    XRAM[13621] = 8'b0;
    XRAM[13622] = 8'b0;
    XRAM[13623] = 8'b0;
    XRAM[13624] = 8'b0;
    XRAM[13625] = 8'b0;
    XRAM[13626] = 8'b0;
    XRAM[13627] = 8'b0;
    XRAM[13628] = 8'b0;
    XRAM[13629] = 8'b0;
    XRAM[13630] = 8'b0;
    XRAM[13631] = 8'b0;
    XRAM[13632] = 8'b0;
    XRAM[13633] = 8'b0;
    XRAM[13634] = 8'b0;
    XRAM[13635] = 8'b0;
    XRAM[13636] = 8'b0;
    XRAM[13637] = 8'b0;
    XRAM[13638] = 8'b0;
    XRAM[13639] = 8'b0;
    XRAM[13640] = 8'b0;
    XRAM[13641] = 8'b0;
    XRAM[13642] = 8'b0;
    XRAM[13643] = 8'b0;
    XRAM[13644] = 8'b0;
    XRAM[13645] = 8'b0;
    XRAM[13646] = 8'b0;
    XRAM[13647] = 8'b0;
    XRAM[13648] = 8'b0;
    XRAM[13649] = 8'b0;
    XRAM[13650] = 8'b0;
    XRAM[13651] = 8'b0;
    XRAM[13652] = 8'b0;
    XRAM[13653] = 8'b0;
    XRAM[13654] = 8'b0;
    XRAM[13655] = 8'b0;
    XRAM[13656] = 8'b0;
    XRAM[13657] = 8'b0;
    XRAM[13658] = 8'b0;
    XRAM[13659] = 8'b0;
    XRAM[13660] = 8'b0;
    XRAM[13661] = 8'b0;
    XRAM[13662] = 8'b0;
    XRAM[13663] = 8'b0;
    XRAM[13664] = 8'b0;
    XRAM[13665] = 8'b0;
    XRAM[13666] = 8'b0;
    XRAM[13667] = 8'b0;
    XRAM[13668] = 8'b0;
    XRAM[13669] = 8'b0;
    XRAM[13670] = 8'b0;
    XRAM[13671] = 8'b0;
    XRAM[13672] = 8'b0;
    XRAM[13673] = 8'b0;
    XRAM[13674] = 8'b0;
    XRAM[13675] = 8'b0;
    XRAM[13676] = 8'b0;
    XRAM[13677] = 8'b0;
    XRAM[13678] = 8'b0;
    XRAM[13679] = 8'b0;
    XRAM[13680] = 8'b0;
    XRAM[13681] = 8'b0;
    XRAM[13682] = 8'b0;
    XRAM[13683] = 8'b0;
    XRAM[13684] = 8'b0;
    XRAM[13685] = 8'b0;
    XRAM[13686] = 8'b0;
    XRAM[13687] = 8'b0;
    XRAM[13688] = 8'b0;
    XRAM[13689] = 8'b0;
    XRAM[13690] = 8'b0;
    XRAM[13691] = 8'b0;
    XRAM[13692] = 8'b0;
    XRAM[13693] = 8'b0;
    XRAM[13694] = 8'b0;
    XRAM[13695] = 8'b0;
    XRAM[13696] = 8'b0;
    XRAM[13697] = 8'b0;
    XRAM[13698] = 8'b0;
    XRAM[13699] = 8'b0;
    XRAM[13700] = 8'b0;
    XRAM[13701] = 8'b0;
    XRAM[13702] = 8'b0;
    XRAM[13703] = 8'b0;
    XRAM[13704] = 8'b0;
    XRAM[13705] = 8'b0;
    XRAM[13706] = 8'b0;
    XRAM[13707] = 8'b0;
    XRAM[13708] = 8'b0;
    XRAM[13709] = 8'b0;
    XRAM[13710] = 8'b0;
    XRAM[13711] = 8'b0;
    XRAM[13712] = 8'b0;
    XRAM[13713] = 8'b0;
    XRAM[13714] = 8'b0;
    XRAM[13715] = 8'b0;
    XRAM[13716] = 8'b0;
    XRAM[13717] = 8'b0;
    XRAM[13718] = 8'b0;
    XRAM[13719] = 8'b0;
    XRAM[13720] = 8'b0;
    XRAM[13721] = 8'b0;
    XRAM[13722] = 8'b0;
    XRAM[13723] = 8'b0;
    XRAM[13724] = 8'b0;
    XRAM[13725] = 8'b0;
    XRAM[13726] = 8'b0;
    XRAM[13727] = 8'b0;
    XRAM[13728] = 8'b0;
    XRAM[13729] = 8'b0;
    XRAM[13730] = 8'b0;
    XRAM[13731] = 8'b0;
    XRAM[13732] = 8'b0;
    XRAM[13733] = 8'b0;
    XRAM[13734] = 8'b0;
    XRAM[13735] = 8'b0;
    XRAM[13736] = 8'b0;
    XRAM[13737] = 8'b0;
    XRAM[13738] = 8'b0;
    XRAM[13739] = 8'b0;
    XRAM[13740] = 8'b0;
    XRAM[13741] = 8'b0;
    XRAM[13742] = 8'b0;
    XRAM[13743] = 8'b0;
    XRAM[13744] = 8'b0;
    XRAM[13745] = 8'b0;
    XRAM[13746] = 8'b0;
    XRAM[13747] = 8'b0;
    XRAM[13748] = 8'b0;
    XRAM[13749] = 8'b0;
    XRAM[13750] = 8'b0;
    XRAM[13751] = 8'b0;
    XRAM[13752] = 8'b0;
    XRAM[13753] = 8'b0;
    XRAM[13754] = 8'b0;
    XRAM[13755] = 8'b0;
    XRAM[13756] = 8'b0;
    XRAM[13757] = 8'b0;
    XRAM[13758] = 8'b0;
    XRAM[13759] = 8'b0;
    XRAM[13760] = 8'b0;
    XRAM[13761] = 8'b0;
    XRAM[13762] = 8'b0;
    XRAM[13763] = 8'b0;
    XRAM[13764] = 8'b0;
    XRAM[13765] = 8'b0;
    XRAM[13766] = 8'b0;
    XRAM[13767] = 8'b0;
    XRAM[13768] = 8'b0;
    XRAM[13769] = 8'b0;
    XRAM[13770] = 8'b0;
    XRAM[13771] = 8'b0;
    XRAM[13772] = 8'b0;
    XRAM[13773] = 8'b0;
    XRAM[13774] = 8'b0;
    XRAM[13775] = 8'b0;
    XRAM[13776] = 8'b0;
    XRAM[13777] = 8'b0;
    XRAM[13778] = 8'b0;
    XRAM[13779] = 8'b0;
    XRAM[13780] = 8'b0;
    XRAM[13781] = 8'b0;
    XRAM[13782] = 8'b0;
    XRAM[13783] = 8'b0;
    XRAM[13784] = 8'b0;
    XRAM[13785] = 8'b0;
    XRAM[13786] = 8'b0;
    XRAM[13787] = 8'b0;
    XRAM[13788] = 8'b0;
    XRAM[13789] = 8'b0;
    XRAM[13790] = 8'b0;
    XRAM[13791] = 8'b0;
    XRAM[13792] = 8'b0;
    XRAM[13793] = 8'b0;
    XRAM[13794] = 8'b0;
    XRAM[13795] = 8'b0;
    XRAM[13796] = 8'b0;
    XRAM[13797] = 8'b0;
    XRAM[13798] = 8'b0;
    XRAM[13799] = 8'b0;
    XRAM[13800] = 8'b0;
    XRAM[13801] = 8'b0;
    XRAM[13802] = 8'b0;
    XRAM[13803] = 8'b0;
    XRAM[13804] = 8'b0;
    XRAM[13805] = 8'b0;
    XRAM[13806] = 8'b0;
    XRAM[13807] = 8'b0;
    XRAM[13808] = 8'b0;
    XRAM[13809] = 8'b0;
    XRAM[13810] = 8'b0;
    XRAM[13811] = 8'b0;
    XRAM[13812] = 8'b0;
    XRAM[13813] = 8'b0;
    XRAM[13814] = 8'b0;
    XRAM[13815] = 8'b0;
    XRAM[13816] = 8'b0;
    XRAM[13817] = 8'b0;
    XRAM[13818] = 8'b0;
    XRAM[13819] = 8'b0;
    XRAM[13820] = 8'b0;
    XRAM[13821] = 8'b0;
    XRAM[13822] = 8'b0;
    XRAM[13823] = 8'b0;
    XRAM[13824] = 8'b0;
    XRAM[13825] = 8'b0;
    XRAM[13826] = 8'b0;
    XRAM[13827] = 8'b0;
    XRAM[13828] = 8'b0;
    XRAM[13829] = 8'b0;
    XRAM[13830] = 8'b0;
    XRAM[13831] = 8'b0;
    XRAM[13832] = 8'b0;
    XRAM[13833] = 8'b0;
    XRAM[13834] = 8'b0;
    XRAM[13835] = 8'b0;
    XRAM[13836] = 8'b0;
    XRAM[13837] = 8'b0;
    XRAM[13838] = 8'b0;
    XRAM[13839] = 8'b0;
    XRAM[13840] = 8'b0;
    XRAM[13841] = 8'b0;
    XRAM[13842] = 8'b0;
    XRAM[13843] = 8'b0;
    XRAM[13844] = 8'b0;
    XRAM[13845] = 8'b0;
    XRAM[13846] = 8'b0;
    XRAM[13847] = 8'b0;
    XRAM[13848] = 8'b0;
    XRAM[13849] = 8'b0;
    XRAM[13850] = 8'b0;
    XRAM[13851] = 8'b0;
    XRAM[13852] = 8'b0;
    XRAM[13853] = 8'b0;
    XRAM[13854] = 8'b0;
    XRAM[13855] = 8'b0;
    XRAM[13856] = 8'b0;
    XRAM[13857] = 8'b0;
    XRAM[13858] = 8'b0;
    XRAM[13859] = 8'b0;
    XRAM[13860] = 8'b0;
    XRAM[13861] = 8'b0;
    XRAM[13862] = 8'b0;
    XRAM[13863] = 8'b0;
    XRAM[13864] = 8'b0;
    XRAM[13865] = 8'b0;
    XRAM[13866] = 8'b0;
    XRAM[13867] = 8'b0;
    XRAM[13868] = 8'b0;
    XRAM[13869] = 8'b0;
    XRAM[13870] = 8'b0;
    XRAM[13871] = 8'b0;
    XRAM[13872] = 8'b0;
    XRAM[13873] = 8'b0;
    XRAM[13874] = 8'b0;
    XRAM[13875] = 8'b0;
    XRAM[13876] = 8'b0;
    XRAM[13877] = 8'b0;
    XRAM[13878] = 8'b0;
    XRAM[13879] = 8'b0;
    XRAM[13880] = 8'b0;
    XRAM[13881] = 8'b0;
    XRAM[13882] = 8'b0;
    XRAM[13883] = 8'b0;
    XRAM[13884] = 8'b0;
    XRAM[13885] = 8'b0;
    XRAM[13886] = 8'b0;
    XRAM[13887] = 8'b0;
    XRAM[13888] = 8'b0;
    XRAM[13889] = 8'b0;
    XRAM[13890] = 8'b0;
    XRAM[13891] = 8'b0;
    XRAM[13892] = 8'b0;
    XRAM[13893] = 8'b0;
    XRAM[13894] = 8'b0;
    XRAM[13895] = 8'b0;
    XRAM[13896] = 8'b0;
    XRAM[13897] = 8'b0;
    XRAM[13898] = 8'b0;
    XRAM[13899] = 8'b0;
    XRAM[13900] = 8'b0;
    XRAM[13901] = 8'b0;
    XRAM[13902] = 8'b0;
    XRAM[13903] = 8'b0;
    XRAM[13904] = 8'b0;
    XRAM[13905] = 8'b0;
    XRAM[13906] = 8'b0;
    XRAM[13907] = 8'b0;
    XRAM[13908] = 8'b0;
    XRAM[13909] = 8'b0;
    XRAM[13910] = 8'b0;
    XRAM[13911] = 8'b0;
    XRAM[13912] = 8'b0;
    XRAM[13913] = 8'b0;
    XRAM[13914] = 8'b0;
    XRAM[13915] = 8'b0;
    XRAM[13916] = 8'b0;
    XRAM[13917] = 8'b0;
    XRAM[13918] = 8'b0;
    XRAM[13919] = 8'b0;
    XRAM[13920] = 8'b0;
    XRAM[13921] = 8'b0;
    XRAM[13922] = 8'b0;
    XRAM[13923] = 8'b0;
    XRAM[13924] = 8'b0;
    XRAM[13925] = 8'b0;
    XRAM[13926] = 8'b0;
    XRAM[13927] = 8'b0;
    XRAM[13928] = 8'b0;
    XRAM[13929] = 8'b0;
    XRAM[13930] = 8'b0;
    XRAM[13931] = 8'b0;
    XRAM[13932] = 8'b0;
    XRAM[13933] = 8'b0;
    XRAM[13934] = 8'b0;
    XRAM[13935] = 8'b0;
    XRAM[13936] = 8'b0;
    XRAM[13937] = 8'b0;
    XRAM[13938] = 8'b0;
    XRAM[13939] = 8'b0;
    XRAM[13940] = 8'b0;
    XRAM[13941] = 8'b0;
    XRAM[13942] = 8'b0;
    XRAM[13943] = 8'b0;
    XRAM[13944] = 8'b0;
    XRAM[13945] = 8'b0;
    XRAM[13946] = 8'b0;
    XRAM[13947] = 8'b0;
    XRAM[13948] = 8'b0;
    XRAM[13949] = 8'b0;
    XRAM[13950] = 8'b0;
    XRAM[13951] = 8'b0;
    XRAM[13952] = 8'b0;
    XRAM[13953] = 8'b0;
    XRAM[13954] = 8'b0;
    XRAM[13955] = 8'b0;
    XRAM[13956] = 8'b0;
    XRAM[13957] = 8'b0;
    XRAM[13958] = 8'b0;
    XRAM[13959] = 8'b0;
    XRAM[13960] = 8'b0;
    XRAM[13961] = 8'b0;
    XRAM[13962] = 8'b0;
    XRAM[13963] = 8'b0;
    XRAM[13964] = 8'b0;
    XRAM[13965] = 8'b0;
    XRAM[13966] = 8'b0;
    XRAM[13967] = 8'b0;
    XRAM[13968] = 8'b0;
    XRAM[13969] = 8'b0;
    XRAM[13970] = 8'b0;
    XRAM[13971] = 8'b0;
    XRAM[13972] = 8'b0;
    XRAM[13973] = 8'b0;
    XRAM[13974] = 8'b0;
    XRAM[13975] = 8'b0;
    XRAM[13976] = 8'b0;
    XRAM[13977] = 8'b0;
    XRAM[13978] = 8'b0;
    XRAM[13979] = 8'b0;
    XRAM[13980] = 8'b0;
    XRAM[13981] = 8'b0;
    XRAM[13982] = 8'b0;
    XRAM[13983] = 8'b0;
    XRAM[13984] = 8'b0;
    XRAM[13985] = 8'b0;
    XRAM[13986] = 8'b0;
    XRAM[13987] = 8'b0;
    XRAM[13988] = 8'b0;
    XRAM[13989] = 8'b0;
    XRAM[13990] = 8'b0;
    XRAM[13991] = 8'b0;
    XRAM[13992] = 8'b0;
    XRAM[13993] = 8'b0;
    XRAM[13994] = 8'b0;
    XRAM[13995] = 8'b0;
    XRAM[13996] = 8'b0;
    XRAM[13997] = 8'b0;
    XRAM[13998] = 8'b0;
    XRAM[13999] = 8'b0;
    XRAM[14000] = 8'b0;
    XRAM[14001] = 8'b0;
    XRAM[14002] = 8'b0;
    XRAM[14003] = 8'b0;
    XRAM[14004] = 8'b0;
    XRAM[14005] = 8'b0;
    XRAM[14006] = 8'b0;
    XRAM[14007] = 8'b0;
    XRAM[14008] = 8'b0;
    XRAM[14009] = 8'b0;
    XRAM[14010] = 8'b0;
    XRAM[14011] = 8'b0;
    XRAM[14012] = 8'b0;
    XRAM[14013] = 8'b0;
    XRAM[14014] = 8'b0;
    XRAM[14015] = 8'b0;
    XRAM[14016] = 8'b0;
    XRAM[14017] = 8'b0;
    XRAM[14018] = 8'b0;
    XRAM[14019] = 8'b0;
    XRAM[14020] = 8'b0;
    XRAM[14021] = 8'b0;
    XRAM[14022] = 8'b0;
    XRAM[14023] = 8'b0;
    XRAM[14024] = 8'b0;
    XRAM[14025] = 8'b0;
    XRAM[14026] = 8'b0;
    XRAM[14027] = 8'b0;
    XRAM[14028] = 8'b0;
    XRAM[14029] = 8'b0;
    XRAM[14030] = 8'b0;
    XRAM[14031] = 8'b0;
    XRAM[14032] = 8'b0;
    XRAM[14033] = 8'b0;
    XRAM[14034] = 8'b0;
    XRAM[14035] = 8'b0;
    XRAM[14036] = 8'b0;
    XRAM[14037] = 8'b0;
    XRAM[14038] = 8'b0;
    XRAM[14039] = 8'b0;
    XRAM[14040] = 8'b0;
    XRAM[14041] = 8'b0;
    XRAM[14042] = 8'b0;
    XRAM[14043] = 8'b0;
    XRAM[14044] = 8'b0;
    XRAM[14045] = 8'b0;
    XRAM[14046] = 8'b0;
    XRAM[14047] = 8'b0;
    XRAM[14048] = 8'b0;
    XRAM[14049] = 8'b0;
    XRAM[14050] = 8'b0;
    XRAM[14051] = 8'b0;
    XRAM[14052] = 8'b0;
    XRAM[14053] = 8'b0;
    XRAM[14054] = 8'b0;
    XRAM[14055] = 8'b0;
    XRAM[14056] = 8'b0;
    XRAM[14057] = 8'b0;
    XRAM[14058] = 8'b0;
    XRAM[14059] = 8'b0;
    XRAM[14060] = 8'b0;
    XRAM[14061] = 8'b0;
    XRAM[14062] = 8'b0;
    XRAM[14063] = 8'b0;
    XRAM[14064] = 8'b0;
    XRAM[14065] = 8'b0;
    XRAM[14066] = 8'b0;
    XRAM[14067] = 8'b0;
    XRAM[14068] = 8'b0;
    XRAM[14069] = 8'b0;
    XRAM[14070] = 8'b0;
    XRAM[14071] = 8'b0;
    XRAM[14072] = 8'b0;
    XRAM[14073] = 8'b0;
    XRAM[14074] = 8'b0;
    XRAM[14075] = 8'b0;
    XRAM[14076] = 8'b0;
    XRAM[14077] = 8'b0;
    XRAM[14078] = 8'b0;
    XRAM[14079] = 8'b0;
    XRAM[14080] = 8'b0;
    XRAM[14081] = 8'b0;
    XRAM[14082] = 8'b0;
    XRAM[14083] = 8'b0;
    XRAM[14084] = 8'b0;
    XRAM[14085] = 8'b0;
    XRAM[14086] = 8'b0;
    XRAM[14087] = 8'b0;
    XRAM[14088] = 8'b0;
    XRAM[14089] = 8'b0;
    XRAM[14090] = 8'b0;
    XRAM[14091] = 8'b0;
    XRAM[14092] = 8'b0;
    XRAM[14093] = 8'b0;
    XRAM[14094] = 8'b0;
    XRAM[14095] = 8'b0;
    XRAM[14096] = 8'b0;
    XRAM[14097] = 8'b0;
    XRAM[14098] = 8'b0;
    XRAM[14099] = 8'b0;
    XRAM[14100] = 8'b0;
    XRAM[14101] = 8'b0;
    XRAM[14102] = 8'b0;
    XRAM[14103] = 8'b0;
    XRAM[14104] = 8'b0;
    XRAM[14105] = 8'b0;
    XRAM[14106] = 8'b0;
    XRAM[14107] = 8'b0;
    XRAM[14108] = 8'b0;
    XRAM[14109] = 8'b0;
    XRAM[14110] = 8'b0;
    XRAM[14111] = 8'b0;
    XRAM[14112] = 8'b0;
    XRAM[14113] = 8'b0;
    XRAM[14114] = 8'b0;
    XRAM[14115] = 8'b0;
    XRAM[14116] = 8'b0;
    XRAM[14117] = 8'b0;
    XRAM[14118] = 8'b0;
    XRAM[14119] = 8'b0;
    XRAM[14120] = 8'b0;
    XRAM[14121] = 8'b0;
    XRAM[14122] = 8'b0;
    XRAM[14123] = 8'b0;
    XRAM[14124] = 8'b0;
    XRAM[14125] = 8'b0;
    XRAM[14126] = 8'b0;
    XRAM[14127] = 8'b0;
    XRAM[14128] = 8'b0;
    XRAM[14129] = 8'b0;
    XRAM[14130] = 8'b0;
    XRAM[14131] = 8'b0;
    XRAM[14132] = 8'b0;
    XRAM[14133] = 8'b0;
    XRAM[14134] = 8'b0;
    XRAM[14135] = 8'b0;
    XRAM[14136] = 8'b0;
    XRAM[14137] = 8'b0;
    XRAM[14138] = 8'b0;
    XRAM[14139] = 8'b0;
    XRAM[14140] = 8'b0;
    XRAM[14141] = 8'b0;
    XRAM[14142] = 8'b0;
    XRAM[14143] = 8'b0;
    XRAM[14144] = 8'b0;
    XRAM[14145] = 8'b0;
    XRAM[14146] = 8'b0;
    XRAM[14147] = 8'b0;
    XRAM[14148] = 8'b0;
    XRAM[14149] = 8'b0;
    XRAM[14150] = 8'b0;
    XRAM[14151] = 8'b0;
    XRAM[14152] = 8'b0;
    XRAM[14153] = 8'b0;
    XRAM[14154] = 8'b0;
    XRAM[14155] = 8'b0;
    XRAM[14156] = 8'b0;
    XRAM[14157] = 8'b0;
    XRAM[14158] = 8'b0;
    XRAM[14159] = 8'b0;
    XRAM[14160] = 8'b0;
    XRAM[14161] = 8'b0;
    XRAM[14162] = 8'b0;
    XRAM[14163] = 8'b0;
    XRAM[14164] = 8'b0;
    XRAM[14165] = 8'b0;
    XRAM[14166] = 8'b0;
    XRAM[14167] = 8'b0;
    XRAM[14168] = 8'b0;
    XRAM[14169] = 8'b0;
    XRAM[14170] = 8'b0;
    XRAM[14171] = 8'b0;
    XRAM[14172] = 8'b0;
    XRAM[14173] = 8'b0;
    XRAM[14174] = 8'b0;
    XRAM[14175] = 8'b0;
    XRAM[14176] = 8'b0;
    XRAM[14177] = 8'b0;
    XRAM[14178] = 8'b0;
    XRAM[14179] = 8'b0;
    XRAM[14180] = 8'b0;
    XRAM[14181] = 8'b0;
    XRAM[14182] = 8'b0;
    XRAM[14183] = 8'b0;
    XRAM[14184] = 8'b0;
    XRAM[14185] = 8'b0;
    XRAM[14186] = 8'b0;
    XRAM[14187] = 8'b0;
    XRAM[14188] = 8'b0;
    XRAM[14189] = 8'b0;
    XRAM[14190] = 8'b0;
    XRAM[14191] = 8'b0;
    XRAM[14192] = 8'b0;
    XRAM[14193] = 8'b0;
    XRAM[14194] = 8'b0;
    XRAM[14195] = 8'b0;
    XRAM[14196] = 8'b0;
    XRAM[14197] = 8'b0;
    XRAM[14198] = 8'b0;
    XRAM[14199] = 8'b0;
    XRAM[14200] = 8'b0;
    XRAM[14201] = 8'b0;
    XRAM[14202] = 8'b0;
    XRAM[14203] = 8'b0;
    XRAM[14204] = 8'b0;
    XRAM[14205] = 8'b0;
    XRAM[14206] = 8'b0;
    XRAM[14207] = 8'b0;
    XRAM[14208] = 8'b0;
    XRAM[14209] = 8'b0;
    XRAM[14210] = 8'b0;
    XRAM[14211] = 8'b0;
    XRAM[14212] = 8'b0;
    XRAM[14213] = 8'b0;
    XRAM[14214] = 8'b0;
    XRAM[14215] = 8'b0;
    XRAM[14216] = 8'b0;
    XRAM[14217] = 8'b0;
    XRAM[14218] = 8'b0;
    XRAM[14219] = 8'b0;
    XRAM[14220] = 8'b0;
    XRAM[14221] = 8'b0;
    XRAM[14222] = 8'b0;
    XRAM[14223] = 8'b0;
    XRAM[14224] = 8'b0;
    XRAM[14225] = 8'b0;
    XRAM[14226] = 8'b0;
    XRAM[14227] = 8'b0;
    XRAM[14228] = 8'b0;
    XRAM[14229] = 8'b0;
    XRAM[14230] = 8'b0;
    XRAM[14231] = 8'b0;
    XRAM[14232] = 8'b0;
    XRAM[14233] = 8'b0;
    XRAM[14234] = 8'b0;
    XRAM[14235] = 8'b0;
    XRAM[14236] = 8'b0;
    XRAM[14237] = 8'b0;
    XRAM[14238] = 8'b0;
    XRAM[14239] = 8'b0;
    XRAM[14240] = 8'b0;
    XRAM[14241] = 8'b0;
    XRAM[14242] = 8'b0;
    XRAM[14243] = 8'b0;
    XRAM[14244] = 8'b0;
    XRAM[14245] = 8'b0;
    XRAM[14246] = 8'b0;
    XRAM[14247] = 8'b0;
    XRAM[14248] = 8'b0;
    XRAM[14249] = 8'b0;
    XRAM[14250] = 8'b0;
    XRAM[14251] = 8'b0;
    XRAM[14252] = 8'b0;
    XRAM[14253] = 8'b0;
    XRAM[14254] = 8'b0;
    XRAM[14255] = 8'b0;
    XRAM[14256] = 8'b0;
    XRAM[14257] = 8'b0;
    XRAM[14258] = 8'b0;
    XRAM[14259] = 8'b0;
    XRAM[14260] = 8'b0;
    XRAM[14261] = 8'b0;
    XRAM[14262] = 8'b0;
    XRAM[14263] = 8'b0;
    XRAM[14264] = 8'b0;
    XRAM[14265] = 8'b0;
    XRAM[14266] = 8'b0;
    XRAM[14267] = 8'b0;
    XRAM[14268] = 8'b0;
    XRAM[14269] = 8'b0;
    XRAM[14270] = 8'b0;
    XRAM[14271] = 8'b0;
    XRAM[14272] = 8'b0;
    XRAM[14273] = 8'b0;
    XRAM[14274] = 8'b0;
    XRAM[14275] = 8'b0;
    XRAM[14276] = 8'b0;
    XRAM[14277] = 8'b0;
    XRAM[14278] = 8'b0;
    XRAM[14279] = 8'b0;
    XRAM[14280] = 8'b0;
    XRAM[14281] = 8'b0;
    XRAM[14282] = 8'b0;
    XRAM[14283] = 8'b0;
    XRAM[14284] = 8'b0;
    XRAM[14285] = 8'b0;
    XRAM[14286] = 8'b0;
    XRAM[14287] = 8'b0;
    XRAM[14288] = 8'b0;
    XRAM[14289] = 8'b0;
    XRAM[14290] = 8'b0;
    XRAM[14291] = 8'b0;
    XRAM[14292] = 8'b0;
    XRAM[14293] = 8'b0;
    XRAM[14294] = 8'b0;
    XRAM[14295] = 8'b0;
    XRAM[14296] = 8'b0;
    XRAM[14297] = 8'b0;
    XRAM[14298] = 8'b0;
    XRAM[14299] = 8'b0;
    XRAM[14300] = 8'b0;
    XRAM[14301] = 8'b0;
    XRAM[14302] = 8'b0;
    XRAM[14303] = 8'b0;
    XRAM[14304] = 8'b0;
    XRAM[14305] = 8'b0;
    XRAM[14306] = 8'b0;
    XRAM[14307] = 8'b0;
    XRAM[14308] = 8'b0;
    XRAM[14309] = 8'b0;
    XRAM[14310] = 8'b0;
    XRAM[14311] = 8'b0;
    XRAM[14312] = 8'b0;
    XRAM[14313] = 8'b0;
    XRAM[14314] = 8'b0;
    XRAM[14315] = 8'b0;
    XRAM[14316] = 8'b0;
    XRAM[14317] = 8'b0;
    XRAM[14318] = 8'b0;
    XRAM[14319] = 8'b0;
    XRAM[14320] = 8'b0;
    XRAM[14321] = 8'b0;
    XRAM[14322] = 8'b0;
    XRAM[14323] = 8'b0;
    XRAM[14324] = 8'b0;
    XRAM[14325] = 8'b0;
    XRAM[14326] = 8'b0;
    XRAM[14327] = 8'b0;
    XRAM[14328] = 8'b0;
    XRAM[14329] = 8'b0;
    XRAM[14330] = 8'b0;
    XRAM[14331] = 8'b0;
    XRAM[14332] = 8'b0;
    XRAM[14333] = 8'b0;
    XRAM[14334] = 8'b0;
    XRAM[14335] = 8'b0;
    XRAM[14336] = 8'b0;
    XRAM[14337] = 8'b0;
    XRAM[14338] = 8'b0;
    XRAM[14339] = 8'b0;
    XRAM[14340] = 8'b0;
    XRAM[14341] = 8'b0;
    XRAM[14342] = 8'b0;
    XRAM[14343] = 8'b0;
    XRAM[14344] = 8'b0;
    XRAM[14345] = 8'b0;
    XRAM[14346] = 8'b0;
    XRAM[14347] = 8'b0;
    XRAM[14348] = 8'b0;
    XRAM[14349] = 8'b0;
    XRAM[14350] = 8'b0;
    XRAM[14351] = 8'b0;
    XRAM[14352] = 8'b0;
    XRAM[14353] = 8'b0;
    XRAM[14354] = 8'b0;
    XRAM[14355] = 8'b0;
    XRAM[14356] = 8'b0;
    XRAM[14357] = 8'b0;
    XRAM[14358] = 8'b0;
    XRAM[14359] = 8'b0;
    XRAM[14360] = 8'b0;
    XRAM[14361] = 8'b0;
    XRAM[14362] = 8'b0;
    XRAM[14363] = 8'b0;
    XRAM[14364] = 8'b0;
    XRAM[14365] = 8'b0;
    XRAM[14366] = 8'b0;
    XRAM[14367] = 8'b0;
    XRAM[14368] = 8'b0;
    XRAM[14369] = 8'b0;
    XRAM[14370] = 8'b0;
    XRAM[14371] = 8'b0;
    XRAM[14372] = 8'b0;
    XRAM[14373] = 8'b0;
    XRAM[14374] = 8'b0;
    XRAM[14375] = 8'b0;
    XRAM[14376] = 8'b0;
    XRAM[14377] = 8'b0;
    XRAM[14378] = 8'b0;
    XRAM[14379] = 8'b0;
    XRAM[14380] = 8'b0;
    XRAM[14381] = 8'b0;
    XRAM[14382] = 8'b0;
    XRAM[14383] = 8'b0;
    XRAM[14384] = 8'b0;
    XRAM[14385] = 8'b0;
    XRAM[14386] = 8'b0;
    XRAM[14387] = 8'b0;
    XRAM[14388] = 8'b0;
    XRAM[14389] = 8'b0;
    XRAM[14390] = 8'b0;
    XRAM[14391] = 8'b0;
    XRAM[14392] = 8'b0;
    XRAM[14393] = 8'b0;
    XRAM[14394] = 8'b0;
    XRAM[14395] = 8'b0;
    XRAM[14396] = 8'b0;
    XRAM[14397] = 8'b0;
    XRAM[14398] = 8'b0;
    XRAM[14399] = 8'b0;
    XRAM[14400] = 8'b0;
    XRAM[14401] = 8'b0;
    XRAM[14402] = 8'b0;
    XRAM[14403] = 8'b0;
    XRAM[14404] = 8'b0;
    XRAM[14405] = 8'b0;
    XRAM[14406] = 8'b0;
    XRAM[14407] = 8'b0;
    XRAM[14408] = 8'b0;
    XRAM[14409] = 8'b0;
    XRAM[14410] = 8'b0;
    XRAM[14411] = 8'b0;
    XRAM[14412] = 8'b0;
    XRAM[14413] = 8'b0;
    XRAM[14414] = 8'b0;
    XRAM[14415] = 8'b0;
    XRAM[14416] = 8'b0;
    XRAM[14417] = 8'b0;
    XRAM[14418] = 8'b0;
    XRAM[14419] = 8'b0;
    XRAM[14420] = 8'b0;
    XRAM[14421] = 8'b0;
    XRAM[14422] = 8'b0;
    XRAM[14423] = 8'b0;
    XRAM[14424] = 8'b0;
    XRAM[14425] = 8'b0;
    XRAM[14426] = 8'b0;
    XRAM[14427] = 8'b0;
    XRAM[14428] = 8'b0;
    XRAM[14429] = 8'b0;
    XRAM[14430] = 8'b0;
    XRAM[14431] = 8'b0;
    XRAM[14432] = 8'b0;
    XRAM[14433] = 8'b0;
    XRAM[14434] = 8'b0;
    XRAM[14435] = 8'b0;
    XRAM[14436] = 8'b0;
    XRAM[14437] = 8'b0;
    XRAM[14438] = 8'b0;
    XRAM[14439] = 8'b0;
    XRAM[14440] = 8'b0;
    XRAM[14441] = 8'b0;
    XRAM[14442] = 8'b0;
    XRAM[14443] = 8'b0;
    XRAM[14444] = 8'b0;
    XRAM[14445] = 8'b0;
    XRAM[14446] = 8'b0;
    XRAM[14447] = 8'b0;
    XRAM[14448] = 8'b0;
    XRAM[14449] = 8'b0;
    XRAM[14450] = 8'b0;
    XRAM[14451] = 8'b0;
    XRAM[14452] = 8'b0;
    XRAM[14453] = 8'b0;
    XRAM[14454] = 8'b0;
    XRAM[14455] = 8'b0;
    XRAM[14456] = 8'b0;
    XRAM[14457] = 8'b0;
    XRAM[14458] = 8'b0;
    XRAM[14459] = 8'b0;
    XRAM[14460] = 8'b0;
    XRAM[14461] = 8'b0;
    XRAM[14462] = 8'b0;
    XRAM[14463] = 8'b0;
    XRAM[14464] = 8'b0;
    XRAM[14465] = 8'b0;
    XRAM[14466] = 8'b0;
    XRAM[14467] = 8'b0;
    XRAM[14468] = 8'b0;
    XRAM[14469] = 8'b0;
    XRAM[14470] = 8'b0;
    XRAM[14471] = 8'b0;
    XRAM[14472] = 8'b0;
    XRAM[14473] = 8'b0;
    XRAM[14474] = 8'b0;
    XRAM[14475] = 8'b0;
    XRAM[14476] = 8'b0;
    XRAM[14477] = 8'b0;
    XRAM[14478] = 8'b0;
    XRAM[14479] = 8'b0;
    XRAM[14480] = 8'b0;
    XRAM[14481] = 8'b0;
    XRAM[14482] = 8'b0;
    XRAM[14483] = 8'b0;
    XRAM[14484] = 8'b0;
    XRAM[14485] = 8'b0;
    XRAM[14486] = 8'b0;
    XRAM[14487] = 8'b0;
    XRAM[14488] = 8'b0;
    XRAM[14489] = 8'b0;
    XRAM[14490] = 8'b0;
    XRAM[14491] = 8'b0;
    XRAM[14492] = 8'b0;
    XRAM[14493] = 8'b0;
    XRAM[14494] = 8'b0;
    XRAM[14495] = 8'b0;
    XRAM[14496] = 8'b0;
    XRAM[14497] = 8'b0;
    XRAM[14498] = 8'b0;
    XRAM[14499] = 8'b0;
    XRAM[14500] = 8'b0;
    XRAM[14501] = 8'b0;
    XRAM[14502] = 8'b0;
    XRAM[14503] = 8'b0;
    XRAM[14504] = 8'b0;
    XRAM[14505] = 8'b0;
    XRAM[14506] = 8'b0;
    XRAM[14507] = 8'b0;
    XRAM[14508] = 8'b0;
    XRAM[14509] = 8'b0;
    XRAM[14510] = 8'b0;
    XRAM[14511] = 8'b0;
    XRAM[14512] = 8'b0;
    XRAM[14513] = 8'b0;
    XRAM[14514] = 8'b0;
    XRAM[14515] = 8'b0;
    XRAM[14516] = 8'b0;
    XRAM[14517] = 8'b0;
    XRAM[14518] = 8'b0;
    XRAM[14519] = 8'b0;
    XRAM[14520] = 8'b0;
    XRAM[14521] = 8'b0;
    XRAM[14522] = 8'b0;
    XRAM[14523] = 8'b0;
    XRAM[14524] = 8'b0;
    XRAM[14525] = 8'b0;
    XRAM[14526] = 8'b0;
    XRAM[14527] = 8'b0;
    XRAM[14528] = 8'b0;
    XRAM[14529] = 8'b0;
    XRAM[14530] = 8'b0;
    XRAM[14531] = 8'b0;
    XRAM[14532] = 8'b0;
    XRAM[14533] = 8'b0;
    XRAM[14534] = 8'b0;
    XRAM[14535] = 8'b0;
    XRAM[14536] = 8'b0;
    XRAM[14537] = 8'b0;
    XRAM[14538] = 8'b0;
    XRAM[14539] = 8'b0;
    XRAM[14540] = 8'b0;
    XRAM[14541] = 8'b0;
    XRAM[14542] = 8'b0;
    XRAM[14543] = 8'b0;
    XRAM[14544] = 8'b0;
    XRAM[14545] = 8'b0;
    XRAM[14546] = 8'b0;
    XRAM[14547] = 8'b0;
    XRAM[14548] = 8'b0;
    XRAM[14549] = 8'b0;
    XRAM[14550] = 8'b0;
    XRAM[14551] = 8'b0;
    XRAM[14552] = 8'b0;
    XRAM[14553] = 8'b0;
    XRAM[14554] = 8'b0;
    XRAM[14555] = 8'b0;
    XRAM[14556] = 8'b0;
    XRAM[14557] = 8'b0;
    XRAM[14558] = 8'b0;
    XRAM[14559] = 8'b0;
    XRAM[14560] = 8'b0;
    XRAM[14561] = 8'b0;
    XRAM[14562] = 8'b0;
    XRAM[14563] = 8'b0;
    XRAM[14564] = 8'b0;
    XRAM[14565] = 8'b0;
    XRAM[14566] = 8'b0;
    XRAM[14567] = 8'b0;
    XRAM[14568] = 8'b0;
    XRAM[14569] = 8'b0;
    XRAM[14570] = 8'b0;
    XRAM[14571] = 8'b0;
    XRAM[14572] = 8'b0;
    XRAM[14573] = 8'b0;
    XRAM[14574] = 8'b0;
    XRAM[14575] = 8'b0;
    XRAM[14576] = 8'b0;
    XRAM[14577] = 8'b0;
    XRAM[14578] = 8'b0;
    XRAM[14579] = 8'b0;
    XRAM[14580] = 8'b0;
    XRAM[14581] = 8'b0;
    XRAM[14582] = 8'b0;
    XRAM[14583] = 8'b0;
    XRAM[14584] = 8'b0;
    XRAM[14585] = 8'b0;
    XRAM[14586] = 8'b0;
    XRAM[14587] = 8'b0;
    XRAM[14588] = 8'b0;
    XRAM[14589] = 8'b0;
    XRAM[14590] = 8'b0;
    XRAM[14591] = 8'b0;
    XRAM[14592] = 8'b0;
    XRAM[14593] = 8'b0;
    XRAM[14594] = 8'b0;
    XRAM[14595] = 8'b0;
    XRAM[14596] = 8'b0;
    XRAM[14597] = 8'b0;
    XRAM[14598] = 8'b0;
    XRAM[14599] = 8'b0;
    XRAM[14600] = 8'b0;
    XRAM[14601] = 8'b0;
    XRAM[14602] = 8'b0;
    XRAM[14603] = 8'b0;
    XRAM[14604] = 8'b0;
    XRAM[14605] = 8'b0;
    XRAM[14606] = 8'b0;
    XRAM[14607] = 8'b0;
    XRAM[14608] = 8'b0;
    XRAM[14609] = 8'b0;
    XRAM[14610] = 8'b0;
    XRAM[14611] = 8'b0;
    XRAM[14612] = 8'b0;
    XRAM[14613] = 8'b0;
    XRAM[14614] = 8'b0;
    XRAM[14615] = 8'b0;
    XRAM[14616] = 8'b0;
    XRAM[14617] = 8'b0;
    XRAM[14618] = 8'b0;
    XRAM[14619] = 8'b0;
    XRAM[14620] = 8'b0;
    XRAM[14621] = 8'b0;
    XRAM[14622] = 8'b0;
    XRAM[14623] = 8'b0;
    XRAM[14624] = 8'b0;
    XRAM[14625] = 8'b0;
    XRAM[14626] = 8'b0;
    XRAM[14627] = 8'b0;
    XRAM[14628] = 8'b0;
    XRAM[14629] = 8'b0;
    XRAM[14630] = 8'b0;
    XRAM[14631] = 8'b0;
    XRAM[14632] = 8'b0;
    XRAM[14633] = 8'b0;
    XRAM[14634] = 8'b0;
    XRAM[14635] = 8'b0;
    XRAM[14636] = 8'b0;
    XRAM[14637] = 8'b0;
    XRAM[14638] = 8'b0;
    XRAM[14639] = 8'b0;
    XRAM[14640] = 8'b0;
    XRAM[14641] = 8'b0;
    XRAM[14642] = 8'b0;
    XRAM[14643] = 8'b0;
    XRAM[14644] = 8'b0;
    XRAM[14645] = 8'b0;
    XRAM[14646] = 8'b0;
    XRAM[14647] = 8'b0;
    XRAM[14648] = 8'b0;
    XRAM[14649] = 8'b0;
    XRAM[14650] = 8'b0;
    XRAM[14651] = 8'b0;
    XRAM[14652] = 8'b0;
    XRAM[14653] = 8'b0;
    XRAM[14654] = 8'b0;
    XRAM[14655] = 8'b0;
    XRAM[14656] = 8'b0;
    XRAM[14657] = 8'b0;
    XRAM[14658] = 8'b0;
    XRAM[14659] = 8'b0;
    XRAM[14660] = 8'b0;
    XRAM[14661] = 8'b0;
    XRAM[14662] = 8'b0;
    XRAM[14663] = 8'b0;
    XRAM[14664] = 8'b0;
    XRAM[14665] = 8'b0;
    XRAM[14666] = 8'b0;
    XRAM[14667] = 8'b0;
    XRAM[14668] = 8'b0;
    XRAM[14669] = 8'b0;
    XRAM[14670] = 8'b0;
    XRAM[14671] = 8'b0;
    XRAM[14672] = 8'b0;
    XRAM[14673] = 8'b0;
    XRAM[14674] = 8'b0;
    XRAM[14675] = 8'b0;
    XRAM[14676] = 8'b0;
    XRAM[14677] = 8'b0;
    XRAM[14678] = 8'b0;
    XRAM[14679] = 8'b0;
    XRAM[14680] = 8'b0;
    XRAM[14681] = 8'b0;
    XRAM[14682] = 8'b0;
    XRAM[14683] = 8'b0;
    XRAM[14684] = 8'b0;
    XRAM[14685] = 8'b0;
    XRAM[14686] = 8'b0;
    XRAM[14687] = 8'b0;
    XRAM[14688] = 8'b0;
    XRAM[14689] = 8'b0;
    XRAM[14690] = 8'b0;
    XRAM[14691] = 8'b0;
    XRAM[14692] = 8'b0;
    XRAM[14693] = 8'b0;
    XRAM[14694] = 8'b0;
    XRAM[14695] = 8'b0;
    XRAM[14696] = 8'b0;
    XRAM[14697] = 8'b0;
    XRAM[14698] = 8'b0;
    XRAM[14699] = 8'b0;
    XRAM[14700] = 8'b0;
    XRAM[14701] = 8'b0;
    XRAM[14702] = 8'b0;
    XRAM[14703] = 8'b0;
    XRAM[14704] = 8'b0;
    XRAM[14705] = 8'b0;
    XRAM[14706] = 8'b0;
    XRAM[14707] = 8'b0;
    XRAM[14708] = 8'b0;
    XRAM[14709] = 8'b0;
    XRAM[14710] = 8'b0;
    XRAM[14711] = 8'b0;
    XRAM[14712] = 8'b0;
    XRAM[14713] = 8'b0;
    XRAM[14714] = 8'b0;
    XRAM[14715] = 8'b0;
    XRAM[14716] = 8'b0;
    XRAM[14717] = 8'b0;
    XRAM[14718] = 8'b0;
    XRAM[14719] = 8'b0;
    XRAM[14720] = 8'b0;
    XRAM[14721] = 8'b0;
    XRAM[14722] = 8'b0;
    XRAM[14723] = 8'b0;
    XRAM[14724] = 8'b0;
    XRAM[14725] = 8'b0;
    XRAM[14726] = 8'b0;
    XRAM[14727] = 8'b0;
    XRAM[14728] = 8'b0;
    XRAM[14729] = 8'b0;
    XRAM[14730] = 8'b0;
    XRAM[14731] = 8'b0;
    XRAM[14732] = 8'b0;
    XRAM[14733] = 8'b0;
    XRAM[14734] = 8'b0;
    XRAM[14735] = 8'b0;
    XRAM[14736] = 8'b0;
    XRAM[14737] = 8'b0;
    XRAM[14738] = 8'b0;
    XRAM[14739] = 8'b0;
    XRAM[14740] = 8'b0;
    XRAM[14741] = 8'b0;
    XRAM[14742] = 8'b0;
    XRAM[14743] = 8'b0;
    XRAM[14744] = 8'b0;
    XRAM[14745] = 8'b0;
    XRAM[14746] = 8'b0;
    XRAM[14747] = 8'b0;
    XRAM[14748] = 8'b0;
    XRAM[14749] = 8'b0;
    XRAM[14750] = 8'b0;
    XRAM[14751] = 8'b0;
    XRAM[14752] = 8'b0;
    XRAM[14753] = 8'b0;
    XRAM[14754] = 8'b0;
    XRAM[14755] = 8'b0;
    XRAM[14756] = 8'b0;
    XRAM[14757] = 8'b0;
    XRAM[14758] = 8'b0;
    XRAM[14759] = 8'b0;
    XRAM[14760] = 8'b0;
    XRAM[14761] = 8'b0;
    XRAM[14762] = 8'b0;
    XRAM[14763] = 8'b0;
    XRAM[14764] = 8'b0;
    XRAM[14765] = 8'b0;
    XRAM[14766] = 8'b0;
    XRAM[14767] = 8'b0;
    XRAM[14768] = 8'b0;
    XRAM[14769] = 8'b0;
    XRAM[14770] = 8'b0;
    XRAM[14771] = 8'b0;
    XRAM[14772] = 8'b0;
    XRAM[14773] = 8'b0;
    XRAM[14774] = 8'b0;
    XRAM[14775] = 8'b0;
    XRAM[14776] = 8'b0;
    XRAM[14777] = 8'b0;
    XRAM[14778] = 8'b0;
    XRAM[14779] = 8'b0;
    XRAM[14780] = 8'b0;
    XRAM[14781] = 8'b0;
    XRAM[14782] = 8'b0;
    XRAM[14783] = 8'b0;
    XRAM[14784] = 8'b0;
    XRAM[14785] = 8'b0;
    XRAM[14786] = 8'b0;
    XRAM[14787] = 8'b0;
    XRAM[14788] = 8'b0;
    XRAM[14789] = 8'b0;
    XRAM[14790] = 8'b0;
    XRAM[14791] = 8'b0;
    XRAM[14792] = 8'b0;
    XRAM[14793] = 8'b0;
    XRAM[14794] = 8'b0;
    XRAM[14795] = 8'b0;
    XRAM[14796] = 8'b0;
    XRAM[14797] = 8'b0;
    XRAM[14798] = 8'b0;
    XRAM[14799] = 8'b0;
    XRAM[14800] = 8'b0;
    XRAM[14801] = 8'b0;
    XRAM[14802] = 8'b0;
    XRAM[14803] = 8'b0;
    XRAM[14804] = 8'b0;
    XRAM[14805] = 8'b0;
    XRAM[14806] = 8'b0;
    XRAM[14807] = 8'b0;
    XRAM[14808] = 8'b0;
    XRAM[14809] = 8'b0;
    XRAM[14810] = 8'b0;
    XRAM[14811] = 8'b0;
    XRAM[14812] = 8'b0;
    XRAM[14813] = 8'b0;
    XRAM[14814] = 8'b0;
    XRAM[14815] = 8'b0;
    XRAM[14816] = 8'b0;
    XRAM[14817] = 8'b0;
    XRAM[14818] = 8'b0;
    XRAM[14819] = 8'b0;
    XRAM[14820] = 8'b0;
    XRAM[14821] = 8'b0;
    XRAM[14822] = 8'b0;
    XRAM[14823] = 8'b0;
    XRAM[14824] = 8'b0;
    XRAM[14825] = 8'b0;
    XRAM[14826] = 8'b0;
    XRAM[14827] = 8'b0;
    XRAM[14828] = 8'b0;
    XRAM[14829] = 8'b0;
    XRAM[14830] = 8'b0;
    XRAM[14831] = 8'b0;
    XRAM[14832] = 8'b0;
    XRAM[14833] = 8'b0;
    XRAM[14834] = 8'b0;
    XRAM[14835] = 8'b0;
    XRAM[14836] = 8'b0;
    XRAM[14837] = 8'b0;
    XRAM[14838] = 8'b0;
    XRAM[14839] = 8'b0;
    XRAM[14840] = 8'b0;
    XRAM[14841] = 8'b0;
    XRAM[14842] = 8'b0;
    XRAM[14843] = 8'b0;
    XRAM[14844] = 8'b0;
    XRAM[14845] = 8'b0;
    XRAM[14846] = 8'b0;
    XRAM[14847] = 8'b0;
    XRAM[14848] = 8'b0;
    XRAM[14849] = 8'b0;
    XRAM[14850] = 8'b0;
    XRAM[14851] = 8'b0;
    XRAM[14852] = 8'b0;
    XRAM[14853] = 8'b0;
    XRAM[14854] = 8'b0;
    XRAM[14855] = 8'b0;
    XRAM[14856] = 8'b0;
    XRAM[14857] = 8'b0;
    XRAM[14858] = 8'b0;
    XRAM[14859] = 8'b0;
    XRAM[14860] = 8'b0;
    XRAM[14861] = 8'b0;
    XRAM[14862] = 8'b0;
    XRAM[14863] = 8'b0;
    XRAM[14864] = 8'b0;
    XRAM[14865] = 8'b0;
    XRAM[14866] = 8'b0;
    XRAM[14867] = 8'b0;
    XRAM[14868] = 8'b0;
    XRAM[14869] = 8'b0;
    XRAM[14870] = 8'b0;
    XRAM[14871] = 8'b0;
    XRAM[14872] = 8'b0;
    XRAM[14873] = 8'b0;
    XRAM[14874] = 8'b0;
    XRAM[14875] = 8'b0;
    XRAM[14876] = 8'b0;
    XRAM[14877] = 8'b0;
    XRAM[14878] = 8'b0;
    XRAM[14879] = 8'b0;
    XRAM[14880] = 8'b0;
    XRAM[14881] = 8'b0;
    XRAM[14882] = 8'b0;
    XRAM[14883] = 8'b0;
    XRAM[14884] = 8'b0;
    XRAM[14885] = 8'b0;
    XRAM[14886] = 8'b0;
    XRAM[14887] = 8'b0;
    XRAM[14888] = 8'b0;
    XRAM[14889] = 8'b0;
    XRAM[14890] = 8'b0;
    XRAM[14891] = 8'b0;
    XRAM[14892] = 8'b0;
    XRAM[14893] = 8'b0;
    XRAM[14894] = 8'b0;
    XRAM[14895] = 8'b0;
    XRAM[14896] = 8'b0;
    XRAM[14897] = 8'b0;
    XRAM[14898] = 8'b0;
    XRAM[14899] = 8'b0;
    XRAM[14900] = 8'b0;
    XRAM[14901] = 8'b0;
    XRAM[14902] = 8'b0;
    XRAM[14903] = 8'b0;
    XRAM[14904] = 8'b0;
    XRAM[14905] = 8'b0;
    XRAM[14906] = 8'b0;
    XRAM[14907] = 8'b0;
    XRAM[14908] = 8'b0;
    XRAM[14909] = 8'b0;
    XRAM[14910] = 8'b0;
    XRAM[14911] = 8'b0;
    XRAM[14912] = 8'b0;
    XRAM[14913] = 8'b0;
    XRAM[14914] = 8'b0;
    XRAM[14915] = 8'b0;
    XRAM[14916] = 8'b0;
    XRAM[14917] = 8'b0;
    XRAM[14918] = 8'b0;
    XRAM[14919] = 8'b0;
    XRAM[14920] = 8'b0;
    XRAM[14921] = 8'b0;
    XRAM[14922] = 8'b0;
    XRAM[14923] = 8'b0;
    XRAM[14924] = 8'b0;
    XRAM[14925] = 8'b0;
    XRAM[14926] = 8'b0;
    XRAM[14927] = 8'b0;
    XRAM[14928] = 8'b0;
    XRAM[14929] = 8'b0;
    XRAM[14930] = 8'b0;
    XRAM[14931] = 8'b0;
    XRAM[14932] = 8'b0;
    XRAM[14933] = 8'b0;
    XRAM[14934] = 8'b0;
    XRAM[14935] = 8'b0;
    XRAM[14936] = 8'b0;
    XRAM[14937] = 8'b0;
    XRAM[14938] = 8'b0;
    XRAM[14939] = 8'b0;
    XRAM[14940] = 8'b0;
    XRAM[14941] = 8'b0;
    XRAM[14942] = 8'b0;
    XRAM[14943] = 8'b0;
    XRAM[14944] = 8'b0;
    XRAM[14945] = 8'b0;
    XRAM[14946] = 8'b0;
    XRAM[14947] = 8'b0;
    XRAM[14948] = 8'b0;
    XRAM[14949] = 8'b0;
    XRAM[14950] = 8'b0;
    XRAM[14951] = 8'b0;
    XRAM[14952] = 8'b0;
    XRAM[14953] = 8'b0;
    XRAM[14954] = 8'b0;
    XRAM[14955] = 8'b0;
    XRAM[14956] = 8'b0;
    XRAM[14957] = 8'b0;
    XRAM[14958] = 8'b0;
    XRAM[14959] = 8'b0;
    XRAM[14960] = 8'b0;
    XRAM[14961] = 8'b0;
    XRAM[14962] = 8'b0;
    XRAM[14963] = 8'b0;
    XRAM[14964] = 8'b0;
    XRAM[14965] = 8'b0;
    XRAM[14966] = 8'b0;
    XRAM[14967] = 8'b0;
    XRAM[14968] = 8'b0;
    XRAM[14969] = 8'b0;
    XRAM[14970] = 8'b0;
    XRAM[14971] = 8'b0;
    XRAM[14972] = 8'b0;
    XRAM[14973] = 8'b0;
    XRAM[14974] = 8'b0;
    XRAM[14975] = 8'b0;
    XRAM[14976] = 8'b0;
    XRAM[14977] = 8'b0;
    XRAM[14978] = 8'b0;
    XRAM[14979] = 8'b0;
    XRAM[14980] = 8'b0;
    XRAM[14981] = 8'b0;
    XRAM[14982] = 8'b0;
    XRAM[14983] = 8'b0;
    XRAM[14984] = 8'b0;
    XRAM[14985] = 8'b0;
    XRAM[14986] = 8'b0;
    XRAM[14987] = 8'b0;
    XRAM[14988] = 8'b0;
    XRAM[14989] = 8'b0;
    XRAM[14990] = 8'b0;
    XRAM[14991] = 8'b0;
    XRAM[14992] = 8'b0;
    XRAM[14993] = 8'b0;
    XRAM[14994] = 8'b0;
    XRAM[14995] = 8'b0;
    XRAM[14996] = 8'b0;
    XRAM[14997] = 8'b0;
    XRAM[14998] = 8'b0;
    XRAM[14999] = 8'b0;
    XRAM[15000] = 8'b0;
    XRAM[15001] = 8'b0;
    XRAM[15002] = 8'b0;
    XRAM[15003] = 8'b0;
    XRAM[15004] = 8'b0;
    XRAM[15005] = 8'b0;
    XRAM[15006] = 8'b0;
    XRAM[15007] = 8'b0;
    XRAM[15008] = 8'b0;
    XRAM[15009] = 8'b0;
    XRAM[15010] = 8'b0;
    XRAM[15011] = 8'b0;
    XRAM[15012] = 8'b0;
    XRAM[15013] = 8'b0;
    XRAM[15014] = 8'b0;
    XRAM[15015] = 8'b0;
    XRAM[15016] = 8'b0;
    XRAM[15017] = 8'b0;
    XRAM[15018] = 8'b0;
    XRAM[15019] = 8'b0;
    XRAM[15020] = 8'b0;
    XRAM[15021] = 8'b0;
    XRAM[15022] = 8'b0;
    XRAM[15023] = 8'b0;
    XRAM[15024] = 8'b0;
    XRAM[15025] = 8'b0;
    XRAM[15026] = 8'b0;
    XRAM[15027] = 8'b0;
    XRAM[15028] = 8'b0;
    XRAM[15029] = 8'b0;
    XRAM[15030] = 8'b0;
    XRAM[15031] = 8'b0;
    XRAM[15032] = 8'b0;
    XRAM[15033] = 8'b0;
    XRAM[15034] = 8'b0;
    XRAM[15035] = 8'b0;
    XRAM[15036] = 8'b0;
    XRAM[15037] = 8'b0;
    XRAM[15038] = 8'b0;
    XRAM[15039] = 8'b0;
    XRAM[15040] = 8'b0;
    XRAM[15041] = 8'b0;
    XRAM[15042] = 8'b0;
    XRAM[15043] = 8'b0;
    XRAM[15044] = 8'b0;
    XRAM[15045] = 8'b0;
    XRAM[15046] = 8'b0;
    XRAM[15047] = 8'b0;
    XRAM[15048] = 8'b0;
    XRAM[15049] = 8'b0;
    XRAM[15050] = 8'b0;
    XRAM[15051] = 8'b0;
    XRAM[15052] = 8'b0;
    XRAM[15053] = 8'b0;
    XRAM[15054] = 8'b0;
    XRAM[15055] = 8'b0;
    XRAM[15056] = 8'b0;
    XRAM[15057] = 8'b0;
    XRAM[15058] = 8'b0;
    XRAM[15059] = 8'b0;
    XRAM[15060] = 8'b0;
    XRAM[15061] = 8'b0;
    XRAM[15062] = 8'b0;
    XRAM[15063] = 8'b0;
    XRAM[15064] = 8'b0;
    XRAM[15065] = 8'b0;
    XRAM[15066] = 8'b0;
    XRAM[15067] = 8'b0;
    XRAM[15068] = 8'b0;
    XRAM[15069] = 8'b0;
    XRAM[15070] = 8'b0;
    XRAM[15071] = 8'b0;
    XRAM[15072] = 8'b0;
    XRAM[15073] = 8'b0;
    XRAM[15074] = 8'b0;
    XRAM[15075] = 8'b0;
    XRAM[15076] = 8'b0;
    XRAM[15077] = 8'b0;
    XRAM[15078] = 8'b0;
    XRAM[15079] = 8'b0;
    XRAM[15080] = 8'b0;
    XRAM[15081] = 8'b0;
    XRAM[15082] = 8'b0;
    XRAM[15083] = 8'b0;
    XRAM[15084] = 8'b0;
    XRAM[15085] = 8'b0;
    XRAM[15086] = 8'b0;
    XRAM[15087] = 8'b0;
    XRAM[15088] = 8'b0;
    XRAM[15089] = 8'b0;
    XRAM[15090] = 8'b0;
    XRAM[15091] = 8'b0;
    XRAM[15092] = 8'b0;
    XRAM[15093] = 8'b0;
    XRAM[15094] = 8'b0;
    XRAM[15095] = 8'b0;
    XRAM[15096] = 8'b0;
    XRAM[15097] = 8'b0;
    XRAM[15098] = 8'b0;
    XRAM[15099] = 8'b0;
    XRAM[15100] = 8'b0;
    XRAM[15101] = 8'b0;
    XRAM[15102] = 8'b0;
    XRAM[15103] = 8'b0;
    XRAM[15104] = 8'b0;
    XRAM[15105] = 8'b0;
    XRAM[15106] = 8'b0;
    XRAM[15107] = 8'b0;
    XRAM[15108] = 8'b0;
    XRAM[15109] = 8'b0;
    XRAM[15110] = 8'b0;
    XRAM[15111] = 8'b0;
    XRAM[15112] = 8'b0;
    XRAM[15113] = 8'b0;
    XRAM[15114] = 8'b0;
    XRAM[15115] = 8'b0;
    XRAM[15116] = 8'b0;
    XRAM[15117] = 8'b0;
    XRAM[15118] = 8'b0;
    XRAM[15119] = 8'b0;
    XRAM[15120] = 8'b0;
    XRAM[15121] = 8'b0;
    XRAM[15122] = 8'b0;
    XRAM[15123] = 8'b0;
    XRAM[15124] = 8'b0;
    XRAM[15125] = 8'b0;
    XRAM[15126] = 8'b0;
    XRAM[15127] = 8'b0;
    XRAM[15128] = 8'b0;
    XRAM[15129] = 8'b0;
    XRAM[15130] = 8'b0;
    XRAM[15131] = 8'b0;
    XRAM[15132] = 8'b0;
    XRAM[15133] = 8'b0;
    XRAM[15134] = 8'b0;
    XRAM[15135] = 8'b0;
    XRAM[15136] = 8'b0;
    XRAM[15137] = 8'b0;
    XRAM[15138] = 8'b0;
    XRAM[15139] = 8'b0;
    XRAM[15140] = 8'b0;
    XRAM[15141] = 8'b0;
    XRAM[15142] = 8'b0;
    XRAM[15143] = 8'b0;
    XRAM[15144] = 8'b0;
    XRAM[15145] = 8'b0;
    XRAM[15146] = 8'b0;
    XRAM[15147] = 8'b0;
    XRAM[15148] = 8'b0;
    XRAM[15149] = 8'b0;
    XRAM[15150] = 8'b0;
    XRAM[15151] = 8'b0;
    XRAM[15152] = 8'b0;
    XRAM[15153] = 8'b0;
    XRAM[15154] = 8'b0;
    XRAM[15155] = 8'b0;
    XRAM[15156] = 8'b0;
    XRAM[15157] = 8'b0;
    XRAM[15158] = 8'b0;
    XRAM[15159] = 8'b0;
    XRAM[15160] = 8'b0;
    XRAM[15161] = 8'b0;
    XRAM[15162] = 8'b0;
    XRAM[15163] = 8'b0;
    XRAM[15164] = 8'b0;
    XRAM[15165] = 8'b0;
    XRAM[15166] = 8'b0;
    XRAM[15167] = 8'b0;
    XRAM[15168] = 8'b0;
    XRAM[15169] = 8'b0;
    XRAM[15170] = 8'b0;
    XRAM[15171] = 8'b0;
    XRAM[15172] = 8'b0;
    XRAM[15173] = 8'b0;
    XRAM[15174] = 8'b0;
    XRAM[15175] = 8'b0;
    XRAM[15176] = 8'b0;
    XRAM[15177] = 8'b0;
    XRAM[15178] = 8'b0;
    XRAM[15179] = 8'b0;
    XRAM[15180] = 8'b0;
    XRAM[15181] = 8'b0;
    XRAM[15182] = 8'b0;
    XRAM[15183] = 8'b0;
    XRAM[15184] = 8'b0;
    XRAM[15185] = 8'b0;
    XRAM[15186] = 8'b0;
    XRAM[15187] = 8'b0;
    XRAM[15188] = 8'b0;
    XRAM[15189] = 8'b0;
    XRAM[15190] = 8'b0;
    XRAM[15191] = 8'b0;
    XRAM[15192] = 8'b0;
    XRAM[15193] = 8'b0;
    XRAM[15194] = 8'b0;
    XRAM[15195] = 8'b0;
    XRAM[15196] = 8'b0;
    XRAM[15197] = 8'b0;
    XRAM[15198] = 8'b0;
    XRAM[15199] = 8'b0;
    XRAM[15200] = 8'b0;
    XRAM[15201] = 8'b0;
    XRAM[15202] = 8'b0;
    XRAM[15203] = 8'b0;
    XRAM[15204] = 8'b0;
    XRAM[15205] = 8'b0;
    XRAM[15206] = 8'b0;
    XRAM[15207] = 8'b0;
    XRAM[15208] = 8'b0;
    XRAM[15209] = 8'b0;
    XRAM[15210] = 8'b0;
    XRAM[15211] = 8'b0;
    XRAM[15212] = 8'b0;
    XRAM[15213] = 8'b0;
    XRAM[15214] = 8'b0;
    XRAM[15215] = 8'b0;
    XRAM[15216] = 8'b0;
    XRAM[15217] = 8'b0;
    XRAM[15218] = 8'b0;
    XRAM[15219] = 8'b0;
    XRAM[15220] = 8'b0;
    XRAM[15221] = 8'b0;
    XRAM[15222] = 8'b0;
    XRAM[15223] = 8'b0;
    XRAM[15224] = 8'b0;
    XRAM[15225] = 8'b0;
    XRAM[15226] = 8'b0;
    XRAM[15227] = 8'b0;
    XRAM[15228] = 8'b0;
    XRAM[15229] = 8'b0;
    XRAM[15230] = 8'b0;
    XRAM[15231] = 8'b0;
    XRAM[15232] = 8'b0;
    XRAM[15233] = 8'b0;
    XRAM[15234] = 8'b0;
    XRAM[15235] = 8'b0;
    XRAM[15236] = 8'b0;
    XRAM[15237] = 8'b0;
    XRAM[15238] = 8'b0;
    XRAM[15239] = 8'b0;
    XRAM[15240] = 8'b0;
    XRAM[15241] = 8'b0;
    XRAM[15242] = 8'b0;
    XRAM[15243] = 8'b0;
    XRAM[15244] = 8'b0;
    XRAM[15245] = 8'b0;
    XRAM[15246] = 8'b0;
    XRAM[15247] = 8'b0;
    XRAM[15248] = 8'b0;
    XRAM[15249] = 8'b0;
    XRAM[15250] = 8'b0;
    XRAM[15251] = 8'b0;
    XRAM[15252] = 8'b0;
    XRAM[15253] = 8'b0;
    XRAM[15254] = 8'b0;
    XRAM[15255] = 8'b0;
    XRAM[15256] = 8'b0;
    XRAM[15257] = 8'b0;
    XRAM[15258] = 8'b0;
    XRAM[15259] = 8'b0;
    XRAM[15260] = 8'b0;
    XRAM[15261] = 8'b0;
    XRAM[15262] = 8'b0;
    XRAM[15263] = 8'b0;
    XRAM[15264] = 8'b0;
    XRAM[15265] = 8'b0;
    XRAM[15266] = 8'b0;
    XRAM[15267] = 8'b0;
    XRAM[15268] = 8'b0;
    XRAM[15269] = 8'b0;
    XRAM[15270] = 8'b0;
    XRAM[15271] = 8'b0;
    XRAM[15272] = 8'b0;
    XRAM[15273] = 8'b0;
    XRAM[15274] = 8'b0;
    XRAM[15275] = 8'b0;
    XRAM[15276] = 8'b0;
    XRAM[15277] = 8'b0;
    XRAM[15278] = 8'b0;
    XRAM[15279] = 8'b0;
    XRAM[15280] = 8'b0;
    XRAM[15281] = 8'b0;
    XRAM[15282] = 8'b0;
    XRAM[15283] = 8'b0;
    XRAM[15284] = 8'b0;
    XRAM[15285] = 8'b0;
    XRAM[15286] = 8'b0;
    XRAM[15287] = 8'b0;
    XRAM[15288] = 8'b0;
    XRAM[15289] = 8'b0;
    XRAM[15290] = 8'b0;
    XRAM[15291] = 8'b0;
    XRAM[15292] = 8'b0;
    XRAM[15293] = 8'b0;
    XRAM[15294] = 8'b0;
    XRAM[15295] = 8'b0;
    XRAM[15296] = 8'b0;
    XRAM[15297] = 8'b0;
    XRAM[15298] = 8'b0;
    XRAM[15299] = 8'b0;
    XRAM[15300] = 8'b0;
    XRAM[15301] = 8'b0;
    XRAM[15302] = 8'b0;
    XRAM[15303] = 8'b0;
    XRAM[15304] = 8'b0;
    XRAM[15305] = 8'b0;
    XRAM[15306] = 8'b0;
    XRAM[15307] = 8'b0;
    XRAM[15308] = 8'b0;
    XRAM[15309] = 8'b0;
    XRAM[15310] = 8'b0;
    XRAM[15311] = 8'b0;
    XRAM[15312] = 8'b0;
    XRAM[15313] = 8'b0;
    XRAM[15314] = 8'b0;
    XRAM[15315] = 8'b0;
    XRAM[15316] = 8'b0;
    XRAM[15317] = 8'b0;
    XRAM[15318] = 8'b0;
    XRAM[15319] = 8'b0;
    XRAM[15320] = 8'b0;
    XRAM[15321] = 8'b0;
    XRAM[15322] = 8'b0;
    XRAM[15323] = 8'b0;
    XRAM[15324] = 8'b0;
    XRAM[15325] = 8'b0;
    XRAM[15326] = 8'b0;
    XRAM[15327] = 8'b0;
    XRAM[15328] = 8'b0;
    XRAM[15329] = 8'b0;
    XRAM[15330] = 8'b0;
    XRAM[15331] = 8'b0;
    XRAM[15332] = 8'b0;
    XRAM[15333] = 8'b0;
    XRAM[15334] = 8'b0;
    XRAM[15335] = 8'b0;
    XRAM[15336] = 8'b0;
    XRAM[15337] = 8'b0;
    XRAM[15338] = 8'b0;
    XRAM[15339] = 8'b0;
    XRAM[15340] = 8'b0;
    XRAM[15341] = 8'b0;
    XRAM[15342] = 8'b0;
    XRAM[15343] = 8'b0;
    XRAM[15344] = 8'b0;
    XRAM[15345] = 8'b0;
    XRAM[15346] = 8'b0;
    XRAM[15347] = 8'b0;
    XRAM[15348] = 8'b0;
    XRAM[15349] = 8'b0;
    XRAM[15350] = 8'b0;
    XRAM[15351] = 8'b0;
    XRAM[15352] = 8'b0;
    XRAM[15353] = 8'b0;
    XRAM[15354] = 8'b0;
    XRAM[15355] = 8'b0;
    XRAM[15356] = 8'b0;
    XRAM[15357] = 8'b0;
    XRAM[15358] = 8'b0;
    XRAM[15359] = 8'b0;
    XRAM[15360] = 8'b0;
    XRAM[15361] = 8'b0;
    XRAM[15362] = 8'b0;
    XRAM[15363] = 8'b0;
    XRAM[15364] = 8'b0;
    XRAM[15365] = 8'b0;
    XRAM[15366] = 8'b0;
    XRAM[15367] = 8'b0;
    XRAM[15368] = 8'b0;
    XRAM[15369] = 8'b0;
    XRAM[15370] = 8'b0;
    XRAM[15371] = 8'b0;
    XRAM[15372] = 8'b0;
    XRAM[15373] = 8'b0;
    XRAM[15374] = 8'b0;
    XRAM[15375] = 8'b0;
    XRAM[15376] = 8'b0;
    XRAM[15377] = 8'b0;
    XRAM[15378] = 8'b0;
    XRAM[15379] = 8'b0;
    XRAM[15380] = 8'b0;
    XRAM[15381] = 8'b0;
    XRAM[15382] = 8'b0;
    XRAM[15383] = 8'b0;
    XRAM[15384] = 8'b0;
    XRAM[15385] = 8'b0;
    XRAM[15386] = 8'b0;
    XRAM[15387] = 8'b0;
    XRAM[15388] = 8'b0;
    XRAM[15389] = 8'b0;
    XRAM[15390] = 8'b0;
    XRAM[15391] = 8'b0;
    XRAM[15392] = 8'b0;
    XRAM[15393] = 8'b0;
    XRAM[15394] = 8'b0;
    XRAM[15395] = 8'b0;
    XRAM[15396] = 8'b0;
    XRAM[15397] = 8'b0;
    XRAM[15398] = 8'b0;
    XRAM[15399] = 8'b0;
    XRAM[15400] = 8'b0;
    XRAM[15401] = 8'b0;
    XRAM[15402] = 8'b0;
    XRAM[15403] = 8'b0;
    XRAM[15404] = 8'b0;
    XRAM[15405] = 8'b0;
    XRAM[15406] = 8'b0;
    XRAM[15407] = 8'b0;
    XRAM[15408] = 8'b0;
    XRAM[15409] = 8'b0;
    XRAM[15410] = 8'b0;
    XRAM[15411] = 8'b0;
    XRAM[15412] = 8'b0;
    XRAM[15413] = 8'b0;
    XRAM[15414] = 8'b0;
    XRAM[15415] = 8'b0;
    XRAM[15416] = 8'b0;
    XRAM[15417] = 8'b0;
    XRAM[15418] = 8'b0;
    XRAM[15419] = 8'b0;
    XRAM[15420] = 8'b0;
    XRAM[15421] = 8'b0;
    XRAM[15422] = 8'b0;
    XRAM[15423] = 8'b0;
    XRAM[15424] = 8'b0;
    XRAM[15425] = 8'b0;
    XRAM[15426] = 8'b0;
    XRAM[15427] = 8'b0;
    XRAM[15428] = 8'b0;
    XRAM[15429] = 8'b0;
    XRAM[15430] = 8'b0;
    XRAM[15431] = 8'b0;
    XRAM[15432] = 8'b0;
    XRAM[15433] = 8'b0;
    XRAM[15434] = 8'b0;
    XRAM[15435] = 8'b0;
    XRAM[15436] = 8'b0;
    XRAM[15437] = 8'b0;
    XRAM[15438] = 8'b0;
    XRAM[15439] = 8'b0;
    XRAM[15440] = 8'b0;
    XRAM[15441] = 8'b0;
    XRAM[15442] = 8'b0;
    XRAM[15443] = 8'b0;
    XRAM[15444] = 8'b0;
    XRAM[15445] = 8'b0;
    XRAM[15446] = 8'b0;
    XRAM[15447] = 8'b0;
    XRAM[15448] = 8'b0;
    XRAM[15449] = 8'b0;
    XRAM[15450] = 8'b0;
    XRAM[15451] = 8'b0;
    XRAM[15452] = 8'b0;
    XRAM[15453] = 8'b0;
    XRAM[15454] = 8'b0;
    XRAM[15455] = 8'b0;
    XRAM[15456] = 8'b0;
    XRAM[15457] = 8'b0;
    XRAM[15458] = 8'b0;
    XRAM[15459] = 8'b0;
    XRAM[15460] = 8'b0;
    XRAM[15461] = 8'b0;
    XRAM[15462] = 8'b0;
    XRAM[15463] = 8'b0;
    XRAM[15464] = 8'b0;
    XRAM[15465] = 8'b0;
    XRAM[15466] = 8'b0;
    XRAM[15467] = 8'b0;
    XRAM[15468] = 8'b0;
    XRAM[15469] = 8'b0;
    XRAM[15470] = 8'b0;
    XRAM[15471] = 8'b0;
    XRAM[15472] = 8'b0;
    XRAM[15473] = 8'b0;
    XRAM[15474] = 8'b0;
    XRAM[15475] = 8'b0;
    XRAM[15476] = 8'b0;
    XRAM[15477] = 8'b0;
    XRAM[15478] = 8'b0;
    XRAM[15479] = 8'b0;
    XRAM[15480] = 8'b0;
    XRAM[15481] = 8'b0;
    XRAM[15482] = 8'b0;
    XRAM[15483] = 8'b0;
    XRAM[15484] = 8'b0;
    XRAM[15485] = 8'b0;
    XRAM[15486] = 8'b0;
    XRAM[15487] = 8'b0;
    XRAM[15488] = 8'b0;
    XRAM[15489] = 8'b0;
    XRAM[15490] = 8'b0;
    XRAM[15491] = 8'b0;
    XRAM[15492] = 8'b0;
    XRAM[15493] = 8'b0;
    XRAM[15494] = 8'b0;
    XRAM[15495] = 8'b0;
    XRAM[15496] = 8'b0;
    XRAM[15497] = 8'b0;
    XRAM[15498] = 8'b0;
    XRAM[15499] = 8'b0;
    XRAM[15500] = 8'b0;
    XRAM[15501] = 8'b0;
    XRAM[15502] = 8'b0;
    XRAM[15503] = 8'b0;
    XRAM[15504] = 8'b0;
    XRAM[15505] = 8'b0;
    XRAM[15506] = 8'b0;
    XRAM[15507] = 8'b0;
    XRAM[15508] = 8'b0;
    XRAM[15509] = 8'b0;
    XRAM[15510] = 8'b0;
    XRAM[15511] = 8'b0;
    XRAM[15512] = 8'b0;
    XRAM[15513] = 8'b0;
    XRAM[15514] = 8'b0;
    XRAM[15515] = 8'b0;
    XRAM[15516] = 8'b0;
    XRAM[15517] = 8'b0;
    XRAM[15518] = 8'b0;
    XRAM[15519] = 8'b0;
    XRAM[15520] = 8'b0;
    XRAM[15521] = 8'b0;
    XRAM[15522] = 8'b0;
    XRAM[15523] = 8'b0;
    XRAM[15524] = 8'b0;
    XRAM[15525] = 8'b0;
    XRAM[15526] = 8'b0;
    XRAM[15527] = 8'b0;
    XRAM[15528] = 8'b0;
    XRAM[15529] = 8'b0;
    XRAM[15530] = 8'b0;
    XRAM[15531] = 8'b0;
    XRAM[15532] = 8'b0;
    XRAM[15533] = 8'b0;
    XRAM[15534] = 8'b0;
    XRAM[15535] = 8'b0;
    XRAM[15536] = 8'b0;
    XRAM[15537] = 8'b0;
    XRAM[15538] = 8'b0;
    XRAM[15539] = 8'b0;
    XRAM[15540] = 8'b0;
    XRAM[15541] = 8'b0;
    XRAM[15542] = 8'b0;
    XRAM[15543] = 8'b0;
    XRAM[15544] = 8'b0;
    XRAM[15545] = 8'b0;
    XRAM[15546] = 8'b0;
    XRAM[15547] = 8'b0;
    XRAM[15548] = 8'b0;
    XRAM[15549] = 8'b0;
    XRAM[15550] = 8'b0;
    XRAM[15551] = 8'b0;
    XRAM[15552] = 8'b0;
    XRAM[15553] = 8'b0;
    XRAM[15554] = 8'b0;
    XRAM[15555] = 8'b0;
    XRAM[15556] = 8'b0;
    XRAM[15557] = 8'b0;
    XRAM[15558] = 8'b0;
    XRAM[15559] = 8'b0;
    XRAM[15560] = 8'b0;
    XRAM[15561] = 8'b0;
    XRAM[15562] = 8'b0;
    XRAM[15563] = 8'b0;
    XRAM[15564] = 8'b0;
    XRAM[15565] = 8'b0;
    XRAM[15566] = 8'b0;
    XRAM[15567] = 8'b0;
    XRAM[15568] = 8'b0;
    XRAM[15569] = 8'b0;
    XRAM[15570] = 8'b0;
    XRAM[15571] = 8'b0;
    XRAM[15572] = 8'b0;
    XRAM[15573] = 8'b0;
    XRAM[15574] = 8'b0;
    XRAM[15575] = 8'b0;
    XRAM[15576] = 8'b0;
    XRAM[15577] = 8'b0;
    XRAM[15578] = 8'b0;
    XRAM[15579] = 8'b0;
    XRAM[15580] = 8'b0;
    XRAM[15581] = 8'b0;
    XRAM[15582] = 8'b0;
    XRAM[15583] = 8'b0;
    XRAM[15584] = 8'b0;
    XRAM[15585] = 8'b0;
    XRAM[15586] = 8'b0;
    XRAM[15587] = 8'b0;
    XRAM[15588] = 8'b0;
    XRAM[15589] = 8'b0;
    XRAM[15590] = 8'b0;
    XRAM[15591] = 8'b0;
    XRAM[15592] = 8'b0;
    XRAM[15593] = 8'b0;
    XRAM[15594] = 8'b0;
    XRAM[15595] = 8'b0;
    XRAM[15596] = 8'b0;
    XRAM[15597] = 8'b0;
    XRAM[15598] = 8'b0;
    XRAM[15599] = 8'b0;
    XRAM[15600] = 8'b0;
    XRAM[15601] = 8'b0;
    XRAM[15602] = 8'b0;
    XRAM[15603] = 8'b0;
    XRAM[15604] = 8'b0;
    XRAM[15605] = 8'b0;
    XRAM[15606] = 8'b0;
    XRAM[15607] = 8'b0;
    XRAM[15608] = 8'b0;
    XRAM[15609] = 8'b0;
    XRAM[15610] = 8'b0;
    XRAM[15611] = 8'b0;
    XRAM[15612] = 8'b0;
    XRAM[15613] = 8'b0;
    XRAM[15614] = 8'b0;
    XRAM[15615] = 8'b0;
    XRAM[15616] = 8'b0;
    XRAM[15617] = 8'b0;
    XRAM[15618] = 8'b0;
    XRAM[15619] = 8'b0;
    XRAM[15620] = 8'b0;
    XRAM[15621] = 8'b0;
    XRAM[15622] = 8'b0;
    XRAM[15623] = 8'b0;
    XRAM[15624] = 8'b0;
    XRAM[15625] = 8'b0;
    XRAM[15626] = 8'b0;
    XRAM[15627] = 8'b0;
    XRAM[15628] = 8'b0;
    XRAM[15629] = 8'b0;
    XRAM[15630] = 8'b0;
    XRAM[15631] = 8'b0;
    XRAM[15632] = 8'b0;
    XRAM[15633] = 8'b0;
    XRAM[15634] = 8'b0;
    XRAM[15635] = 8'b0;
    XRAM[15636] = 8'b0;
    XRAM[15637] = 8'b0;
    XRAM[15638] = 8'b0;
    XRAM[15639] = 8'b0;
    XRAM[15640] = 8'b0;
    XRAM[15641] = 8'b0;
    XRAM[15642] = 8'b0;
    XRAM[15643] = 8'b0;
    XRAM[15644] = 8'b0;
    XRAM[15645] = 8'b0;
    XRAM[15646] = 8'b0;
    XRAM[15647] = 8'b0;
    XRAM[15648] = 8'b0;
    XRAM[15649] = 8'b0;
    XRAM[15650] = 8'b0;
    XRAM[15651] = 8'b0;
    XRAM[15652] = 8'b0;
    XRAM[15653] = 8'b0;
    XRAM[15654] = 8'b0;
    XRAM[15655] = 8'b0;
    XRAM[15656] = 8'b0;
    XRAM[15657] = 8'b0;
    XRAM[15658] = 8'b0;
    XRAM[15659] = 8'b0;
    XRAM[15660] = 8'b0;
    XRAM[15661] = 8'b0;
    XRAM[15662] = 8'b0;
    XRAM[15663] = 8'b0;
    XRAM[15664] = 8'b0;
    XRAM[15665] = 8'b0;
    XRAM[15666] = 8'b0;
    XRAM[15667] = 8'b0;
    XRAM[15668] = 8'b0;
    XRAM[15669] = 8'b0;
    XRAM[15670] = 8'b0;
    XRAM[15671] = 8'b0;
    XRAM[15672] = 8'b0;
    XRAM[15673] = 8'b0;
    XRAM[15674] = 8'b0;
    XRAM[15675] = 8'b0;
    XRAM[15676] = 8'b0;
    XRAM[15677] = 8'b0;
    XRAM[15678] = 8'b0;
    XRAM[15679] = 8'b0;
    XRAM[15680] = 8'b0;
    XRAM[15681] = 8'b0;
    XRAM[15682] = 8'b0;
    XRAM[15683] = 8'b0;
    XRAM[15684] = 8'b0;
    XRAM[15685] = 8'b0;
    XRAM[15686] = 8'b0;
    XRAM[15687] = 8'b0;
    XRAM[15688] = 8'b0;
    XRAM[15689] = 8'b0;
    XRAM[15690] = 8'b0;
    XRAM[15691] = 8'b0;
    XRAM[15692] = 8'b0;
    XRAM[15693] = 8'b0;
    XRAM[15694] = 8'b0;
    XRAM[15695] = 8'b0;
    XRAM[15696] = 8'b0;
    XRAM[15697] = 8'b0;
    XRAM[15698] = 8'b0;
    XRAM[15699] = 8'b0;
    XRAM[15700] = 8'b0;
    XRAM[15701] = 8'b0;
    XRAM[15702] = 8'b0;
    XRAM[15703] = 8'b0;
    XRAM[15704] = 8'b0;
    XRAM[15705] = 8'b0;
    XRAM[15706] = 8'b0;
    XRAM[15707] = 8'b0;
    XRAM[15708] = 8'b0;
    XRAM[15709] = 8'b0;
    XRAM[15710] = 8'b0;
    XRAM[15711] = 8'b0;
    XRAM[15712] = 8'b0;
    XRAM[15713] = 8'b0;
    XRAM[15714] = 8'b0;
    XRAM[15715] = 8'b0;
    XRAM[15716] = 8'b0;
    XRAM[15717] = 8'b0;
    XRAM[15718] = 8'b0;
    XRAM[15719] = 8'b0;
    XRAM[15720] = 8'b0;
    XRAM[15721] = 8'b0;
    XRAM[15722] = 8'b0;
    XRAM[15723] = 8'b0;
    XRAM[15724] = 8'b0;
    XRAM[15725] = 8'b0;
    XRAM[15726] = 8'b0;
    XRAM[15727] = 8'b0;
    XRAM[15728] = 8'b0;
    XRAM[15729] = 8'b0;
    XRAM[15730] = 8'b0;
    XRAM[15731] = 8'b0;
    XRAM[15732] = 8'b0;
    XRAM[15733] = 8'b0;
    XRAM[15734] = 8'b0;
    XRAM[15735] = 8'b0;
    XRAM[15736] = 8'b0;
    XRAM[15737] = 8'b0;
    XRAM[15738] = 8'b0;
    XRAM[15739] = 8'b0;
    XRAM[15740] = 8'b0;
    XRAM[15741] = 8'b0;
    XRAM[15742] = 8'b0;
    XRAM[15743] = 8'b0;
    XRAM[15744] = 8'b0;
    XRAM[15745] = 8'b0;
    XRAM[15746] = 8'b0;
    XRAM[15747] = 8'b0;
    XRAM[15748] = 8'b0;
    XRAM[15749] = 8'b0;
    XRAM[15750] = 8'b0;
    XRAM[15751] = 8'b0;
    XRAM[15752] = 8'b0;
    XRAM[15753] = 8'b0;
    XRAM[15754] = 8'b0;
    XRAM[15755] = 8'b0;
    XRAM[15756] = 8'b0;
    XRAM[15757] = 8'b0;
    XRAM[15758] = 8'b0;
    XRAM[15759] = 8'b0;
    XRAM[15760] = 8'b0;
    XRAM[15761] = 8'b0;
    XRAM[15762] = 8'b0;
    XRAM[15763] = 8'b0;
    XRAM[15764] = 8'b0;
    XRAM[15765] = 8'b0;
    XRAM[15766] = 8'b0;
    XRAM[15767] = 8'b0;
    XRAM[15768] = 8'b0;
    XRAM[15769] = 8'b0;
    XRAM[15770] = 8'b0;
    XRAM[15771] = 8'b0;
    XRAM[15772] = 8'b0;
    XRAM[15773] = 8'b0;
    XRAM[15774] = 8'b0;
    XRAM[15775] = 8'b0;
    XRAM[15776] = 8'b0;
    XRAM[15777] = 8'b0;
    XRAM[15778] = 8'b0;
    XRAM[15779] = 8'b0;
    XRAM[15780] = 8'b0;
    XRAM[15781] = 8'b0;
    XRAM[15782] = 8'b0;
    XRAM[15783] = 8'b0;
    XRAM[15784] = 8'b0;
    XRAM[15785] = 8'b0;
    XRAM[15786] = 8'b0;
    XRAM[15787] = 8'b0;
    XRAM[15788] = 8'b0;
    XRAM[15789] = 8'b0;
    XRAM[15790] = 8'b0;
    XRAM[15791] = 8'b0;
    XRAM[15792] = 8'b0;
    XRAM[15793] = 8'b0;
    XRAM[15794] = 8'b0;
    XRAM[15795] = 8'b0;
    XRAM[15796] = 8'b0;
    XRAM[15797] = 8'b0;
    XRAM[15798] = 8'b0;
    XRAM[15799] = 8'b0;
    XRAM[15800] = 8'b0;
    XRAM[15801] = 8'b0;
    XRAM[15802] = 8'b0;
    XRAM[15803] = 8'b0;
    XRAM[15804] = 8'b0;
    XRAM[15805] = 8'b0;
    XRAM[15806] = 8'b0;
    XRAM[15807] = 8'b0;
    XRAM[15808] = 8'b0;
    XRAM[15809] = 8'b0;
    XRAM[15810] = 8'b0;
    XRAM[15811] = 8'b0;
    XRAM[15812] = 8'b0;
    XRAM[15813] = 8'b0;
    XRAM[15814] = 8'b0;
    XRAM[15815] = 8'b0;
    XRAM[15816] = 8'b0;
    XRAM[15817] = 8'b0;
    XRAM[15818] = 8'b0;
    XRAM[15819] = 8'b0;
    XRAM[15820] = 8'b0;
    XRAM[15821] = 8'b0;
    XRAM[15822] = 8'b0;
    XRAM[15823] = 8'b0;
    XRAM[15824] = 8'b0;
    XRAM[15825] = 8'b0;
    XRAM[15826] = 8'b0;
    XRAM[15827] = 8'b0;
    XRAM[15828] = 8'b0;
    XRAM[15829] = 8'b0;
    XRAM[15830] = 8'b0;
    XRAM[15831] = 8'b0;
    XRAM[15832] = 8'b0;
    XRAM[15833] = 8'b0;
    XRAM[15834] = 8'b0;
    XRAM[15835] = 8'b0;
    XRAM[15836] = 8'b0;
    XRAM[15837] = 8'b0;
    XRAM[15838] = 8'b0;
    XRAM[15839] = 8'b0;
    XRAM[15840] = 8'b0;
    XRAM[15841] = 8'b0;
    XRAM[15842] = 8'b0;
    XRAM[15843] = 8'b0;
    XRAM[15844] = 8'b0;
    XRAM[15845] = 8'b0;
    XRAM[15846] = 8'b0;
    XRAM[15847] = 8'b0;
    XRAM[15848] = 8'b0;
    XRAM[15849] = 8'b0;
    XRAM[15850] = 8'b0;
    XRAM[15851] = 8'b0;
    XRAM[15852] = 8'b0;
    XRAM[15853] = 8'b0;
    XRAM[15854] = 8'b0;
    XRAM[15855] = 8'b0;
    XRAM[15856] = 8'b0;
    XRAM[15857] = 8'b0;
    XRAM[15858] = 8'b0;
    XRAM[15859] = 8'b0;
    XRAM[15860] = 8'b0;
    XRAM[15861] = 8'b0;
    XRAM[15862] = 8'b0;
    XRAM[15863] = 8'b0;
    XRAM[15864] = 8'b0;
    XRAM[15865] = 8'b0;
    XRAM[15866] = 8'b0;
    XRAM[15867] = 8'b0;
    XRAM[15868] = 8'b0;
    XRAM[15869] = 8'b0;
    XRAM[15870] = 8'b0;
    XRAM[15871] = 8'b0;
    XRAM[15872] = 8'b0;
    XRAM[15873] = 8'b0;
    XRAM[15874] = 8'b0;
    XRAM[15875] = 8'b0;
    XRAM[15876] = 8'b0;
    XRAM[15877] = 8'b0;
    XRAM[15878] = 8'b0;
    XRAM[15879] = 8'b0;
    XRAM[15880] = 8'b0;
    XRAM[15881] = 8'b0;
    XRAM[15882] = 8'b0;
    XRAM[15883] = 8'b0;
    XRAM[15884] = 8'b0;
    XRAM[15885] = 8'b0;
    XRAM[15886] = 8'b0;
    XRAM[15887] = 8'b0;
    XRAM[15888] = 8'b0;
    XRAM[15889] = 8'b0;
    XRAM[15890] = 8'b0;
    XRAM[15891] = 8'b0;
    XRAM[15892] = 8'b0;
    XRAM[15893] = 8'b0;
    XRAM[15894] = 8'b0;
    XRAM[15895] = 8'b0;
    XRAM[15896] = 8'b0;
    XRAM[15897] = 8'b0;
    XRAM[15898] = 8'b0;
    XRAM[15899] = 8'b0;
    XRAM[15900] = 8'b0;
    XRAM[15901] = 8'b0;
    XRAM[15902] = 8'b0;
    XRAM[15903] = 8'b0;
    XRAM[15904] = 8'b0;
    XRAM[15905] = 8'b0;
    XRAM[15906] = 8'b0;
    XRAM[15907] = 8'b0;
    XRAM[15908] = 8'b0;
    XRAM[15909] = 8'b0;
    XRAM[15910] = 8'b0;
    XRAM[15911] = 8'b0;
    XRAM[15912] = 8'b0;
    XRAM[15913] = 8'b0;
    XRAM[15914] = 8'b0;
    XRAM[15915] = 8'b0;
    XRAM[15916] = 8'b0;
    XRAM[15917] = 8'b0;
    XRAM[15918] = 8'b0;
    XRAM[15919] = 8'b0;
    XRAM[15920] = 8'b0;
    XRAM[15921] = 8'b0;
    XRAM[15922] = 8'b0;
    XRAM[15923] = 8'b0;
    XRAM[15924] = 8'b0;
    XRAM[15925] = 8'b0;
    XRAM[15926] = 8'b0;
    XRAM[15927] = 8'b0;
    XRAM[15928] = 8'b0;
    XRAM[15929] = 8'b0;
    XRAM[15930] = 8'b0;
    XRAM[15931] = 8'b0;
    XRAM[15932] = 8'b0;
    XRAM[15933] = 8'b0;
    XRAM[15934] = 8'b0;
    XRAM[15935] = 8'b0;
    XRAM[15936] = 8'b0;
    XRAM[15937] = 8'b0;
    XRAM[15938] = 8'b0;
    XRAM[15939] = 8'b0;
    XRAM[15940] = 8'b0;
    XRAM[15941] = 8'b0;
    XRAM[15942] = 8'b0;
    XRAM[15943] = 8'b0;
    XRAM[15944] = 8'b0;
    XRAM[15945] = 8'b0;
    XRAM[15946] = 8'b0;
    XRAM[15947] = 8'b0;
    XRAM[15948] = 8'b0;
    XRAM[15949] = 8'b0;
    XRAM[15950] = 8'b0;
    XRAM[15951] = 8'b0;
    XRAM[15952] = 8'b0;
    XRAM[15953] = 8'b0;
    XRAM[15954] = 8'b0;
    XRAM[15955] = 8'b0;
    XRAM[15956] = 8'b0;
    XRAM[15957] = 8'b0;
    XRAM[15958] = 8'b0;
    XRAM[15959] = 8'b0;
    XRAM[15960] = 8'b0;
    XRAM[15961] = 8'b0;
    XRAM[15962] = 8'b0;
    XRAM[15963] = 8'b0;
    XRAM[15964] = 8'b0;
    XRAM[15965] = 8'b0;
    XRAM[15966] = 8'b0;
    XRAM[15967] = 8'b0;
    XRAM[15968] = 8'b0;
    XRAM[15969] = 8'b0;
    XRAM[15970] = 8'b0;
    XRAM[15971] = 8'b0;
    XRAM[15972] = 8'b0;
    XRAM[15973] = 8'b0;
    XRAM[15974] = 8'b0;
    XRAM[15975] = 8'b0;
    XRAM[15976] = 8'b0;
    XRAM[15977] = 8'b0;
    XRAM[15978] = 8'b0;
    XRAM[15979] = 8'b0;
    XRAM[15980] = 8'b0;
    XRAM[15981] = 8'b0;
    XRAM[15982] = 8'b0;
    XRAM[15983] = 8'b0;
    XRAM[15984] = 8'b0;
    XRAM[15985] = 8'b0;
    XRAM[15986] = 8'b0;
    XRAM[15987] = 8'b0;
    XRAM[15988] = 8'b0;
    XRAM[15989] = 8'b0;
    XRAM[15990] = 8'b0;
    XRAM[15991] = 8'b0;
    XRAM[15992] = 8'b0;
    XRAM[15993] = 8'b0;
    XRAM[15994] = 8'b0;
    XRAM[15995] = 8'b0;
    XRAM[15996] = 8'b0;
    XRAM[15997] = 8'b0;
    XRAM[15998] = 8'b0;
    XRAM[15999] = 8'b0;
    XRAM[16000] = 8'b0;
    XRAM[16001] = 8'b0;
    XRAM[16002] = 8'b0;
    XRAM[16003] = 8'b0;
    XRAM[16004] = 8'b0;
    XRAM[16005] = 8'b0;
    XRAM[16006] = 8'b0;
    XRAM[16007] = 8'b0;
    XRAM[16008] = 8'b0;
    XRAM[16009] = 8'b0;
    XRAM[16010] = 8'b0;
    XRAM[16011] = 8'b0;
    XRAM[16012] = 8'b0;
    XRAM[16013] = 8'b0;
    XRAM[16014] = 8'b0;
    XRAM[16015] = 8'b0;
    XRAM[16016] = 8'b0;
    XRAM[16017] = 8'b0;
    XRAM[16018] = 8'b0;
    XRAM[16019] = 8'b0;
    XRAM[16020] = 8'b0;
    XRAM[16021] = 8'b0;
    XRAM[16022] = 8'b0;
    XRAM[16023] = 8'b0;
    XRAM[16024] = 8'b0;
    XRAM[16025] = 8'b0;
    XRAM[16026] = 8'b0;
    XRAM[16027] = 8'b0;
    XRAM[16028] = 8'b0;
    XRAM[16029] = 8'b0;
    XRAM[16030] = 8'b0;
    XRAM[16031] = 8'b0;
    XRAM[16032] = 8'b0;
    XRAM[16033] = 8'b0;
    XRAM[16034] = 8'b0;
    XRAM[16035] = 8'b0;
    XRAM[16036] = 8'b0;
    XRAM[16037] = 8'b0;
    XRAM[16038] = 8'b0;
    XRAM[16039] = 8'b0;
    XRAM[16040] = 8'b0;
    XRAM[16041] = 8'b0;
    XRAM[16042] = 8'b0;
    XRAM[16043] = 8'b0;
    XRAM[16044] = 8'b0;
    XRAM[16045] = 8'b0;
    XRAM[16046] = 8'b0;
    XRAM[16047] = 8'b0;
    XRAM[16048] = 8'b0;
    XRAM[16049] = 8'b0;
    XRAM[16050] = 8'b0;
    XRAM[16051] = 8'b0;
    XRAM[16052] = 8'b0;
    XRAM[16053] = 8'b0;
    XRAM[16054] = 8'b0;
    XRAM[16055] = 8'b0;
    XRAM[16056] = 8'b0;
    XRAM[16057] = 8'b0;
    XRAM[16058] = 8'b0;
    XRAM[16059] = 8'b0;
    XRAM[16060] = 8'b0;
    XRAM[16061] = 8'b0;
    XRAM[16062] = 8'b0;
    XRAM[16063] = 8'b0;
    XRAM[16064] = 8'b0;
    XRAM[16065] = 8'b0;
    XRAM[16066] = 8'b0;
    XRAM[16067] = 8'b0;
    XRAM[16068] = 8'b0;
    XRAM[16069] = 8'b0;
    XRAM[16070] = 8'b0;
    XRAM[16071] = 8'b0;
    XRAM[16072] = 8'b0;
    XRAM[16073] = 8'b0;
    XRAM[16074] = 8'b0;
    XRAM[16075] = 8'b0;
    XRAM[16076] = 8'b0;
    XRAM[16077] = 8'b0;
    XRAM[16078] = 8'b0;
    XRAM[16079] = 8'b0;
    XRAM[16080] = 8'b0;
    XRAM[16081] = 8'b0;
    XRAM[16082] = 8'b0;
    XRAM[16083] = 8'b0;
    XRAM[16084] = 8'b0;
    XRAM[16085] = 8'b0;
    XRAM[16086] = 8'b0;
    XRAM[16087] = 8'b0;
    XRAM[16088] = 8'b0;
    XRAM[16089] = 8'b0;
    XRAM[16090] = 8'b0;
    XRAM[16091] = 8'b0;
    XRAM[16092] = 8'b0;
    XRAM[16093] = 8'b0;
    XRAM[16094] = 8'b0;
    XRAM[16095] = 8'b0;
    XRAM[16096] = 8'b0;
    XRAM[16097] = 8'b0;
    XRAM[16098] = 8'b0;
    XRAM[16099] = 8'b0;
    XRAM[16100] = 8'b0;
    XRAM[16101] = 8'b0;
    XRAM[16102] = 8'b0;
    XRAM[16103] = 8'b0;
    XRAM[16104] = 8'b0;
    XRAM[16105] = 8'b0;
    XRAM[16106] = 8'b0;
    XRAM[16107] = 8'b0;
    XRAM[16108] = 8'b0;
    XRAM[16109] = 8'b0;
    XRAM[16110] = 8'b0;
    XRAM[16111] = 8'b0;
    XRAM[16112] = 8'b0;
    XRAM[16113] = 8'b0;
    XRAM[16114] = 8'b0;
    XRAM[16115] = 8'b0;
    XRAM[16116] = 8'b0;
    XRAM[16117] = 8'b0;
    XRAM[16118] = 8'b0;
    XRAM[16119] = 8'b0;
    XRAM[16120] = 8'b0;
    XRAM[16121] = 8'b0;
    XRAM[16122] = 8'b0;
    XRAM[16123] = 8'b0;
    XRAM[16124] = 8'b0;
    XRAM[16125] = 8'b0;
    XRAM[16126] = 8'b0;
    XRAM[16127] = 8'b0;
    XRAM[16128] = 8'b0;
    XRAM[16129] = 8'b0;
    XRAM[16130] = 8'b0;
    XRAM[16131] = 8'b0;
    XRAM[16132] = 8'b0;
    XRAM[16133] = 8'b0;
    XRAM[16134] = 8'b0;
    XRAM[16135] = 8'b0;
    XRAM[16136] = 8'b0;
    XRAM[16137] = 8'b0;
    XRAM[16138] = 8'b0;
    XRAM[16139] = 8'b0;
    XRAM[16140] = 8'b0;
    XRAM[16141] = 8'b0;
    XRAM[16142] = 8'b0;
    XRAM[16143] = 8'b0;
    XRAM[16144] = 8'b0;
    XRAM[16145] = 8'b0;
    XRAM[16146] = 8'b0;
    XRAM[16147] = 8'b0;
    XRAM[16148] = 8'b0;
    XRAM[16149] = 8'b0;
    XRAM[16150] = 8'b0;
    XRAM[16151] = 8'b0;
    XRAM[16152] = 8'b0;
    XRAM[16153] = 8'b0;
    XRAM[16154] = 8'b0;
    XRAM[16155] = 8'b0;
    XRAM[16156] = 8'b0;
    XRAM[16157] = 8'b0;
    XRAM[16158] = 8'b0;
    XRAM[16159] = 8'b0;
    XRAM[16160] = 8'b0;
    XRAM[16161] = 8'b0;
    XRAM[16162] = 8'b0;
    XRAM[16163] = 8'b0;
    XRAM[16164] = 8'b0;
    XRAM[16165] = 8'b0;
    XRAM[16166] = 8'b0;
    XRAM[16167] = 8'b0;
    XRAM[16168] = 8'b0;
    XRAM[16169] = 8'b0;
    XRAM[16170] = 8'b0;
    XRAM[16171] = 8'b0;
    XRAM[16172] = 8'b0;
    XRAM[16173] = 8'b0;
    XRAM[16174] = 8'b0;
    XRAM[16175] = 8'b0;
    XRAM[16176] = 8'b0;
    XRAM[16177] = 8'b0;
    XRAM[16178] = 8'b0;
    XRAM[16179] = 8'b0;
    XRAM[16180] = 8'b0;
    XRAM[16181] = 8'b0;
    XRAM[16182] = 8'b0;
    XRAM[16183] = 8'b0;
    XRAM[16184] = 8'b0;
    XRAM[16185] = 8'b0;
    XRAM[16186] = 8'b0;
    XRAM[16187] = 8'b0;
    XRAM[16188] = 8'b0;
    XRAM[16189] = 8'b0;
    XRAM[16190] = 8'b0;
    XRAM[16191] = 8'b0;
    XRAM[16192] = 8'b0;
    XRAM[16193] = 8'b0;
    XRAM[16194] = 8'b0;
    XRAM[16195] = 8'b0;
    XRAM[16196] = 8'b0;
    XRAM[16197] = 8'b0;
    XRAM[16198] = 8'b0;
    XRAM[16199] = 8'b0;
    XRAM[16200] = 8'b0;
    XRAM[16201] = 8'b0;
    XRAM[16202] = 8'b0;
    XRAM[16203] = 8'b0;
    XRAM[16204] = 8'b0;
    XRAM[16205] = 8'b0;
    XRAM[16206] = 8'b0;
    XRAM[16207] = 8'b0;
    XRAM[16208] = 8'b0;
    XRAM[16209] = 8'b0;
    XRAM[16210] = 8'b0;
    XRAM[16211] = 8'b0;
    XRAM[16212] = 8'b0;
    XRAM[16213] = 8'b0;
    XRAM[16214] = 8'b0;
    XRAM[16215] = 8'b0;
    XRAM[16216] = 8'b0;
    XRAM[16217] = 8'b0;
    XRAM[16218] = 8'b0;
    XRAM[16219] = 8'b0;
    XRAM[16220] = 8'b0;
    XRAM[16221] = 8'b0;
    XRAM[16222] = 8'b0;
    XRAM[16223] = 8'b0;
    XRAM[16224] = 8'b0;
    XRAM[16225] = 8'b0;
    XRAM[16226] = 8'b0;
    XRAM[16227] = 8'b0;
    XRAM[16228] = 8'b0;
    XRAM[16229] = 8'b0;
    XRAM[16230] = 8'b0;
    XRAM[16231] = 8'b0;
    XRAM[16232] = 8'b0;
    XRAM[16233] = 8'b0;
    XRAM[16234] = 8'b0;
    XRAM[16235] = 8'b0;
    XRAM[16236] = 8'b0;
    XRAM[16237] = 8'b0;
    XRAM[16238] = 8'b0;
    XRAM[16239] = 8'b0;
    XRAM[16240] = 8'b0;
    XRAM[16241] = 8'b0;
    XRAM[16242] = 8'b0;
    XRAM[16243] = 8'b0;
    XRAM[16244] = 8'b0;
    XRAM[16245] = 8'b0;
    XRAM[16246] = 8'b0;
    XRAM[16247] = 8'b0;
    XRAM[16248] = 8'b0;
    XRAM[16249] = 8'b0;
    XRAM[16250] = 8'b0;
    XRAM[16251] = 8'b0;
    XRAM[16252] = 8'b0;
    XRAM[16253] = 8'b0;
    XRAM[16254] = 8'b0;
    XRAM[16255] = 8'b0;
    XRAM[16256] = 8'b0;
    XRAM[16257] = 8'b0;
    XRAM[16258] = 8'b0;
    XRAM[16259] = 8'b0;
    XRAM[16260] = 8'b0;
    XRAM[16261] = 8'b0;
    XRAM[16262] = 8'b0;
    XRAM[16263] = 8'b0;
    XRAM[16264] = 8'b0;
    XRAM[16265] = 8'b0;
    XRAM[16266] = 8'b0;
    XRAM[16267] = 8'b0;
    XRAM[16268] = 8'b0;
    XRAM[16269] = 8'b0;
    XRAM[16270] = 8'b0;
    XRAM[16271] = 8'b0;
    XRAM[16272] = 8'b0;
    XRAM[16273] = 8'b0;
    XRAM[16274] = 8'b0;
    XRAM[16275] = 8'b0;
    XRAM[16276] = 8'b0;
    XRAM[16277] = 8'b0;
    XRAM[16278] = 8'b0;
    XRAM[16279] = 8'b0;
    XRAM[16280] = 8'b0;
    XRAM[16281] = 8'b0;
    XRAM[16282] = 8'b0;
    XRAM[16283] = 8'b0;
    XRAM[16284] = 8'b0;
    XRAM[16285] = 8'b0;
    XRAM[16286] = 8'b0;
    XRAM[16287] = 8'b0;
    XRAM[16288] = 8'b0;
    XRAM[16289] = 8'b0;
    XRAM[16290] = 8'b0;
    XRAM[16291] = 8'b0;
    XRAM[16292] = 8'b0;
    XRAM[16293] = 8'b0;
    XRAM[16294] = 8'b0;
    XRAM[16295] = 8'b0;
    XRAM[16296] = 8'b0;
    XRAM[16297] = 8'b0;
    XRAM[16298] = 8'b0;
    XRAM[16299] = 8'b0;
    XRAM[16300] = 8'b0;
    XRAM[16301] = 8'b0;
    XRAM[16302] = 8'b0;
    XRAM[16303] = 8'b0;
    XRAM[16304] = 8'b0;
    XRAM[16305] = 8'b0;
    XRAM[16306] = 8'b0;
    XRAM[16307] = 8'b0;
    XRAM[16308] = 8'b0;
    XRAM[16309] = 8'b0;
    XRAM[16310] = 8'b0;
    XRAM[16311] = 8'b0;
    XRAM[16312] = 8'b0;
    XRAM[16313] = 8'b0;
    XRAM[16314] = 8'b0;
    XRAM[16315] = 8'b0;
    XRAM[16316] = 8'b0;
    XRAM[16317] = 8'b0;
    XRAM[16318] = 8'b0;
    XRAM[16319] = 8'b0;
    XRAM[16320] = 8'b0;
    XRAM[16321] = 8'b0;
    XRAM[16322] = 8'b0;
    XRAM[16323] = 8'b0;
    XRAM[16324] = 8'b0;
    XRAM[16325] = 8'b0;
    XRAM[16326] = 8'b0;
    XRAM[16327] = 8'b0;
    XRAM[16328] = 8'b0;
    XRAM[16329] = 8'b0;
    XRAM[16330] = 8'b0;
    XRAM[16331] = 8'b0;
    XRAM[16332] = 8'b0;
    XRAM[16333] = 8'b0;
    XRAM[16334] = 8'b0;
    XRAM[16335] = 8'b0;
    XRAM[16336] = 8'b0;
    XRAM[16337] = 8'b0;
    XRAM[16338] = 8'b0;
    XRAM[16339] = 8'b0;
    XRAM[16340] = 8'b0;
    XRAM[16341] = 8'b0;
    XRAM[16342] = 8'b0;
    XRAM[16343] = 8'b0;
    XRAM[16344] = 8'b0;
    XRAM[16345] = 8'b0;
    XRAM[16346] = 8'b0;
    XRAM[16347] = 8'b0;
    XRAM[16348] = 8'b0;
    XRAM[16349] = 8'b0;
    XRAM[16350] = 8'b0;
    XRAM[16351] = 8'b0;
    XRAM[16352] = 8'b0;
    XRAM[16353] = 8'b0;
    XRAM[16354] = 8'b0;
    XRAM[16355] = 8'b0;
    XRAM[16356] = 8'b0;
    XRAM[16357] = 8'b0;
    XRAM[16358] = 8'b0;
    XRAM[16359] = 8'b0;
    XRAM[16360] = 8'b0;
    XRAM[16361] = 8'b0;
    XRAM[16362] = 8'b0;
    XRAM[16363] = 8'b0;
    XRAM[16364] = 8'b0;
    XRAM[16365] = 8'b0;
    XRAM[16366] = 8'b0;
    XRAM[16367] = 8'b0;
    XRAM[16368] = 8'b0;
    XRAM[16369] = 8'b0;
    XRAM[16370] = 8'b0;
    XRAM[16371] = 8'b0;
    XRAM[16372] = 8'b0;
    XRAM[16373] = 8'b0;
    XRAM[16374] = 8'b0;
    XRAM[16375] = 8'b0;
    XRAM[16376] = 8'b0;
    XRAM[16377] = 8'b0;
    XRAM[16378] = 8'b0;
    XRAM[16379] = 8'b0;
    XRAM[16380] = 8'b0;
    XRAM[16381] = 8'b0;
    XRAM[16382] = 8'b0;
    XRAM[16383] = 8'b0;
    XRAM[16384] = 8'b0;
    XRAM[16385] = 8'b0;
    XRAM[16386] = 8'b0;
    XRAM[16387] = 8'b0;
    XRAM[16388] = 8'b0;
    XRAM[16389] = 8'b0;
    XRAM[16390] = 8'b0;
    XRAM[16391] = 8'b0;
    XRAM[16392] = 8'b0;
    XRAM[16393] = 8'b0;
    XRAM[16394] = 8'b0;
    XRAM[16395] = 8'b0;
    XRAM[16396] = 8'b0;
    XRAM[16397] = 8'b0;
    XRAM[16398] = 8'b0;
    XRAM[16399] = 8'b0;
    XRAM[16400] = 8'b0;
    XRAM[16401] = 8'b0;
    XRAM[16402] = 8'b0;
    XRAM[16403] = 8'b0;
    XRAM[16404] = 8'b0;
    XRAM[16405] = 8'b0;
    XRAM[16406] = 8'b0;
    XRAM[16407] = 8'b0;
    XRAM[16408] = 8'b0;
    XRAM[16409] = 8'b0;
    XRAM[16410] = 8'b0;
    XRAM[16411] = 8'b0;
    XRAM[16412] = 8'b0;
    XRAM[16413] = 8'b0;
    XRAM[16414] = 8'b0;
    XRAM[16415] = 8'b0;
    XRAM[16416] = 8'b0;
    XRAM[16417] = 8'b0;
    XRAM[16418] = 8'b0;
    XRAM[16419] = 8'b0;
    XRAM[16420] = 8'b0;
    XRAM[16421] = 8'b0;
    XRAM[16422] = 8'b0;
    XRAM[16423] = 8'b0;
    XRAM[16424] = 8'b0;
    XRAM[16425] = 8'b0;
    XRAM[16426] = 8'b0;
    XRAM[16427] = 8'b0;
    XRAM[16428] = 8'b0;
    XRAM[16429] = 8'b0;
    XRAM[16430] = 8'b0;
    XRAM[16431] = 8'b0;
    XRAM[16432] = 8'b0;
    XRAM[16433] = 8'b0;
    XRAM[16434] = 8'b0;
    XRAM[16435] = 8'b0;
    XRAM[16436] = 8'b0;
    XRAM[16437] = 8'b0;
    XRAM[16438] = 8'b0;
    XRAM[16439] = 8'b0;
    XRAM[16440] = 8'b0;
    XRAM[16441] = 8'b0;
    XRAM[16442] = 8'b0;
    XRAM[16443] = 8'b0;
    XRAM[16444] = 8'b0;
    XRAM[16445] = 8'b0;
    XRAM[16446] = 8'b0;
    XRAM[16447] = 8'b0;
    XRAM[16448] = 8'b0;
    XRAM[16449] = 8'b0;
    XRAM[16450] = 8'b0;
    XRAM[16451] = 8'b0;
    XRAM[16452] = 8'b0;
    XRAM[16453] = 8'b0;
    XRAM[16454] = 8'b0;
    XRAM[16455] = 8'b0;
    XRAM[16456] = 8'b0;
    XRAM[16457] = 8'b0;
    XRAM[16458] = 8'b0;
    XRAM[16459] = 8'b0;
    XRAM[16460] = 8'b0;
    XRAM[16461] = 8'b0;
    XRAM[16462] = 8'b0;
    XRAM[16463] = 8'b0;
    XRAM[16464] = 8'b0;
    XRAM[16465] = 8'b0;
    XRAM[16466] = 8'b0;
    XRAM[16467] = 8'b0;
    XRAM[16468] = 8'b0;
    XRAM[16469] = 8'b0;
    XRAM[16470] = 8'b0;
    XRAM[16471] = 8'b0;
    XRAM[16472] = 8'b0;
    XRAM[16473] = 8'b0;
    XRAM[16474] = 8'b0;
    XRAM[16475] = 8'b0;
    XRAM[16476] = 8'b0;
    XRAM[16477] = 8'b0;
    XRAM[16478] = 8'b0;
    XRAM[16479] = 8'b0;
    XRAM[16480] = 8'b0;
    XRAM[16481] = 8'b0;
    XRAM[16482] = 8'b0;
    XRAM[16483] = 8'b0;
    XRAM[16484] = 8'b0;
    XRAM[16485] = 8'b0;
    XRAM[16486] = 8'b0;
    XRAM[16487] = 8'b0;
    XRAM[16488] = 8'b0;
    XRAM[16489] = 8'b0;
    XRAM[16490] = 8'b0;
    XRAM[16491] = 8'b0;
    XRAM[16492] = 8'b0;
    XRAM[16493] = 8'b0;
    XRAM[16494] = 8'b0;
    XRAM[16495] = 8'b0;
    XRAM[16496] = 8'b0;
    XRAM[16497] = 8'b0;
    XRAM[16498] = 8'b0;
    XRAM[16499] = 8'b0;
    XRAM[16500] = 8'b0;
    XRAM[16501] = 8'b0;
    XRAM[16502] = 8'b0;
    XRAM[16503] = 8'b0;
    XRAM[16504] = 8'b0;
    XRAM[16505] = 8'b0;
    XRAM[16506] = 8'b0;
    XRAM[16507] = 8'b0;
    XRAM[16508] = 8'b0;
    XRAM[16509] = 8'b0;
    XRAM[16510] = 8'b0;
    XRAM[16511] = 8'b0;
    XRAM[16512] = 8'b0;
    XRAM[16513] = 8'b0;
    XRAM[16514] = 8'b0;
    XRAM[16515] = 8'b0;
    XRAM[16516] = 8'b0;
    XRAM[16517] = 8'b0;
    XRAM[16518] = 8'b0;
    XRAM[16519] = 8'b0;
    XRAM[16520] = 8'b0;
    XRAM[16521] = 8'b0;
    XRAM[16522] = 8'b0;
    XRAM[16523] = 8'b0;
    XRAM[16524] = 8'b0;
    XRAM[16525] = 8'b0;
    XRAM[16526] = 8'b0;
    XRAM[16527] = 8'b0;
    XRAM[16528] = 8'b0;
    XRAM[16529] = 8'b0;
    XRAM[16530] = 8'b0;
    XRAM[16531] = 8'b0;
    XRAM[16532] = 8'b0;
    XRAM[16533] = 8'b0;
    XRAM[16534] = 8'b0;
    XRAM[16535] = 8'b0;
    XRAM[16536] = 8'b0;
    XRAM[16537] = 8'b0;
    XRAM[16538] = 8'b0;
    XRAM[16539] = 8'b0;
    XRAM[16540] = 8'b0;
    XRAM[16541] = 8'b0;
    XRAM[16542] = 8'b0;
    XRAM[16543] = 8'b0;
    XRAM[16544] = 8'b0;
    XRAM[16545] = 8'b0;
    XRAM[16546] = 8'b0;
    XRAM[16547] = 8'b0;
    XRAM[16548] = 8'b0;
    XRAM[16549] = 8'b0;
    XRAM[16550] = 8'b0;
    XRAM[16551] = 8'b0;
    XRAM[16552] = 8'b0;
    XRAM[16553] = 8'b0;
    XRAM[16554] = 8'b0;
    XRAM[16555] = 8'b0;
    XRAM[16556] = 8'b0;
    XRAM[16557] = 8'b0;
    XRAM[16558] = 8'b0;
    XRAM[16559] = 8'b0;
    XRAM[16560] = 8'b0;
    XRAM[16561] = 8'b0;
    XRAM[16562] = 8'b0;
    XRAM[16563] = 8'b0;
    XRAM[16564] = 8'b0;
    XRAM[16565] = 8'b0;
    XRAM[16566] = 8'b0;
    XRAM[16567] = 8'b0;
    XRAM[16568] = 8'b0;
    XRAM[16569] = 8'b0;
    XRAM[16570] = 8'b0;
    XRAM[16571] = 8'b0;
    XRAM[16572] = 8'b0;
    XRAM[16573] = 8'b0;
    XRAM[16574] = 8'b0;
    XRAM[16575] = 8'b0;
    XRAM[16576] = 8'b0;
    XRAM[16577] = 8'b0;
    XRAM[16578] = 8'b0;
    XRAM[16579] = 8'b0;
    XRAM[16580] = 8'b0;
    XRAM[16581] = 8'b0;
    XRAM[16582] = 8'b0;
    XRAM[16583] = 8'b0;
    XRAM[16584] = 8'b0;
    XRAM[16585] = 8'b0;
    XRAM[16586] = 8'b0;
    XRAM[16587] = 8'b0;
    XRAM[16588] = 8'b0;
    XRAM[16589] = 8'b0;
    XRAM[16590] = 8'b0;
    XRAM[16591] = 8'b0;
    XRAM[16592] = 8'b0;
    XRAM[16593] = 8'b0;
    XRAM[16594] = 8'b0;
    XRAM[16595] = 8'b0;
    XRAM[16596] = 8'b0;
    XRAM[16597] = 8'b0;
    XRAM[16598] = 8'b0;
    XRAM[16599] = 8'b0;
    XRAM[16600] = 8'b0;
    XRAM[16601] = 8'b0;
    XRAM[16602] = 8'b0;
    XRAM[16603] = 8'b0;
    XRAM[16604] = 8'b0;
    XRAM[16605] = 8'b0;
    XRAM[16606] = 8'b0;
    XRAM[16607] = 8'b0;
    XRAM[16608] = 8'b0;
    XRAM[16609] = 8'b0;
    XRAM[16610] = 8'b0;
    XRAM[16611] = 8'b0;
    XRAM[16612] = 8'b0;
    XRAM[16613] = 8'b0;
    XRAM[16614] = 8'b0;
    XRAM[16615] = 8'b0;
    XRAM[16616] = 8'b0;
    XRAM[16617] = 8'b0;
    XRAM[16618] = 8'b0;
    XRAM[16619] = 8'b0;
    XRAM[16620] = 8'b0;
    XRAM[16621] = 8'b0;
    XRAM[16622] = 8'b0;
    XRAM[16623] = 8'b0;
    XRAM[16624] = 8'b0;
    XRAM[16625] = 8'b0;
    XRAM[16626] = 8'b0;
    XRAM[16627] = 8'b0;
    XRAM[16628] = 8'b0;
    XRAM[16629] = 8'b0;
    XRAM[16630] = 8'b0;
    XRAM[16631] = 8'b0;
    XRAM[16632] = 8'b0;
    XRAM[16633] = 8'b0;
    XRAM[16634] = 8'b0;
    XRAM[16635] = 8'b0;
    XRAM[16636] = 8'b0;
    XRAM[16637] = 8'b0;
    XRAM[16638] = 8'b0;
    XRAM[16639] = 8'b0;
    XRAM[16640] = 8'b0;
    XRAM[16641] = 8'b0;
    XRAM[16642] = 8'b0;
    XRAM[16643] = 8'b0;
    XRAM[16644] = 8'b0;
    XRAM[16645] = 8'b0;
    XRAM[16646] = 8'b0;
    XRAM[16647] = 8'b0;
    XRAM[16648] = 8'b0;
    XRAM[16649] = 8'b0;
    XRAM[16650] = 8'b0;
    XRAM[16651] = 8'b0;
    XRAM[16652] = 8'b0;
    XRAM[16653] = 8'b0;
    XRAM[16654] = 8'b0;
    XRAM[16655] = 8'b0;
    XRAM[16656] = 8'b0;
    XRAM[16657] = 8'b0;
    XRAM[16658] = 8'b0;
    XRAM[16659] = 8'b0;
    XRAM[16660] = 8'b0;
    XRAM[16661] = 8'b0;
    XRAM[16662] = 8'b0;
    XRAM[16663] = 8'b0;
    XRAM[16664] = 8'b0;
    XRAM[16665] = 8'b0;
    XRAM[16666] = 8'b0;
    XRAM[16667] = 8'b0;
    XRAM[16668] = 8'b0;
    XRAM[16669] = 8'b0;
    XRAM[16670] = 8'b0;
    XRAM[16671] = 8'b0;
    XRAM[16672] = 8'b0;
    XRAM[16673] = 8'b0;
    XRAM[16674] = 8'b0;
    XRAM[16675] = 8'b0;
    XRAM[16676] = 8'b0;
    XRAM[16677] = 8'b0;
    XRAM[16678] = 8'b0;
    XRAM[16679] = 8'b0;
    XRAM[16680] = 8'b0;
    XRAM[16681] = 8'b0;
    XRAM[16682] = 8'b0;
    XRAM[16683] = 8'b0;
    XRAM[16684] = 8'b0;
    XRAM[16685] = 8'b0;
    XRAM[16686] = 8'b0;
    XRAM[16687] = 8'b0;
    XRAM[16688] = 8'b0;
    XRAM[16689] = 8'b0;
    XRAM[16690] = 8'b0;
    XRAM[16691] = 8'b0;
    XRAM[16692] = 8'b0;
    XRAM[16693] = 8'b0;
    XRAM[16694] = 8'b0;
    XRAM[16695] = 8'b0;
    XRAM[16696] = 8'b0;
    XRAM[16697] = 8'b0;
    XRAM[16698] = 8'b0;
    XRAM[16699] = 8'b0;
    XRAM[16700] = 8'b0;
    XRAM[16701] = 8'b0;
    XRAM[16702] = 8'b0;
    XRAM[16703] = 8'b0;
    XRAM[16704] = 8'b0;
    XRAM[16705] = 8'b0;
    XRAM[16706] = 8'b0;
    XRAM[16707] = 8'b0;
    XRAM[16708] = 8'b0;
    XRAM[16709] = 8'b0;
    XRAM[16710] = 8'b0;
    XRAM[16711] = 8'b0;
    XRAM[16712] = 8'b0;
    XRAM[16713] = 8'b0;
    XRAM[16714] = 8'b0;
    XRAM[16715] = 8'b0;
    XRAM[16716] = 8'b0;
    XRAM[16717] = 8'b0;
    XRAM[16718] = 8'b0;
    XRAM[16719] = 8'b0;
    XRAM[16720] = 8'b0;
    XRAM[16721] = 8'b0;
    XRAM[16722] = 8'b0;
    XRAM[16723] = 8'b0;
    XRAM[16724] = 8'b0;
    XRAM[16725] = 8'b0;
    XRAM[16726] = 8'b0;
    XRAM[16727] = 8'b0;
    XRAM[16728] = 8'b0;
    XRAM[16729] = 8'b0;
    XRAM[16730] = 8'b0;
    XRAM[16731] = 8'b0;
    XRAM[16732] = 8'b0;
    XRAM[16733] = 8'b0;
    XRAM[16734] = 8'b0;
    XRAM[16735] = 8'b0;
    XRAM[16736] = 8'b0;
    XRAM[16737] = 8'b0;
    XRAM[16738] = 8'b0;
    XRAM[16739] = 8'b0;
    XRAM[16740] = 8'b0;
    XRAM[16741] = 8'b0;
    XRAM[16742] = 8'b0;
    XRAM[16743] = 8'b0;
    XRAM[16744] = 8'b0;
    XRAM[16745] = 8'b0;
    XRAM[16746] = 8'b0;
    XRAM[16747] = 8'b0;
    XRAM[16748] = 8'b0;
    XRAM[16749] = 8'b0;
    XRAM[16750] = 8'b0;
    XRAM[16751] = 8'b0;
    XRAM[16752] = 8'b0;
    XRAM[16753] = 8'b0;
    XRAM[16754] = 8'b0;
    XRAM[16755] = 8'b0;
    XRAM[16756] = 8'b0;
    XRAM[16757] = 8'b0;
    XRAM[16758] = 8'b0;
    XRAM[16759] = 8'b0;
    XRAM[16760] = 8'b0;
    XRAM[16761] = 8'b0;
    XRAM[16762] = 8'b0;
    XRAM[16763] = 8'b0;
    XRAM[16764] = 8'b0;
    XRAM[16765] = 8'b0;
    XRAM[16766] = 8'b0;
    XRAM[16767] = 8'b0;
    XRAM[16768] = 8'b0;
    XRAM[16769] = 8'b0;
    XRAM[16770] = 8'b0;
    XRAM[16771] = 8'b0;
    XRAM[16772] = 8'b0;
    XRAM[16773] = 8'b0;
    XRAM[16774] = 8'b0;
    XRAM[16775] = 8'b0;
    XRAM[16776] = 8'b0;
    XRAM[16777] = 8'b0;
    XRAM[16778] = 8'b0;
    XRAM[16779] = 8'b0;
    XRAM[16780] = 8'b0;
    XRAM[16781] = 8'b0;
    XRAM[16782] = 8'b0;
    XRAM[16783] = 8'b0;
    XRAM[16784] = 8'b0;
    XRAM[16785] = 8'b0;
    XRAM[16786] = 8'b0;
    XRAM[16787] = 8'b0;
    XRAM[16788] = 8'b0;
    XRAM[16789] = 8'b0;
    XRAM[16790] = 8'b0;
    XRAM[16791] = 8'b0;
    XRAM[16792] = 8'b0;
    XRAM[16793] = 8'b0;
    XRAM[16794] = 8'b0;
    XRAM[16795] = 8'b0;
    XRAM[16796] = 8'b0;
    XRAM[16797] = 8'b0;
    XRAM[16798] = 8'b0;
    XRAM[16799] = 8'b0;
    XRAM[16800] = 8'b0;
    XRAM[16801] = 8'b0;
    XRAM[16802] = 8'b0;
    XRAM[16803] = 8'b0;
    XRAM[16804] = 8'b0;
    XRAM[16805] = 8'b0;
    XRAM[16806] = 8'b0;
    XRAM[16807] = 8'b0;
    XRAM[16808] = 8'b0;
    XRAM[16809] = 8'b0;
    XRAM[16810] = 8'b0;
    XRAM[16811] = 8'b0;
    XRAM[16812] = 8'b0;
    XRAM[16813] = 8'b0;
    XRAM[16814] = 8'b0;
    XRAM[16815] = 8'b0;
    XRAM[16816] = 8'b0;
    XRAM[16817] = 8'b0;
    XRAM[16818] = 8'b0;
    XRAM[16819] = 8'b0;
    XRAM[16820] = 8'b0;
    XRAM[16821] = 8'b0;
    XRAM[16822] = 8'b0;
    XRAM[16823] = 8'b0;
    XRAM[16824] = 8'b0;
    XRAM[16825] = 8'b0;
    XRAM[16826] = 8'b0;
    XRAM[16827] = 8'b0;
    XRAM[16828] = 8'b0;
    XRAM[16829] = 8'b0;
    XRAM[16830] = 8'b0;
    XRAM[16831] = 8'b0;
    XRAM[16832] = 8'b0;
    XRAM[16833] = 8'b0;
    XRAM[16834] = 8'b0;
    XRAM[16835] = 8'b0;
    XRAM[16836] = 8'b0;
    XRAM[16837] = 8'b0;
    XRAM[16838] = 8'b0;
    XRAM[16839] = 8'b0;
    XRAM[16840] = 8'b0;
    XRAM[16841] = 8'b0;
    XRAM[16842] = 8'b0;
    XRAM[16843] = 8'b0;
    XRAM[16844] = 8'b0;
    XRAM[16845] = 8'b0;
    XRAM[16846] = 8'b0;
    XRAM[16847] = 8'b0;
    XRAM[16848] = 8'b0;
    XRAM[16849] = 8'b0;
    XRAM[16850] = 8'b0;
    XRAM[16851] = 8'b0;
    XRAM[16852] = 8'b0;
    XRAM[16853] = 8'b0;
    XRAM[16854] = 8'b0;
    XRAM[16855] = 8'b0;
    XRAM[16856] = 8'b0;
    XRAM[16857] = 8'b0;
    XRAM[16858] = 8'b0;
    XRAM[16859] = 8'b0;
    XRAM[16860] = 8'b0;
    XRAM[16861] = 8'b0;
    XRAM[16862] = 8'b0;
    XRAM[16863] = 8'b0;
    XRAM[16864] = 8'b0;
    XRAM[16865] = 8'b0;
    XRAM[16866] = 8'b0;
    XRAM[16867] = 8'b0;
    XRAM[16868] = 8'b0;
    XRAM[16869] = 8'b0;
    XRAM[16870] = 8'b0;
    XRAM[16871] = 8'b0;
    XRAM[16872] = 8'b0;
    XRAM[16873] = 8'b0;
    XRAM[16874] = 8'b0;
    XRAM[16875] = 8'b0;
    XRAM[16876] = 8'b0;
    XRAM[16877] = 8'b0;
    XRAM[16878] = 8'b0;
    XRAM[16879] = 8'b0;
    XRAM[16880] = 8'b0;
    XRAM[16881] = 8'b0;
    XRAM[16882] = 8'b0;
    XRAM[16883] = 8'b0;
    XRAM[16884] = 8'b0;
    XRAM[16885] = 8'b0;
    XRAM[16886] = 8'b0;
    XRAM[16887] = 8'b0;
    XRAM[16888] = 8'b0;
    XRAM[16889] = 8'b0;
    XRAM[16890] = 8'b0;
    XRAM[16891] = 8'b0;
    XRAM[16892] = 8'b0;
    XRAM[16893] = 8'b0;
    XRAM[16894] = 8'b0;
    XRAM[16895] = 8'b0;
    XRAM[16896] = 8'b0;
    XRAM[16897] = 8'b0;
    XRAM[16898] = 8'b0;
    XRAM[16899] = 8'b0;
    XRAM[16900] = 8'b0;
    XRAM[16901] = 8'b0;
    XRAM[16902] = 8'b0;
    XRAM[16903] = 8'b0;
    XRAM[16904] = 8'b0;
    XRAM[16905] = 8'b0;
    XRAM[16906] = 8'b0;
    XRAM[16907] = 8'b0;
    XRAM[16908] = 8'b0;
    XRAM[16909] = 8'b0;
    XRAM[16910] = 8'b0;
    XRAM[16911] = 8'b0;
    XRAM[16912] = 8'b0;
    XRAM[16913] = 8'b0;
    XRAM[16914] = 8'b0;
    XRAM[16915] = 8'b0;
    XRAM[16916] = 8'b0;
    XRAM[16917] = 8'b0;
    XRAM[16918] = 8'b0;
    XRAM[16919] = 8'b0;
    XRAM[16920] = 8'b0;
    XRAM[16921] = 8'b0;
    XRAM[16922] = 8'b0;
    XRAM[16923] = 8'b0;
    XRAM[16924] = 8'b0;
    XRAM[16925] = 8'b0;
    XRAM[16926] = 8'b0;
    XRAM[16927] = 8'b0;
    XRAM[16928] = 8'b0;
    XRAM[16929] = 8'b0;
    XRAM[16930] = 8'b0;
    XRAM[16931] = 8'b0;
    XRAM[16932] = 8'b0;
    XRAM[16933] = 8'b0;
    XRAM[16934] = 8'b0;
    XRAM[16935] = 8'b0;
    XRAM[16936] = 8'b0;
    XRAM[16937] = 8'b0;
    XRAM[16938] = 8'b0;
    XRAM[16939] = 8'b0;
    XRAM[16940] = 8'b0;
    XRAM[16941] = 8'b0;
    XRAM[16942] = 8'b0;
    XRAM[16943] = 8'b0;
    XRAM[16944] = 8'b0;
    XRAM[16945] = 8'b0;
    XRAM[16946] = 8'b0;
    XRAM[16947] = 8'b0;
    XRAM[16948] = 8'b0;
    XRAM[16949] = 8'b0;
    XRAM[16950] = 8'b0;
    XRAM[16951] = 8'b0;
    XRAM[16952] = 8'b0;
    XRAM[16953] = 8'b0;
    XRAM[16954] = 8'b0;
    XRAM[16955] = 8'b0;
    XRAM[16956] = 8'b0;
    XRAM[16957] = 8'b0;
    XRAM[16958] = 8'b0;
    XRAM[16959] = 8'b0;
    XRAM[16960] = 8'b0;
    XRAM[16961] = 8'b0;
    XRAM[16962] = 8'b0;
    XRAM[16963] = 8'b0;
    XRAM[16964] = 8'b0;
    XRAM[16965] = 8'b0;
    XRAM[16966] = 8'b0;
    XRAM[16967] = 8'b0;
    XRAM[16968] = 8'b0;
    XRAM[16969] = 8'b0;
    XRAM[16970] = 8'b0;
    XRAM[16971] = 8'b0;
    XRAM[16972] = 8'b0;
    XRAM[16973] = 8'b0;
    XRAM[16974] = 8'b0;
    XRAM[16975] = 8'b0;
    XRAM[16976] = 8'b0;
    XRAM[16977] = 8'b0;
    XRAM[16978] = 8'b0;
    XRAM[16979] = 8'b0;
    XRAM[16980] = 8'b0;
    XRAM[16981] = 8'b0;
    XRAM[16982] = 8'b0;
    XRAM[16983] = 8'b0;
    XRAM[16984] = 8'b0;
    XRAM[16985] = 8'b0;
    XRAM[16986] = 8'b0;
    XRAM[16987] = 8'b0;
    XRAM[16988] = 8'b0;
    XRAM[16989] = 8'b0;
    XRAM[16990] = 8'b0;
    XRAM[16991] = 8'b0;
    XRAM[16992] = 8'b0;
    XRAM[16993] = 8'b0;
    XRAM[16994] = 8'b0;
    XRAM[16995] = 8'b0;
    XRAM[16996] = 8'b0;
    XRAM[16997] = 8'b0;
    XRAM[16998] = 8'b0;
    XRAM[16999] = 8'b0;
    XRAM[17000] = 8'b0;
    XRAM[17001] = 8'b0;
    XRAM[17002] = 8'b0;
    XRAM[17003] = 8'b0;
    XRAM[17004] = 8'b0;
    XRAM[17005] = 8'b0;
    XRAM[17006] = 8'b0;
    XRAM[17007] = 8'b0;
    XRAM[17008] = 8'b0;
    XRAM[17009] = 8'b0;
    XRAM[17010] = 8'b0;
    XRAM[17011] = 8'b0;
    XRAM[17012] = 8'b0;
    XRAM[17013] = 8'b0;
    XRAM[17014] = 8'b0;
    XRAM[17015] = 8'b0;
    XRAM[17016] = 8'b0;
    XRAM[17017] = 8'b0;
    XRAM[17018] = 8'b0;
    XRAM[17019] = 8'b0;
    XRAM[17020] = 8'b0;
    XRAM[17021] = 8'b0;
    XRAM[17022] = 8'b0;
    XRAM[17023] = 8'b0;
    XRAM[17024] = 8'b0;
    XRAM[17025] = 8'b0;
    XRAM[17026] = 8'b0;
    XRAM[17027] = 8'b0;
    XRAM[17028] = 8'b0;
    XRAM[17029] = 8'b0;
    XRAM[17030] = 8'b0;
    XRAM[17031] = 8'b0;
    XRAM[17032] = 8'b0;
    XRAM[17033] = 8'b0;
    XRAM[17034] = 8'b0;
    XRAM[17035] = 8'b0;
    XRAM[17036] = 8'b0;
    XRAM[17037] = 8'b0;
    XRAM[17038] = 8'b0;
    XRAM[17039] = 8'b0;
    XRAM[17040] = 8'b0;
    XRAM[17041] = 8'b0;
    XRAM[17042] = 8'b0;
    XRAM[17043] = 8'b0;
    XRAM[17044] = 8'b0;
    XRAM[17045] = 8'b0;
    XRAM[17046] = 8'b0;
    XRAM[17047] = 8'b0;
    XRAM[17048] = 8'b0;
    XRAM[17049] = 8'b0;
    XRAM[17050] = 8'b0;
    XRAM[17051] = 8'b0;
    XRAM[17052] = 8'b0;
    XRAM[17053] = 8'b0;
    XRAM[17054] = 8'b0;
    XRAM[17055] = 8'b0;
    XRAM[17056] = 8'b0;
    XRAM[17057] = 8'b0;
    XRAM[17058] = 8'b0;
    XRAM[17059] = 8'b0;
    XRAM[17060] = 8'b0;
    XRAM[17061] = 8'b0;
    XRAM[17062] = 8'b0;
    XRAM[17063] = 8'b0;
    XRAM[17064] = 8'b0;
    XRAM[17065] = 8'b0;
    XRAM[17066] = 8'b0;
    XRAM[17067] = 8'b0;
    XRAM[17068] = 8'b0;
    XRAM[17069] = 8'b0;
    XRAM[17070] = 8'b0;
    XRAM[17071] = 8'b0;
    XRAM[17072] = 8'b0;
    XRAM[17073] = 8'b0;
    XRAM[17074] = 8'b0;
    XRAM[17075] = 8'b0;
    XRAM[17076] = 8'b0;
    XRAM[17077] = 8'b0;
    XRAM[17078] = 8'b0;
    XRAM[17079] = 8'b0;
    XRAM[17080] = 8'b0;
    XRAM[17081] = 8'b0;
    XRAM[17082] = 8'b0;
    XRAM[17083] = 8'b0;
    XRAM[17084] = 8'b0;
    XRAM[17085] = 8'b0;
    XRAM[17086] = 8'b0;
    XRAM[17087] = 8'b0;
    XRAM[17088] = 8'b0;
    XRAM[17089] = 8'b0;
    XRAM[17090] = 8'b0;
    XRAM[17091] = 8'b0;
    XRAM[17092] = 8'b0;
    XRAM[17093] = 8'b0;
    XRAM[17094] = 8'b0;
    XRAM[17095] = 8'b0;
    XRAM[17096] = 8'b0;
    XRAM[17097] = 8'b0;
    XRAM[17098] = 8'b0;
    XRAM[17099] = 8'b0;
    XRAM[17100] = 8'b0;
    XRAM[17101] = 8'b0;
    XRAM[17102] = 8'b0;
    XRAM[17103] = 8'b0;
    XRAM[17104] = 8'b0;
    XRAM[17105] = 8'b0;
    XRAM[17106] = 8'b0;
    XRAM[17107] = 8'b0;
    XRAM[17108] = 8'b0;
    XRAM[17109] = 8'b0;
    XRAM[17110] = 8'b0;
    XRAM[17111] = 8'b0;
    XRAM[17112] = 8'b0;
    XRAM[17113] = 8'b0;
    XRAM[17114] = 8'b0;
    XRAM[17115] = 8'b0;
    XRAM[17116] = 8'b0;
    XRAM[17117] = 8'b0;
    XRAM[17118] = 8'b0;
    XRAM[17119] = 8'b0;
    XRAM[17120] = 8'b0;
    XRAM[17121] = 8'b0;
    XRAM[17122] = 8'b0;
    XRAM[17123] = 8'b0;
    XRAM[17124] = 8'b0;
    XRAM[17125] = 8'b0;
    XRAM[17126] = 8'b0;
    XRAM[17127] = 8'b0;
    XRAM[17128] = 8'b0;
    XRAM[17129] = 8'b0;
    XRAM[17130] = 8'b0;
    XRAM[17131] = 8'b0;
    XRAM[17132] = 8'b0;
    XRAM[17133] = 8'b0;
    XRAM[17134] = 8'b0;
    XRAM[17135] = 8'b0;
    XRAM[17136] = 8'b0;
    XRAM[17137] = 8'b0;
    XRAM[17138] = 8'b0;
    XRAM[17139] = 8'b0;
    XRAM[17140] = 8'b0;
    XRAM[17141] = 8'b0;
    XRAM[17142] = 8'b0;
    XRAM[17143] = 8'b0;
    XRAM[17144] = 8'b0;
    XRAM[17145] = 8'b0;
    XRAM[17146] = 8'b0;
    XRAM[17147] = 8'b0;
    XRAM[17148] = 8'b0;
    XRAM[17149] = 8'b0;
    XRAM[17150] = 8'b0;
    XRAM[17151] = 8'b0;
    XRAM[17152] = 8'b0;
    XRAM[17153] = 8'b0;
    XRAM[17154] = 8'b0;
    XRAM[17155] = 8'b0;
    XRAM[17156] = 8'b0;
    XRAM[17157] = 8'b0;
    XRAM[17158] = 8'b0;
    XRAM[17159] = 8'b0;
    XRAM[17160] = 8'b0;
    XRAM[17161] = 8'b0;
    XRAM[17162] = 8'b0;
    XRAM[17163] = 8'b0;
    XRAM[17164] = 8'b0;
    XRAM[17165] = 8'b0;
    XRAM[17166] = 8'b0;
    XRAM[17167] = 8'b0;
    XRAM[17168] = 8'b0;
    XRAM[17169] = 8'b0;
    XRAM[17170] = 8'b0;
    XRAM[17171] = 8'b0;
    XRAM[17172] = 8'b0;
    XRAM[17173] = 8'b0;
    XRAM[17174] = 8'b0;
    XRAM[17175] = 8'b0;
    XRAM[17176] = 8'b0;
    XRAM[17177] = 8'b0;
    XRAM[17178] = 8'b0;
    XRAM[17179] = 8'b0;
    XRAM[17180] = 8'b0;
    XRAM[17181] = 8'b0;
    XRAM[17182] = 8'b0;
    XRAM[17183] = 8'b0;
    XRAM[17184] = 8'b0;
    XRAM[17185] = 8'b0;
    XRAM[17186] = 8'b0;
    XRAM[17187] = 8'b0;
    XRAM[17188] = 8'b0;
    XRAM[17189] = 8'b0;
    XRAM[17190] = 8'b0;
    XRAM[17191] = 8'b0;
    XRAM[17192] = 8'b0;
    XRAM[17193] = 8'b0;
    XRAM[17194] = 8'b0;
    XRAM[17195] = 8'b0;
    XRAM[17196] = 8'b0;
    XRAM[17197] = 8'b0;
    XRAM[17198] = 8'b0;
    XRAM[17199] = 8'b0;
    XRAM[17200] = 8'b0;
    XRAM[17201] = 8'b0;
    XRAM[17202] = 8'b0;
    XRAM[17203] = 8'b0;
    XRAM[17204] = 8'b0;
    XRAM[17205] = 8'b0;
    XRAM[17206] = 8'b0;
    XRAM[17207] = 8'b0;
    XRAM[17208] = 8'b0;
    XRAM[17209] = 8'b0;
    XRAM[17210] = 8'b0;
    XRAM[17211] = 8'b0;
    XRAM[17212] = 8'b0;
    XRAM[17213] = 8'b0;
    XRAM[17214] = 8'b0;
    XRAM[17215] = 8'b0;
    XRAM[17216] = 8'b0;
    XRAM[17217] = 8'b0;
    XRAM[17218] = 8'b0;
    XRAM[17219] = 8'b0;
    XRAM[17220] = 8'b0;
    XRAM[17221] = 8'b0;
    XRAM[17222] = 8'b0;
    XRAM[17223] = 8'b0;
    XRAM[17224] = 8'b0;
    XRAM[17225] = 8'b0;
    XRAM[17226] = 8'b0;
    XRAM[17227] = 8'b0;
    XRAM[17228] = 8'b0;
    XRAM[17229] = 8'b0;
    XRAM[17230] = 8'b0;
    XRAM[17231] = 8'b0;
    XRAM[17232] = 8'b0;
    XRAM[17233] = 8'b0;
    XRAM[17234] = 8'b0;
    XRAM[17235] = 8'b0;
    XRAM[17236] = 8'b0;
    XRAM[17237] = 8'b0;
    XRAM[17238] = 8'b0;
    XRAM[17239] = 8'b0;
    XRAM[17240] = 8'b0;
    XRAM[17241] = 8'b0;
    XRAM[17242] = 8'b0;
    XRAM[17243] = 8'b0;
    XRAM[17244] = 8'b0;
    XRAM[17245] = 8'b0;
    XRAM[17246] = 8'b0;
    XRAM[17247] = 8'b0;
    XRAM[17248] = 8'b0;
    XRAM[17249] = 8'b0;
    XRAM[17250] = 8'b0;
    XRAM[17251] = 8'b0;
    XRAM[17252] = 8'b0;
    XRAM[17253] = 8'b0;
    XRAM[17254] = 8'b0;
    XRAM[17255] = 8'b0;
    XRAM[17256] = 8'b0;
    XRAM[17257] = 8'b0;
    XRAM[17258] = 8'b0;
    XRAM[17259] = 8'b0;
    XRAM[17260] = 8'b0;
    XRAM[17261] = 8'b0;
    XRAM[17262] = 8'b0;
    XRAM[17263] = 8'b0;
    XRAM[17264] = 8'b0;
    XRAM[17265] = 8'b0;
    XRAM[17266] = 8'b0;
    XRAM[17267] = 8'b0;
    XRAM[17268] = 8'b0;
    XRAM[17269] = 8'b0;
    XRAM[17270] = 8'b0;
    XRAM[17271] = 8'b0;
    XRAM[17272] = 8'b0;
    XRAM[17273] = 8'b0;
    XRAM[17274] = 8'b0;
    XRAM[17275] = 8'b0;
    XRAM[17276] = 8'b0;
    XRAM[17277] = 8'b0;
    XRAM[17278] = 8'b0;
    XRAM[17279] = 8'b0;
    XRAM[17280] = 8'b0;
    XRAM[17281] = 8'b0;
    XRAM[17282] = 8'b0;
    XRAM[17283] = 8'b0;
    XRAM[17284] = 8'b0;
    XRAM[17285] = 8'b0;
    XRAM[17286] = 8'b0;
    XRAM[17287] = 8'b0;
    XRAM[17288] = 8'b0;
    XRAM[17289] = 8'b0;
    XRAM[17290] = 8'b0;
    XRAM[17291] = 8'b0;
    XRAM[17292] = 8'b0;
    XRAM[17293] = 8'b0;
    XRAM[17294] = 8'b0;
    XRAM[17295] = 8'b0;
    XRAM[17296] = 8'b0;
    XRAM[17297] = 8'b0;
    XRAM[17298] = 8'b0;
    XRAM[17299] = 8'b0;
    XRAM[17300] = 8'b0;
    XRAM[17301] = 8'b0;
    XRAM[17302] = 8'b0;
    XRAM[17303] = 8'b0;
    XRAM[17304] = 8'b0;
    XRAM[17305] = 8'b0;
    XRAM[17306] = 8'b0;
    XRAM[17307] = 8'b0;
    XRAM[17308] = 8'b0;
    XRAM[17309] = 8'b0;
    XRAM[17310] = 8'b0;
    XRAM[17311] = 8'b0;
    XRAM[17312] = 8'b0;
    XRAM[17313] = 8'b0;
    XRAM[17314] = 8'b0;
    XRAM[17315] = 8'b0;
    XRAM[17316] = 8'b0;
    XRAM[17317] = 8'b0;
    XRAM[17318] = 8'b0;
    XRAM[17319] = 8'b0;
    XRAM[17320] = 8'b0;
    XRAM[17321] = 8'b0;
    XRAM[17322] = 8'b0;
    XRAM[17323] = 8'b0;
    XRAM[17324] = 8'b0;
    XRAM[17325] = 8'b0;
    XRAM[17326] = 8'b0;
    XRAM[17327] = 8'b0;
    XRAM[17328] = 8'b0;
    XRAM[17329] = 8'b0;
    XRAM[17330] = 8'b0;
    XRAM[17331] = 8'b0;
    XRAM[17332] = 8'b0;
    XRAM[17333] = 8'b0;
    XRAM[17334] = 8'b0;
    XRAM[17335] = 8'b0;
    XRAM[17336] = 8'b0;
    XRAM[17337] = 8'b0;
    XRAM[17338] = 8'b0;
    XRAM[17339] = 8'b0;
    XRAM[17340] = 8'b0;
    XRAM[17341] = 8'b0;
    XRAM[17342] = 8'b0;
    XRAM[17343] = 8'b0;
    XRAM[17344] = 8'b0;
    XRAM[17345] = 8'b0;
    XRAM[17346] = 8'b0;
    XRAM[17347] = 8'b0;
    XRAM[17348] = 8'b0;
    XRAM[17349] = 8'b0;
    XRAM[17350] = 8'b0;
    XRAM[17351] = 8'b0;
    XRAM[17352] = 8'b0;
    XRAM[17353] = 8'b0;
    XRAM[17354] = 8'b0;
    XRAM[17355] = 8'b0;
    XRAM[17356] = 8'b0;
    XRAM[17357] = 8'b0;
    XRAM[17358] = 8'b0;
    XRAM[17359] = 8'b0;
    XRAM[17360] = 8'b0;
    XRAM[17361] = 8'b0;
    XRAM[17362] = 8'b0;
    XRAM[17363] = 8'b0;
    XRAM[17364] = 8'b0;
    XRAM[17365] = 8'b0;
    XRAM[17366] = 8'b0;
    XRAM[17367] = 8'b0;
    XRAM[17368] = 8'b0;
    XRAM[17369] = 8'b0;
    XRAM[17370] = 8'b0;
    XRAM[17371] = 8'b0;
    XRAM[17372] = 8'b0;
    XRAM[17373] = 8'b0;
    XRAM[17374] = 8'b0;
    XRAM[17375] = 8'b0;
    XRAM[17376] = 8'b0;
    XRAM[17377] = 8'b0;
    XRAM[17378] = 8'b0;
    XRAM[17379] = 8'b0;
    XRAM[17380] = 8'b0;
    XRAM[17381] = 8'b0;
    XRAM[17382] = 8'b0;
    XRAM[17383] = 8'b0;
    XRAM[17384] = 8'b0;
    XRAM[17385] = 8'b0;
    XRAM[17386] = 8'b0;
    XRAM[17387] = 8'b0;
    XRAM[17388] = 8'b0;
    XRAM[17389] = 8'b0;
    XRAM[17390] = 8'b0;
    XRAM[17391] = 8'b0;
    XRAM[17392] = 8'b0;
    XRAM[17393] = 8'b0;
    XRAM[17394] = 8'b0;
    XRAM[17395] = 8'b0;
    XRAM[17396] = 8'b0;
    XRAM[17397] = 8'b0;
    XRAM[17398] = 8'b0;
    XRAM[17399] = 8'b0;
    XRAM[17400] = 8'b0;
    XRAM[17401] = 8'b0;
    XRAM[17402] = 8'b0;
    XRAM[17403] = 8'b0;
    XRAM[17404] = 8'b0;
    XRAM[17405] = 8'b0;
    XRAM[17406] = 8'b0;
    XRAM[17407] = 8'b0;
    XRAM[17408] = 8'b0;
    XRAM[17409] = 8'b0;
    XRAM[17410] = 8'b0;
    XRAM[17411] = 8'b0;
    XRAM[17412] = 8'b0;
    XRAM[17413] = 8'b0;
    XRAM[17414] = 8'b0;
    XRAM[17415] = 8'b0;
    XRAM[17416] = 8'b0;
    XRAM[17417] = 8'b0;
    XRAM[17418] = 8'b0;
    XRAM[17419] = 8'b0;
    XRAM[17420] = 8'b0;
    XRAM[17421] = 8'b0;
    XRAM[17422] = 8'b0;
    XRAM[17423] = 8'b0;
    XRAM[17424] = 8'b0;
    XRAM[17425] = 8'b0;
    XRAM[17426] = 8'b0;
    XRAM[17427] = 8'b0;
    XRAM[17428] = 8'b0;
    XRAM[17429] = 8'b0;
    XRAM[17430] = 8'b0;
    XRAM[17431] = 8'b0;
    XRAM[17432] = 8'b0;
    XRAM[17433] = 8'b0;
    XRAM[17434] = 8'b0;
    XRAM[17435] = 8'b0;
    XRAM[17436] = 8'b0;
    XRAM[17437] = 8'b0;
    XRAM[17438] = 8'b0;
    XRAM[17439] = 8'b0;
    XRAM[17440] = 8'b0;
    XRAM[17441] = 8'b0;
    XRAM[17442] = 8'b0;
    XRAM[17443] = 8'b0;
    XRAM[17444] = 8'b0;
    XRAM[17445] = 8'b0;
    XRAM[17446] = 8'b0;
    XRAM[17447] = 8'b0;
    XRAM[17448] = 8'b0;
    XRAM[17449] = 8'b0;
    XRAM[17450] = 8'b0;
    XRAM[17451] = 8'b0;
    XRAM[17452] = 8'b0;
    XRAM[17453] = 8'b0;
    XRAM[17454] = 8'b0;
    XRAM[17455] = 8'b0;
    XRAM[17456] = 8'b0;
    XRAM[17457] = 8'b0;
    XRAM[17458] = 8'b0;
    XRAM[17459] = 8'b0;
    XRAM[17460] = 8'b0;
    XRAM[17461] = 8'b0;
    XRAM[17462] = 8'b0;
    XRAM[17463] = 8'b0;
    XRAM[17464] = 8'b0;
    XRAM[17465] = 8'b0;
    XRAM[17466] = 8'b0;
    XRAM[17467] = 8'b0;
    XRAM[17468] = 8'b0;
    XRAM[17469] = 8'b0;
    XRAM[17470] = 8'b0;
    XRAM[17471] = 8'b0;
    XRAM[17472] = 8'b0;
    XRAM[17473] = 8'b0;
    XRAM[17474] = 8'b0;
    XRAM[17475] = 8'b0;
    XRAM[17476] = 8'b0;
    XRAM[17477] = 8'b0;
    XRAM[17478] = 8'b0;
    XRAM[17479] = 8'b0;
    XRAM[17480] = 8'b0;
    XRAM[17481] = 8'b0;
    XRAM[17482] = 8'b0;
    XRAM[17483] = 8'b0;
    XRAM[17484] = 8'b0;
    XRAM[17485] = 8'b0;
    XRAM[17486] = 8'b0;
    XRAM[17487] = 8'b0;
    XRAM[17488] = 8'b0;
    XRAM[17489] = 8'b0;
    XRAM[17490] = 8'b0;
    XRAM[17491] = 8'b0;
    XRAM[17492] = 8'b0;
    XRAM[17493] = 8'b0;
    XRAM[17494] = 8'b0;
    XRAM[17495] = 8'b0;
    XRAM[17496] = 8'b0;
    XRAM[17497] = 8'b0;
    XRAM[17498] = 8'b0;
    XRAM[17499] = 8'b0;
    XRAM[17500] = 8'b0;
    XRAM[17501] = 8'b0;
    XRAM[17502] = 8'b0;
    XRAM[17503] = 8'b0;
    XRAM[17504] = 8'b0;
    XRAM[17505] = 8'b0;
    XRAM[17506] = 8'b0;
    XRAM[17507] = 8'b0;
    XRAM[17508] = 8'b0;
    XRAM[17509] = 8'b0;
    XRAM[17510] = 8'b0;
    XRAM[17511] = 8'b0;
    XRAM[17512] = 8'b0;
    XRAM[17513] = 8'b0;
    XRAM[17514] = 8'b0;
    XRAM[17515] = 8'b0;
    XRAM[17516] = 8'b0;
    XRAM[17517] = 8'b0;
    XRAM[17518] = 8'b0;
    XRAM[17519] = 8'b0;
    XRAM[17520] = 8'b0;
    XRAM[17521] = 8'b0;
    XRAM[17522] = 8'b0;
    XRAM[17523] = 8'b0;
    XRAM[17524] = 8'b0;
    XRAM[17525] = 8'b0;
    XRAM[17526] = 8'b0;
    XRAM[17527] = 8'b0;
    XRAM[17528] = 8'b0;
    XRAM[17529] = 8'b0;
    XRAM[17530] = 8'b0;
    XRAM[17531] = 8'b0;
    XRAM[17532] = 8'b0;
    XRAM[17533] = 8'b0;
    XRAM[17534] = 8'b0;
    XRAM[17535] = 8'b0;
    XRAM[17536] = 8'b0;
    XRAM[17537] = 8'b0;
    XRAM[17538] = 8'b0;
    XRAM[17539] = 8'b0;
    XRAM[17540] = 8'b0;
    XRAM[17541] = 8'b0;
    XRAM[17542] = 8'b0;
    XRAM[17543] = 8'b0;
    XRAM[17544] = 8'b0;
    XRAM[17545] = 8'b0;
    XRAM[17546] = 8'b0;
    XRAM[17547] = 8'b0;
    XRAM[17548] = 8'b0;
    XRAM[17549] = 8'b0;
    XRAM[17550] = 8'b0;
    XRAM[17551] = 8'b0;
    XRAM[17552] = 8'b0;
    XRAM[17553] = 8'b0;
    XRAM[17554] = 8'b0;
    XRAM[17555] = 8'b0;
    XRAM[17556] = 8'b0;
    XRAM[17557] = 8'b0;
    XRAM[17558] = 8'b0;
    XRAM[17559] = 8'b0;
    XRAM[17560] = 8'b0;
    XRAM[17561] = 8'b0;
    XRAM[17562] = 8'b0;
    XRAM[17563] = 8'b0;
    XRAM[17564] = 8'b0;
    XRAM[17565] = 8'b0;
    XRAM[17566] = 8'b0;
    XRAM[17567] = 8'b0;
    XRAM[17568] = 8'b0;
    XRAM[17569] = 8'b0;
    XRAM[17570] = 8'b0;
    XRAM[17571] = 8'b0;
    XRAM[17572] = 8'b0;
    XRAM[17573] = 8'b0;
    XRAM[17574] = 8'b0;
    XRAM[17575] = 8'b0;
    XRAM[17576] = 8'b0;
    XRAM[17577] = 8'b0;
    XRAM[17578] = 8'b0;
    XRAM[17579] = 8'b0;
    XRAM[17580] = 8'b0;
    XRAM[17581] = 8'b0;
    XRAM[17582] = 8'b0;
    XRAM[17583] = 8'b0;
    XRAM[17584] = 8'b0;
    XRAM[17585] = 8'b0;
    XRAM[17586] = 8'b0;
    XRAM[17587] = 8'b0;
    XRAM[17588] = 8'b0;
    XRAM[17589] = 8'b0;
    XRAM[17590] = 8'b0;
    XRAM[17591] = 8'b0;
    XRAM[17592] = 8'b0;
    XRAM[17593] = 8'b0;
    XRAM[17594] = 8'b0;
    XRAM[17595] = 8'b0;
    XRAM[17596] = 8'b0;
    XRAM[17597] = 8'b0;
    XRAM[17598] = 8'b0;
    XRAM[17599] = 8'b0;
    XRAM[17600] = 8'b0;
    XRAM[17601] = 8'b0;
    XRAM[17602] = 8'b0;
    XRAM[17603] = 8'b0;
    XRAM[17604] = 8'b0;
    XRAM[17605] = 8'b0;
    XRAM[17606] = 8'b0;
    XRAM[17607] = 8'b0;
    XRAM[17608] = 8'b0;
    XRAM[17609] = 8'b0;
    XRAM[17610] = 8'b0;
    XRAM[17611] = 8'b0;
    XRAM[17612] = 8'b0;
    XRAM[17613] = 8'b0;
    XRAM[17614] = 8'b0;
    XRAM[17615] = 8'b0;
    XRAM[17616] = 8'b0;
    XRAM[17617] = 8'b0;
    XRAM[17618] = 8'b0;
    XRAM[17619] = 8'b0;
    XRAM[17620] = 8'b0;
    XRAM[17621] = 8'b0;
    XRAM[17622] = 8'b0;
    XRAM[17623] = 8'b0;
    XRAM[17624] = 8'b0;
    XRAM[17625] = 8'b0;
    XRAM[17626] = 8'b0;
    XRAM[17627] = 8'b0;
    XRAM[17628] = 8'b0;
    XRAM[17629] = 8'b0;
    XRAM[17630] = 8'b0;
    XRAM[17631] = 8'b0;
    XRAM[17632] = 8'b0;
    XRAM[17633] = 8'b0;
    XRAM[17634] = 8'b0;
    XRAM[17635] = 8'b0;
    XRAM[17636] = 8'b0;
    XRAM[17637] = 8'b0;
    XRAM[17638] = 8'b0;
    XRAM[17639] = 8'b0;
    XRAM[17640] = 8'b0;
    XRAM[17641] = 8'b0;
    XRAM[17642] = 8'b0;
    XRAM[17643] = 8'b0;
    XRAM[17644] = 8'b0;
    XRAM[17645] = 8'b0;
    XRAM[17646] = 8'b0;
    XRAM[17647] = 8'b0;
    XRAM[17648] = 8'b0;
    XRAM[17649] = 8'b0;
    XRAM[17650] = 8'b0;
    XRAM[17651] = 8'b0;
    XRAM[17652] = 8'b0;
    XRAM[17653] = 8'b0;
    XRAM[17654] = 8'b0;
    XRAM[17655] = 8'b0;
    XRAM[17656] = 8'b0;
    XRAM[17657] = 8'b0;
    XRAM[17658] = 8'b0;
    XRAM[17659] = 8'b0;
    XRAM[17660] = 8'b0;
    XRAM[17661] = 8'b0;
    XRAM[17662] = 8'b0;
    XRAM[17663] = 8'b0;
    XRAM[17664] = 8'b0;
    XRAM[17665] = 8'b0;
    XRAM[17666] = 8'b0;
    XRAM[17667] = 8'b0;
    XRAM[17668] = 8'b0;
    XRAM[17669] = 8'b0;
    XRAM[17670] = 8'b0;
    XRAM[17671] = 8'b0;
    XRAM[17672] = 8'b0;
    XRAM[17673] = 8'b0;
    XRAM[17674] = 8'b0;
    XRAM[17675] = 8'b0;
    XRAM[17676] = 8'b0;
    XRAM[17677] = 8'b0;
    XRAM[17678] = 8'b0;
    XRAM[17679] = 8'b0;
    XRAM[17680] = 8'b0;
    XRAM[17681] = 8'b0;
    XRAM[17682] = 8'b0;
    XRAM[17683] = 8'b0;
    XRAM[17684] = 8'b0;
    XRAM[17685] = 8'b0;
    XRAM[17686] = 8'b0;
    XRAM[17687] = 8'b0;
    XRAM[17688] = 8'b0;
    XRAM[17689] = 8'b0;
    XRAM[17690] = 8'b0;
    XRAM[17691] = 8'b0;
    XRAM[17692] = 8'b0;
    XRAM[17693] = 8'b0;
    XRAM[17694] = 8'b0;
    XRAM[17695] = 8'b0;
    XRAM[17696] = 8'b0;
    XRAM[17697] = 8'b0;
    XRAM[17698] = 8'b0;
    XRAM[17699] = 8'b0;
    XRAM[17700] = 8'b0;
    XRAM[17701] = 8'b0;
    XRAM[17702] = 8'b0;
    XRAM[17703] = 8'b0;
    XRAM[17704] = 8'b0;
    XRAM[17705] = 8'b0;
    XRAM[17706] = 8'b0;
    XRAM[17707] = 8'b0;
    XRAM[17708] = 8'b0;
    XRAM[17709] = 8'b0;
    XRAM[17710] = 8'b0;
    XRAM[17711] = 8'b0;
    XRAM[17712] = 8'b0;
    XRAM[17713] = 8'b0;
    XRAM[17714] = 8'b0;
    XRAM[17715] = 8'b0;
    XRAM[17716] = 8'b0;
    XRAM[17717] = 8'b0;
    XRAM[17718] = 8'b0;
    XRAM[17719] = 8'b0;
    XRAM[17720] = 8'b0;
    XRAM[17721] = 8'b0;
    XRAM[17722] = 8'b0;
    XRAM[17723] = 8'b0;
    XRAM[17724] = 8'b0;
    XRAM[17725] = 8'b0;
    XRAM[17726] = 8'b0;
    XRAM[17727] = 8'b0;
    XRAM[17728] = 8'b0;
    XRAM[17729] = 8'b0;
    XRAM[17730] = 8'b0;
    XRAM[17731] = 8'b0;
    XRAM[17732] = 8'b0;
    XRAM[17733] = 8'b0;
    XRAM[17734] = 8'b0;
    XRAM[17735] = 8'b0;
    XRAM[17736] = 8'b0;
    XRAM[17737] = 8'b0;
    XRAM[17738] = 8'b0;
    XRAM[17739] = 8'b0;
    XRAM[17740] = 8'b0;
    XRAM[17741] = 8'b0;
    XRAM[17742] = 8'b0;
    XRAM[17743] = 8'b0;
    XRAM[17744] = 8'b0;
    XRAM[17745] = 8'b0;
    XRAM[17746] = 8'b0;
    XRAM[17747] = 8'b0;
    XRAM[17748] = 8'b0;
    XRAM[17749] = 8'b0;
    XRAM[17750] = 8'b0;
    XRAM[17751] = 8'b0;
    XRAM[17752] = 8'b0;
    XRAM[17753] = 8'b0;
    XRAM[17754] = 8'b0;
    XRAM[17755] = 8'b0;
    XRAM[17756] = 8'b0;
    XRAM[17757] = 8'b0;
    XRAM[17758] = 8'b0;
    XRAM[17759] = 8'b0;
    XRAM[17760] = 8'b0;
    XRAM[17761] = 8'b0;
    XRAM[17762] = 8'b0;
    XRAM[17763] = 8'b0;
    XRAM[17764] = 8'b0;
    XRAM[17765] = 8'b0;
    XRAM[17766] = 8'b0;
    XRAM[17767] = 8'b0;
    XRAM[17768] = 8'b0;
    XRAM[17769] = 8'b0;
    XRAM[17770] = 8'b0;
    XRAM[17771] = 8'b0;
    XRAM[17772] = 8'b0;
    XRAM[17773] = 8'b0;
    XRAM[17774] = 8'b0;
    XRAM[17775] = 8'b0;
    XRAM[17776] = 8'b0;
    XRAM[17777] = 8'b0;
    XRAM[17778] = 8'b0;
    XRAM[17779] = 8'b0;
    XRAM[17780] = 8'b0;
    XRAM[17781] = 8'b0;
    XRAM[17782] = 8'b0;
    XRAM[17783] = 8'b0;
    XRAM[17784] = 8'b0;
    XRAM[17785] = 8'b0;
    XRAM[17786] = 8'b0;
    XRAM[17787] = 8'b0;
    XRAM[17788] = 8'b0;
    XRAM[17789] = 8'b0;
    XRAM[17790] = 8'b0;
    XRAM[17791] = 8'b0;
    XRAM[17792] = 8'b0;
    XRAM[17793] = 8'b0;
    XRAM[17794] = 8'b0;
    XRAM[17795] = 8'b0;
    XRAM[17796] = 8'b0;
    XRAM[17797] = 8'b0;
    XRAM[17798] = 8'b0;
    XRAM[17799] = 8'b0;
    XRAM[17800] = 8'b0;
    XRAM[17801] = 8'b0;
    XRAM[17802] = 8'b0;
    XRAM[17803] = 8'b0;
    XRAM[17804] = 8'b0;
    XRAM[17805] = 8'b0;
    XRAM[17806] = 8'b0;
    XRAM[17807] = 8'b0;
    XRAM[17808] = 8'b0;
    XRAM[17809] = 8'b0;
    XRAM[17810] = 8'b0;
    XRAM[17811] = 8'b0;
    XRAM[17812] = 8'b0;
    XRAM[17813] = 8'b0;
    XRAM[17814] = 8'b0;
    XRAM[17815] = 8'b0;
    XRAM[17816] = 8'b0;
    XRAM[17817] = 8'b0;
    XRAM[17818] = 8'b0;
    XRAM[17819] = 8'b0;
    XRAM[17820] = 8'b0;
    XRAM[17821] = 8'b0;
    XRAM[17822] = 8'b0;
    XRAM[17823] = 8'b0;
    XRAM[17824] = 8'b0;
    XRAM[17825] = 8'b0;
    XRAM[17826] = 8'b0;
    XRAM[17827] = 8'b0;
    XRAM[17828] = 8'b0;
    XRAM[17829] = 8'b0;
    XRAM[17830] = 8'b0;
    XRAM[17831] = 8'b0;
    XRAM[17832] = 8'b0;
    XRAM[17833] = 8'b0;
    XRAM[17834] = 8'b0;
    XRAM[17835] = 8'b0;
    XRAM[17836] = 8'b0;
    XRAM[17837] = 8'b0;
    XRAM[17838] = 8'b0;
    XRAM[17839] = 8'b0;
    XRAM[17840] = 8'b0;
    XRAM[17841] = 8'b0;
    XRAM[17842] = 8'b0;
    XRAM[17843] = 8'b0;
    XRAM[17844] = 8'b0;
    XRAM[17845] = 8'b0;
    XRAM[17846] = 8'b0;
    XRAM[17847] = 8'b0;
    XRAM[17848] = 8'b0;
    XRAM[17849] = 8'b0;
    XRAM[17850] = 8'b0;
    XRAM[17851] = 8'b0;
    XRAM[17852] = 8'b0;
    XRAM[17853] = 8'b0;
    XRAM[17854] = 8'b0;
    XRAM[17855] = 8'b0;
    XRAM[17856] = 8'b0;
    XRAM[17857] = 8'b0;
    XRAM[17858] = 8'b0;
    XRAM[17859] = 8'b0;
    XRAM[17860] = 8'b0;
    XRAM[17861] = 8'b0;
    XRAM[17862] = 8'b0;
    XRAM[17863] = 8'b0;
    XRAM[17864] = 8'b0;
    XRAM[17865] = 8'b0;
    XRAM[17866] = 8'b0;
    XRAM[17867] = 8'b0;
    XRAM[17868] = 8'b0;
    XRAM[17869] = 8'b0;
    XRAM[17870] = 8'b0;
    XRAM[17871] = 8'b0;
    XRAM[17872] = 8'b0;
    XRAM[17873] = 8'b0;
    XRAM[17874] = 8'b0;
    XRAM[17875] = 8'b0;
    XRAM[17876] = 8'b0;
    XRAM[17877] = 8'b0;
    XRAM[17878] = 8'b0;
    XRAM[17879] = 8'b0;
    XRAM[17880] = 8'b0;
    XRAM[17881] = 8'b0;
    XRAM[17882] = 8'b0;
    XRAM[17883] = 8'b0;
    XRAM[17884] = 8'b0;
    XRAM[17885] = 8'b0;
    XRAM[17886] = 8'b0;
    XRAM[17887] = 8'b0;
    XRAM[17888] = 8'b0;
    XRAM[17889] = 8'b0;
    XRAM[17890] = 8'b0;
    XRAM[17891] = 8'b0;
    XRAM[17892] = 8'b0;
    XRAM[17893] = 8'b0;
    XRAM[17894] = 8'b0;
    XRAM[17895] = 8'b0;
    XRAM[17896] = 8'b0;
    XRAM[17897] = 8'b0;
    XRAM[17898] = 8'b0;
    XRAM[17899] = 8'b0;
    XRAM[17900] = 8'b0;
    XRAM[17901] = 8'b0;
    XRAM[17902] = 8'b0;
    XRAM[17903] = 8'b0;
    XRAM[17904] = 8'b0;
    XRAM[17905] = 8'b0;
    XRAM[17906] = 8'b0;
    XRAM[17907] = 8'b0;
    XRAM[17908] = 8'b0;
    XRAM[17909] = 8'b0;
    XRAM[17910] = 8'b0;
    XRAM[17911] = 8'b0;
    XRAM[17912] = 8'b0;
    XRAM[17913] = 8'b0;
    XRAM[17914] = 8'b0;
    XRAM[17915] = 8'b0;
    XRAM[17916] = 8'b0;
    XRAM[17917] = 8'b0;
    XRAM[17918] = 8'b0;
    XRAM[17919] = 8'b0;
    XRAM[17920] = 8'b0;
    XRAM[17921] = 8'b0;
    XRAM[17922] = 8'b0;
    XRAM[17923] = 8'b0;
    XRAM[17924] = 8'b0;
    XRAM[17925] = 8'b0;
    XRAM[17926] = 8'b0;
    XRAM[17927] = 8'b0;
    XRAM[17928] = 8'b0;
    XRAM[17929] = 8'b0;
    XRAM[17930] = 8'b0;
    XRAM[17931] = 8'b0;
    XRAM[17932] = 8'b0;
    XRAM[17933] = 8'b0;
    XRAM[17934] = 8'b0;
    XRAM[17935] = 8'b0;
    XRAM[17936] = 8'b0;
    XRAM[17937] = 8'b0;
    XRAM[17938] = 8'b0;
    XRAM[17939] = 8'b0;
    XRAM[17940] = 8'b0;
    XRAM[17941] = 8'b0;
    XRAM[17942] = 8'b0;
    XRAM[17943] = 8'b0;
    XRAM[17944] = 8'b0;
    XRAM[17945] = 8'b0;
    XRAM[17946] = 8'b0;
    XRAM[17947] = 8'b0;
    XRAM[17948] = 8'b0;
    XRAM[17949] = 8'b0;
    XRAM[17950] = 8'b0;
    XRAM[17951] = 8'b0;
    XRAM[17952] = 8'b0;
    XRAM[17953] = 8'b0;
    XRAM[17954] = 8'b0;
    XRAM[17955] = 8'b0;
    XRAM[17956] = 8'b0;
    XRAM[17957] = 8'b0;
    XRAM[17958] = 8'b0;
    XRAM[17959] = 8'b0;
    XRAM[17960] = 8'b0;
    XRAM[17961] = 8'b0;
    XRAM[17962] = 8'b0;
    XRAM[17963] = 8'b0;
    XRAM[17964] = 8'b0;
    XRAM[17965] = 8'b0;
    XRAM[17966] = 8'b0;
    XRAM[17967] = 8'b0;
    XRAM[17968] = 8'b0;
    XRAM[17969] = 8'b0;
    XRAM[17970] = 8'b0;
    XRAM[17971] = 8'b0;
    XRAM[17972] = 8'b0;
    XRAM[17973] = 8'b0;
    XRAM[17974] = 8'b0;
    XRAM[17975] = 8'b0;
    XRAM[17976] = 8'b0;
    XRAM[17977] = 8'b0;
    XRAM[17978] = 8'b0;
    XRAM[17979] = 8'b0;
    XRAM[17980] = 8'b0;
    XRAM[17981] = 8'b0;
    XRAM[17982] = 8'b0;
    XRAM[17983] = 8'b0;
    XRAM[17984] = 8'b0;
    XRAM[17985] = 8'b0;
    XRAM[17986] = 8'b0;
    XRAM[17987] = 8'b0;
    XRAM[17988] = 8'b0;
    XRAM[17989] = 8'b0;
    XRAM[17990] = 8'b0;
    XRAM[17991] = 8'b0;
    XRAM[17992] = 8'b0;
    XRAM[17993] = 8'b0;
    XRAM[17994] = 8'b0;
    XRAM[17995] = 8'b0;
    XRAM[17996] = 8'b0;
    XRAM[17997] = 8'b0;
    XRAM[17998] = 8'b0;
    XRAM[17999] = 8'b0;
    XRAM[18000] = 8'b0;
    XRAM[18001] = 8'b0;
    XRAM[18002] = 8'b0;
    XRAM[18003] = 8'b0;
    XRAM[18004] = 8'b0;
    XRAM[18005] = 8'b0;
    XRAM[18006] = 8'b0;
    XRAM[18007] = 8'b0;
    XRAM[18008] = 8'b0;
    XRAM[18009] = 8'b0;
    XRAM[18010] = 8'b0;
    XRAM[18011] = 8'b0;
    XRAM[18012] = 8'b0;
    XRAM[18013] = 8'b0;
    XRAM[18014] = 8'b0;
    XRAM[18015] = 8'b0;
    XRAM[18016] = 8'b0;
    XRAM[18017] = 8'b0;
    XRAM[18018] = 8'b0;
    XRAM[18019] = 8'b0;
    XRAM[18020] = 8'b0;
    XRAM[18021] = 8'b0;
    XRAM[18022] = 8'b0;
    XRAM[18023] = 8'b0;
    XRAM[18024] = 8'b0;
    XRAM[18025] = 8'b0;
    XRAM[18026] = 8'b0;
    XRAM[18027] = 8'b0;
    XRAM[18028] = 8'b0;
    XRAM[18029] = 8'b0;
    XRAM[18030] = 8'b0;
    XRAM[18031] = 8'b0;
    XRAM[18032] = 8'b0;
    XRAM[18033] = 8'b0;
    XRAM[18034] = 8'b0;
    XRAM[18035] = 8'b0;
    XRAM[18036] = 8'b0;
    XRAM[18037] = 8'b0;
    XRAM[18038] = 8'b0;
    XRAM[18039] = 8'b0;
    XRAM[18040] = 8'b0;
    XRAM[18041] = 8'b0;
    XRAM[18042] = 8'b0;
    XRAM[18043] = 8'b0;
    XRAM[18044] = 8'b0;
    XRAM[18045] = 8'b0;
    XRAM[18046] = 8'b0;
    XRAM[18047] = 8'b0;
    XRAM[18048] = 8'b0;
    XRAM[18049] = 8'b0;
    XRAM[18050] = 8'b0;
    XRAM[18051] = 8'b0;
    XRAM[18052] = 8'b0;
    XRAM[18053] = 8'b0;
    XRAM[18054] = 8'b0;
    XRAM[18055] = 8'b0;
    XRAM[18056] = 8'b0;
    XRAM[18057] = 8'b0;
    XRAM[18058] = 8'b0;
    XRAM[18059] = 8'b0;
    XRAM[18060] = 8'b0;
    XRAM[18061] = 8'b0;
    XRAM[18062] = 8'b0;
    XRAM[18063] = 8'b0;
    XRAM[18064] = 8'b0;
    XRAM[18065] = 8'b0;
    XRAM[18066] = 8'b0;
    XRAM[18067] = 8'b0;
    XRAM[18068] = 8'b0;
    XRAM[18069] = 8'b0;
    XRAM[18070] = 8'b0;
    XRAM[18071] = 8'b0;
    XRAM[18072] = 8'b0;
    XRAM[18073] = 8'b0;
    XRAM[18074] = 8'b0;
    XRAM[18075] = 8'b0;
    XRAM[18076] = 8'b0;
    XRAM[18077] = 8'b0;
    XRAM[18078] = 8'b0;
    XRAM[18079] = 8'b0;
    XRAM[18080] = 8'b0;
    XRAM[18081] = 8'b0;
    XRAM[18082] = 8'b0;
    XRAM[18083] = 8'b0;
    XRAM[18084] = 8'b0;
    XRAM[18085] = 8'b0;
    XRAM[18086] = 8'b0;
    XRAM[18087] = 8'b0;
    XRAM[18088] = 8'b0;
    XRAM[18089] = 8'b0;
    XRAM[18090] = 8'b0;
    XRAM[18091] = 8'b0;
    XRAM[18092] = 8'b0;
    XRAM[18093] = 8'b0;
    XRAM[18094] = 8'b0;
    XRAM[18095] = 8'b0;
    XRAM[18096] = 8'b0;
    XRAM[18097] = 8'b0;
    XRAM[18098] = 8'b0;
    XRAM[18099] = 8'b0;
    XRAM[18100] = 8'b0;
    XRAM[18101] = 8'b0;
    XRAM[18102] = 8'b0;
    XRAM[18103] = 8'b0;
    XRAM[18104] = 8'b0;
    XRAM[18105] = 8'b0;
    XRAM[18106] = 8'b0;
    XRAM[18107] = 8'b0;
    XRAM[18108] = 8'b0;
    XRAM[18109] = 8'b0;
    XRAM[18110] = 8'b0;
    XRAM[18111] = 8'b0;
    XRAM[18112] = 8'b0;
    XRAM[18113] = 8'b0;
    XRAM[18114] = 8'b0;
    XRAM[18115] = 8'b0;
    XRAM[18116] = 8'b0;
    XRAM[18117] = 8'b0;
    XRAM[18118] = 8'b0;
    XRAM[18119] = 8'b0;
    XRAM[18120] = 8'b0;
    XRAM[18121] = 8'b0;
    XRAM[18122] = 8'b0;
    XRAM[18123] = 8'b0;
    XRAM[18124] = 8'b0;
    XRAM[18125] = 8'b0;
    XRAM[18126] = 8'b0;
    XRAM[18127] = 8'b0;
    XRAM[18128] = 8'b0;
    XRAM[18129] = 8'b0;
    XRAM[18130] = 8'b0;
    XRAM[18131] = 8'b0;
    XRAM[18132] = 8'b0;
    XRAM[18133] = 8'b0;
    XRAM[18134] = 8'b0;
    XRAM[18135] = 8'b0;
    XRAM[18136] = 8'b0;
    XRAM[18137] = 8'b0;
    XRAM[18138] = 8'b0;
    XRAM[18139] = 8'b0;
    XRAM[18140] = 8'b0;
    XRAM[18141] = 8'b0;
    XRAM[18142] = 8'b0;
    XRAM[18143] = 8'b0;
    XRAM[18144] = 8'b0;
    XRAM[18145] = 8'b0;
    XRAM[18146] = 8'b0;
    XRAM[18147] = 8'b0;
    XRAM[18148] = 8'b0;
    XRAM[18149] = 8'b0;
    XRAM[18150] = 8'b0;
    XRAM[18151] = 8'b0;
    XRAM[18152] = 8'b0;
    XRAM[18153] = 8'b0;
    XRAM[18154] = 8'b0;
    XRAM[18155] = 8'b0;
    XRAM[18156] = 8'b0;
    XRAM[18157] = 8'b0;
    XRAM[18158] = 8'b0;
    XRAM[18159] = 8'b0;
    XRAM[18160] = 8'b0;
    XRAM[18161] = 8'b0;
    XRAM[18162] = 8'b0;
    XRAM[18163] = 8'b0;
    XRAM[18164] = 8'b0;
    XRAM[18165] = 8'b0;
    XRAM[18166] = 8'b0;
    XRAM[18167] = 8'b0;
    XRAM[18168] = 8'b0;
    XRAM[18169] = 8'b0;
    XRAM[18170] = 8'b0;
    XRAM[18171] = 8'b0;
    XRAM[18172] = 8'b0;
    XRAM[18173] = 8'b0;
    XRAM[18174] = 8'b0;
    XRAM[18175] = 8'b0;
    XRAM[18176] = 8'b0;
    XRAM[18177] = 8'b0;
    XRAM[18178] = 8'b0;
    XRAM[18179] = 8'b0;
    XRAM[18180] = 8'b0;
    XRAM[18181] = 8'b0;
    XRAM[18182] = 8'b0;
    XRAM[18183] = 8'b0;
    XRAM[18184] = 8'b0;
    XRAM[18185] = 8'b0;
    XRAM[18186] = 8'b0;
    XRAM[18187] = 8'b0;
    XRAM[18188] = 8'b0;
    XRAM[18189] = 8'b0;
    XRAM[18190] = 8'b0;
    XRAM[18191] = 8'b0;
    XRAM[18192] = 8'b0;
    XRAM[18193] = 8'b0;
    XRAM[18194] = 8'b0;
    XRAM[18195] = 8'b0;
    XRAM[18196] = 8'b0;
    XRAM[18197] = 8'b0;
    XRAM[18198] = 8'b0;
    XRAM[18199] = 8'b0;
    XRAM[18200] = 8'b0;
    XRAM[18201] = 8'b0;
    XRAM[18202] = 8'b0;
    XRAM[18203] = 8'b0;
    XRAM[18204] = 8'b0;
    XRAM[18205] = 8'b0;
    XRAM[18206] = 8'b0;
    XRAM[18207] = 8'b0;
    XRAM[18208] = 8'b0;
    XRAM[18209] = 8'b0;
    XRAM[18210] = 8'b0;
    XRAM[18211] = 8'b0;
    XRAM[18212] = 8'b0;
    XRAM[18213] = 8'b0;
    XRAM[18214] = 8'b0;
    XRAM[18215] = 8'b0;
    XRAM[18216] = 8'b0;
    XRAM[18217] = 8'b0;
    XRAM[18218] = 8'b0;
    XRAM[18219] = 8'b0;
    XRAM[18220] = 8'b0;
    XRAM[18221] = 8'b0;
    XRAM[18222] = 8'b0;
    XRAM[18223] = 8'b0;
    XRAM[18224] = 8'b0;
    XRAM[18225] = 8'b0;
    XRAM[18226] = 8'b0;
    XRAM[18227] = 8'b0;
    XRAM[18228] = 8'b0;
    XRAM[18229] = 8'b0;
    XRAM[18230] = 8'b0;
    XRAM[18231] = 8'b0;
    XRAM[18232] = 8'b0;
    XRAM[18233] = 8'b0;
    XRAM[18234] = 8'b0;
    XRAM[18235] = 8'b0;
    XRAM[18236] = 8'b0;
    XRAM[18237] = 8'b0;
    XRAM[18238] = 8'b0;
    XRAM[18239] = 8'b0;
    XRAM[18240] = 8'b0;
    XRAM[18241] = 8'b0;
    XRAM[18242] = 8'b0;
    XRAM[18243] = 8'b0;
    XRAM[18244] = 8'b0;
    XRAM[18245] = 8'b0;
    XRAM[18246] = 8'b0;
    XRAM[18247] = 8'b0;
    XRAM[18248] = 8'b0;
    XRAM[18249] = 8'b0;
    XRAM[18250] = 8'b0;
    XRAM[18251] = 8'b0;
    XRAM[18252] = 8'b0;
    XRAM[18253] = 8'b0;
    XRAM[18254] = 8'b0;
    XRAM[18255] = 8'b0;
    XRAM[18256] = 8'b0;
    XRAM[18257] = 8'b0;
    XRAM[18258] = 8'b0;
    XRAM[18259] = 8'b0;
    XRAM[18260] = 8'b0;
    XRAM[18261] = 8'b0;
    XRAM[18262] = 8'b0;
    XRAM[18263] = 8'b0;
    XRAM[18264] = 8'b0;
    XRAM[18265] = 8'b0;
    XRAM[18266] = 8'b0;
    XRAM[18267] = 8'b0;
    XRAM[18268] = 8'b0;
    XRAM[18269] = 8'b0;
    XRAM[18270] = 8'b0;
    XRAM[18271] = 8'b0;
    XRAM[18272] = 8'b0;
    XRAM[18273] = 8'b0;
    XRAM[18274] = 8'b0;
    XRAM[18275] = 8'b0;
    XRAM[18276] = 8'b0;
    XRAM[18277] = 8'b0;
    XRAM[18278] = 8'b0;
    XRAM[18279] = 8'b0;
    XRAM[18280] = 8'b0;
    XRAM[18281] = 8'b0;
    XRAM[18282] = 8'b0;
    XRAM[18283] = 8'b0;
    XRAM[18284] = 8'b0;
    XRAM[18285] = 8'b0;
    XRAM[18286] = 8'b0;
    XRAM[18287] = 8'b0;
    XRAM[18288] = 8'b0;
    XRAM[18289] = 8'b0;
    XRAM[18290] = 8'b0;
    XRAM[18291] = 8'b0;
    XRAM[18292] = 8'b0;
    XRAM[18293] = 8'b0;
    XRAM[18294] = 8'b0;
    XRAM[18295] = 8'b0;
    XRAM[18296] = 8'b0;
    XRAM[18297] = 8'b0;
    XRAM[18298] = 8'b0;
    XRAM[18299] = 8'b0;
    XRAM[18300] = 8'b0;
    XRAM[18301] = 8'b0;
    XRAM[18302] = 8'b0;
    XRAM[18303] = 8'b0;
    XRAM[18304] = 8'b0;
    XRAM[18305] = 8'b0;
    XRAM[18306] = 8'b0;
    XRAM[18307] = 8'b0;
    XRAM[18308] = 8'b0;
    XRAM[18309] = 8'b0;
    XRAM[18310] = 8'b0;
    XRAM[18311] = 8'b0;
    XRAM[18312] = 8'b0;
    XRAM[18313] = 8'b0;
    XRAM[18314] = 8'b0;
    XRAM[18315] = 8'b0;
    XRAM[18316] = 8'b0;
    XRAM[18317] = 8'b0;
    XRAM[18318] = 8'b0;
    XRAM[18319] = 8'b0;
    XRAM[18320] = 8'b0;
    XRAM[18321] = 8'b0;
    XRAM[18322] = 8'b0;
    XRAM[18323] = 8'b0;
    XRAM[18324] = 8'b0;
    XRAM[18325] = 8'b0;
    XRAM[18326] = 8'b0;
    XRAM[18327] = 8'b0;
    XRAM[18328] = 8'b0;
    XRAM[18329] = 8'b0;
    XRAM[18330] = 8'b0;
    XRAM[18331] = 8'b0;
    XRAM[18332] = 8'b0;
    XRAM[18333] = 8'b0;
    XRAM[18334] = 8'b0;
    XRAM[18335] = 8'b0;
    XRAM[18336] = 8'b0;
    XRAM[18337] = 8'b0;
    XRAM[18338] = 8'b0;
    XRAM[18339] = 8'b0;
    XRAM[18340] = 8'b0;
    XRAM[18341] = 8'b0;
    XRAM[18342] = 8'b0;
    XRAM[18343] = 8'b0;
    XRAM[18344] = 8'b0;
    XRAM[18345] = 8'b0;
    XRAM[18346] = 8'b0;
    XRAM[18347] = 8'b0;
    XRAM[18348] = 8'b0;
    XRAM[18349] = 8'b0;
    XRAM[18350] = 8'b0;
    XRAM[18351] = 8'b0;
    XRAM[18352] = 8'b0;
    XRAM[18353] = 8'b0;
    XRAM[18354] = 8'b0;
    XRAM[18355] = 8'b0;
    XRAM[18356] = 8'b0;
    XRAM[18357] = 8'b0;
    XRAM[18358] = 8'b0;
    XRAM[18359] = 8'b0;
    XRAM[18360] = 8'b0;
    XRAM[18361] = 8'b0;
    XRAM[18362] = 8'b0;
    XRAM[18363] = 8'b0;
    XRAM[18364] = 8'b0;
    XRAM[18365] = 8'b0;
    XRAM[18366] = 8'b0;
    XRAM[18367] = 8'b0;
    XRAM[18368] = 8'b0;
    XRAM[18369] = 8'b0;
    XRAM[18370] = 8'b0;
    XRAM[18371] = 8'b0;
    XRAM[18372] = 8'b0;
    XRAM[18373] = 8'b0;
    XRAM[18374] = 8'b0;
    XRAM[18375] = 8'b0;
    XRAM[18376] = 8'b0;
    XRAM[18377] = 8'b0;
    XRAM[18378] = 8'b0;
    XRAM[18379] = 8'b0;
    XRAM[18380] = 8'b0;
    XRAM[18381] = 8'b0;
    XRAM[18382] = 8'b0;
    XRAM[18383] = 8'b0;
    XRAM[18384] = 8'b0;
    XRAM[18385] = 8'b0;
    XRAM[18386] = 8'b0;
    XRAM[18387] = 8'b0;
    XRAM[18388] = 8'b0;
    XRAM[18389] = 8'b0;
    XRAM[18390] = 8'b0;
    XRAM[18391] = 8'b0;
    XRAM[18392] = 8'b0;
    XRAM[18393] = 8'b0;
    XRAM[18394] = 8'b0;
    XRAM[18395] = 8'b0;
    XRAM[18396] = 8'b0;
    XRAM[18397] = 8'b0;
    XRAM[18398] = 8'b0;
    XRAM[18399] = 8'b0;
    XRAM[18400] = 8'b0;
    XRAM[18401] = 8'b0;
    XRAM[18402] = 8'b0;
    XRAM[18403] = 8'b0;
    XRAM[18404] = 8'b0;
    XRAM[18405] = 8'b0;
    XRAM[18406] = 8'b0;
    XRAM[18407] = 8'b0;
    XRAM[18408] = 8'b0;
    XRAM[18409] = 8'b0;
    XRAM[18410] = 8'b0;
    XRAM[18411] = 8'b0;
    XRAM[18412] = 8'b0;
    XRAM[18413] = 8'b0;
    XRAM[18414] = 8'b0;
    XRAM[18415] = 8'b0;
    XRAM[18416] = 8'b0;
    XRAM[18417] = 8'b0;
    XRAM[18418] = 8'b0;
    XRAM[18419] = 8'b0;
    XRAM[18420] = 8'b0;
    XRAM[18421] = 8'b0;
    XRAM[18422] = 8'b0;
    XRAM[18423] = 8'b0;
    XRAM[18424] = 8'b0;
    XRAM[18425] = 8'b0;
    XRAM[18426] = 8'b0;
    XRAM[18427] = 8'b0;
    XRAM[18428] = 8'b0;
    XRAM[18429] = 8'b0;
    XRAM[18430] = 8'b0;
    XRAM[18431] = 8'b0;
    XRAM[18432] = 8'b0;
    XRAM[18433] = 8'b0;
    XRAM[18434] = 8'b0;
    XRAM[18435] = 8'b0;
    XRAM[18436] = 8'b0;
    XRAM[18437] = 8'b0;
    XRAM[18438] = 8'b0;
    XRAM[18439] = 8'b0;
    XRAM[18440] = 8'b0;
    XRAM[18441] = 8'b0;
    XRAM[18442] = 8'b0;
    XRAM[18443] = 8'b0;
    XRAM[18444] = 8'b0;
    XRAM[18445] = 8'b0;
    XRAM[18446] = 8'b0;
    XRAM[18447] = 8'b0;
    XRAM[18448] = 8'b0;
    XRAM[18449] = 8'b0;
    XRAM[18450] = 8'b0;
    XRAM[18451] = 8'b0;
    XRAM[18452] = 8'b0;
    XRAM[18453] = 8'b0;
    XRAM[18454] = 8'b0;
    XRAM[18455] = 8'b0;
    XRAM[18456] = 8'b0;
    XRAM[18457] = 8'b0;
    XRAM[18458] = 8'b0;
    XRAM[18459] = 8'b0;
    XRAM[18460] = 8'b0;
    XRAM[18461] = 8'b0;
    XRAM[18462] = 8'b0;
    XRAM[18463] = 8'b0;
    XRAM[18464] = 8'b0;
    XRAM[18465] = 8'b0;
    XRAM[18466] = 8'b0;
    XRAM[18467] = 8'b0;
    XRAM[18468] = 8'b0;
    XRAM[18469] = 8'b0;
    XRAM[18470] = 8'b0;
    XRAM[18471] = 8'b0;
    XRAM[18472] = 8'b0;
    XRAM[18473] = 8'b0;
    XRAM[18474] = 8'b0;
    XRAM[18475] = 8'b0;
    XRAM[18476] = 8'b0;
    XRAM[18477] = 8'b0;
    XRAM[18478] = 8'b0;
    XRAM[18479] = 8'b0;
    XRAM[18480] = 8'b0;
    XRAM[18481] = 8'b0;
    XRAM[18482] = 8'b0;
    XRAM[18483] = 8'b0;
    XRAM[18484] = 8'b0;
    XRAM[18485] = 8'b0;
    XRAM[18486] = 8'b0;
    XRAM[18487] = 8'b0;
    XRAM[18488] = 8'b0;
    XRAM[18489] = 8'b0;
    XRAM[18490] = 8'b0;
    XRAM[18491] = 8'b0;
    XRAM[18492] = 8'b0;
    XRAM[18493] = 8'b0;
    XRAM[18494] = 8'b0;
    XRAM[18495] = 8'b0;
    XRAM[18496] = 8'b0;
    XRAM[18497] = 8'b0;
    XRAM[18498] = 8'b0;
    XRAM[18499] = 8'b0;
    XRAM[18500] = 8'b0;
    XRAM[18501] = 8'b0;
    XRAM[18502] = 8'b0;
    XRAM[18503] = 8'b0;
    XRAM[18504] = 8'b0;
    XRAM[18505] = 8'b0;
    XRAM[18506] = 8'b0;
    XRAM[18507] = 8'b0;
    XRAM[18508] = 8'b0;
    XRAM[18509] = 8'b0;
    XRAM[18510] = 8'b0;
    XRAM[18511] = 8'b0;
    XRAM[18512] = 8'b0;
    XRAM[18513] = 8'b0;
    XRAM[18514] = 8'b0;
    XRAM[18515] = 8'b0;
    XRAM[18516] = 8'b0;
    XRAM[18517] = 8'b0;
    XRAM[18518] = 8'b0;
    XRAM[18519] = 8'b0;
    XRAM[18520] = 8'b0;
    XRAM[18521] = 8'b0;
    XRAM[18522] = 8'b0;
    XRAM[18523] = 8'b0;
    XRAM[18524] = 8'b0;
    XRAM[18525] = 8'b0;
    XRAM[18526] = 8'b0;
    XRAM[18527] = 8'b0;
    XRAM[18528] = 8'b0;
    XRAM[18529] = 8'b0;
    XRAM[18530] = 8'b0;
    XRAM[18531] = 8'b0;
    XRAM[18532] = 8'b0;
    XRAM[18533] = 8'b0;
    XRAM[18534] = 8'b0;
    XRAM[18535] = 8'b0;
    XRAM[18536] = 8'b0;
    XRAM[18537] = 8'b0;
    XRAM[18538] = 8'b0;
    XRAM[18539] = 8'b0;
    XRAM[18540] = 8'b0;
    XRAM[18541] = 8'b0;
    XRAM[18542] = 8'b0;
    XRAM[18543] = 8'b0;
    XRAM[18544] = 8'b0;
    XRAM[18545] = 8'b0;
    XRAM[18546] = 8'b0;
    XRAM[18547] = 8'b0;
    XRAM[18548] = 8'b0;
    XRAM[18549] = 8'b0;
    XRAM[18550] = 8'b0;
    XRAM[18551] = 8'b0;
    XRAM[18552] = 8'b0;
    XRAM[18553] = 8'b0;
    XRAM[18554] = 8'b0;
    XRAM[18555] = 8'b0;
    XRAM[18556] = 8'b0;
    XRAM[18557] = 8'b0;
    XRAM[18558] = 8'b0;
    XRAM[18559] = 8'b0;
    XRAM[18560] = 8'b0;
    XRAM[18561] = 8'b0;
    XRAM[18562] = 8'b0;
    XRAM[18563] = 8'b0;
    XRAM[18564] = 8'b0;
    XRAM[18565] = 8'b0;
    XRAM[18566] = 8'b0;
    XRAM[18567] = 8'b0;
    XRAM[18568] = 8'b0;
    XRAM[18569] = 8'b0;
    XRAM[18570] = 8'b0;
    XRAM[18571] = 8'b0;
    XRAM[18572] = 8'b0;
    XRAM[18573] = 8'b0;
    XRAM[18574] = 8'b0;
    XRAM[18575] = 8'b0;
    XRAM[18576] = 8'b0;
    XRAM[18577] = 8'b0;
    XRAM[18578] = 8'b0;
    XRAM[18579] = 8'b0;
    XRAM[18580] = 8'b0;
    XRAM[18581] = 8'b0;
    XRAM[18582] = 8'b0;
    XRAM[18583] = 8'b0;
    XRAM[18584] = 8'b0;
    XRAM[18585] = 8'b0;
    XRAM[18586] = 8'b0;
    XRAM[18587] = 8'b0;
    XRAM[18588] = 8'b0;
    XRAM[18589] = 8'b0;
    XRAM[18590] = 8'b0;
    XRAM[18591] = 8'b0;
    XRAM[18592] = 8'b0;
    XRAM[18593] = 8'b0;
    XRAM[18594] = 8'b0;
    XRAM[18595] = 8'b0;
    XRAM[18596] = 8'b0;
    XRAM[18597] = 8'b0;
    XRAM[18598] = 8'b0;
    XRAM[18599] = 8'b0;
    XRAM[18600] = 8'b0;
    XRAM[18601] = 8'b0;
    XRAM[18602] = 8'b0;
    XRAM[18603] = 8'b0;
    XRAM[18604] = 8'b0;
    XRAM[18605] = 8'b0;
    XRAM[18606] = 8'b0;
    XRAM[18607] = 8'b0;
    XRAM[18608] = 8'b0;
    XRAM[18609] = 8'b0;
    XRAM[18610] = 8'b0;
    XRAM[18611] = 8'b0;
    XRAM[18612] = 8'b0;
    XRAM[18613] = 8'b0;
    XRAM[18614] = 8'b0;
    XRAM[18615] = 8'b0;
    XRAM[18616] = 8'b0;
    XRAM[18617] = 8'b0;
    XRAM[18618] = 8'b0;
    XRAM[18619] = 8'b0;
    XRAM[18620] = 8'b0;
    XRAM[18621] = 8'b0;
    XRAM[18622] = 8'b0;
    XRAM[18623] = 8'b0;
    XRAM[18624] = 8'b0;
    XRAM[18625] = 8'b0;
    XRAM[18626] = 8'b0;
    XRAM[18627] = 8'b0;
    XRAM[18628] = 8'b0;
    XRAM[18629] = 8'b0;
    XRAM[18630] = 8'b0;
    XRAM[18631] = 8'b0;
    XRAM[18632] = 8'b0;
    XRAM[18633] = 8'b0;
    XRAM[18634] = 8'b0;
    XRAM[18635] = 8'b0;
    XRAM[18636] = 8'b0;
    XRAM[18637] = 8'b0;
    XRAM[18638] = 8'b0;
    XRAM[18639] = 8'b0;
    XRAM[18640] = 8'b0;
    XRAM[18641] = 8'b0;
    XRAM[18642] = 8'b0;
    XRAM[18643] = 8'b0;
    XRAM[18644] = 8'b0;
    XRAM[18645] = 8'b0;
    XRAM[18646] = 8'b0;
    XRAM[18647] = 8'b0;
    XRAM[18648] = 8'b0;
    XRAM[18649] = 8'b0;
    XRAM[18650] = 8'b0;
    XRAM[18651] = 8'b0;
    XRAM[18652] = 8'b0;
    XRAM[18653] = 8'b0;
    XRAM[18654] = 8'b0;
    XRAM[18655] = 8'b0;
    XRAM[18656] = 8'b0;
    XRAM[18657] = 8'b0;
    XRAM[18658] = 8'b0;
    XRAM[18659] = 8'b0;
    XRAM[18660] = 8'b0;
    XRAM[18661] = 8'b0;
    XRAM[18662] = 8'b0;
    XRAM[18663] = 8'b0;
    XRAM[18664] = 8'b0;
    XRAM[18665] = 8'b0;
    XRAM[18666] = 8'b0;
    XRAM[18667] = 8'b0;
    XRAM[18668] = 8'b0;
    XRAM[18669] = 8'b0;
    XRAM[18670] = 8'b0;
    XRAM[18671] = 8'b0;
    XRAM[18672] = 8'b0;
    XRAM[18673] = 8'b0;
    XRAM[18674] = 8'b0;
    XRAM[18675] = 8'b0;
    XRAM[18676] = 8'b0;
    XRAM[18677] = 8'b0;
    XRAM[18678] = 8'b0;
    XRAM[18679] = 8'b0;
    XRAM[18680] = 8'b0;
    XRAM[18681] = 8'b0;
    XRAM[18682] = 8'b0;
    XRAM[18683] = 8'b0;
    XRAM[18684] = 8'b0;
    XRAM[18685] = 8'b0;
    XRAM[18686] = 8'b0;
    XRAM[18687] = 8'b0;
    XRAM[18688] = 8'b0;
    XRAM[18689] = 8'b0;
    XRAM[18690] = 8'b0;
    XRAM[18691] = 8'b0;
    XRAM[18692] = 8'b0;
    XRAM[18693] = 8'b0;
    XRAM[18694] = 8'b0;
    XRAM[18695] = 8'b0;
    XRAM[18696] = 8'b0;
    XRAM[18697] = 8'b0;
    XRAM[18698] = 8'b0;
    XRAM[18699] = 8'b0;
    XRAM[18700] = 8'b0;
    XRAM[18701] = 8'b0;
    XRAM[18702] = 8'b0;
    XRAM[18703] = 8'b0;
    XRAM[18704] = 8'b0;
    XRAM[18705] = 8'b0;
    XRAM[18706] = 8'b0;
    XRAM[18707] = 8'b0;
    XRAM[18708] = 8'b0;
    XRAM[18709] = 8'b0;
    XRAM[18710] = 8'b0;
    XRAM[18711] = 8'b0;
    XRAM[18712] = 8'b0;
    XRAM[18713] = 8'b0;
    XRAM[18714] = 8'b0;
    XRAM[18715] = 8'b0;
    XRAM[18716] = 8'b0;
    XRAM[18717] = 8'b0;
    XRAM[18718] = 8'b0;
    XRAM[18719] = 8'b0;
    XRAM[18720] = 8'b0;
    XRAM[18721] = 8'b0;
    XRAM[18722] = 8'b0;
    XRAM[18723] = 8'b0;
    XRAM[18724] = 8'b0;
    XRAM[18725] = 8'b0;
    XRAM[18726] = 8'b0;
    XRAM[18727] = 8'b0;
    XRAM[18728] = 8'b0;
    XRAM[18729] = 8'b0;
    XRAM[18730] = 8'b0;
    XRAM[18731] = 8'b0;
    XRAM[18732] = 8'b0;
    XRAM[18733] = 8'b0;
    XRAM[18734] = 8'b0;
    XRAM[18735] = 8'b0;
    XRAM[18736] = 8'b0;
    XRAM[18737] = 8'b0;
    XRAM[18738] = 8'b0;
    XRAM[18739] = 8'b0;
    XRAM[18740] = 8'b0;
    XRAM[18741] = 8'b0;
    XRAM[18742] = 8'b0;
    XRAM[18743] = 8'b0;
    XRAM[18744] = 8'b0;
    XRAM[18745] = 8'b0;
    XRAM[18746] = 8'b0;
    XRAM[18747] = 8'b0;
    XRAM[18748] = 8'b0;
    XRAM[18749] = 8'b0;
    XRAM[18750] = 8'b0;
    XRAM[18751] = 8'b0;
    XRAM[18752] = 8'b0;
    XRAM[18753] = 8'b0;
    XRAM[18754] = 8'b0;
    XRAM[18755] = 8'b0;
    XRAM[18756] = 8'b0;
    XRAM[18757] = 8'b0;
    XRAM[18758] = 8'b0;
    XRAM[18759] = 8'b0;
    XRAM[18760] = 8'b0;
    XRAM[18761] = 8'b0;
    XRAM[18762] = 8'b0;
    XRAM[18763] = 8'b0;
    XRAM[18764] = 8'b0;
    XRAM[18765] = 8'b0;
    XRAM[18766] = 8'b0;
    XRAM[18767] = 8'b0;
    XRAM[18768] = 8'b0;
    XRAM[18769] = 8'b0;
    XRAM[18770] = 8'b0;
    XRAM[18771] = 8'b0;
    XRAM[18772] = 8'b0;
    XRAM[18773] = 8'b0;
    XRAM[18774] = 8'b0;
    XRAM[18775] = 8'b0;
    XRAM[18776] = 8'b0;
    XRAM[18777] = 8'b0;
    XRAM[18778] = 8'b0;
    XRAM[18779] = 8'b0;
    XRAM[18780] = 8'b0;
    XRAM[18781] = 8'b0;
    XRAM[18782] = 8'b0;
    XRAM[18783] = 8'b0;
    XRAM[18784] = 8'b0;
    XRAM[18785] = 8'b0;
    XRAM[18786] = 8'b0;
    XRAM[18787] = 8'b0;
    XRAM[18788] = 8'b0;
    XRAM[18789] = 8'b0;
    XRAM[18790] = 8'b0;
    XRAM[18791] = 8'b0;
    XRAM[18792] = 8'b0;
    XRAM[18793] = 8'b0;
    XRAM[18794] = 8'b0;
    XRAM[18795] = 8'b0;
    XRAM[18796] = 8'b0;
    XRAM[18797] = 8'b0;
    XRAM[18798] = 8'b0;
    XRAM[18799] = 8'b0;
    XRAM[18800] = 8'b0;
    XRAM[18801] = 8'b0;
    XRAM[18802] = 8'b0;
    XRAM[18803] = 8'b0;
    XRAM[18804] = 8'b0;
    XRAM[18805] = 8'b0;
    XRAM[18806] = 8'b0;
    XRAM[18807] = 8'b0;
    XRAM[18808] = 8'b0;
    XRAM[18809] = 8'b0;
    XRAM[18810] = 8'b0;
    XRAM[18811] = 8'b0;
    XRAM[18812] = 8'b0;
    XRAM[18813] = 8'b0;
    XRAM[18814] = 8'b0;
    XRAM[18815] = 8'b0;
    XRAM[18816] = 8'b0;
    XRAM[18817] = 8'b0;
    XRAM[18818] = 8'b0;
    XRAM[18819] = 8'b0;
    XRAM[18820] = 8'b0;
    XRAM[18821] = 8'b0;
    XRAM[18822] = 8'b0;
    XRAM[18823] = 8'b0;
    XRAM[18824] = 8'b0;
    XRAM[18825] = 8'b0;
    XRAM[18826] = 8'b0;
    XRAM[18827] = 8'b0;
    XRAM[18828] = 8'b0;
    XRAM[18829] = 8'b0;
    XRAM[18830] = 8'b0;
    XRAM[18831] = 8'b0;
    XRAM[18832] = 8'b0;
    XRAM[18833] = 8'b0;
    XRAM[18834] = 8'b0;
    XRAM[18835] = 8'b0;
    XRAM[18836] = 8'b0;
    XRAM[18837] = 8'b0;
    XRAM[18838] = 8'b0;
    XRAM[18839] = 8'b0;
    XRAM[18840] = 8'b0;
    XRAM[18841] = 8'b0;
    XRAM[18842] = 8'b0;
    XRAM[18843] = 8'b0;
    XRAM[18844] = 8'b0;
    XRAM[18845] = 8'b0;
    XRAM[18846] = 8'b0;
    XRAM[18847] = 8'b0;
    XRAM[18848] = 8'b0;
    XRAM[18849] = 8'b0;
    XRAM[18850] = 8'b0;
    XRAM[18851] = 8'b0;
    XRAM[18852] = 8'b0;
    XRAM[18853] = 8'b0;
    XRAM[18854] = 8'b0;
    XRAM[18855] = 8'b0;
    XRAM[18856] = 8'b0;
    XRAM[18857] = 8'b0;
    XRAM[18858] = 8'b0;
    XRAM[18859] = 8'b0;
    XRAM[18860] = 8'b0;
    XRAM[18861] = 8'b0;
    XRAM[18862] = 8'b0;
    XRAM[18863] = 8'b0;
    XRAM[18864] = 8'b0;
    XRAM[18865] = 8'b0;
    XRAM[18866] = 8'b0;
    XRAM[18867] = 8'b0;
    XRAM[18868] = 8'b0;
    XRAM[18869] = 8'b0;
    XRAM[18870] = 8'b0;
    XRAM[18871] = 8'b0;
    XRAM[18872] = 8'b0;
    XRAM[18873] = 8'b0;
    XRAM[18874] = 8'b0;
    XRAM[18875] = 8'b0;
    XRAM[18876] = 8'b0;
    XRAM[18877] = 8'b0;
    XRAM[18878] = 8'b0;
    XRAM[18879] = 8'b0;
    XRAM[18880] = 8'b0;
    XRAM[18881] = 8'b0;
    XRAM[18882] = 8'b0;
    XRAM[18883] = 8'b0;
    XRAM[18884] = 8'b0;
    XRAM[18885] = 8'b0;
    XRAM[18886] = 8'b0;
    XRAM[18887] = 8'b0;
    XRAM[18888] = 8'b0;
    XRAM[18889] = 8'b0;
    XRAM[18890] = 8'b0;
    XRAM[18891] = 8'b0;
    XRAM[18892] = 8'b0;
    XRAM[18893] = 8'b0;
    XRAM[18894] = 8'b0;
    XRAM[18895] = 8'b0;
    XRAM[18896] = 8'b0;
    XRAM[18897] = 8'b0;
    XRAM[18898] = 8'b0;
    XRAM[18899] = 8'b0;
    XRAM[18900] = 8'b0;
    XRAM[18901] = 8'b0;
    XRAM[18902] = 8'b0;
    XRAM[18903] = 8'b0;
    XRAM[18904] = 8'b0;
    XRAM[18905] = 8'b0;
    XRAM[18906] = 8'b0;
    XRAM[18907] = 8'b0;
    XRAM[18908] = 8'b0;
    XRAM[18909] = 8'b0;
    XRAM[18910] = 8'b0;
    XRAM[18911] = 8'b0;
    XRAM[18912] = 8'b0;
    XRAM[18913] = 8'b0;
    XRAM[18914] = 8'b0;
    XRAM[18915] = 8'b0;
    XRAM[18916] = 8'b0;
    XRAM[18917] = 8'b0;
    XRAM[18918] = 8'b0;
    XRAM[18919] = 8'b0;
    XRAM[18920] = 8'b0;
    XRAM[18921] = 8'b0;
    XRAM[18922] = 8'b0;
    XRAM[18923] = 8'b0;
    XRAM[18924] = 8'b0;
    XRAM[18925] = 8'b0;
    XRAM[18926] = 8'b0;
    XRAM[18927] = 8'b0;
    XRAM[18928] = 8'b0;
    XRAM[18929] = 8'b0;
    XRAM[18930] = 8'b0;
    XRAM[18931] = 8'b0;
    XRAM[18932] = 8'b0;
    XRAM[18933] = 8'b0;
    XRAM[18934] = 8'b0;
    XRAM[18935] = 8'b0;
    XRAM[18936] = 8'b0;
    XRAM[18937] = 8'b0;
    XRAM[18938] = 8'b0;
    XRAM[18939] = 8'b0;
    XRAM[18940] = 8'b0;
    XRAM[18941] = 8'b0;
    XRAM[18942] = 8'b0;
    XRAM[18943] = 8'b0;
    XRAM[18944] = 8'b0;
    XRAM[18945] = 8'b0;
    XRAM[18946] = 8'b0;
    XRAM[18947] = 8'b0;
    XRAM[18948] = 8'b0;
    XRAM[18949] = 8'b0;
    XRAM[18950] = 8'b0;
    XRAM[18951] = 8'b0;
    XRAM[18952] = 8'b0;
    XRAM[18953] = 8'b0;
    XRAM[18954] = 8'b0;
    XRAM[18955] = 8'b0;
    XRAM[18956] = 8'b0;
    XRAM[18957] = 8'b0;
    XRAM[18958] = 8'b0;
    XRAM[18959] = 8'b0;
    XRAM[18960] = 8'b0;
    XRAM[18961] = 8'b0;
    XRAM[18962] = 8'b0;
    XRAM[18963] = 8'b0;
    XRAM[18964] = 8'b0;
    XRAM[18965] = 8'b0;
    XRAM[18966] = 8'b0;
    XRAM[18967] = 8'b0;
    XRAM[18968] = 8'b0;
    XRAM[18969] = 8'b0;
    XRAM[18970] = 8'b0;
    XRAM[18971] = 8'b0;
    XRAM[18972] = 8'b0;
    XRAM[18973] = 8'b0;
    XRAM[18974] = 8'b0;
    XRAM[18975] = 8'b0;
    XRAM[18976] = 8'b0;
    XRAM[18977] = 8'b0;
    XRAM[18978] = 8'b0;
    XRAM[18979] = 8'b0;
    XRAM[18980] = 8'b0;
    XRAM[18981] = 8'b0;
    XRAM[18982] = 8'b0;
    XRAM[18983] = 8'b0;
    XRAM[18984] = 8'b0;
    XRAM[18985] = 8'b0;
    XRAM[18986] = 8'b0;
    XRAM[18987] = 8'b0;
    XRAM[18988] = 8'b0;
    XRAM[18989] = 8'b0;
    XRAM[18990] = 8'b0;
    XRAM[18991] = 8'b0;
    XRAM[18992] = 8'b0;
    XRAM[18993] = 8'b0;
    XRAM[18994] = 8'b0;
    XRAM[18995] = 8'b0;
    XRAM[18996] = 8'b0;
    XRAM[18997] = 8'b0;
    XRAM[18998] = 8'b0;
    XRAM[18999] = 8'b0;
    XRAM[19000] = 8'b0;
    XRAM[19001] = 8'b0;
    XRAM[19002] = 8'b0;
    XRAM[19003] = 8'b0;
    XRAM[19004] = 8'b0;
    XRAM[19005] = 8'b0;
    XRAM[19006] = 8'b0;
    XRAM[19007] = 8'b0;
    XRAM[19008] = 8'b0;
    XRAM[19009] = 8'b0;
    XRAM[19010] = 8'b0;
    XRAM[19011] = 8'b0;
    XRAM[19012] = 8'b0;
    XRAM[19013] = 8'b0;
    XRAM[19014] = 8'b0;
    XRAM[19015] = 8'b0;
    XRAM[19016] = 8'b0;
    XRAM[19017] = 8'b0;
    XRAM[19018] = 8'b0;
    XRAM[19019] = 8'b0;
    XRAM[19020] = 8'b0;
    XRAM[19021] = 8'b0;
    XRAM[19022] = 8'b0;
    XRAM[19023] = 8'b0;
    XRAM[19024] = 8'b0;
    XRAM[19025] = 8'b0;
    XRAM[19026] = 8'b0;
    XRAM[19027] = 8'b0;
    XRAM[19028] = 8'b0;
    XRAM[19029] = 8'b0;
    XRAM[19030] = 8'b0;
    XRAM[19031] = 8'b0;
    XRAM[19032] = 8'b0;
    XRAM[19033] = 8'b0;
    XRAM[19034] = 8'b0;
    XRAM[19035] = 8'b0;
    XRAM[19036] = 8'b0;
    XRAM[19037] = 8'b0;
    XRAM[19038] = 8'b0;
    XRAM[19039] = 8'b0;
    XRAM[19040] = 8'b0;
    XRAM[19041] = 8'b0;
    XRAM[19042] = 8'b0;
    XRAM[19043] = 8'b0;
    XRAM[19044] = 8'b0;
    XRAM[19045] = 8'b0;
    XRAM[19046] = 8'b0;
    XRAM[19047] = 8'b0;
    XRAM[19048] = 8'b0;
    XRAM[19049] = 8'b0;
    XRAM[19050] = 8'b0;
    XRAM[19051] = 8'b0;
    XRAM[19052] = 8'b0;
    XRAM[19053] = 8'b0;
    XRAM[19054] = 8'b0;
    XRAM[19055] = 8'b0;
    XRAM[19056] = 8'b0;
    XRAM[19057] = 8'b0;
    XRAM[19058] = 8'b0;
    XRAM[19059] = 8'b0;
    XRAM[19060] = 8'b0;
    XRAM[19061] = 8'b0;
    XRAM[19062] = 8'b0;
    XRAM[19063] = 8'b0;
    XRAM[19064] = 8'b0;
    XRAM[19065] = 8'b0;
    XRAM[19066] = 8'b0;
    XRAM[19067] = 8'b0;
    XRAM[19068] = 8'b0;
    XRAM[19069] = 8'b0;
    XRAM[19070] = 8'b0;
    XRAM[19071] = 8'b0;
    XRAM[19072] = 8'b0;
    XRAM[19073] = 8'b0;
    XRAM[19074] = 8'b0;
    XRAM[19075] = 8'b0;
    XRAM[19076] = 8'b0;
    XRAM[19077] = 8'b0;
    XRAM[19078] = 8'b0;
    XRAM[19079] = 8'b0;
    XRAM[19080] = 8'b0;
    XRAM[19081] = 8'b0;
    XRAM[19082] = 8'b0;
    XRAM[19083] = 8'b0;
    XRAM[19084] = 8'b0;
    XRAM[19085] = 8'b0;
    XRAM[19086] = 8'b0;
    XRAM[19087] = 8'b0;
    XRAM[19088] = 8'b0;
    XRAM[19089] = 8'b0;
    XRAM[19090] = 8'b0;
    XRAM[19091] = 8'b0;
    XRAM[19092] = 8'b0;
    XRAM[19093] = 8'b0;
    XRAM[19094] = 8'b0;
    XRAM[19095] = 8'b0;
    XRAM[19096] = 8'b0;
    XRAM[19097] = 8'b0;
    XRAM[19098] = 8'b0;
    XRAM[19099] = 8'b0;
    XRAM[19100] = 8'b0;
    XRAM[19101] = 8'b0;
    XRAM[19102] = 8'b0;
    XRAM[19103] = 8'b0;
    XRAM[19104] = 8'b0;
    XRAM[19105] = 8'b0;
    XRAM[19106] = 8'b0;
    XRAM[19107] = 8'b0;
    XRAM[19108] = 8'b0;
    XRAM[19109] = 8'b0;
    XRAM[19110] = 8'b0;
    XRAM[19111] = 8'b0;
    XRAM[19112] = 8'b0;
    XRAM[19113] = 8'b0;
    XRAM[19114] = 8'b0;
    XRAM[19115] = 8'b0;
    XRAM[19116] = 8'b0;
    XRAM[19117] = 8'b0;
    XRAM[19118] = 8'b0;
    XRAM[19119] = 8'b0;
    XRAM[19120] = 8'b0;
    XRAM[19121] = 8'b0;
    XRAM[19122] = 8'b0;
    XRAM[19123] = 8'b0;
    XRAM[19124] = 8'b0;
    XRAM[19125] = 8'b0;
    XRAM[19126] = 8'b0;
    XRAM[19127] = 8'b0;
    XRAM[19128] = 8'b0;
    XRAM[19129] = 8'b0;
    XRAM[19130] = 8'b0;
    XRAM[19131] = 8'b0;
    XRAM[19132] = 8'b0;
    XRAM[19133] = 8'b0;
    XRAM[19134] = 8'b0;
    XRAM[19135] = 8'b0;
    XRAM[19136] = 8'b0;
    XRAM[19137] = 8'b0;
    XRAM[19138] = 8'b0;
    XRAM[19139] = 8'b0;
    XRAM[19140] = 8'b0;
    XRAM[19141] = 8'b0;
    XRAM[19142] = 8'b0;
    XRAM[19143] = 8'b0;
    XRAM[19144] = 8'b0;
    XRAM[19145] = 8'b0;
    XRAM[19146] = 8'b0;
    XRAM[19147] = 8'b0;
    XRAM[19148] = 8'b0;
    XRAM[19149] = 8'b0;
    XRAM[19150] = 8'b0;
    XRAM[19151] = 8'b0;
    XRAM[19152] = 8'b0;
    XRAM[19153] = 8'b0;
    XRAM[19154] = 8'b0;
    XRAM[19155] = 8'b0;
    XRAM[19156] = 8'b0;
    XRAM[19157] = 8'b0;
    XRAM[19158] = 8'b0;
    XRAM[19159] = 8'b0;
    XRAM[19160] = 8'b0;
    XRAM[19161] = 8'b0;
    XRAM[19162] = 8'b0;
    XRAM[19163] = 8'b0;
    XRAM[19164] = 8'b0;
    XRAM[19165] = 8'b0;
    XRAM[19166] = 8'b0;
    XRAM[19167] = 8'b0;
    XRAM[19168] = 8'b0;
    XRAM[19169] = 8'b0;
    XRAM[19170] = 8'b0;
    XRAM[19171] = 8'b0;
    XRAM[19172] = 8'b0;
    XRAM[19173] = 8'b0;
    XRAM[19174] = 8'b0;
    XRAM[19175] = 8'b0;
    XRAM[19176] = 8'b0;
    XRAM[19177] = 8'b0;
    XRAM[19178] = 8'b0;
    XRAM[19179] = 8'b0;
    XRAM[19180] = 8'b0;
    XRAM[19181] = 8'b0;
    XRAM[19182] = 8'b0;
    XRAM[19183] = 8'b0;
    XRAM[19184] = 8'b0;
    XRAM[19185] = 8'b0;
    XRAM[19186] = 8'b0;
    XRAM[19187] = 8'b0;
    XRAM[19188] = 8'b0;
    XRAM[19189] = 8'b0;
    XRAM[19190] = 8'b0;
    XRAM[19191] = 8'b0;
    XRAM[19192] = 8'b0;
    XRAM[19193] = 8'b0;
    XRAM[19194] = 8'b0;
    XRAM[19195] = 8'b0;
    XRAM[19196] = 8'b0;
    XRAM[19197] = 8'b0;
    XRAM[19198] = 8'b0;
    XRAM[19199] = 8'b0;
    XRAM[19200] = 8'b0;
    XRAM[19201] = 8'b0;
    XRAM[19202] = 8'b0;
    XRAM[19203] = 8'b0;
    XRAM[19204] = 8'b0;
    XRAM[19205] = 8'b0;
    XRAM[19206] = 8'b0;
    XRAM[19207] = 8'b0;
    XRAM[19208] = 8'b0;
    XRAM[19209] = 8'b0;
    XRAM[19210] = 8'b0;
    XRAM[19211] = 8'b0;
    XRAM[19212] = 8'b0;
    XRAM[19213] = 8'b0;
    XRAM[19214] = 8'b0;
    XRAM[19215] = 8'b0;
    XRAM[19216] = 8'b0;
    XRAM[19217] = 8'b0;
    XRAM[19218] = 8'b0;
    XRAM[19219] = 8'b0;
    XRAM[19220] = 8'b0;
    XRAM[19221] = 8'b0;
    XRAM[19222] = 8'b0;
    XRAM[19223] = 8'b0;
    XRAM[19224] = 8'b0;
    XRAM[19225] = 8'b0;
    XRAM[19226] = 8'b0;
    XRAM[19227] = 8'b0;
    XRAM[19228] = 8'b0;
    XRAM[19229] = 8'b0;
    XRAM[19230] = 8'b0;
    XRAM[19231] = 8'b0;
    XRAM[19232] = 8'b0;
    XRAM[19233] = 8'b0;
    XRAM[19234] = 8'b0;
    XRAM[19235] = 8'b0;
    XRAM[19236] = 8'b0;
    XRAM[19237] = 8'b0;
    XRAM[19238] = 8'b0;
    XRAM[19239] = 8'b0;
    XRAM[19240] = 8'b0;
    XRAM[19241] = 8'b0;
    XRAM[19242] = 8'b0;
    XRAM[19243] = 8'b0;
    XRAM[19244] = 8'b0;
    XRAM[19245] = 8'b0;
    XRAM[19246] = 8'b0;
    XRAM[19247] = 8'b0;
    XRAM[19248] = 8'b0;
    XRAM[19249] = 8'b0;
    XRAM[19250] = 8'b0;
    XRAM[19251] = 8'b0;
    XRAM[19252] = 8'b0;
    XRAM[19253] = 8'b0;
    XRAM[19254] = 8'b0;
    XRAM[19255] = 8'b0;
    XRAM[19256] = 8'b0;
    XRAM[19257] = 8'b0;
    XRAM[19258] = 8'b0;
    XRAM[19259] = 8'b0;
    XRAM[19260] = 8'b0;
    XRAM[19261] = 8'b0;
    XRAM[19262] = 8'b0;
    XRAM[19263] = 8'b0;
    XRAM[19264] = 8'b0;
    XRAM[19265] = 8'b0;
    XRAM[19266] = 8'b0;
    XRAM[19267] = 8'b0;
    XRAM[19268] = 8'b0;
    XRAM[19269] = 8'b0;
    XRAM[19270] = 8'b0;
    XRAM[19271] = 8'b0;
    XRAM[19272] = 8'b0;
    XRAM[19273] = 8'b0;
    XRAM[19274] = 8'b0;
    XRAM[19275] = 8'b0;
    XRAM[19276] = 8'b0;
    XRAM[19277] = 8'b0;
    XRAM[19278] = 8'b0;
    XRAM[19279] = 8'b0;
    XRAM[19280] = 8'b0;
    XRAM[19281] = 8'b0;
    XRAM[19282] = 8'b0;
    XRAM[19283] = 8'b0;
    XRAM[19284] = 8'b0;
    XRAM[19285] = 8'b0;
    XRAM[19286] = 8'b0;
    XRAM[19287] = 8'b0;
    XRAM[19288] = 8'b0;
    XRAM[19289] = 8'b0;
    XRAM[19290] = 8'b0;
    XRAM[19291] = 8'b0;
    XRAM[19292] = 8'b0;
    XRAM[19293] = 8'b0;
    XRAM[19294] = 8'b0;
    XRAM[19295] = 8'b0;
    XRAM[19296] = 8'b0;
    XRAM[19297] = 8'b0;
    XRAM[19298] = 8'b0;
    XRAM[19299] = 8'b0;
    XRAM[19300] = 8'b0;
    XRAM[19301] = 8'b0;
    XRAM[19302] = 8'b0;
    XRAM[19303] = 8'b0;
    XRAM[19304] = 8'b0;
    XRAM[19305] = 8'b0;
    XRAM[19306] = 8'b0;
    XRAM[19307] = 8'b0;
    XRAM[19308] = 8'b0;
    XRAM[19309] = 8'b0;
    XRAM[19310] = 8'b0;
    XRAM[19311] = 8'b0;
    XRAM[19312] = 8'b0;
    XRAM[19313] = 8'b0;
    XRAM[19314] = 8'b0;
    XRAM[19315] = 8'b0;
    XRAM[19316] = 8'b0;
    XRAM[19317] = 8'b0;
    XRAM[19318] = 8'b0;
    XRAM[19319] = 8'b0;
    XRAM[19320] = 8'b0;
    XRAM[19321] = 8'b0;
    XRAM[19322] = 8'b0;
    XRAM[19323] = 8'b0;
    XRAM[19324] = 8'b0;
    XRAM[19325] = 8'b0;
    XRAM[19326] = 8'b0;
    XRAM[19327] = 8'b0;
    XRAM[19328] = 8'b0;
    XRAM[19329] = 8'b0;
    XRAM[19330] = 8'b0;
    XRAM[19331] = 8'b0;
    XRAM[19332] = 8'b0;
    XRAM[19333] = 8'b0;
    XRAM[19334] = 8'b0;
    XRAM[19335] = 8'b0;
    XRAM[19336] = 8'b0;
    XRAM[19337] = 8'b0;
    XRAM[19338] = 8'b0;
    XRAM[19339] = 8'b0;
    XRAM[19340] = 8'b0;
    XRAM[19341] = 8'b0;
    XRAM[19342] = 8'b0;
    XRAM[19343] = 8'b0;
    XRAM[19344] = 8'b0;
    XRAM[19345] = 8'b0;
    XRAM[19346] = 8'b0;
    XRAM[19347] = 8'b0;
    XRAM[19348] = 8'b0;
    XRAM[19349] = 8'b0;
    XRAM[19350] = 8'b0;
    XRAM[19351] = 8'b0;
    XRAM[19352] = 8'b0;
    XRAM[19353] = 8'b0;
    XRAM[19354] = 8'b0;
    XRAM[19355] = 8'b0;
    XRAM[19356] = 8'b0;
    XRAM[19357] = 8'b0;
    XRAM[19358] = 8'b0;
    XRAM[19359] = 8'b0;
    XRAM[19360] = 8'b0;
    XRAM[19361] = 8'b0;
    XRAM[19362] = 8'b0;
    XRAM[19363] = 8'b0;
    XRAM[19364] = 8'b0;
    XRAM[19365] = 8'b0;
    XRAM[19366] = 8'b0;
    XRAM[19367] = 8'b0;
    XRAM[19368] = 8'b0;
    XRAM[19369] = 8'b0;
    XRAM[19370] = 8'b0;
    XRAM[19371] = 8'b0;
    XRAM[19372] = 8'b0;
    XRAM[19373] = 8'b0;
    XRAM[19374] = 8'b0;
    XRAM[19375] = 8'b0;
    XRAM[19376] = 8'b0;
    XRAM[19377] = 8'b0;
    XRAM[19378] = 8'b0;
    XRAM[19379] = 8'b0;
    XRAM[19380] = 8'b0;
    XRAM[19381] = 8'b0;
    XRAM[19382] = 8'b0;
    XRAM[19383] = 8'b0;
    XRAM[19384] = 8'b0;
    XRAM[19385] = 8'b0;
    XRAM[19386] = 8'b0;
    XRAM[19387] = 8'b0;
    XRAM[19388] = 8'b0;
    XRAM[19389] = 8'b0;
    XRAM[19390] = 8'b0;
    XRAM[19391] = 8'b0;
    XRAM[19392] = 8'b0;
    XRAM[19393] = 8'b0;
    XRAM[19394] = 8'b0;
    XRAM[19395] = 8'b0;
    XRAM[19396] = 8'b0;
    XRAM[19397] = 8'b0;
    XRAM[19398] = 8'b0;
    XRAM[19399] = 8'b0;
    XRAM[19400] = 8'b0;
    XRAM[19401] = 8'b0;
    XRAM[19402] = 8'b0;
    XRAM[19403] = 8'b0;
    XRAM[19404] = 8'b0;
    XRAM[19405] = 8'b0;
    XRAM[19406] = 8'b0;
    XRAM[19407] = 8'b0;
    XRAM[19408] = 8'b0;
    XRAM[19409] = 8'b0;
    XRAM[19410] = 8'b0;
    XRAM[19411] = 8'b0;
    XRAM[19412] = 8'b0;
    XRAM[19413] = 8'b0;
    XRAM[19414] = 8'b0;
    XRAM[19415] = 8'b0;
    XRAM[19416] = 8'b0;
    XRAM[19417] = 8'b0;
    XRAM[19418] = 8'b0;
    XRAM[19419] = 8'b0;
    XRAM[19420] = 8'b0;
    XRAM[19421] = 8'b0;
    XRAM[19422] = 8'b0;
    XRAM[19423] = 8'b0;
    XRAM[19424] = 8'b0;
    XRAM[19425] = 8'b0;
    XRAM[19426] = 8'b0;
    XRAM[19427] = 8'b0;
    XRAM[19428] = 8'b0;
    XRAM[19429] = 8'b0;
    XRAM[19430] = 8'b0;
    XRAM[19431] = 8'b0;
    XRAM[19432] = 8'b0;
    XRAM[19433] = 8'b0;
    XRAM[19434] = 8'b0;
    XRAM[19435] = 8'b0;
    XRAM[19436] = 8'b0;
    XRAM[19437] = 8'b0;
    XRAM[19438] = 8'b0;
    XRAM[19439] = 8'b0;
    XRAM[19440] = 8'b0;
    XRAM[19441] = 8'b0;
    XRAM[19442] = 8'b0;
    XRAM[19443] = 8'b0;
    XRAM[19444] = 8'b0;
    XRAM[19445] = 8'b0;
    XRAM[19446] = 8'b0;
    XRAM[19447] = 8'b0;
    XRAM[19448] = 8'b0;
    XRAM[19449] = 8'b0;
    XRAM[19450] = 8'b0;
    XRAM[19451] = 8'b0;
    XRAM[19452] = 8'b0;
    XRAM[19453] = 8'b0;
    XRAM[19454] = 8'b0;
    XRAM[19455] = 8'b0;
    XRAM[19456] = 8'b0;
    XRAM[19457] = 8'b0;
    XRAM[19458] = 8'b0;
    XRAM[19459] = 8'b0;
    XRAM[19460] = 8'b0;
    XRAM[19461] = 8'b0;
    XRAM[19462] = 8'b0;
    XRAM[19463] = 8'b0;
    XRAM[19464] = 8'b0;
    XRAM[19465] = 8'b0;
    XRAM[19466] = 8'b0;
    XRAM[19467] = 8'b0;
    XRAM[19468] = 8'b0;
    XRAM[19469] = 8'b0;
    XRAM[19470] = 8'b0;
    XRAM[19471] = 8'b0;
    XRAM[19472] = 8'b0;
    XRAM[19473] = 8'b0;
    XRAM[19474] = 8'b0;
    XRAM[19475] = 8'b0;
    XRAM[19476] = 8'b0;
    XRAM[19477] = 8'b0;
    XRAM[19478] = 8'b0;
    XRAM[19479] = 8'b0;
    XRAM[19480] = 8'b0;
    XRAM[19481] = 8'b0;
    XRAM[19482] = 8'b0;
    XRAM[19483] = 8'b0;
    XRAM[19484] = 8'b0;
    XRAM[19485] = 8'b0;
    XRAM[19486] = 8'b0;
    XRAM[19487] = 8'b0;
    XRAM[19488] = 8'b0;
    XRAM[19489] = 8'b0;
    XRAM[19490] = 8'b0;
    XRAM[19491] = 8'b0;
    XRAM[19492] = 8'b0;
    XRAM[19493] = 8'b0;
    XRAM[19494] = 8'b0;
    XRAM[19495] = 8'b0;
    XRAM[19496] = 8'b0;
    XRAM[19497] = 8'b0;
    XRAM[19498] = 8'b0;
    XRAM[19499] = 8'b0;
    XRAM[19500] = 8'b0;
    XRAM[19501] = 8'b0;
    XRAM[19502] = 8'b0;
    XRAM[19503] = 8'b0;
    XRAM[19504] = 8'b0;
    XRAM[19505] = 8'b0;
    XRAM[19506] = 8'b0;
    XRAM[19507] = 8'b0;
    XRAM[19508] = 8'b0;
    XRAM[19509] = 8'b0;
    XRAM[19510] = 8'b0;
    XRAM[19511] = 8'b0;
    XRAM[19512] = 8'b0;
    XRAM[19513] = 8'b0;
    XRAM[19514] = 8'b0;
    XRAM[19515] = 8'b0;
    XRAM[19516] = 8'b0;
    XRAM[19517] = 8'b0;
    XRAM[19518] = 8'b0;
    XRAM[19519] = 8'b0;
    XRAM[19520] = 8'b0;
    XRAM[19521] = 8'b0;
    XRAM[19522] = 8'b0;
    XRAM[19523] = 8'b0;
    XRAM[19524] = 8'b0;
    XRAM[19525] = 8'b0;
    XRAM[19526] = 8'b0;
    XRAM[19527] = 8'b0;
    XRAM[19528] = 8'b0;
    XRAM[19529] = 8'b0;
    XRAM[19530] = 8'b0;
    XRAM[19531] = 8'b0;
    XRAM[19532] = 8'b0;
    XRAM[19533] = 8'b0;
    XRAM[19534] = 8'b0;
    XRAM[19535] = 8'b0;
    XRAM[19536] = 8'b0;
    XRAM[19537] = 8'b0;
    XRAM[19538] = 8'b0;
    XRAM[19539] = 8'b0;
    XRAM[19540] = 8'b0;
    XRAM[19541] = 8'b0;
    XRAM[19542] = 8'b0;
    XRAM[19543] = 8'b0;
    XRAM[19544] = 8'b0;
    XRAM[19545] = 8'b0;
    XRAM[19546] = 8'b0;
    XRAM[19547] = 8'b0;
    XRAM[19548] = 8'b0;
    XRAM[19549] = 8'b0;
    XRAM[19550] = 8'b0;
    XRAM[19551] = 8'b0;
    XRAM[19552] = 8'b0;
    XRAM[19553] = 8'b0;
    XRAM[19554] = 8'b0;
    XRAM[19555] = 8'b0;
    XRAM[19556] = 8'b0;
    XRAM[19557] = 8'b0;
    XRAM[19558] = 8'b0;
    XRAM[19559] = 8'b0;
    XRAM[19560] = 8'b0;
    XRAM[19561] = 8'b0;
    XRAM[19562] = 8'b0;
    XRAM[19563] = 8'b0;
    XRAM[19564] = 8'b0;
    XRAM[19565] = 8'b0;
    XRAM[19566] = 8'b0;
    XRAM[19567] = 8'b0;
    XRAM[19568] = 8'b0;
    XRAM[19569] = 8'b0;
    XRAM[19570] = 8'b0;
    XRAM[19571] = 8'b0;
    XRAM[19572] = 8'b0;
    XRAM[19573] = 8'b0;
    XRAM[19574] = 8'b0;
    XRAM[19575] = 8'b0;
    XRAM[19576] = 8'b0;
    XRAM[19577] = 8'b0;
    XRAM[19578] = 8'b0;
    XRAM[19579] = 8'b0;
    XRAM[19580] = 8'b0;
    XRAM[19581] = 8'b0;
    XRAM[19582] = 8'b0;
    XRAM[19583] = 8'b0;
    XRAM[19584] = 8'b0;
    XRAM[19585] = 8'b0;
    XRAM[19586] = 8'b0;
    XRAM[19587] = 8'b0;
    XRAM[19588] = 8'b0;
    XRAM[19589] = 8'b0;
    XRAM[19590] = 8'b0;
    XRAM[19591] = 8'b0;
    XRAM[19592] = 8'b0;
    XRAM[19593] = 8'b0;
    XRAM[19594] = 8'b0;
    XRAM[19595] = 8'b0;
    XRAM[19596] = 8'b0;
    XRAM[19597] = 8'b0;
    XRAM[19598] = 8'b0;
    XRAM[19599] = 8'b0;
    XRAM[19600] = 8'b0;
    XRAM[19601] = 8'b0;
    XRAM[19602] = 8'b0;
    XRAM[19603] = 8'b0;
    XRAM[19604] = 8'b0;
    XRAM[19605] = 8'b0;
    XRAM[19606] = 8'b0;
    XRAM[19607] = 8'b0;
    XRAM[19608] = 8'b0;
    XRAM[19609] = 8'b0;
    XRAM[19610] = 8'b0;
    XRAM[19611] = 8'b0;
    XRAM[19612] = 8'b0;
    XRAM[19613] = 8'b0;
    XRAM[19614] = 8'b0;
    XRAM[19615] = 8'b0;
    XRAM[19616] = 8'b0;
    XRAM[19617] = 8'b0;
    XRAM[19618] = 8'b0;
    XRAM[19619] = 8'b0;
    XRAM[19620] = 8'b0;
    XRAM[19621] = 8'b0;
    XRAM[19622] = 8'b0;
    XRAM[19623] = 8'b0;
    XRAM[19624] = 8'b0;
    XRAM[19625] = 8'b0;
    XRAM[19626] = 8'b0;
    XRAM[19627] = 8'b0;
    XRAM[19628] = 8'b0;
    XRAM[19629] = 8'b0;
    XRAM[19630] = 8'b0;
    XRAM[19631] = 8'b0;
    XRAM[19632] = 8'b0;
    XRAM[19633] = 8'b0;
    XRAM[19634] = 8'b0;
    XRAM[19635] = 8'b0;
    XRAM[19636] = 8'b0;
    XRAM[19637] = 8'b0;
    XRAM[19638] = 8'b0;
    XRAM[19639] = 8'b0;
    XRAM[19640] = 8'b0;
    XRAM[19641] = 8'b0;
    XRAM[19642] = 8'b0;
    XRAM[19643] = 8'b0;
    XRAM[19644] = 8'b0;
    XRAM[19645] = 8'b0;
    XRAM[19646] = 8'b0;
    XRAM[19647] = 8'b0;
    XRAM[19648] = 8'b0;
    XRAM[19649] = 8'b0;
    XRAM[19650] = 8'b0;
    XRAM[19651] = 8'b0;
    XRAM[19652] = 8'b0;
    XRAM[19653] = 8'b0;
    XRAM[19654] = 8'b0;
    XRAM[19655] = 8'b0;
    XRAM[19656] = 8'b0;
    XRAM[19657] = 8'b0;
    XRAM[19658] = 8'b0;
    XRAM[19659] = 8'b0;
    XRAM[19660] = 8'b0;
    XRAM[19661] = 8'b0;
    XRAM[19662] = 8'b0;
    XRAM[19663] = 8'b0;
    XRAM[19664] = 8'b0;
    XRAM[19665] = 8'b0;
    XRAM[19666] = 8'b0;
    XRAM[19667] = 8'b0;
    XRAM[19668] = 8'b0;
    XRAM[19669] = 8'b0;
    XRAM[19670] = 8'b0;
    XRAM[19671] = 8'b0;
    XRAM[19672] = 8'b0;
    XRAM[19673] = 8'b0;
    XRAM[19674] = 8'b0;
    XRAM[19675] = 8'b0;
    XRAM[19676] = 8'b0;
    XRAM[19677] = 8'b0;
    XRAM[19678] = 8'b0;
    XRAM[19679] = 8'b0;
    XRAM[19680] = 8'b0;
    XRAM[19681] = 8'b0;
    XRAM[19682] = 8'b0;
    XRAM[19683] = 8'b0;
    XRAM[19684] = 8'b0;
    XRAM[19685] = 8'b0;
    XRAM[19686] = 8'b0;
    XRAM[19687] = 8'b0;
    XRAM[19688] = 8'b0;
    XRAM[19689] = 8'b0;
    XRAM[19690] = 8'b0;
    XRAM[19691] = 8'b0;
    XRAM[19692] = 8'b0;
    XRAM[19693] = 8'b0;
    XRAM[19694] = 8'b0;
    XRAM[19695] = 8'b0;
    XRAM[19696] = 8'b0;
    XRAM[19697] = 8'b0;
    XRAM[19698] = 8'b0;
    XRAM[19699] = 8'b0;
    XRAM[19700] = 8'b0;
    XRAM[19701] = 8'b0;
    XRAM[19702] = 8'b0;
    XRAM[19703] = 8'b0;
    XRAM[19704] = 8'b0;
    XRAM[19705] = 8'b0;
    XRAM[19706] = 8'b0;
    XRAM[19707] = 8'b0;
    XRAM[19708] = 8'b0;
    XRAM[19709] = 8'b0;
    XRAM[19710] = 8'b0;
    XRAM[19711] = 8'b0;
    XRAM[19712] = 8'b0;
    XRAM[19713] = 8'b0;
    XRAM[19714] = 8'b0;
    XRAM[19715] = 8'b0;
    XRAM[19716] = 8'b0;
    XRAM[19717] = 8'b0;
    XRAM[19718] = 8'b0;
    XRAM[19719] = 8'b0;
    XRAM[19720] = 8'b0;
    XRAM[19721] = 8'b0;
    XRAM[19722] = 8'b0;
    XRAM[19723] = 8'b0;
    XRAM[19724] = 8'b0;
    XRAM[19725] = 8'b0;
    XRAM[19726] = 8'b0;
    XRAM[19727] = 8'b0;
    XRAM[19728] = 8'b0;
    XRAM[19729] = 8'b0;
    XRAM[19730] = 8'b0;
    XRAM[19731] = 8'b0;
    XRAM[19732] = 8'b0;
    XRAM[19733] = 8'b0;
    XRAM[19734] = 8'b0;
    XRAM[19735] = 8'b0;
    XRAM[19736] = 8'b0;
    XRAM[19737] = 8'b0;
    XRAM[19738] = 8'b0;
    XRAM[19739] = 8'b0;
    XRAM[19740] = 8'b0;
    XRAM[19741] = 8'b0;
    XRAM[19742] = 8'b0;
    XRAM[19743] = 8'b0;
    XRAM[19744] = 8'b0;
    XRAM[19745] = 8'b0;
    XRAM[19746] = 8'b0;
    XRAM[19747] = 8'b0;
    XRAM[19748] = 8'b0;
    XRAM[19749] = 8'b0;
    XRAM[19750] = 8'b0;
    XRAM[19751] = 8'b0;
    XRAM[19752] = 8'b0;
    XRAM[19753] = 8'b0;
    XRAM[19754] = 8'b0;
    XRAM[19755] = 8'b0;
    XRAM[19756] = 8'b0;
    XRAM[19757] = 8'b0;
    XRAM[19758] = 8'b0;
    XRAM[19759] = 8'b0;
    XRAM[19760] = 8'b0;
    XRAM[19761] = 8'b0;
    XRAM[19762] = 8'b0;
    XRAM[19763] = 8'b0;
    XRAM[19764] = 8'b0;
    XRAM[19765] = 8'b0;
    XRAM[19766] = 8'b0;
    XRAM[19767] = 8'b0;
    XRAM[19768] = 8'b0;
    XRAM[19769] = 8'b0;
    XRAM[19770] = 8'b0;
    XRAM[19771] = 8'b0;
    XRAM[19772] = 8'b0;
    XRAM[19773] = 8'b0;
    XRAM[19774] = 8'b0;
    XRAM[19775] = 8'b0;
    XRAM[19776] = 8'b0;
    XRAM[19777] = 8'b0;
    XRAM[19778] = 8'b0;
    XRAM[19779] = 8'b0;
    XRAM[19780] = 8'b0;
    XRAM[19781] = 8'b0;
    XRAM[19782] = 8'b0;
    XRAM[19783] = 8'b0;
    XRAM[19784] = 8'b0;
    XRAM[19785] = 8'b0;
    XRAM[19786] = 8'b0;
    XRAM[19787] = 8'b0;
    XRAM[19788] = 8'b0;
    XRAM[19789] = 8'b0;
    XRAM[19790] = 8'b0;
    XRAM[19791] = 8'b0;
    XRAM[19792] = 8'b0;
    XRAM[19793] = 8'b0;
    XRAM[19794] = 8'b0;
    XRAM[19795] = 8'b0;
    XRAM[19796] = 8'b0;
    XRAM[19797] = 8'b0;
    XRAM[19798] = 8'b0;
    XRAM[19799] = 8'b0;
    XRAM[19800] = 8'b0;
    XRAM[19801] = 8'b0;
    XRAM[19802] = 8'b0;
    XRAM[19803] = 8'b0;
    XRAM[19804] = 8'b0;
    XRAM[19805] = 8'b0;
    XRAM[19806] = 8'b0;
    XRAM[19807] = 8'b0;
    XRAM[19808] = 8'b0;
    XRAM[19809] = 8'b0;
    XRAM[19810] = 8'b0;
    XRAM[19811] = 8'b0;
    XRAM[19812] = 8'b0;
    XRAM[19813] = 8'b0;
    XRAM[19814] = 8'b0;
    XRAM[19815] = 8'b0;
    XRAM[19816] = 8'b0;
    XRAM[19817] = 8'b0;
    XRAM[19818] = 8'b0;
    XRAM[19819] = 8'b0;
    XRAM[19820] = 8'b0;
    XRAM[19821] = 8'b0;
    XRAM[19822] = 8'b0;
    XRAM[19823] = 8'b0;
    XRAM[19824] = 8'b0;
    XRAM[19825] = 8'b0;
    XRAM[19826] = 8'b0;
    XRAM[19827] = 8'b0;
    XRAM[19828] = 8'b0;
    XRAM[19829] = 8'b0;
    XRAM[19830] = 8'b0;
    XRAM[19831] = 8'b0;
    XRAM[19832] = 8'b0;
    XRAM[19833] = 8'b0;
    XRAM[19834] = 8'b0;
    XRAM[19835] = 8'b0;
    XRAM[19836] = 8'b0;
    XRAM[19837] = 8'b0;
    XRAM[19838] = 8'b0;
    XRAM[19839] = 8'b0;
    XRAM[19840] = 8'b0;
    XRAM[19841] = 8'b0;
    XRAM[19842] = 8'b0;
    XRAM[19843] = 8'b0;
    XRAM[19844] = 8'b0;
    XRAM[19845] = 8'b0;
    XRAM[19846] = 8'b0;
    XRAM[19847] = 8'b0;
    XRAM[19848] = 8'b0;
    XRAM[19849] = 8'b0;
    XRAM[19850] = 8'b0;
    XRAM[19851] = 8'b0;
    XRAM[19852] = 8'b0;
    XRAM[19853] = 8'b0;
    XRAM[19854] = 8'b0;
    XRAM[19855] = 8'b0;
    XRAM[19856] = 8'b0;
    XRAM[19857] = 8'b0;
    XRAM[19858] = 8'b0;
    XRAM[19859] = 8'b0;
    XRAM[19860] = 8'b0;
    XRAM[19861] = 8'b0;
    XRAM[19862] = 8'b0;
    XRAM[19863] = 8'b0;
    XRAM[19864] = 8'b0;
    XRAM[19865] = 8'b0;
    XRAM[19866] = 8'b0;
    XRAM[19867] = 8'b0;
    XRAM[19868] = 8'b0;
    XRAM[19869] = 8'b0;
    XRAM[19870] = 8'b0;
    XRAM[19871] = 8'b0;
    XRAM[19872] = 8'b0;
    XRAM[19873] = 8'b0;
    XRAM[19874] = 8'b0;
    XRAM[19875] = 8'b0;
    XRAM[19876] = 8'b0;
    XRAM[19877] = 8'b0;
    XRAM[19878] = 8'b0;
    XRAM[19879] = 8'b0;
    XRAM[19880] = 8'b0;
    XRAM[19881] = 8'b0;
    XRAM[19882] = 8'b0;
    XRAM[19883] = 8'b0;
    XRAM[19884] = 8'b0;
    XRAM[19885] = 8'b0;
    XRAM[19886] = 8'b0;
    XRAM[19887] = 8'b0;
    XRAM[19888] = 8'b0;
    XRAM[19889] = 8'b0;
    XRAM[19890] = 8'b0;
    XRAM[19891] = 8'b0;
    XRAM[19892] = 8'b0;
    XRAM[19893] = 8'b0;
    XRAM[19894] = 8'b0;
    XRAM[19895] = 8'b0;
    XRAM[19896] = 8'b0;
    XRAM[19897] = 8'b0;
    XRAM[19898] = 8'b0;
    XRAM[19899] = 8'b0;
    XRAM[19900] = 8'b0;
    XRAM[19901] = 8'b0;
    XRAM[19902] = 8'b0;
    XRAM[19903] = 8'b0;
    XRAM[19904] = 8'b0;
    XRAM[19905] = 8'b0;
    XRAM[19906] = 8'b0;
    XRAM[19907] = 8'b0;
    XRAM[19908] = 8'b0;
    XRAM[19909] = 8'b0;
    XRAM[19910] = 8'b0;
    XRAM[19911] = 8'b0;
    XRAM[19912] = 8'b0;
    XRAM[19913] = 8'b0;
    XRAM[19914] = 8'b0;
    XRAM[19915] = 8'b0;
    XRAM[19916] = 8'b0;
    XRAM[19917] = 8'b0;
    XRAM[19918] = 8'b0;
    XRAM[19919] = 8'b0;
    XRAM[19920] = 8'b0;
    XRAM[19921] = 8'b0;
    XRAM[19922] = 8'b0;
    XRAM[19923] = 8'b0;
    XRAM[19924] = 8'b0;
    XRAM[19925] = 8'b0;
    XRAM[19926] = 8'b0;
    XRAM[19927] = 8'b0;
    XRAM[19928] = 8'b0;
    XRAM[19929] = 8'b0;
    XRAM[19930] = 8'b0;
    XRAM[19931] = 8'b0;
    XRAM[19932] = 8'b0;
    XRAM[19933] = 8'b0;
    XRAM[19934] = 8'b0;
    XRAM[19935] = 8'b0;
    XRAM[19936] = 8'b0;
    XRAM[19937] = 8'b0;
    XRAM[19938] = 8'b0;
    XRAM[19939] = 8'b0;
    XRAM[19940] = 8'b0;
    XRAM[19941] = 8'b0;
    XRAM[19942] = 8'b0;
    XRAM[19943] = 8'b0;
    XRAM[19944] = 8'b0;
    XRAM[19945] = 8'b0;
    XRAM[19946] = 8'b0;
    XRAM[19947] = 8'b0;
    XRAM[19948] = 8'b0;
    XRAM[19949] = 8'b0;
    XRAM[19950] = 8'b0;
    XRAM[19951] = 8'b0;
    XRAM[19952] = 8'b0;
    XRAM[19953] = 8'b0;
    XRAM[19954] = 8'b0;
    XRAM[19955] = 8'b0;
    XRAM[19956] = 8'b0;
    XRAM[19957] = 8'b0;
    XRAM[19958] = 8'b0;
    XRAM[19959] = 8'b0;
    XRAM[19960] = 8'b0;
    XRAM[19961] = 8'b0;
    XRAM[19962] = 8'b0;
    XRAM[19963] = 8'b0;
    XRAM[19964] = 8'b0;
    XRAM[19965] = 8'b0;
    XRAM[19966] = 8'b0;
    XRAM[19967] = 8'b0;
    XRAM[19968] = 8'b0;
    XRAM[19969] = 8'b0;
    XRAM[19970] = 8'b0;
    XRAM[19971] = 8'b0;
    XRAM[19972] = 8'b0;
    XRAM[19973] = 8'b0;
    XRAM[19974] = 8'b0;
    XRAM[19975] = 8'b0;
    XRAM[19976] = 8'b0;
    XRAM[19977] = 8'b0;
    XRAM[19978] = 8'b0;
    XRAM[19979] = 8'b0;
    XRAM[19980] = 8'b0;
    XRAM[19981] = 8'b0;
    XRAM[19982] = 8'b0;
    XRAM[19983] = 8'b0;
    XRAM[19984] = 8'b0;
    XRAM[19985] = 8'b0;
    XRAM[19986] = 8'b0;
    XRAM[19987] = 8'b0;
    XRAM[19988] = 8'b0;
    XRAM[19989] = 8'b0;
    XRAM[19990] = 8'b0;
    XRAM[19991] = 8'b0;
    XRAM[19992] = 8'b0;
    XRAM[19993] = 8'b0;
    XRAM[19994] = 8'b0;
    XRAM[19995] = 8'b0;
    XRAM[19996] = 8'b0;
    XRAM[19997] = 8'b0;
    XRAM[19998] = 8'b0;
    XRAM[19999] = 8'b0;
    XRAM[20000] = 8'b0;
    XRAM[20001] = 8'b0;
    XRAM[20002] = 8'b0;
    XRAM[20003] = 8'b0;
    XRAM[20004] = 8'b0;
    XRAM[20005] = 8'b0;
    XRAM[20006] = 8'b0;
    XRAM[20007] = 8'b0;
    XRAM[20008] = 8'b0;
    XRAM[20009] = 8'b0;
    XRAM[20010] = 8'b0;
    XRAM[20011] = 8'b0;
    XRAM[20012] = 8'b0;
    XRAM[20013] = 8'b0;
    XRAM[20014] = 8'b0;
    XRAM[20015] = 8'b0;
    XRAM[20016] = 8'b0;
    XRAM[20017] = 8'b0;
    XRAM[20018] = 8'b0;
    XRAM[20019] = 8'b0;
    XRAM[20020] = 8'b0;
    XRAM[20021] = 8'b0;
    XRAM[20022] = 8'b0;
    XRAM[20023] = 8'b0;
    XRAM[20024] = 8'b0;
    XRAM[20025] = 8'b0;
    XRAM[20026] = 8'b0;
    XRAM[20027] = 8'b0;
    XRAM[20028] = 8'b0;
    XRAM[20029] = 8'b0;
    XRAM[20030] = 8'b0;
    XRAM[20031] = 8'b0;
    XRAM[20032] = 8'b0;
    XRAM[20033] = 8'b0;
    XRAM[20034] = 8'b0;
    XRAM[20035] = 8'b0;
    XRAM[20036] = 8'b0;
    XRAM[20037] = 8'b0;
    XRAM[20038] = 8'b0;
    XRAM[20039] = 8'b0;
    XRAM[20040] = 8'b0;
    XRAM[20041] = 8'b0;
    XRAM[20042] = 8'b0;
    XRAM[20043] = 8'b0;
    XRAM[20044] = 8'b0;
    XRAM[20045] = 8'b0;
    XRAM[20046] = 8'b0;
    XRAM[20047] = 8'b0;
    XRAM[20048] = 8'b0;
    XRAM[20049] = 8'b0;
    XRAM[20050] = 8'b0;
    XRAM[20051] = 8'b0;
    XRAM[20052] = 8'b0;
    XRAM[20053] = 8'b0;
    XRAM[20054] = 8'b0;
    XRAM[20055] = 8'b0;
    XRAM[20056] = 8'b0;
    XRAM[20057] = 8'b0;
    XRAM[20058] = 8'b0;
    XRAM[20059] = 8'b0;
    XRAM[20060] = 8'b0;
    XRAM[20061] = 8'b0;
    XRAM[20062] = 8'b0;
    XRAM[20063] = 8'b0;
    XRAM[20064] = 8'b0;
    XRAM[20065] = 8'b0;
    XRAM[20066] = 8'b0;
    XRAM[20067] = 8'b0;
    XRAM[20068] = 8'b0;
    XRAM[20069] = 8'b0;
    XRAM[20070] = 8'b0;
    XRAM[20071] = 8'b0;
    XRAM[20072] = 8'b0;
    XRAM[20073] = 8'b0;
    XRAM[20074] = 8'b0;
    XRAM[20075] = 8'b0;
    XRAM[20076] = 8'b0;
    XRAM[20077] = 8'b0;
    XRAM[20078] = 8'b0;
    XRAM[20079] = 8'b0;
    XRAM[20080] = 8'b0;
    XRAM[20081] = 8'b0;
    XRAM[20082] = 8'b0;
    XRAM[20083] = 8'b0;
    XRAM[20084] = 8'b0;
    XRAM[20085] = 8'b0;
    XRAM[20086] = 8'b0;
    XRAM[20087] = 8'b0;
    XRAM[20088] = 8'b0;
    XRAM[20089] = 8'b0;
    XRAM[20090] = 8'b0;
    XRAM[20091] = 8'b0;
    XRAM[20092] = 8'b0;
    XRAM[20093] = 8'b0;
    XRAM[20094] = 8'b0;
    XRAM[20095] = 8'b0;
    XRAM[20096] = 8'b0;
    XRAM[20097] = 8'b0;
    XRAM[20098] = 8'b0;
    XRAM[20099] = 8'b0;
    XRAM[20100] = 8'b0;
    XRAM[20101] = 8'b0;
    XRAM[20102] = 8'b0;
    XRAM[20103] = 8'b0;
    XRAM[20104] = 8'b0;
    XRAM[20105] = 8'b0;
    XRAM[20106] = 8'b0;
    XRAM[20107] = 8'b0;
    XRAM[20108] = 8'b0;
    XRAM[20109] = 8'b0;
    XRAM[20110] = 8'b0;
    XRAM[20111] = 8'b0;
    XRAM[20112] = 8'b0;
    XRAM[20113] = 8'b0;
    XRAM[20114] = 8'b0;
    XRAM[20115] = 8'b0;
    XRAM[20116] = 8'b0;
    XRAM[20117] = 8'b0;
    XRAM[20118] = 8'b0;
    XRAM[20119] = 8'b0;
    XRAM[20120] = 8'b0;
    XRAM[20121] = 8'b0;
    XRAM[20122] = 8'b0;
    XRAM[20123] = 8'b0;
    XRAM[20124] = 8'b0;
    XRAM[20125] = 8'b0;
    XRAM[20126] = 8'b0;
    XRAM[20127] = 8'b0;
    XRAM[20128] = 8'b0;
    XRAM[20129] = 8'b0;
    XRAM[20130] = 8'b0;
    XRAM[20131] = 8'b0;
    XRAM[20132] = 8'b0;
    XRAM[20133] = 8'b0;
    XRAM[20134] = 8'b0;
    XRAM[20135] = 8'b0;
    XRAM[20136] = 8'b0;
    XRAM[20137] = 8'b0;
    XRAM[20138] = 8'b0;
    XRAM[20139] = 8'b0;
    XRAM[20140] = 8'b0;
    XRAM[20141] = 8'b0;
    XRAM[20142] = 8'b0;
    XRAM[20143] = 8'b0;
    XRAM[20144] = 8'b0;
    XRAM[20145] = 8'b0;
    XRAM[20146] = 8'b0;
    XRAM[20147] = 8'b0;
    XRAM[20148] = 8'b0;
    XRAM[20149] = 8'b0;
    XRAM[20150] = 8'b0;
    XRAM[20151] = 8'b0;
    XRAM[20152] = 8'b0;
    XRAM[20153] = 8'b0;
    XRAM[20154] = 8'b0;
    XRAM[20155] = 8'b0;
    XRAM[20156] = 8'b0;
    XRAM[20157] = 8'b0;
    XRAM[20158] = 8'b0;
    XRAM[20159] = 8'b0;
    XRAM[20160] = 8'b0;
    XRAM[20161] = 8'b0;
    XRAM[20162] = 8'b0;
    XRAM[20163] = 8'b0;
    XRAM[20164] = 8'b0;
    XRAM[20165] = 8'b0;
    XRAM[20166] = 8'b0;
    XRAM[20167] = 8'b0;
    XRAM[20168] = 8'b0;
    XRAM[20169] = 8'b0;
    XRAM[20170] = 8'b0;
    XRAM[20171] = 8'b0;
    XRAM[20172] = 8'b0;
    XRAM[20173] = 8'b0;
    XRAM[20174] = 8'b0;
    XRAM[20175] = 8'b0;
    XRAM[20176] = 8'b0;
    XRAM[20177] = 8'b0;
    XRAM[20178] = 8'b0;
    XRAM[20179] = 8'b0;
    XRAM[20180] = 8'b0;
    XRAM[20181] = 8'b0;
    XRAM[20182] = 8'b0;
    XRAM[20183] = 8'b0;
    XRAM[20184] = 8'b0;
    XRAM[20185] = 8'b0;
    XRAM[20186] = 8'b0;
    XRAM[20187] = 8'b0;
    XRAM[20188] = 8'b0;
    XRAM[20189] = 8'b0;
    XRAM[20190] = 8'b0;
    XRAM[20191] = 8'b0;
    XRAM[20192] = 8'b0;
    XRAM[20193] = 8'b0;
    XRAM[20194] = 8'b0;
    XRAM[20195] = 8'b0;
    XRAM[20196] = 8'b0;
    XRAM[20197] = 8'b0;
    XRAM[20198] = 8'b0;
    XRAM[20199] = 8'b0;
    XRAM[20200] = 8'b0;
    XRAM[20201] = 8'b0;
    XRAM[20202] = 8'b0;
    XRAM[20203] = 8'b0;
    XRAM[20204] = 8'b0;
    XRAM[20205] = 8'b0;
    XRAM[20206] = 8'b0;
    XRAM[20207] = 8'b0;
    XRAM[20208] = 8'b0;
    XRAM[20209] = 8'b0;
    XRAM[20210] = 8'b0;
    XRAM[20211] = 8'b0;
    XRAM[20212] = 8'b0;
    XRAM[20213] = 8'b0;
    XRAM[20214] = 8'b0;
    XRAM[20215] = 8'b0;
    XRAM[20216] = 8'b0;
    XRAM[20217] = 8'b0;
    XRAM[20218] = 8'b0;
    XRAM[20219] = 8'b0;
    XRAM[20220] = 8'b0;
    XRAM[20221] = 8'b0;
    XRAM[20222] = 8'b0;
    XRAM[20223] = 8'b0;
    XRAM[20224] = 8'b0;
    XRAM[20225] = 8'b0;
    XRAM[20226] = 8'b0;
    XRAM[20227] = 8'b0;
    XRAM[20228] = 8'b0;
    XRAM[20229] = 8'b0;
    XRAM[20230] = 8'b0;
    XRAM[20231] = 8'b0;
    XRAM[20232] = 8'b0;
    XRAM[20233] = 8'b0;
    XRAM[20234] = 8'b0;
    XRAM[20235] = 8'b0;
    XRAM[20236] = 8'b0;
    XRAM[20237] = 8'b0;
    XRAM[20238] = 8'b0;
    XRAM[20239] = 8'b0;
    XRAM[20240] = 8'b0;
    XRAM[20241] = 8'b0;
    XRAM[20242] = 8'b0;
    XRAM[20243] = 8'b0;
    XRAM[20244] = 8'b0;
    XRAM[20245] = 8'b0;
    XRAM[20246] = 8'b0;
    XRAM[20247] = 8'b0;
    XRAM[20248] = 8'b0;
    XRAM[20249] = 8'b0;
    XRAM[20250] = 8'b0;
    XRAM[20251] = 8'b0;
    XRAM[20252] = 8'b0;
    XRAM[20253] = 8'b0;
    XRAM[20254] = 8'b0;
    XRAM[20255] = 8'b0;
    XRAM[20256] = 8'b0;
    XRAM[20257] = 8'b0;
    XRAM[20258] = 8'b0;
    XRAM[20259] = 8'b0;
    XRAM[20260] = 8'b0;
    XRAM[20261] = 8'b0;
    XRAM[20262] = 8'b0;
    XRAM[20263] = 8'b0;
    XRAM[20264] = 8'b0;
    XRAM[20265] = 8'b0;
    XRAM[20266] = 8'b0;
    XRAM[20267] = 8'b0;
    XRAM[20268] = 8'b0;
    XRAM[20269] = 8'b0;
    XRAM[20270] = 8'b0;
    XRAM[20271] = 8'b0;
    XRAM[20272] = 8'b0;
    XRAM[20273] = 8'b0;
    XRAM[20274] = 8'b0;
    XRAM[20275] = 8'b0;
    XRAM[20276] = 8'b0;
    XRAM[20277] = 8'b0;
    XRAM[20278] = 8'b0;
    XRAM[20279] = 8'b0;
    XRAM[20280] = 8'b0;
    XRAM[20281] = 8'b0;
    XRAM[20282] = 8'b0;
    XRAM[20283] = 8'b0;
    XRAM[20284] = 8'b0;
    XRAM[20285] = 8'b0;
    XRAM[20286] = 8'b0;
    XRAM[20287] = 8'b0;
    XRAM[20288] = 8'b0;
    XRAM[20289] = 8'b0;
    XRAM[20290] = 8'b0;
    XRAM[20291] = 8'b0;
    XRAM[20292] = 8'b0;
    XRAM[20293] = 8'b0;
    XRAM[20294] = 8'b0;
    XRAM[20295] = 8'b0;
    XRAM[20296] = 8'b0;
    XRAM[20297] = 8'b0;
    XRAM[20298] = 8'b0;
    XRAM[20299] = 8'b0;
    XRAM[20300] = 8'b0;
    XRAM[20301] = 8'b0;
    XRAM[20302] = 8'b0;
    XRAM[20303] = 8'b0;
    XRAM[20304] = 8'b0;
    XRAM[20305] = 8'b0;
    XRAM[20306] = 8'b0;
    XRAM[20307] = 8'b0;
    XRAM[20308] = 8'b0;
    XRAM[20309] = 8'b0;
    XRAM[20310] = 8'b0;
    XRAM[20311] = 8'b0;
    XRAM[20312] = 8'b0;
    XRAM[20313] = 8'b0;
    XRAM[20314] = 8'b0;
    XRAM[20315] = 8'b0;
    XRAM[20316] = 8'b0;
    XRAM[20317] = 8'b0;
    XRAM[20318] = 8'b0;
    XRAM[20319] = 8'b0;
    XRAM[20320] = 8'b0;
    XRAM[20321] = 8'b0;
    XRAM[20322] = 8'b0;
    XRAM[20323] = 8'b0;
    XRAM[20324] = 8'b0;
    XRAM[20325] = 8'b0;
    XRAM[20326] = 8'b0;
    XRAM[20327] = 8'b0;
    XRAM[20328] = 8'b0;
    XRAM[20329] = 8'b0;
    XRAM[20330] = 8'b0;
    XRAM[20331] = 8'b0;
    XRAM[20332] = 8'b0;
    XRAM[20333] = 8'b0;
    XRAM[20334] = 8'b0;
    XRAM[20335] = 8'b0;
    XRAM[20336] = 8'b0;
    XRAM[20337] = 8'b0;
    XRAM[20338] = 8'b0;
    XRAM[20339] = 8'b0;
    XRAM[20340] = 8'b0;
    XRAM[20341] = 8'b0;
    XRAM[20342] = 8'b0;
    XRAM[20343] = 8'b0;
    XRAM[20344] = 8'b0;
    XRAM[20345] = 8'b0;
    XRAM[20346] = 8'b0;
    XRAM[20347] = 8'b0;
    XRAM[20348] = 8'b0;
    XRAM[20349] = 8'b0;
    XRAM[20350] = 8'b0;
    XRAM[20351] = 8'b0;
    XRAM[20352] = 8'b0;
    XRAM[20353] = 8'b0;
    XRAM[20354] = 8'b0;
    XRAM[20355] = 8'b0;
    XRAM[20356] = 8'b0;
    XRAM[20357] = 8'b0;
    XRAM[20358] = 8'b0;
    XRAM[20359] = 8'b0;
    XRAM[20360] = 8'b0;
    XRAM[20361] = 8'b0;
    XRAM[20362] = 8'b0;
    XRAM[20363] = 8'b0;
    XRAM[20364] = 8'b0;
    XRAM[20365] = 8'b0;
    XRAM[20366] = 8'b0;
    XRAM[20367] = 8'b0;
    XRAM[20368] = 8'b0;
    XRAM[20369] = 8'b0;
    XRAM[20370] = 8'b0;
    XRAM[20371] = 8'b0;
    XRAM[20372] = 8'b0;
    XRAM[20373] = 8'b0;
    XRAM[20374] = 8'b0;
    XRAM[20375] = 8'b0;
    XRAM[20376] = 8'b0;
    XRAM[20377] = 8'b0;
    XRAM[20378] = 8'b0;
    XRAM[20379] = 8'b0;
    XRAM[20380] = 8'b0;
    XRAM[20381] = 8'b0;
    XRAM[20382] = 8'b0;
    XRAM[20383] = 8'b0;
    XRAM[20384] = 8'b0;
    XRAM[20385] = 8'b0;
    XRAM[20386] = 8'b0;
    XRAM[20387] = 8'b0;
    XRAM[20388] = 8'b0;
    XRAM[20389] = 8'b0;
    XRAM[20390] = 8'b0;
    XRAM[20391] = 8'b0;
    XRAM[20392] = 8'b0;
    XRAM[20393] = 8'b0;
    XRAM[20394] = 8'b0;
    XRAM[20395] = 8'b0;
    XRAM[20396] = 8'b0;
    XRAM[20397] = 8'b0;
    XRAM[20398] = 8'b0;
    XRAM[20399] = 8'b0;
    XRAM[20400] = 8'b0;
    XRAM[20401] = 8'b0;
    XRAM[20402] = 8'b0;
    XRAM[20403] = 8'b0;
    XRAM[20404] = 8'b0;
    XRAM[20405] = 8'b0;
    XRAM[20406] = 8'b0;
    XRAM[20407] = 8'b0;
    XRAM[20408] = 8'b0;
    XRAM[20409] = 8'b0;
    XRAM[20410] = 8'b0;
    XRAM[20411] = 8'b0;
    XRAM[20412] = 8'b0;
    XRAM[20413] = 8'b0;
    XRAM[20414] = 8'b0;
    XRAM[20415] = 8'b0;
    XRAM[20416] = 8'b0;
    XRAM[20417] = 8'b0;
    XRAM[20418] = 8'b0;
    XRAM[20419] = 8'b0;
    XRAM[20420] = 8'b0;
    XRAM[20421] = 8'b0;
    XRAM[20422] = 8'b0;
    XRAM[20423] = 8'b0;
    XRAM[20424] = 8'b0;
    XRAM[20425] = 8'b0;
    XRAM[20426] = 8'b0;
    XRAM[20427] = 8'b0;
    XRAM[20428] = 8'b0;
    XRAM[20429] = 8'b0;
    XRAM[20430] = 8'b0;
    XRAM[20431] = 8'b0;
    XRAM[20432] = 8'b0;
    XRAM[20433] = 8'b0;
    XRAM[20434] = 8'b0;
    XRAM[20435] = 8'b0;
    XRAM[20436] = 8'b0;
    XRAM[20437] = 8'b0;
    XRAM[20438] = 8'b0;
    XRAM[20439] = 8'b0;
    XRAM[20440] = 8'b0;
    XRAM[20441] = 8'b0;
    XRAM[20442] = 8'b0;
    XRAM[20443] = 8'b0;
    XRAM[20444] = 8'b0;
    XRAM[20445] = 8'b0;
    XRAM[20446] = 8'b0;
    XRAM[20447] = 8'b0;
    XRAM[20448] = 8'b0;
    XRAM[20449] = 8'b0;
    XRAM[20450] = 8'b0;
    XRAM[20451] = 8'b0;
    XRAM[20452] = 8'b0;
    XRAM[20453] = 8'b0;
    XRAM[20454] = 8'b0;
    XRAM[20455] = 8'b0;
    XRAM[20456] = 8'b0;
    XRAM[20457] = 8'b0;
    XRAM[20458] = 8'b0;
    XRAM[20459] = 8'b0;
    XRAM[20460] = 8'b0;
    XRAM[20461] = 8'b0;
    XRAM[20462] = 8'b0;
    XRAM[20463] = 8'b0;
    XRAM[20464] = 8'b0;
    XRAM[20465] = 8'b0;
    XRAM[20466] = 8'b0;
    XRAM[20467] = 8'b0;
    XRAM[20468] = 8'b0;
    XRAM[20469] = 8'b0;
    XRAM[20470] = 8'b0;
    XRAM[20471] = 8'b0;
    XRAM[20472] = 8'b0;
    XRAM[20473] = 8'b0;
    XRAM[20474] = 8'b0;
    XRAM[20475] = 8'b0;
    XRAM[20476] = 8'b0;
    XRAM[20477] = 8'b0;
    XRAM[20478] = 8'b0;
    XRAM[20479] = 8'b0;
    XRAM[20480] = 8'b0;
    XRAM[20481] = 8'b0;
    XRAM[20482] = 8'b0;
    XRAM[20483] = 8'b0;
    XRAM[20484] = 8'b0;
    XRAM[20485] = 8'b0;
    XRAM[20486] = 8'b0;
    XRAM[20487] = 8'b0;
    XRAM[20488] = 8'b0;
    XRAM[20489] = 8'b0;
    XRAM[20490] = 8'b0;
    XRAM[20491] = 8'b0;
    XRAM[20492] = 8'b0;
    XRAM[20493] = 8'b0;
    XRAM[20494] = 8'b0;
    XRAM[20495] = 8'b0;
    XRAM[20496] = 8'b0;
    XRAM[20497] = 8'b0;
    XRAM[20498] = 8'b0;
    XRAM[20499] = 8'b0;
    XRAM[20500] = 8'b0;
    XRAM[20501] = 8'b0;
    XRAM[20502] = 8'b0;
    XRAM[20503] = 8'b0;
    XRAM[20504] = 8'b0;
    XRAM[20505] = 8'b0;
    XRAM[20506] = 8'b0;
    XRAM[20507] = 8'b0;
    XRAM[20508] = 8'b0;
    XRAM[20509] = 8'b0;
    XRAM[20510] = 8'b0;
    XRAM[20511] = 8'b0;
    XRAM[20512] = 8'b0;
    XRAM[20513] = 8'b0;
    XRAM[20514] = 8'b0;
    XRAM[20515] = 8'b0;
    XRAM[20516] = 8'b0;
    XRAM[20517] = 8'b0;
    XRAM[20518] = 8'b0;
    XRAM[20519] = 8'b0;
    XRAM[20520] = 8'b0;
    XRAM[20521] = 8'b0;
    XRAM[20522] = 8'b0;
    XRAM[20523] = 8'b0;
    XRAM[20524] = 8'b0;
    XRAM[20525] = 8'b0;
    XRAM[20526] = 8'b0;
    XRAM[20527] = 8'b0;
    XRAM[20528] = 8'b0;
    XRAM[20529] = 8'b0;
    XRAM[20530] = 8'b0;
    XRAM[20531] = 8'b0;
    XRAM[20532] = 8'b0;
    XRAM[20533] = 8'b0;
    XRAM[20534] = 8'b0;
    XRAM[20535] = 8'b0;
    XRAM[20536] = 8'b0;
    XRAM[20537] = 8'b0;
    XRAM[20538] = 8'b0;
    XRAM[20539] = 8'b0;
    XRAM[20540] = 8'b0;
    XRAM[20541] = 8'b0;
    XRAM[20542] = 8'b0;
    XRAM[20543] = 8'b0;
    XRAM[20544] = 8'b0;
    XRAM[20545] = 8'b0;
    XRAM[20546] = 8'b0;
    XRAM[20547] = 8'b0;
    XRAM[20548] = 8'b0;
    XRAM[20549] = 8'b0;
    XRAM[20550] = 8'b0;
    XRAM[20551] = 8'b0;
    XRAM[20552] = 8'b0;
    XRAM[20553] = 8'b0;
    XRAM[20554] = 8'b0;
    XRAM[20555] = 8'b0;
    XRAM[20556] = 8'b0;
    XRAM[20557] = 8'b0;
    XRAM[20558] = 8'b0;
    XRAM[20559] = 8'b0;
    XRAM[20560] = 8'b0;
    XRAM[20561] = 8'b0;
    XRAM[20562] = 8'b0;
    XRAM[20563] = 8'b0;
    XRAM[20564] = 8'b0;
    XRAM[20565] = 8'b0;
    XRAM[20566] = 8'b0;
    XRAM[20567] = 8'b0;
    XRAM[20568] = 8'b0;
    XRAM[20569] = 8'b0;
    XRAM[20570] = 8'b0;
    XRAM[20571] = 8'b0;
    XRAM[20572] = 8'b0;
    XRAM[20573] = 8'b0;
    XRAM[20574] = 8'b0;
    XRAM[20575] = 8'b0;
    XRAM[20576] = 8'b0;
    XRAM[20577] = 8'b0;
    XRAM[20578] = 8'b0;
    XRAM[20579] = 8'b0;
    XRAM[20580] = 8'b0;
    XRAM[20581] = 8'b0;
    XRAM[20582] = 8'b0;
    XRAM[20583] = 8'b0;
    XRAM[20584] = 8'b0;
    XRAM[20585] = 8'b0;
    XRAM[20586] = 8'b0;
    XRAM[20587] = 8'b0;
    XRAM[20588] = 8'b0;
    XRAM[20589] = 8'b0;
    XRAM[20590] = 8'b0;
    XRAM[20591] = 8'b0;
    XRAM[20592] = 8'b0;
    XRAM[20593] = 8'b0;
    XRAM[20594] = 8'b0;
    XRAM[20595] = 8'b0;
    XRAM[20596] = 8'b0;
    XRAM[20597] = 8'b0;
    XRAM[20598] = 8'b0;
    XRAM[20599] = 8'b0;
    XRAM[20600] = 8'b0;
    XRAM[20601] = 8'b0;
    XRAM[20602] = 8'b0;
    XRAM[20603] = 8'b0;
    XRAM[20604] = 8'b0;
    XRAM[20605] = 8'b0;
    XRAM[20606] = 8'b0;
    XRAM[20607] = 8'b0;
    XRAM[20608] = 8'b0;
    XRAM[20609] = 8'b0;
    XRAM[20610] = 8'b0;
    XRAM[20611] = 8'b0;
    XRAM[20612] = 8'b0;
    XRAM[20613] = 8'b0;
    XRAM[20614] = 8'b0;
    XRAM[20615] = 8'b0;
    XRAM[20616] = 8'b0;
    XRAM[20617] = 8'b0;
    XRAM[20618] = 8'b0;
    XRAM[20619] = 8'b0;
    XRAM[20620] = 8'b0;
    XRAM[20621] = 8'b0;
    XRAM[20622] = 8'b0;
    XRAM[20623] = 8'b0;
    XRAM[20624] = 8'b0;
    XRAM[20625] = 8'b0;
    XRAM[20626] = 8'b0;
    XRAM[20627] = 8'b0;
    XRAM[20628] = 8'b0;
    XRAM[20629] = 8'b0;
    XRAM[20630] = 8'b0;
    XRAM[20631] = 8'b0;
    XRAM[20632] = 8'b0;
    XRAM[20633] = 8'b0;
    XRAM[20634] = 8'b0;
    XRAM[20635] = 8'b0;
    XRAM[20636] = 8'b0;
    XRAM[20637] = 8'b0;
    XRAM[20638] = 8'b0;
    XRAM[20639] = 8'b0;
    XRAM[20640] = 8'b0;
    XRAM[20641] = 8'b0;
    XRAM[20642] = 8'b0;
    XRAM[20643] = 8'b0;
    XRAM[20644] = 8'b0;
    XRAM[20645] = 8'b0;
    XRAM[20646] = 8'b0;
    XRAM[20647] = 8'b0;
    XRAM[20648] = 8'b0;
    XRAM[20649] = 8'b0;
    XRAM[20650] = 8'b0;
    XRAM[20651] = 8'b0;
    XRAM[20652] = 8'b0;
    XRAM[20653] = 8'b0;
    XRAM[20654] = 8'b0;
    XRAM[20655] = 8'b0;
    XRAM[20656] = 8'b0;
    XRAM[20657] = 8'b0;
    XRAM[20658] = 8'b0;
    XRAM[20659] = 8'b0;
    XRAM[20660] = 8'b0;
    XRAM[20661] = 8'b0;
    XRAM[20662] = 8'b0;
    XRAM[20663] = 8'b0;
    XRAM[20664] = 8'b0;
    XRAM[20665] = 8'b0;
    XRAM[20666] = 8'b0;
    XRAM[20667] = 8'b0;
    XRAM[20668] = 8'b0;
    XRAM[20669] = 8'b0;
    XRAM[20670] = 8'b0;
    XRAM[20671] = 8'b0;
    XRAM[20672] = 8'b0;
    XRAM[20673] = 8'b0;
    XRAM[20674] = 8'b0;
    XRAM[20675] = 8'b0;
    XRAM[20676] = 8'b0;
    XRAM[20677] = 8'b0;
    XRAM[20678] = 8'b0;
    XRAM[20679] = 8'b0;
    XRAM[20680] = 8'b0;
    XRAM[20681] = 8'b0;
    XRAM[20682] = 8'b0;
    XRAM[20683] = 8'b0;
    XRAM[20684] = 8'b0;
    XRAM[20685] = 8'b0;
    XRAM[20686] = 8'b0;
    XRAM[20687] = 8'b0;
    XRAM[20688] = 8'b0;
    XRAM[20689] = 8'b0;
    XRAM[20690] = 8'b0;
    XRAM[20691] = 8'b0;
    XRAM[20692] = 8'b0;
    XRAM[20693] = 8'b0;
    XRAM[20694] = 8'b0;
    XRAM[20695] = 8'b0;
    XRAM[20696] = 8'b0;
    XRAM[20697] = 8'b0;
    XRAM[20698] = 8'b0;
    XRAM[20699] = 8'b0;
    XRAM[20700] = 8'b0;
    XRAM[20701] = 8'b0;
    XRAM[20702] = 8'b0;
    XRAM[20703] = 8'b0;
    XRAM[20704] = 8'b0;
    XRAM[20705] = 8'b0;
    XRAM[20706] = 8'b0;
    XRAM[20707] = 8'b0;
    XRAM[20708] = 8'b0;
    XRAM[20709] = 8'b0;
    XRAM[20710] = 8'b0;
    XRAM[20711] = 8'b0;
    XRAM[20712] = 8'b0;
    XRAM[20713] = 8'b0;
    XRAM[20714] = 8'b0;
    XRAM[20715] = 8'b0;
    XRAM[20716] = 8'b0;
    XRAM[20717] = 8'b0;
    XRAM[20718] = 8'b0;
    XRAM[20719] = 8'b0;
    XRAM[20720] = 8'b0;
    XRAM[20721] = 8'b0;
    XRAM[20722] = 8'b0;
    XRAM[20723] = 8'b0;
    XRAM[20724] = 8'b0;
    XRAM[20725] = 8'b0;
    XRAM[20726] = 8'b0;
    XRAM[20727] = 8'b0;
    XRAM[20728] = 8'b0;
    XRAM[20729] = 8'b0;
    XRAM[20730] = 8'b0;
    XRAM[20731] = 8'b0;
    XRAM[20732] = 8'b0;
    XRAM[20733] = 8'b0;
    XRAM[20734] = 8'b0;
    XRAM[20735] = 8'b0;
    XRAM[20736] = 8'b0;
    XRAM[20737] = 8'b0;
    XRAM[20738] = 8'b0;
    XRAM[20739] = 8'b0;
    XRAM[20740] = 8'b0;
    XRAM[20741] = 8'b0;
    XRAM[20742] = 8'b0;
    XRAM[20743] = 8'b0;
    XRAM[20744] = 8'b0;
    XRAM[20745] = 8'b0;
    XRAM[20746] = 8'b0;
    XRAM[20747] = 8'b0;
    XRAM[20748] = 8'b0;
    XRAM[20749] = 8'b0;
    XRAM[20750] = 8'b0;
    XRAM[20751] = 8'b0;
    XRAM[20752] = 8'b0;
    XRAM[20753] = 8'b0;
    XRAM[20754] = 8'b0;
    XRAM[20755] = 8'b0;
    XRAM[20756] = 8'b0;
    XRAM[20757] = 8'b0;
    XRAM[20758] = 8'b0;
    XRAM[20759] = 8'b0;
    XRAM[20760] = 8'b0;
    XRAM[20761] = 8'b0;
    XRAM[20762] = 8'b0;
    XRAM[20763] = 8'b0;
    XRAM[20764] = 8'b0;
    XRAM[20765] = 8'b0;
    XRAM[20766] = 8'b0;
    XRAM[20767] = 8'b0;
    XRAM[20768] = 8'b0;
    XRAM[20769] = 8'b0;
    XRAM[20770] = 8'b0;
    XRAM[20771] = 8'b0;
    XRAM[20772] = 8'b0;
    XRAM[20773] = 8'b0;
    XRAM[20774] = 8'b0;
    XRAM[20775] = 8'b0;
    XRAM[20776] = 8'b0;
    XRAM[20777] = 8'b0;
    XRAM[20778] = 8'b0;
    XRAM[20779] = 8'b0;
    XRAM[20780] = 8'b0;
    XRAM[20781] = 8'b0;
    XRAM[20782] = 8'b0;
    XRAM[20783] = 8'b0;
    XRAM[20784] = 8'b0;
    XRAM[20785] = 8'b0;
    XRAM[20786] = 8'b0;
    XRAM[20787] = 8'b0;
    XRAM[20788] = 8'b0;
    XRAM[20789] = 8'b0;
    XRAM[20790] = 8'b0;
    XRAM[20791] = 8'b0;
    XRAM[20792] = 8'b0;
    XRAM[20793] = 8'b0;
    XRAM[20794] = 8'b0;
    XRAM[20795] = 8'b0;
    XRAM[20796] = 8'b0;
    XRAM[20797] = 8'b0;
    XRAM[20798] = 8'b0;
    XRAM[20799] = 8'b0;
    XRAM[20800] = 8'b0;
    XRAM[20801] = 8'b0;
    XRAM[20802] = 8'b0;
    XRAM[20803] = 8'b0;
    XRAM[20804] = 8'b0;
    XRAM[20805] = 8'b0;
    XRAM[20806] = 8'b0;
    XRAM[20807] = 8'b0;
    XRAM[20808] = 8'b0;
    XRAM[20809] = 8'b0;
    XRAM[20810] = 8'b0;
    XRAM[20811] = 8'b0;
    XRAM[20812] = 8'b0;
    XRAM[20813] = 8'b0;
    XRAM[20814] = 8'b0;
    XRAM[20815] = 8'b0;
    XRAM[20816] = 8'b0;
    XRAM[20817] = 8'b0;
    XRAM[20818] = 8'b0;
    XRAM[20819] = 8'b0;
    XRAM[20820] = 8'b0;
    XRAM[20821] = 8'b0;
    XRAM[20822] = 8'b0;
    XRAM[20823] = 8'b0;
    XRAM[20824] = 8'b0;
    XRAM[20825] = 8'b0;
    XRAM[20826] = 8'b0;
    XRAM[20827] = 8'b0;
    XRAM[20828] = 8'b0;
    XRAM[20829] = 8'b0;
    XRAM[20830] = 8'b0;
    XRAM[20831] = 8'b0;
    XRAM[20832] = 8'b0;
    XRAM[20833] = 8'b0;
    XRAM[20834] = 8'b0;
    XRAM[20835] = 8'b0;
    XRAM[20836] = 8'b0;
    XRAM[20837] = 8'b0;
    XRAM[20838] = 8'b0;
    XRAM[20839] = 8'b0;
    XRAM[20840] = 8'b0;
    XRAM[20841] = 8'b0;
    XRAM[20842] = 8'b0;
    XRAM[20843] = 8'b0;
    XRAM[20844] = 8'b0;
    XRAM[20845] = 8'b0;
    XRAM[20846] = 8'b0;
    XRAM[20847] = 8'b0;
    XRAM[20848] = 8'b0;
    XRAM[20849] = 8'b0;
    XRAM[20850] = 8'b0;
    XRAM[20851] = 8'b0;
    XRAM[20852] = 8'b0;
    XRAM[20853] = 8'b0;
    XRAM[20854] = 8'b0;
    XRAM[20855] = 8'b0;
    XRAM[20856] = 8'b0;
    XRAM[20857] = 8'b0;
    XRAM[20858] = 8'b0;
    XRAM[20859] = 8'b0;
    XRAM[20860] = 8'b0;
    XRAM[20861] = 8'b0;
    XRAM[20862] = 8'b0;
    XRAM[20863] = 8'b0;
    XRAM[20864] = 8'b0;
    XRAM[20865] = 8'b0;
    XRAM[20866] = 8'b0;
    XRAM[20867] = 8'b0;
    XRAM[20868] = 8'b0;
    XRAM[20869] = 8'b0;
    XRAM[20870] = 8'b0;
    XRAM[20871] = 8'b0;
    XRAM[20872] = 8'b0;
    XRAM[20873] = 8'b0;
    XRAM[20874] = 8'b0;
    XRAM[20875] = 8'b0;
    XRAM[20876] = 8'b0;
    XRAM[20877] = 8'b0;
    XRAM[20878] = 8'b0;
    XRAM[20879] = 8'b0;
    XRAM[20880] = 8'b0;
    XRAM[20881] = 8'b0;
    XRAM[20882] = 8'b0;
    XRAM[20883] = 8'b0;
    XRAM[20884] = 8'b0;
    XRAM[20885] = 8'b0;
    XRAM[20886] = 8'b0;
    XRAM[20887] = 8'b0;
    XRAM[20888] = 8'b0;
    XRAM[20889] = 8'b0;
    XRAM[20890] = 8'b0;
    XRAM[20891] = 8'b0;
    XRAM[20892] = 8'b0;
    XRAM[20893] = 8'b0;
    XRAM[20894] = 8'b0;
    XRAM[20895] = 8'b0;
    XRAM[20896] = 8'b0;
    XRAM[20897] = 8'b0;
    XRAM[20898] = 8'b0;
    XRAM[20899] = 8'b0;
    XRAM[20900] = 8'b0;
    XRAM[20901] = 8'b0;
    XRAM[20902] = 8'b0;
    XRAM[20903] = 8'b0;
    XRAM[20904] = 8'b0;
    XRAM[20905] = 8'b0;
    XRAM[20906] = 8'b0;
    XRAM[20907] = 8'b0;
    XRAM[20908] = 8'b0;
    XRAM[20909] = 8'b0;
    XRAM[20910] = 8'b0;
    XRAM[20911] = 8'b0;
    XRAM[20912] = 8'b0;
    XRAM[20913] = 8'b0;
    XRAM[20914] = 8'b0;
    XRAM[20915] = 8'b0;
    XRAM[20916] = 8'b0;
    XRAM[20917] = 8'b0;
    XRAM[20918] = 8'b0;
    XRAM[20919] = 8'b0;
    XRAM[20920] = 8'b0;
    XRAM[20921] = 8'b0;
    XRAM[20922] = 8'b0;
    XRAM[20923] = 8'b0;
    XRAM[20924] = 8'b0;
    XRAM[20925] = 8'b0;
    XRAM[20926] = 8'b0;
    XRAM[20927] = 8'b0;
    XRAM[20928] = 8'b0;
    XRAM[20929] = 8'b0;
    XRAM[20930] = 8'b0;
    XRAM[20931] = 8'b0;
    XRAM[20932] = 8'b0;
    XRAM[20933] = 8'b0;
    XRAM[20934] = 8'b0;
    XRAM[20935] = 8'b0;
    XRAM[20936] = 8'b0;
    XRAM[20937] = 8'b0;
    XRAM[20938] = 8'b0;
    XRAM[20939] = 8'b0;
    XRAM[20940] = 8'b0;
    XRAM[20941] = 8'b0;
    XRAM[20942] = 8'b0;
    XRAM[20943] = 8'b0;
    XRAM[20944] = 8'b0;
    XRAM[20945] = 8'b0;
    XRAM[20946] = 8'b0;
    XRAM[20947] = 8'b0;
    XRAM[20948] = 8'b0;
    XRAM[20949] = 8'b0;
    XRAM[20950] = 8'b0;
    XRAM[20951] = 8'b0;
    XRAM[20952] = 8'b0;
    XRAM[20953] = 8'b0;
    XRAM[20954] = 8'b0;
    XRAM[20955] = 8'b0;
    XRAM[20956] = 8'b0;
    XRAM[20957] = 8'b0;
    XRAM[20958] = 8'b0;
    XRAM[20959] = 8'b0;
    XRAM[20960] = 8'b0;
    XRAM[20961] = 8'b0;
    XRAM[20962] = 8'b0;
    XRAM[20963] = 8'b0;
    XRAM[20964] = 8'b0;
    XRAM[20965] = 8'b0;
    XRAM[20966] = 8'b0;
    XRAM[20967] = 8'b0;
    XRAM[20968] = 8'b0;
    XRAM[20969] = 8'b0;
    XRAM[20970] = 8'b0;
    XRAM[20971] = 8'b0;
    XRAM[20972] = 8'b0;
    XRAM[20973] = 8'b0;
    XRAM[20974] = 8'b0;
    XRAM[20975] = 8'b0;
    XRAM[20976] = 8'b0;
    XRAM[20977] = 8'b0;
    XRAM[20978] = 8'b0;
    XRAM[20979] = 8'b0;
    XRAM[20980] = 8'b0;
    XRAM[20981] = 8'b0;
    XRAM[20982] = 8'b0;
    XRAM[20983] = 8'b0;
    XRAM[20984] = 8'b0;
    XRAM[20985] = 8'b0;
    XRAM[20986] = 8'b0;
    XRAM[20987] = 8'b0;
    XRAM[20988] = 8'b0;
    XRAM[20989] = 8'b0;
    XRAM[20990] = 8'b0;
    XRAM[20991] = 8'b0;
    XRAM[20992] = 8'b0;
    XRAM[20993] = 8'b0;
    XRAM[20994] = 8'b0;
    XRAM[20995] = 8'b0;
    XRAM[20996] = 8'b0;
    XRAM[20997] = 8'b0;
    XRAM[20998] = 8'b0;
    XRAM[20999] = 8'b0;
    XRAM[21000] = 8'b0;
    XRAM[21001] = 8'b0;
    XRAM[21002] = 8'b0;
    XRAM[21003] = 8'b0;
    XRAM[21004] = 8'b0;
    XRAM[21005] = 8'b0;
    XRAM[21006] = 8'b0;
    XRAM[21007] = 8'b0;
    XRAM[21008] = 8'b0;
    XRAM[21009] = 8'b0;
    XRAM[21010] = 8'b0;
    XRAM[21011] = 8'b0;
    XRAM[21012] = 8'b0;
    XRAM[21013] = 8'b0;
    XRAM[21014] = 8'b0;
    XRAM[21015] = 8'b0;
    XRAM[21016] = 8'b0;
    XRAM[21017] = 8'b0;
    XRAM[21018] = 8'b0;
    XRAM[21019] = 8'b0;
    XRAM[21020] = 8'b0;
    XRAM[21021] = 8'b0;
    XRAM[21022] = 8'b0;
    XRAM[21023] = 8'b0;
    XRAM[21024] = 8'b0;
    XRAM[21025] = 8'b0;
    XRAM[21026] = 8'b0;
    XRAM[21027] = 8'b0;
    XRAM[21028] = 8'b0;
    XRAM[21029] = 8'b0;
    XRAM[21030] = 8'b0;
    XRAM[21031] = 8'b0;
    XRAM[21032] = 8'b0;
    XRAM[21033] = 8'b0;
    XRAM[21034] = 8'b0;
    XRAM[21035] = 8'b0;
    XRAM[21036] = 8'b0;
    XRAM[21037] = 8'b0;
    XRAM[21038] = 8'b0;
    XRAM[21039] = 8'b0;
    XRAM[21040] = 8'b0;
    XRAM[21041] = 8'b0;
    XRAM[21042] = 8'b0;
    XRAM[21043] = 8'b0;
    XRAM[21044] = 8'b0;
    XRAM[21045] = 8'b0;
    XRAM[21046] = 8'b0;
    XRAM[21047] = 8'b0;
    XRAM[21048] = 8'b0;
    XRAM[21049] = 8'b0;
    XRAM[21050] = 8'b0;
    XRAM[21051] = 8'b0;
    XRAM[21052] = 8'b0;
    XRAM[21053] = 8'b0;
    XRAM[21054] = 8'b0;
    XRAM[21055] = 8'b0;
    XRAM[21056] = 8'b0;
    XRAM[21057] = 8'b0;
    XRAM[21058] = 8'b0;
    XRAM[21059] = 8'b0;
    XRAM[21060] = 8'b0;
    XRAM[21061] = 8'b0;
    XRAM[21062] = 8'b0;
    XRAM[21063] = 8'b0;
    XRAM[21064] = 8'b0;
    XRAM[21065] = 8'b0;
    XRAM[21066] = 8'b0;
    XRAM[21067] = 8'b0;
    XRAM[21068] = 8'b0;
    XRAM[21069] = 8'b0;
    XRAM[21070] = 8'b0;
    XRAM[21071] = 8'b0;
    XRAM[21072] = 8'b0;
    XRAM[21073] = 8'b0;
    XRAM[21074] = 8'b0;
    XRAM[21075] = 8'b0;
    XRAM[21076] = 8'b0;
    XRAM[21077] = 8'b0;
    XRAM[21078] = 8'b0;
    XRAM[21079] = 8'b0;
    XRAM[21080] = 8'b0;
    XRAM[21081] = 8'b0;
    XRAM[21082] = 8'b0;
    XRAM[21083] = 8'b0;
    XRAM[21084] = 8'b0;
    XRAM[21085] = 8'b0;
    XRAM[21086] = 8'b0;
    XRAM[21087] = 8'b0;
    XRAM[21088] = 8'b0;
    XRAM[21089] = 8'b0;
    XRAM[21090] = 8'b0;
    XRAM[21091] = 8'b0;
    XRAM[21092] = 8'b0;
    XRAM[21093] = 8'b0;
    XRAM[21094] = 8'b0;
    XRAM[21095] = 8'b0;
    XRAM[21096] = 8'b0;
    XRAM[21097] = 8'b0;
    XRAM[21098] = 8'b0;
    XRAM[21099] = 8'b0;
    XRAM[21100] = 8'b0;
    XRAM[21101] = 8'b0;
    XRAM[21102] = 8'b0;
    XRAM[21103] = 8'b0;
    XRAM[21104] = 8'b0;
    XRAM[21105] = 8'b0;
    XRAM[21106] = 8'b0;
    XRAM[21107] = 8'b0;
    XRAM[21108] = 8'b0;
    XRAM[21109] = 8'b0;
    XRAM[21110] = 8'b0;
    XRAM[21111] = 8'b0;
    XRAM[21112] = 8'b0;
    XRAM[21113] = 8'b0;
    XRAM[21114] = 8'b0;
    XRAM[21115] = 8'b0;
    XRAM[21116] = 8'b0;
    XRAM[21117] = 8'b0;
    XRAM[21118] = 8'b0;
    XRAM[21119] = 8'b0;
    XRAM[21120] = 8'b0;
    XRAM[21121] = 8'b0;
    XRAM[21122] = 8'b0;
    XRAM[21123] = 8'b0;
    XRAM[21124] = 8'b0;
    XRAM[21125] = 8'b0;
    XRAM[21126] = 8'b0;
    XRAM[21127] = 8'b0;
    XRAM[21128] = 8'b0;
    XRAM[21129] = 8'b0;
    XRAM[21130] = 8'b0;
    XRAM[21131] = 8'b0;
    XRAM[21132] = 8'b0;
    XRAM[21133] = 8'b0;
    XRAM[21134] = 8'b0;
    XRAM[21135] = 8'b0;
    XRAM[21136] = 8'b0;
    XRAM[21137] = 8'b0;
    XRAM[21138] = 8'b0;
    XRAM[21139] = 8'b0;
    XRAM[21140] = 8'b0;
    XRAM[21141] = 8'b0;
    XRAM[21142] = 8'b0;
    XRAM[21143] = 8'b0;
    XRAM[21144] = 8'b0;
    XRAM[21145] = 8'b0;
    XRAM[21146] = 8'b0;
    XRAM[21147] = 8'b0;
    XRAM[21148] = 8'b0;
    XRAM[21149] = 8'b0;
    XRAM[21150] = 8'b0;
    XRAM[21151] = 8'b0;
    XRAM[21152] = 8'b0;
    XRAM[21153] = 8'b0;
    XRAM[21154] = 8'b0;
    XRAM[21155] = 8'b0;
    XRAM[21156] = 8'b0;
    XRAM[21157] = 8'b0;
    XRAM[21158] = 8'b0;
    XRAM[21159] = 8'b0;
    XRAM[21160] = 8'b0;
    XRAM[21161] = 8'b0;
    XRAM[21162] = 8'b0;
    XRAM[21163] = 8'b0;
    XRAM[21164] = 8'b0;
    XRAM[21165] = 8'b0;
    XRAM[21166] = 8'b0;
    XRAM[21167] = 8'b0;
    XRAM[21168] = 8'b0;
    XRAM[21169] = 8'b0;
    XRAM[21170] = 8'b0;
    XRAM[21171] = 8'b0;
    XRAM[21172] = 8'b0;
    XRAM[21173] = 8'b0;
    XRAM[21174] = 8'b0;
    XRAM[21175] = 8'b0;
    XRAM[21176] = 8'b0;
    XRAM[21177] = 8'b0;
    XRAM[21178] = 8'b0;
    XRAM[21179] = 8'b0;
    XRAM[21180] = 8'b0;
    XRAM[21181] = 8'b0;
    XRAM[21182] = 8'b0;
    XRAM[21183] = 8'b0;
    XRAM[21184] = 8'b0;
    XRAM[21185] = 8'b0;
    XRAM[21186] = 8'b0;
    XRAM[21187] = 8'b0;
    XRAM[21188] = 8'b0;
    XRAM[21189] = 8'b0;
    XRAM[21190] = 8'b0;
    XRAM[21191] = 8'b0;
    XRAM[21192] = 8'b0;
    XRAM[21193] = 8'b0;
    XRAM[21194] = 8'b0;
    XRAM[21195] = 8'b0;
    XRAM[21196] = 8'b0;
    XRAM[21197] = 8'b0;
    XRAM[21198] = 8'b0;
    XRAM[21199] = 8'b0;
    XRAM[21200] = 8'b0;
    XRAM[21201] = 8'b0;
    XRAM[21202] = 8'b0;
    XRAM[21203] = 8'b0;
    XRAM[21204] = 8'b0;
    XRAM[21205] = 8'b0;
    XRAM[21206] = 8'b0;
    XRAM[21207] = 8'b0;
    XRAM[21208] = 8'b0;
    XRAM[21209] = 8'b0;
    XRAM[21210] = 8'b0;
    XRAM[21211] = 8'b0;
    XRAM[21212] = 8'b0;
    XRAM[21213] = 8'b0;
    XRAM[21214] = 8'b0;
    XRAM[21215] = 8'b0;
    XRAM[21216] = 8'b0;
    XRAM[21217] = 8'b0;
    XRAM[21218] = 8'b0;
    XRAM[21219] = 8'b0;
    XRAM[21220] = 8'b0;
    XRAM[21221] = 8'b0;
    XRAM[21222] = 8'b0;
    XRAM[21223] = 8'b0;
    XRAM[21224] = 8'b0;
    XRAM[21225] = 8'b0;
    XRAM[21226] = 8'b0;
    XRAM[21227] = 8'b0;
    XRAM[21228] = 8'b0;
    XRAM[21229] = 8'b0;
    XRAM[21230] = 8'b0;
    XRAM[21231] = 8'b0;
    XRAM[21232] = 8'b0;
    XRAM[21233] = 8'b0;
    XRAM[21234] = 8'b0;
    XRAM[21235] = 8'b0;
    XRAM[21236] = 8'b0;
    XRAM[21237] = 8'b0;
    XRAM[21238] = 8'b0;
    XRAM[21239] = 8'b0;
    XRAM[21240] = 8'b0;
    XRAM[21241] = 8'b0;
    XRAM[21242] = 8'b0;
    XRAM[21243] = 8'b0;
    XRAM[21244] = 8'b0;
    XRAM[21245] = 8'b0;
    XRAM[21246] = 8'b0;
    XRAM[21247] = 8'b0;
    XRAM[21248] = 8'b0;
    XRAM[21249] = 8'b0;
    XRAM[21250] = 8'b0;
    XRAM[21251] = 8'b0;
    XRAM[21252] = 8'b0;
    XRAM[21253] = 8'b0;
    XRAM[21254] = 8'b0;
    XRAM[21255] = 8'b0;
    XRAM[21256] = 8'b0;
    XRAM[21257] = 8'b0;
    XRAM[21258] = 8'b0;
    XRAM[21259] = 8'b0;
    XRAM[21260] = 8'b0;
    XRAM[21261] = 8'b0;
    XRAM[21262] = 8'b0;
    XRAM[21263] = 8'b0;
    XRAM[21264] = 8'b0;
    XRAM[21265] = 8'b0;
    XRAM[21266] = 8'b0;
    XRAM[21267] = 8'b0;
    XRAM[21268] = 8'b0;
    XRAM[21269] = 8'b0;
    XRAM[21270] = 8'b0;
    XRAM[21271] = 8'b0;
    XRAM[21272] = 8'b0;
    XRAM[21273] = 8'b0;
    XRAM[21274] = 8'b0;
    XRAM[21275] = 8'b0;
    XRAM[21276] = 8'b0;
    XRAM[21277] = 8'b0;
    XRAM[21278] = 8'b0;
    XRAM[21279] = 8'b0;
    XRAM[21280] = 8'b0;
    XRAM[21281] = 8'b0;
    XRAM[21282] = 8'b0;
    XRAM[21283] = 8'b0;
    XRAM[21284] = 8'b0;
    XRAM[21285] = 8'b0;
    XRAM[21286] = 8'b0;
    XRAM[21287] = 8'b0;
    XRAM[21288] = 8'b0;
    XRAM[21289] = 8'b0;
    XRAM[21290] = 8'b0;
    XRAM[21291] = 8'b0;
    XRAM[21292] = 8'b0;
    XRAM[21293] = 8'b0;
    XRAM[21294] = 8'b0;
    XRAM[21295] = 8'b0;
    XRAM[21296] = 8'b0;
    XRAM[21297] = 8'b0;
    XRAM[21298] = 8'b0;
    XRAM[21299] = 8'b0;
    XRAM[21300] = 8'b0;
    XRAM[21301] = 8'b0;
    XRAM[21302] = 8'b0;
    XRAM[21303] = 8'b0;
    XRAM[21304] = 8'b0;
    XRAM[21305] = 8'b0;
    XRAM[21306] = 8'b0;
    XRAM[21307] = 8'b0;
    XRAM[21308] = 8'b0;
    XRAM[21309] = 8'b0;
    XRAM[21310] = 8'b0;
    XRAM[21311] = 8'b0;
    XRAM[21312] = 8'b0;
    XRAM[21313] = 8'b0;
    XRAM[21314] = 8'b0;
    XRAM[21315] = 8'b0;
    XRAM[21316] = 8'b0;
    XRAM[21317] = 8'b0;
    XRAM[21318] = 8'b0;
    XRAM[21319] = 8'b0;
    XRAM[21320] = 8'b0;
    XRAM[21321] = 8'b0;
    XRAM[21322] = 8'b0;
    XRAM[21323] = 8'b0;
    XRAM[21324] = 8'b0;
    XRAM[21325] = 8'b0;
    XRAM[21326] = 8'b0;
    XRAM[21327] = 8'b0;
    XRAM[21328] = 8'b0;
    XRAM[21329] = 8'b0;
    XRAM[21330] = 8'b0;
    XRAM[21331] = 8'b0;
    XRAM[21332] = 8'b0;
    XRAM[21333] = 8'b0;
    XRAM[21334] = 8'b0;
    XRAM[21335] = 8'b0;
    XRAM[21336] = 8'b0;
    XRAM[21337] = 8'b0;
    XRAM[21338] = 8'b0;
    XRAM[21339] = 8'b0;
    XRAM[21340] = 8'b0;
    XRAM[21341] = 8'b0;
    XRAM[21342] = 8'b0;
    XRAM[21343] = 8'b0;
    XRAM[21344] = 8'b0;
    XRAM[21345] = 8'b0;
    XRAM[21346] = 8'b0;
    XRAM[21347] = 8'b0;
    XRAM[21348] = 8'b0;
    XRAM[21349] = 8'b0;
    XRAM[21350] = 8'b0;
    XRAM[21351] = 8'b0;
    XRAM[21352] = 8'b0;
    XRAM[21353] = 8'b0;
    XRAM[21354] = 8'b0;
    XRAM[21355] = 8'b0;
    XRAM[21356] = 8'b0;
    XRAM[21357] = 8'b0;
    XRAM[21358] = 8'b0;
    XRAM[21359] = 8'b0;
    XRAM[21360] = 8'b0;
    XRAM[21361] = 8'b0;
    XRAM[21362] = 8'b0;
    XRAM[21363] = 8'b0;
    XRAM[21364] = 8'b0;
    XRAM[21365] = 8'b0;
    XRAM[21366] = 8'b0;
    XRAM[21367] = 8'b0;
    XRAM[21368] = 8'b0;
    XRAM[21369] = 8'b0;
    XRAM[21370] = 8'b0;
    XRAM[21371] = 8'b0;
    XRAM[21372] = 8'b0;
    XRAM[21373] = 8'b0;
    XRAM[21374] = 8'b0;
    XRAM[21375] = 8'b0;
    XRAM[21376] = 8'b0;
    XRAM[21377] = 8'b0;
    XRAM[21378] = 8'b0;
    XRAM[21379] = 8'b0;
    XRAM[21380] = 8'b0;
    XRAM[21381] = 8'b0;
    XRAM[21382] = 8'b0;
    XRAM[21383] = 8'b0;
    XRAM[21384] = 8'b0;
    XRAM[21385] = 8'b0;
    XRAM[21386] = 8'b0;
    XRAM[21387] = 8'b0;
    XRAM[21388] = 8'b0;
    XRAM[21389] = 8'b0;
    XRAM[21390] = 8'b0;
    XRAM[21391] = 8'b0;
    XRAM[21392] = 8'b0;
    XRAM[21393] = 8'b0;
    XRAM[21394] = 8'b0;
    XRAM[21395] = 8'b0;
    XRAM[21396] = 8'b0;
    XRAM[21397] = 8'b0;
    XRAM[21398] = 8'b0;
    XRAM[21399] = 8'b0;
    XRAM[21400] = 8'b0;
    XRAM[21401] = 8'b0;
    XRAM[21402] = 8'b0;
    XRAM[21403] = 8'b0;
    XRAM[21404] = 8'b0;
    XRAM[21405] = 8'b0;
    XRAM[21406] = 8'b0;
    XRAM[21407] = 8'b0;
    XRAM[21408] = 8'b0;
    XRAM[21409] = 8'b0;
    XRAM[21410] = 8'b0;
    XRAM[21411] = 8'b0;
    XRAM[21412] = 8'b0;
    XRAM[21413] = 8'b0;
    XRAM[21414] = 8'b0;
    XRAM[21415] = 8'b0;
    XRAM[21416] = 8'b0;
    XRAM[21417] = 8'b0;
    XRAM[21418] = 8'b0;
    XRAM[21419] = 8'b0;
    XRAM[21420] = 8'b0;
    XRAM[21421] = 8'b0;
    XRAM[21422] = 8'b0;
    XRAM[21423] = 8'b0;
    XRAM[21424] = 8'b0;
    XRAM[21425] = 8'b0;
    XRAM[21426] = 8'b0;
    XRAM[21427] = 8'b0;
    XRAM[21428] = 8'b0;
    XRAM[21429] = 8'b0;
    XRAM[21430] = 8'b0;
    XRAM[21431] = 8'b0;
    XRAM[21432] = 8'b0;
    XRAM[21433] = 8'b0;
    XRAM[21434] = 8'b0;
    XRAM[21435] = 8'b0;
    XRAM[21436] = 8'b0;
    XRAM[21437] = 8'b0;
    XRAM[21438] = 8'b0;
    XRAM[21439] = 8'b0;
    XRAM[21440] = 8'b0;
    XRAM[21441] = 8'b0;
    XRAM[21442] = 8'b0;
    XRAM[21443] = 8'b0;
    XRAM[21444] = 8'b0;
    XRAM[21445] = 8'b0;
    XRAM[21446] = 8'b0;
    XRAM[21447] = 8'b0;
    XRAM[21448] = 8'b0;
    XRAM[21449] = 8'b0;
    XRAM[21450] = 8'b0;
    XRAM[21451] = 8'b0;
    XRAM[21452] = 8'b0;
    XRAM[21453] = 8'b0;
    XRAM[21454] = 8'b0;
    XRAM[21455] = 8'b0;
    XRAM[21456] = 8'b0;
    XRAM[21457] = 8'b0;
    XRAM[21458] = 8'b0;
    XRAM[21459] = 8'b0;
    XRAM[21460] = 8'b0;
    XRAM[21461] = 8'b0;
    XRAM[21462] = 8'b0;
    XRAM[21463] = 8'b0;
    XRAM[21464] = 8'b0;
    XRAM[21465] = 8'b0;
    XRAM[21466] = 8'b0;
    XRAM[21467] = 8'b0;
    XRAM[21468] = 8'b0;
    XRAM[21469] = 8'b0;
    XRAM[21470] = 8'b0;
    XRAM[21471] = 8'b0;
    XRAM[21472] = 8'b0;
    XRAM[21473] = 8'b0;
    XRAM[21474] = 8'b0;
    XRAM[21475] = 8'b0;
    XRAM[21476] = 8'b0;
    XRAM[21477] = 8'b0;
    XRAM[21478] = 8'b0;
    XRAM[21479] = 8'b0;
    XRAM[21480] = 8'b0;
    XRAM[21481] = 8'b0;
    XRAM[21482] = 8'b0;
    XRAM[21483] = 8'b0;
    XRAM[21484] = 8'b0;
    XRAM[21485] = 8'b0;
    XRAM[21486] = 8'b0;
    XRAM[21487] = 8'b0;
    XRAM[21488] = 8'b0;
    XRAM[21489] = 8'b0;
    XRAM[21490] = 8'b0;
    XRAM[21491] = 8'b0;
    XRAM[21492] = 8'b0;
    XRAM[21493] = 8'b0;
    XRAM[21494] = 8'b0;
    XRAM[21495] = 8'b0;
    XRAM[21496] = 8'b0;
    XRAM[21497] = 8'b0;
    XRAM[21498] = 8'b0;
    XRAM[21499] = 8'b0;
    XRAM[21500] = 8'b0;
    XRAM[21501] = 8'b0;
    XRAM[21502] = 8'b0;
    XRAM[21503] = 8'b0;
    XRAM[21504] = 8'b0;
    XRAM[21505] = 8'b0;
    XRAM[21506] = 8'b0;
    XRAM[21507] = 8'b0;
    XRAM[21508] = 8'b0;
    XRAM[21509] = 8'b0;
    XRAM[21510] = 8'b0;
    XRAM[21511] = 8'b0;
    XRAM[21512] = 8'b0;
    XRAM[21513] = 8'b0;
    XRAM[21514] = 8'b0;
    XRAM[21515] = 8'b0;
    XRAM[21516] = 8'b0;
    XRAM[21517] = 8'b0;
    XRAM[21518] = 8'b0;
    XRAM[21519] = 8'b0;
    XRAM[21520] = 8'b0;
    XRAM[21521] = 8'b0;
    XRAM[21522] = 8'b0;
    XRAM[21523] = 8'b0;
    XRAM[21524] = 8'b0;
    XRAM[21525] = 8'b0;
    XRAM[21526] = 8'b0;
    XRAM[21527] = 8'b0;
    XRAM[21528] = 8'b0;
    XRAM[21529] = 8'b0;
    XRAM[21530] = 8'b0;
    XRAM[21531] = 8'b0;
    XRAM[21532] = 8'b0;
    XRAM[21533] = 8'b0;
    XRAM[21534] = 8'b0;
    XRAM[21535] = 8'b0;
    XRAM[21536] = 8'b0;
    XRAM[21537] = 8'b0;
    XRAM[21538] = 8'b0;
    XRAM[21539] = 8'b0;
    XRAM[21540] = 8'b0;
    XRAM[21541] = 8'b0;
    XRAM[21542] = 8'b0;
    XRAM[21543] = 8'b0;
    XRAM[21544] = 8'b0;
    XRAM[21545] = 8'b0;
    XRAM[21546] = 8'b0;
    XRAM[21547] = 8'b0;
    XRAM[21548] = 8'b0;
    XRAM[21549] = 8'b0;
    XRAM[21550] = 8'b0;
    XRAM[21551] = 8'b0;
    XRAM[21552] = 8'b0;
    XRAM[21553] = 8'b0;
    XRAM[21554] = 8'b0;
    XRAM[21555] = 8'b0;
    XRAM[21556] = 8'b0;
    XRAM[21557] = 8'b0;
    XRAM[21558] = 8'b0;
    XRAM[21559] = 8'b0;
    XRAM[21560] = 8'b0;
    XRAM[21561] = 8'b0;
    XRAM[21562] = 8'b0;
    XRAM[21563] = 8'b0;
    XRAM[21564] = 8'b0;
    XRAM[21565] = 8'b0;
    XRAM[21566] = 8'b0;
    XRAM[21567] = 8'b0;
    XRAM[21568] = 8'b0;
    XRAM[21569] = 8'b0;
    XRAM[21570] = 8'b0;
    XRAM[21571] = 8'b0;
    XRAM[21572] = 8'b0;
    XRAM[21573] = 8'b0;
    XRAM[21574] = 8'b0;
    XRAM[21575] = 8'b0;
    XRAM[21576] = 8'b0;
    XRAM[21577] = 8'b0;
    XRAM[21578] = 8'b0;
    XRAM[21579] = 8'b0;
    XRAM[21580] = 8'b0;
    XRAM[21581] = 8'b0;
    XRAM[21582] = 8'b0;
    XRAM[21583] = 8'b0;
    XRAM[21584] = 8'b0;
    XRAM[21585] = 8'b0;
    XRAM[21586] = 8'b0;
    XRAM[21587] = 8'b0;
    XRAM[21588] = 8'b0;
    XRAM[21589] = 8'b0;
    XRAM[21590] = 8'b0;
    XRAM[21591] = 8'b0;
    XRAM[21592] = 8'b0;
    XRAM[21593] = 8'b0;
    XRAM[21594] = 8'b0;
    XRAM[21595] = 8'b0;
    XRAM[21596] = 8'b0;
    XRAM[21597] = 8'b0;
    XRAM[21598] = 8'b0;
    XRAM[21599] = 8'b0;
    XRAM[21600] = 8'b0;
    XRAM[21601] = 8'b0;
    XRAM[21602] = 8'b0;
    XRAM[21603] = 8'b0;
    XRAM[21604] = 8'b0;
    XRAM[21605] = 8'b0;
    XRAM[21606] = 8'b0;
    XRAM[21607] = 8'b0;
    XRAM[21608] = 8'b0;
    XRAM[21609] = 8'b0;
    XRAM[21610] = 8'b0;
    XRAM[21611] = 8'b0;
    XRAM[21612] = 8'b0;
    XRAM[21613] = 8'b0;
    XRAM[21614] = 8'b0;
    XRAM[21615] = 8'b0;
    XRAM[21616] = 8'b0;
    XRAM[21617] = 8'b0;
    XRAM[21618] = 8'b0;
    XRAM[21619] = 8'b0;
    XRAM[21620] = 8'b0;
    XRAM[21621] = 8'b0;
    XRAM[21622] = 8'b0;
    XRAM[21623] = 8'b0;
    XRAM[21624] = 8'b0;
    XRAM[21625] = 8'b0;
    XRAM[21626] = 8'b0;
    XRAM[21627] = 8'b0;
    XRAM[21628] = 8'b0;
    XRAM[21629] = 8'b0;
    XRAM[21630] = 8'b0;
    XRAM[21631] = 8'b0;
    XRAM[21632] = 8'b0;
    XRAM[21633] = 8'b0;
    XRAM[21634] = 8'b0;
    XRAM[21635] = 8'b0;
    XRAM[21636] = 8'b0;
    XRAM[21637] = 8'b0;
    XRAM[21638] = 8'b0;
    XRAM[21639] = 8'b0;
    XRAM[21640] = 8'b0;
    XRAM[21641] = 8'b0;
    XRAM[21642] = 8'b0;
    XRAM[21643] = 8'b0;
    XRAM[21644] = 8'b0;
    XRAM[21645] = 8'b0;
    XRAM[21646] = 8'b0;
    XRAM[21647] = 8'b0;
    XRAM[21648] = 8'b0;
    XRAM[21649] = 8'b0;
    XRAM[21650] = 8'b0;
    XRAM[21651] = 8'b0;
    XRAM[21652] = 8'b0;
    XRAM[21653] = 8'b0;
    XRAM[21654] = 8'b0;
    XRAM[21655] = 8'b0;
    XRAM[21656] = 8'b0;
    XRAM[21657] = 8'b0;
    XRAM[21658] = 8'b0;
    XRAM[21659] = 8'b0;
    XRAM[21660] = 8'b0;
    XRAM[21661] = 8'b0;
    XRAM[21662] = 8'b0;
    XRAM[21663] = 8'b0;
    XRAM[21664] = 8'b0;
    XRAM[21665] = 8'b0;
    XRAM[21666] = 8'b0;
    XRAM[21667] = 8'b0;
    XRAM[21668] = 8'b0;
    XRAM[21669] = 8'b0;
    XRAM[21670] = 8'b0;
    XRAM[21671] = 8'b0;
    XRAM[21672] = 8'b0;
    XRAM[21673] = 8'b0;
    XRAM[21674] = 8'b0;
    XRAM[21675] = 8'b0;
    XRAM[21676] = 8'b0;
    XRAM[21677] = 8'b0;
    XRAM[21678] = 8'b0;
    XRAM[21679] = 8'b0;
    XRAM[21680] = 8'b0;
    XRAM[21681] = 8'b0;
    XRAM[21682] = 8'b0;
    XRAM[21683] = 8'b0;
    XRAM[21684] = 8'b0;
    XRAM[21685] = 8'b0;
    XRAM[21686] = 8'b0;
    XRAM[21687] = 8'b0;
    XRAM[21688] = 8'b0;
    XRAM[21689] = 8'b0;
    XRAM[21690] = 8'b0;
    XRAM[21691] = 8'b0;
    XRAM[21692] = 8'b0;
    XRAM[21693] = 8'b0;
    XRAM[21694] = 8'b0;
    XRAM[21695] = 8'b0;
    XRAM[21696] = 8'b0;
    XRAM[21697] = 8'b0;
    XRAM[21698] = 8'b0;
    XRAM[21699] = 8'b0;
    XRAM[21700] = 8'b0;
    XRAM[21701] = 8'b0;
    XRAM[21702] = 8'b0;
    XRAM[21703] = 8'b0;
    XRAM[21704] = 8'b0;
    XRAM[21705] = 8'b0;
    XRAM[21706] = 8'b0;
    XRAM[21707] = 8'b0;
    XRAM[21708] = 8'b0;
    XRAM[21709] = 8'b0;
    XRAM[21710] = 8'b0;
    XRAM[21711] = 8'b0;
    XRAM[21712] = 8'b0;
    XRAM[21713] = 8'b0;
    XRAM[21714] = 8'b0;
    XRAM[21715] = 8'b0;
    XRAM[21716] = 8'b0;
    XRAM[21717] = 8'b0;
    XRAM[21718] = 8'b0;
    XRAM[21719] = 8'b0;
    XRAM[21720] = 8'b0;
    XRAM[21721] = 8'b0;
    XRAM[21722] = 8'b0;
    XRAM[21723] = 8'b0;
    XRAM[21724] = 8'b0;
    XRAM[21725] = 8'b0;
    XRAM[21726] = 8'b0;
    XRAM[21727] = 8'b0;
    XRAM[21728] = 8'b0;
    XRAM[21729] = 8'b0;
    XRAM[21730] = 8'b0;
    XRAM[21731] = 8'b0;
    XRAM[21732] = 8'b0;
    XRAM[21733] = 8'b0;
    XRAM[21734] = 8'b0;
    XRAM[21735] = 8'b0;
    XRAM[21736] = 8'b0;
    XRAM[21737] = 8'b0;
    XRAM[21738] = 8'b0;
    XRAM[21739] = 8'b0;
    XRAM[21740] = 8'b0;
    XRAM[21741] = 8'b0;
    XRAM[21742] = 8'b0;
    XRAM[21743] = 8'b0;
    XRAM[21744] = 8'b0;
    XRAM[21745] = 8'b0;
    XRAM[21746] = 8'b0;
    XRAM[21747] = 8'b0;
    XRAM[21748] = 8'b0;
    XRAM[21749] = 8'b0;
    XRAM[21750] = 8'b0;
    XRAM[21751] = 8'b0;
    XRAM[21752] = 8'b0;
    XRAM[21753] = 8'b0;
    XRAM[21754] = 8'b0;
    XRAM[21755] = 8'b0;
    XRAM[21756] = 8'b0;
    XRAM[21757] = 8'b0;
    XRAM[21758] = 8'b0;
    XRAM[21759] = 8'b0;
    XRAM[21760] = 8'b0;
    XRAM[21761] = 8'b0;
    XRAM[21762] = 8'b0;
    XRAM[21763] = 8'b0;
    XRAM[21764] = 8'b0;
    XRAM[21765] = 8'b0;
    XRAM[21766] = 8'b0;
    XRAM[21767] = 8'b0;
    XRAM[21768] = 8'b0;
    XRAM[21769] = 8'b0;
    XRAM[21770] = 8'b0;
    XRAM[21771] = 8'b0;
    XRAM[21772] = 8'b0;
    XRAM[21773] = 8'b0;
    XRAM[21774] = 8'b0;
    XRAM[21775] = 8'b0;
    XRAM[21776] = 8'b0;
    XRAM[21777] = 8'b0;
    XRAM[21778] = 8'b0;
    XRAM[21779] = 8'b0;
    XRAM[21780] = 8'b0;
    XRAM[21781] = 8'b0;
    XRAM[21782] = 8'b0;
    XRAM[21783] = 8'b0;
    XRAM[21784] = 8'b0;
    XRAM[21785] = 8'b0;
    XRAM[21786] = 8'b0;
    XRAM[21787] = 8'b0;
    XRAM[21788] = 8'b0;
    XRAM[21789] = 8'b0;
    XRAM[21790] = 8'b0;
    XRAM[21791] = 8'b0;
    XRAM[21792] = 8'b0;
    XRAM[21793] = 8'b0;
    XRAM[21794] = 8'b0;
    XRAM[21795] = 8'b0;
    XRAM[21796] = 8'b0;
    XRAM[21797] = 8'b0;
    XRAM[21798] = 8'b0;
    XRAM[21799] = 8'b0;
    XRAM[21800] = 8'b0;
    XRAM[21801] = 8'b0;
    XRAM[21802] = 8'b0;
    XRAM[21803] = 8'b0;
    XRAM[21804] = 8'b0;
    XRAM[21805] = 8'b0;
    XRAM[21806] = 8'b0;
    XRAM[21807] = 8'b0;
    XRAM[21808] = 8'b0;
    XRAM[21809] = 8'b0;
    XRAM[21810] = 8'b0;
    XRAM[21811] = 8'b0;
    XRAM[21812] = 8'b0;
    XRAM[21813] = 8'b0;
    XRAM[21814] = 8'b0;
    XRAM[21815] = 8'b0;
    XRAM[21816] = 8'b0;
    XRAM[21817] = 8'b0;
    XRAM[21818] = 8'b0;
    XRAM[21819] = 8'b0;
    XRAM[21820] = 8'b0;
    XRAM[21821] = 8'b0;
    XRAM[21822] = 8'b0;
    XRAM[21823] = 8'b0;
    XRAM[21824] = 8'b0;
    XRAM[21825] = 8'b0;
    XRAM[21826] = 8'b0;
    XRAM[21827] = 8'b0;
    XRAM[21828] = 8'b0;
    XRAM[21829] = 8'b0;
    XRAM[21830] = 8'b0;
    XRAM[21831] = 8'b0;
    XRAM[21832] = 8'b0;
    XRAM[21833] = 8'b0;
    XRAM[21834] = 8'b0;
    XRAM[21835] = 8'b0;
    XRAM[21836] = 8'b0;
    XRAM[21837] = 8'b0;
    XRAM[21838] = 8'b0;
    XRAM[21839] = 8'b0;
    XRAM[21840] = 8'b0;
    XRAM[21841] = 8'b0;
    XRAM[21842] = 8'b0;
    XRAM[21843] = 8'b0;
    XRAM[21844] = 8'b0;
    XRAM[21845] = 8'b0;
    XRAM[21846] = 8'b0;
    XRAM[21847] = 8'b0;
    XRAM[21848] = 8'b0;
    XRAM[21849] = 8'b0;
    XRAM[21850] = 8'b0;
    XRAM[21851] = 8'b0;
    XRAM[21852] = 8'b0;
    XRAM[21853] = 8'b0;
    XRAM[21854] = 8'b0;
    XRAM[21855] = 8'b0;
    XRAM[21856] = 8'b0;
    XRAM[21857] = 8'b0;
    XRAM[21858] = 8'b0;
    XRAM[21859] = 8'b0;
    XRAM[21860] = 8'b0;
    XRAM[21861] = 8'b0;
    XRAM[21862] = 8'b0;
    XRAM[21863] = 8'b0;
    XRAM[21864] = 8'b0;
    XRAM[21865] = 8'b0;
    XRAM[21866] = 8'b0;
    XRAM[21867] = 8'b0;
    XRAM[21868] = 8'b0;
    XRAM[21869] = 8'b0;
    XRAM[21870] = 8'b0;
    XRAM[21871] = 8'b0;
    XRAM[21872] = 8'b0;
    XRAM[21873] = 8'b0;
    XRAM[21874] = 8'b0;
    XRAM[21875] = 8'b0;
    XRAM[21876] = 8'b0;
    XRAM[21877] = 8'b0;
    XRAM[21878] = 8'b0;
    XRAM[21879] = 8'b0;
    XRAM[21880] = 8'b0;
    XRAM[21881] = 8'b0;
    XRAM[21882] = 8'b0;
    XRAM[21883] = 8'b0;
    XRAM[21884] = 8'b0;
    XRAM[21885] = 8'b0;
    XRAM[21886] = 8'b0;
    XRAM[21887] = 8'b0;
    XRAM[21888] = 8'b0;
    XRAM[21889] = 8'b0;
    XRAM[21890] = 8'b0;
    XRAM[21891] = 8'b0;
    XRAM[21892] = 8'b0;
    XRAM[21893] = 8'b0;
    XRAM[21894] = 8'b0;
    XRAM[21895] = 8'b0;
    XRAM[21896] = 8'b0;
    XRAM[21897] = 8'b0;
    XRAM[21898] = 8'b0;
    XRAM[21899] = 8'b0;
    XRAM[21900] = 8'b0;
    XRAM[21901] = 8'b0;
    XRAM[21902] = 8'b0;
    XRAM[21903] = 8'b0;
    XRAM[21904] = 8'b0;
    XRAM[21905] = 8'b0;
    XRAM[21906] = 8'b0;
    XRAM[21907] = 8'b0;
    XRAM[21908] = 8'b0;
    XRAM[21909] = 8'b0;
    XRAM[21910] = 8'b0;
    XRAM[21911] = 8'b0;
    XRAM[21912] = 8'b0;
    XRAM[21913] = 8'b0;
    XRAM[21914] = 8'b0;
    XRAM[21915] = 8'b0;
    XRAM[21916] = 8'b0;
    XRAM[21917] = 8'b0;
    XRAM[21918] = 8'b0;
    XRAM[21919] = 8'b0;
    XRAM[21920] = 8'b0;
    XRAM[21921] = 8'b0;
    XRAM[21922] = 8'b0;
    XRAM[21923] = 8'b0;
    XRAM[21924] = 8'b0;
    XRAM[21925] = 8'b0;
    XRAM[21926] = 8'b0;
    XRAM[21927] = 8'b0;
    XRAM[21928] = 8'b0;
    XRAM[21929] = 8'b0;
    XRAM[21930] = 8'b0;
    XRAM[21931] = 8'b0;
    XRAM[21932] = 8'b0;
    XRAM[21933] = 8'b0;
    XRAM[21934] = 8'b0;
    XRAM[21935] = 8'b0;
    XRAM[21936] = 8'b0;
    XRAM[21937] = 8'b0;
    XRAM[21938] = 8'b0;
    XRAM[21939] = 8'b0;
    XRAM[21940] = 8'b0;
    XRAM[21941] = 8'b0;
    XRAM[21942] = 8'b0;
    XRAM[21943] = 8'b0;
    XRAM[21944] = 8'b0;
    XRAM[21945] = 8'b0;
    XRAM[21946] = 8'b0;
    XRAM[21947] = 8'b0;
    XRAM[21948] = 8'b0;
    XRAM[21949] = 8'b0;
    XRAM[21950] = 8'b0;
    XRAM[21951] = 8'b0;
    XRAM[21952] = 8'b0;
    XRAM[21953] = 8'b0;
    XRAM[21954] = 8'b0;
    XRAM[21955] = 8'b0;
    XRAM[21956] = 8'b0;
    XRAM[21957] = 8'b0;
    XRAM[21958] = 8'b0;
    XRAM[21959] = 8'b0;
    XRAM[21960] = 8'b0;
    XRAM[21961] = 8'b0;
    XRAM[21962] = 8'b0;
    XRAM[21963] = 8'b0;
    XRAM[21964] = 8'b0;
    XRAM[21965] = 8'b0;
    XRAM[21966] = 8'b0;
    XRAM[21967] = 8'b0;
    XRAM[21968] = 8'b0;
    XRAM[21969] = 8'b0;
    XRAM[21970] = 8'b0;
    XRAM[21971] = 8'b0;
    XRAM[21972] = 8'b0;
    XRAM[21973] = 8'b0;
    XRAM[21974] = 8'b0;
    XRAM[21975] = 8'b0;
    XRAM[21976] = 8'b0;
    XRAM[21977] = 8'b0;
    XRAM[21978] = 8'b0;
    XRAM[21979] = 8'b0;
    XRAM[21980] = 8'b0;
    XRAM[21981] = 8'b0;
    XRAM[21982] = 8'b0;
    XRAM[21983] = 8'b0;
    XRAM[21984] = 8'b0;
    XRAM[21985] = 8'b0;
    XRAM[21986] = 8'b0;
    XRAM[21987] = 8'b0;
    XRAM[21988] = 8'b0;
    XRAM[21989] = 8'b0;
    XRAM[21990] = 8'b0;
    XRAM[21991] = 8'b0;
    XRAM[21992] = 8'b0;
    XRAM[21993] = 8'b0;
    XRAM[21994] = 8'b0;
    XRAM[21995] = 8'b0;
    XRAM[21996] = 8'b0;
    XRAM[21997] = 8'b0;
    XRAM[21998] = 8'b0;
    XRAM[21999] = 8'b0;
    XRAM[22000] = 8'b0;
    XRAM[22001] = 8'b0;
    XRAM[22002] = 8'b0;
    XRAM[22003] = 8'b0;
    XRAM[22004] = 8'b0;
    XRAM[22005] = 8'b0;
    XRAM[22006] = 8'b0;
    XRAM[22007] = 8'b0;
    XRAM[22008] = 8'b0;
    XRAM[22009] = 8'b0;
    XRAM[22010] = 8'b0;
    XRAM[22011] = 8'b0;
    XRAM[22012] = 8'b0;
    XRAM[22013] = 8'b0;
    XRAM[22014] = 8'b0;
    XRAM[22015] = 8'b0;
    XRAM[22016] = 8'b0;
    XRAM[22017] = 8'b0;
    XRAM[22018] = 8'b0;
    XRAM[22019] = 8'b0;
    XRAM[22020] = 8'b0;
    XRAM[22021] = 8'b0;
    XRAM[22022] = 8'b0;
    XRAM[22023] = 8'b0;
    XRAM[22024] = 8'b0;
    XRAM[22025] = 8'b0;
    XRAM[22026] = 8'b0;
    XRAM[22027] = 8'b0;
    XRAM[22028] = 8'b0;
    XRAM[22029] = 8'b0;
    XRAM[22030] = 8'b0;
    XRAM[22031] = 8'b0;
    XRAM[22032] = 8'b0;
    XRAM[22033] = 8'b0;
    XRAM[22034] = 8'b0;
    XRAM[22035] = 8'b0;
    XRAM[22036] = 8'b0;
    XRAM[22037] = 8'b0;
    XRAM[22038] = 8'b0;
    XRAM[22039] = 8'b0;
    XRAM[22040] = 8'b0;
    XRAM[22041] = 8'b0;
    XRAM[22042] = 8'b0;
    XRAM[22043] = 8'b0;
    XRAM[22044] = 8'b0;
    XRAM[22045] = 8'b0;
    XRAM[22046] = 8'b0;
    XRAM[22047] = 8'b0;
    XRAM[22048] = 8'b0;
    XRAM[22049] = 8'b0;
    XRAM[22050] = 8'b0;
    XRAM[22051] = 8'b0;
    XRAM[22052] = 8'b0;
    XRAM[22053] = 8'b0;
    XRAM[22054] = 8'b0;
    XRAM[22055] = 8'b0;
    XRAM[22056] = 8'b0;
    XRAM[22057] = 8'b0;
    XRAM[22058] = 8'b0;
    XRAM[22059] = 8'b0;
    XRAM[22060] = 8'b0;
    XRAM[22061] = 8'b0;
    XRAM[22062] = 8'b0;
    XRAM[22063] = 8'b0;
    XRAM[22064] = 8'b0;
    XRAM[22065] = 8'b0;
    XRAM[22066] = 8'b0;
    XRAM[22067] = 8'b0;
    XRAM[22068] = 8'b0;
    XRAM[22069] = 8'b0;
    XRAM[22070] = 8'b0;
    XRAM[22071] = 8'b0;
    XRAM[22072] = 8'b0;
    XRAM[22073] = 8'b0;
    XRAM[22074] = 8'b0;
    XRAM[22075] = 8'b0;
    XRAM[22076] = 8'b0;
    XRAM[22077] = 8'b0;
    XRAM[22078] = 8'b0;
    XRAM[22079] = 8'b0;
    XRAM[22080] = 8'b0;
    XRAM[22081] = 8'b0;
    XRAM[22082] = 8'b0;
    XRAM[22083] = 8'b0;
    XRAM[22084] = 8'b0;
    XRAM[22085] = 8'b0;
    XRAM[22086] = 8'b0;
    XRAM[22087] = 8'b0;
    XRAM[22088] = 8'b0;
    XRAM[22089] = 8'b0;
    XRAM[22090] = 8'b0;
    XRAM[22091] = 8'b0;
    XRAM[22092] = 8'b0;
    XRAM[22093] = 8'b0;
    XRAM[22094] = 8'b0;
    XRAM[22095] = 8'b0;
    XRAM[22096] = 8'b0;
    XRAM[22097] = 8'b0;
    XRAM[22098] = 8'b0;
    XRAM[22099] = 8'b0;
    XRAM[22100] = 8'b0;
    XRAM[22101] = 8'b0;
    XRAM[22102] = 8'b0;
    XRAM[22103] = 8'b0;
    XRAM[22104] = 8'b0;
    XRAM[22105] = 8'b0;
    XRAM[22106] = 8'b0;
    XRAM[22107] = 8'b0;
    XRAM[22108] = 8'b0;
    XRAM[22109] = 8'b0;
    XRAM[22110] = 8'b0;
    XRAM[22111] = 8'b0;
    XRAM[22112] = 8'b0;
    XRAM[22113] = 8'b0;
    XRAM[22114] = 8'b0;
    XRAM[22115] = 8'b0;
    XRAM[22116] = 8'b0;
    XRAM[22117] = 8'b0;
    XRAM[22118] = 8'b0;
    XRAM[22119] = 8'b0;
    XRAM[22120] = 8'b0;
    XRAM[22121] = 8'b0;
    XRAM[22122] = 8'b0;
    XRAM[22123] = 8'b0;
    XRAM[22124] = 8'b0;
    XRAM[22125] = 8'b0;
    XRAM[22126] = 8'b0;
    XRAM[22127] = 8'b0;
    XRAM[22128] = 8'b0;
    XRAM[22129] = 8'b0;
    XRAM[22130] = 8'b0;
    XRAM[22131] = 8'b0;
    XRAM[22132] = 8'b0;
    XRAM[22133] = 8'b0;
    XRAM[22134] = 8'b0;
    XRAM[22135] = 8'b0;
    XRAM[22136] = 8'b0;
    XRAM[22137] = 8'b0;
    XRAM[22138] = 8'b0;
    XRAM[22139] = 8'b0;
    XRAM[22140] = 8'b0;
    XRAM[22141] = 8'b0;
    XRAM[22142] = 8'b0;
    XRAM[22143] = 8'b0;
    XRAM[22144] = 8'b0;
    XRAM[22145] = 8'b0;
    XRAM[22146] = 8'b0;
    XRAM[22147] = 8'b0;
    XRAM[22148] = 8'b0;
    XRAM[22149] = 8'b0;
    XRAM[22150] = 8'b0;
    XRAM[22151] = 8'b0;
    XRAM[22152] = 8'b0;
    XRAM[22153] = 8'b0;
    XRAM[22154] = 8'b0;
    XRAM[22155] = 8'b0;
    XRAM[22156] = 8'b0;
    XRAM[22157] = 8'b0;
    XRAM[22158] = 8'b0;
    XRAM[22159] = 8'b0;
    XRAM[22160] = 8'b0;
    XRAM[22161] = 8'b0;
    XRAM[22162] = 8'b0;
    XRAM[22163] = 8'b0;
    XRAM[22164] = 8'b0;
    XRAM[22165] = 8'b0;
    XRAM[22166] = 8'b0;
    XRAM[22167] = 8'b0;
    XRAM[22168] = 8'b0;
    XRAM[22169] = 8'b0;
    XRAM[22170] = 8'b0;
    XRAM[22171] = 8'b0;
    XRAM[22172] = 8'b0;
    XRAM[22173] = 8'b0;
    XRAM[22174] = 8'b0;
    XRAM[22175] = 8'b0;
    XRAM[22176] = 8'b0;
    XRAM[22177] = 8'b0;
    XRAM[22178] = 8'b0;
    XRAM[22179] = 8'b0;
    XRAM[22180] = 8'b0;
    XRAM[22181] = 8'b0;
    XRAM[22182] = 8'b0;
    XRAM[22183] = 8'b0;
    XRAM[22184] = 8'b0;
    XRAM[22185] = 8'b0;
    XRAM[22186] = 8'b0;
    XRAM[22187] = 8'b0;
    XRAM[22188] = 8'b0;
    XRAM[22189] = 8'b0;
    XRAM[22190] = 8'b0;
    XRAM[22191] = 8'b0;
    XRAM[22192] = 8'b0;
    XRAM[22193] = 8'b0;
    XRAM[22194] = 8'b0;
    XRAM[22195] = 8'b0;
    XRAM[22196] = 8'b0;
    XRAM[22197] = 8'b0;
    XRAM[22198] = 8'b0;
    XRAM[22199] = 8'b0;
    XRAM[22200] = 8'b0;
    XRAM[22201] = 8'b0;
    XRAM[22202] = 8'b0;
    XRAM[22203] = 8'b0;
    XRAM[22204] = 8'b0;
    XRAM[22205] = 8'b0;
    XRAM[22206] = 8'b0;
    XRAM[22207] = 8'b0;
    XRAM[22208] = 8'b0;
    XRAM[22209] = 8'b0;
    XRAM[22210] = 8'b0;
    XRAM[22211] = 8'b0;
    XRAM[22212] = 8'b0;
    XRAM[22213] = 8'b0;
    XRAM[22214] = 8'b0;
    XRAM[22215] = 8'b0;
    XRAM[22216] = 8'b0;
    XRAM[22217] = 8'b0;
    XRAM[22218] = 8'b0;
    XRAM[22219] = 8'b0;
    XRAM[22220] = 8'b0;
    XRAM[22221] = 8'b0;
    XRAM[22222] = 8'b0;
    XRAM[22223] = 8'b0;
    XRAM[22224] = 8'b0;
    XRAM[22225] = 8'b0;
    XRAM[22226] = 8'b0;
    XRAM[22227] = 8'b0;
    XRAM[22228] = 8'b0;
    XRAM[22229] = 8'b0;
    XRAM[22230] = 8'b0;
    XRAM[22231] = 8'b0;
    XRAM[22232] = 8'b0;
    XRAM[22233] = 8'b0;
    XRAM[22234] = 8'b0;
    XRAM[22235] = 8'b0;
    XRAM[22236] = 8'b0;
    XRAM[22237] = 8'b0;
    XRAM[22238] = 8'b0;
    XRAM[22239] = 8'b0;
    XRAM[22240] = 8'b0;
    XRAM[22241] = 8'b0;
    XRAM[22242] = 8'b0;
    XRAM[22243] = 8'b0;
    XRAM[22244] = 8'b0;
    XRAM[22245] = 8'b0;
    XRAM[22246] = 8'b0;
    XRAM[22247] = 8'b0;
    XRAM[22248] = 8'b0;
    XRAM[22249] = 8'b0;
    XRAM[22250] = 8'b0;
    XRAM[22251] = 8'b0;
    XRAM[22252] = 8'b0;
    XRAM[22253] = 8'b0;
    XRAM[22254] = 8'b0;
    XRAM[22255] = 8'b0;
    XRAM[22256] = 8'b0;
    XRAM[22257] = 8'b0;
    XRAM[22258] = 8'b0;
    XRAM[22259] = 8'b0;
    XRAM[22260] = 8'b0;
    XRAM[22261] = 8'b0;
    XRAM[22262] = 8'b0;
    XRAM[22263] = 8'b0;
    XRAM[22264] = 8'b0;
    XRAM[22265] = 8'b0;
    XRAM[22266] = 8'b0;
    XRAM[22267] = 8'b0;
    XRAM[22268] = 8'b0;
    XRAM[22269] = 8'b0;
    XRAM[22270] = 8'b0;
    XRAM[22271] = 8'b0;
    XRAM[22272] = 8'b0;
    XRAM[22273] = 8'b0;
    XRAM[22274] = 8'b0;
    XRAM[22275] = 8'b0;
    XRAM[22276] = 8'b0;
    XRAM[22277] = 8'b0;
    XRAM[22278] = 8'b0;
    XRAM[22279] = 8'b0;
    XRAM[22280] = 8'b0;
    XRAM[22281] = 8'b0;
    XRAM[22282] = 8'b0;
    XRAM[22283] = 8'b0;
    XRAM[22284] = 8'b0;
    XRAM[22285] = 8'b0;
    XRAM[22286] = 8'b0;
    XRAM[22287] = 8'b0;
    XRAM[22288] = 8'b0;
    XRAM[22289] = 8'b0;
    XRAM[22290] = 8'b0;
    XRAM[22291] = 8'b0;
    XRAM[22292] = 8'b0;
    XRAM[22293] = 8'b0;
    XRAM[22294] = 8'b0;
    XRAM[22295] = 8'b0;
    XRAM[22296] = 8'b0;
    XRAM[22297] = 8'b0;
    XRAM[22298] = 8'b0;
    XRAM[22299] = 8'b0;
    XRAM[22300] = 8'b0;
    XRAM[22301] = 8'b0;
    XRAM[22302] = 8'b0;
    XRAM[22303] = 8'b0;
    XRAM[22304] = 8'b0;
    XRAM[22305] = 8'b0;
    XRAM[22306] = 8'b0;
    XRAM[22307] = 8'b0;
    XRAM[22308] = 8'b0;
    XRAM[22309] = 8'b0;
    XRAM[22310] = 8'b0;
    XRAM[22311] = 8'b0;
    XRAM[22312] = 8'b0;
    XRAM[22313] = 8'b0;
    XRAM[22314] = 8'b0;
    XRAM[22315] = 8'b0;
    XRAM[22316] = 8'b0;
    XRAM[22317] = 8'b0;
    XRAM[22318] = 8'b0;
    XRAM[22319] = 8'b0;
    XRAM[22320] = 8'b0;
    XRAM[22321] = 8'b0;
    XRAM[22322] = 8'b0;
    XRAM[22323] = 8'b0;
    XRAM[22324] = 8'b0;
    XRAM[22325] = 8'b0;
    XRAM[22326] = 8'b0;
    XRAM[22327] = 8'b0;
    XRAM[22328] = 8'b0;
    XRAM[22329] = 8'b0;
    XRAM[22330] = 8'b0;
    XRAM[22331] = 8'b0;
    XRAM[22332] = 8'b0;
    XRAM[22333] = 8'b0;
    XRAM[22334] = 8'b0;
    XRAM[22335] = 8'b0;
    XRAM[22336] = 8'b0;
    XRAM[22337] = 8'b0;
    XRAM[22338] = 8'b0;
    XRAM[22339] = 8'b0;
    XRAM[22340] = 8'b0;
    XRAM[22341] = 8'b0;
    XRAM[22342] = 8'b0;
    XRAM[22343] = 8'b0;
    XRAM[22344] = 8'b0;
    XRAM[22345] = 8'b0;
    XRAM[22346] = 8'b0;
    XRAM[22347] = 8'b0;
    XRAM[22348] = 8'b0;
    XRAM[22349] = 8'b0;
    XRAM[22350] = 8'b0;
    XRAM[22351] = 8'b0;
    XRAM[22352] = 8'b0;
    XRAM[22353] = 8'b0;
    XRAM[22354] = 8'b0;
    XRAM[22355] = 8'b0;
    XRAM[22356] = 8'b0;
    XRAM[22357] = 8'b0;
    XRAM[22358] = 8'b0;
    XRAM[22359] = 8'b0;
    XRAM[22360] = 8'b0;
    XRAM[22361] = 8'b0;
    XRAM[22362] = 8'b0;
    XRAM[22363] = 8'b0;
    XRAM[22364] = 8'b0;
    XRAM[22365] = 8'b0;
    XRAM[22366] = 8'b0;
    XRAM[22367] = 8'b0;
    XRAM[22368] = 8'b0;
    XRAM[22369] = 8'b0;
    XRAM[22370] = 8'b0;
    XRAM[22371] = 8'b0;
    XRAM[22372] = 8'b0;
    XRAM[22373] = 8'b0;
    XRAM[22374] = 8'b0;
    XRAM[22375] = 8'b0;
    XRAM[22376] = 8'b0;
    XRAM[22377] = 8'b0;
    XRAM[22378] = 8'b0;
    XRAM[22379] = 8'b0;
    XRAM[22380] = 8'b0;
    XRAM[22381] = 8'b0;
    XRAM[22382] = 8'b0;
    XRAM[22383] = 8'b0;
    XRAM[22384] = 8'b0;
    XRAM[22385] = 8'b0;
    XRAM[22386] = 8'b0;
    XRAM[22387] = 8'b0;
    XRAM[22388] = 8'b0;
    XRAM[22389] = 8'b0;
    XRAM[22390] = 8'b0;
    XRAM[22391] = 8'b0;
    XRAM[22392] = 8'b0;
    XRAM[22393] = 8'b0;
    XRAM[22394] = 8'b0;
    XRAM[22395] = 8'b0;
    XRAM[22396] = 8'b0;
    XRAM[22397] = 8'b0;
    XRAM[22398] = 8'b0;
    XRAM[22399] = 8'b0;
    XRAM[22400] = 8'b0;
    XRAM[22401] = 8'b0;
    XRAM[22402] = 8'b0;
    XRAM[22403] = 8'b0;
    XRAM[22404] = 8'b0;
    XRAM[22405] = 8'b0;
    XRAM[22406] = 8'b0;
    XRAM[22407] = 8'b0;
    XRAM[22408] = 8'b0;
    XRAM[22409] = 8'b0;
    XRAM[22410] = 8'b0;
    XRAM[22411] = 8'b0;
    XRAM[22412] = 8'b0;
    XRAM[22413] = 8'b0;
    XRAM[22414] = 8'b0;
    XRAM[22415] = 8'b0;
    XRAM[22416] = 8'b0;
    XRAM[22417] = 8'b0;
    XRAM[22418] = 8'b0;
    XRAM[22419] = 8'b0;
    XRAM[22420] = 8'b0;
    XRAM[22421] = 8'b0;
    XRAM[22422] = 8'b0;
    XRAM[22423] = 8'b0;
    XRAM[22424] = 8'b0;
    XRAM[22425] = 8'b0;
    XRAM[22426] = 8'b0;
    XRAM[22427] = 8'b0;
    XRAM[22428] = 8'b0;
    XRAM[22429] = 8'b0;
    XRAM[22430] = 8'b0;
    XRAM[22431] = 8'b0;
    XRAM[22432] = 8'b0;
    XRAM[22433] = 8'b0;
    XRAM[22434] = 8'b0;
    XRAM[22435] = 8'b0;
    XRAM[22436] = 8'b0;
    XRAM[22437] = 8'b0;
    XRAM[22438] = 8'b0;
    XRAM[22439] = 8'b0;
    XRAM[22440] = 8'b0;
    XRAM[22441] = 8'b0;
    XRAM[22442] = 8'b0;
    XRAM[22443] = 8'b0;
    XRAM[22444] = 8'b0;
    XRAM[22445] = 8'b0;
    XRAM[22446] = 8'b0;
    XRAM[22447] = 8'b0;
    XRAM[22448] = 8'b0;
    XRAM[22449] = 8'b0;
    XRAM[22450] = 8'b0;
    XRAM[22451] = 8'b0;
    XRAM[22452] = 8'b0;
    XRAM[22453] = 8'b0;
    XRAM[22454] = 8'b0;
    XRAM[22455] = 8'b0;
    XRAM[22456] = 8'b0;
    XRAM[22457] = 8'b0;
    XRAM[22458] = 8'b0;
    XRAM[22459] = 8'b0;
    XRAM[22460] = 8'b0;
    XRAM[22461] = 8'b0;
    XRAM[22462] = 8'b0;
    XRAM[22463] = 8'b0;
    XRAM[22464] = 8'b0;
    XRAM[22465] = 8'b0;
    XRAM[22466] = 8'b0;
    XRAM[22467] = 8'b0;
    XRAM[22468] = 8'b0;
    XRAM[22469] = 8'b0;
    XRAM[22470] = 8'b0;
    XRAM[22471] = 8'b0;
    XRAM[22472] = 8'b0;
    XRAM[22473] = 8'b0;
    XRAM[22474] = 8'b0;
    XRAM[22475] = 8'b0;
    XRAM[22476] = 8'b0;
    XRAM[22477] = 8'b0;
    XRAM[22478] = 8'b0;
    XRAM[22479] = 8'b0;
    XRAM[22480] = 8'b0;
    XRAM[22481] = 8'b0;
    XRAM[22482] = 8'b0;
    XRAM[22483] = 8'b0;
    XRAM[22484] = 8'b0;
    XRAM[22485] = 8'b0;
    XRAM[22486] = 8'b0;
    XRAM[22487] = 8'b0;
    XRAM[22488] = 8'b0;
    XRAM[22489] = 8'b0;
    XRAM[22490] = 8'b0;
    XRAM[22491] = 8'b0;
    XRAM[22492] = 8'b0;
    XRAM[22493] = 8'b0;
    XRAM[22494] = 8'b0;
    XRAM[22495] = 8'b0;
    XRAM[22496] = 8'b0;
    XRAM[22497] = 8'b0;
    XRAM[22498] = 8'b0;
    XRAM[22499] = 8'b0;
    XRAM[22500] = 8'b0;
    XRAM[22501] = 8'b0;
    XRAM[22502] = 8'b0;
    XRAM[22503] = 8'b0;
    XRAM[22504] = 8'b0;
    XRAM[22505] = 8'b0;
    XRAM[22506] = 8'b0;
    XRAM[22507] = 8'b0;
    XRAM[22508] = 8'b0;
    XRAM[22509] = 8'b0;
    XRAM[22510] = 8'b0;
    XRAM[22511] = 8'b0;
    XRAM[22512] = 8'b0;
    XRAM[22513] = 8'b0;
    XRAM[22514] = 8'b0;
    XRAM[22515] = 8'b0;
    XRAM[22516] = 8'b0;
    XRAM[22517] = 8'b0;
    XRAM[22518] = 8'b0;
    XRAM[22519] = 8'b0;
    XRAM[22520] = 8'b0;
    XRAM[22521] = 8'b0;
    XRAM[22522] = 8'b0;
    XRAM[22523] = 8'b0;
    XRAM[22524] = 8'b0;
    XRAM[22525] = 8'b0;
    XRAM[22526] = 8'b0;
    XRAM[22527] = 8'b0;
    XRAM[22528] = 8'b0;
    XRAM[22529] = 8'b0;
    XRAM[22530] = 8'b0;
    XRAM[22531] = 8'b0;
    XRAM[22532] = 8'b0;
    XRAM[22533] = 8'b0;
    XRAM[22534] = 8'b0;
    XRAM[22535] = 8'b0;
    XRAM[22536] = 8'b0;
    XRAM[22537] = 8'b0;
    XRAM[22538] = 8'b0;
    XRAM[22539] = 8'b0;
    XRAM[22540] = 8'b0;
    XRAM[22541] = 8'b0;
    XRAM[22542] = 8'b0;
    XRAM[22543] = 8'b0;
    XRAM[22544] = 8'b0;
    XRAM[22545] = 8'b0;
    XRAM[22546] = 8'b0;
    XRAM[22547] = 8'b0;
    XRAM[22548] = 8'b0;
    XRAM[22549] = 8'b0;
    XRAM[22550] = 8'b0;
    XRAM[22551] = 8'b0;
    XRAM[22552] = 8'b0;
    XRAM[22553] = 8'b0;
    XRAM[22554] = 8'b0;
    XRAM[22555] = 8'b0;
    XRAM[22556] = 8'b0;
    XRAM[22557] = 8'b0;
    XRAM[22558] = 8'b0;
    XRAM[22559] = 8'b0;
    XRAM[22560] = 8'b0;
    XRAM[22561] = 8'b0;
    XRAM[22562] = 8'b0;
    XRAM[22563] = 8'b0;
    XRAM[22564] = 8'b0;
    XRAM[22565] = 8'b0;
    XRAM[22566] = 8'b0;
    XRAM[22567] = 8'b0;
    XRAM[22568] = 8'b0;
    XRAM[22569] = 8'b0;
    XRAM[22570] = 8'b0;
    XRAM[22571] = 8'b0;
    XRAM[22572] = 8'b0;
    XRAM[22573] = 8'b0;
    XRAM[22574] = 8'b0;
    XRAM[22575] = 8'b0;
    XRAM[22576] = 8'b0;
    XRAM[22577] = 8'b0;
    XRAM[22578] = 8'b0;
    XRAM[22579] = 8'b0;
    XRAM[22580] = 8'b0;
    XRAM[22581] = 8'b0;
    XRAM[22582] = 8'b0;
    XRAM[22583] = 8'b0;
    XRAM[22584] = 8'b0;
    XRAM[22585] = 8'b0;
    XRAM[22586] = 8'b0;
    XRAM[22587] = 8'b0;
    XRAM[22588] = 8'b0;
    XRAM[22589] = 8'b0;
    XRAM[22590] = 8'b0;
    XRAM[22591] = 8'b0;
    XRAM[22592] = 8'b0;
    XRAM[22593] = 8'b0;
    XRAM[22594] = 8'b0;
    XRAM[22595] = 8'b0;
    XRAM[22596] = 8'b0;
    XRAM[22597] = 8'b0;
    XRAM[22598] = 8'b0;
    XRAM[22599] = 8'b0;
    XRAM[22600] = 8'b0;
    XRAM[22601] = 8'b0;
    XRAM[22602] = 8'b0;
    XRAM[22603] = 8'b0;
    XRAM[22604] = 8'b0;
    XRAM[22605] = 8'b0;
    XRAM[22606] = 8'b0;
    XRAM[22607] = 8'b0;
    XRAM[22608] = 8'b0;
    XRAM[22609] = 8'b0;
    XRAM[22610] = 8'b0;
    XRAM[22611] = 8'b0;
    XRAM[22612] = 8'b0;
    XRAM[22613] = 8'b0;
    XRAM[22614] = 8'b0;
    XRAM[22615] = 8'b0;
    XRAM[22616] = 8'b0;
    XRAM[22617] = 8'b0;
    XRAM[22618] = 8'b0;
    XRAM[22619] = 8'b0;
    XRAM[22620] = 8'b0;
    XRAM[22621] = 8'b0;
    XRAM[22622] = 8'b0;
    XRAM[22623] = 8'b0;
    XRAM[22624] = 8'b0;
    XRAM[22625] = 8'b0;
    XRAM[22626] = 8'b0;
    XRAM[22627] = 8'b0;
    XRAM[22628] = 8'b0;
    XRAM[22629] = 8'b0;
    XRAM[22630] = 8'b0;
    XRAM[22631] = 8'b0;
    XRAM[22632] = 8'b0;
    XRAM[22633] = 8'b0;
    XRAM[22634] = 8'b0;
    XRAM[22635] = 8'b0;
    XRAM[22636] = 8'b0;
    XRAM[22637] = 8'b0;
    XRAM[22638] = 8'b0;
    XRAM[22639] = 8'b0;
    XRAM[22640] = 8'b0;
    XRAM[22641] = 8'b0;
    XRAM[22642] = 8'b0;
    XRAM[22643] = 8'b0;
    XRAM[22644] = 8'b0;
    XRAM[22645] = 8'b0;
    XRAM[22646] = 8'b0;
    XRAM[22647] = 8'b0;
    XRAM[22648] = 8'b0;
    XRAM[22649] = 8'b0;
    XRAM[22650] = 8'b0;
    XRAM[22651] = 8'b0;
    XRAM[22652] = 8'b0;
    XRAM[22653] = 8'b0;
    XRAM[22654] = 8'b0;
    XRAM[22655] = 8'b0;
    XRAM[22656] = 8'b0;
    XRAM[22657] = 8'b0;
    XRAM[22658] = 8'b0;
    XRAM[22659] = 8'b0;
    XRAM[22660] = 8'b0;
    XRAM[22661] = 8'b0;
    XRAM[22662] = 8'b0;
    XRAM[22663] = 8'b0;
    XRAM[22664] = 8'b0;
    XRAM[22665] = 8'b0;
    XRAM[22666] = 8'b0;
    XRAM[22667] = 8'b0;
    XRAM[22668] = 8'b0;
    XRAM[22669] = 8'b0;
    XRAM[22670] = 8'b0;
    XRAM[22671] = 8'b0;
    XRAM[22672] = 8'b0;
    XRAM[22673] = 8'b0;
    XRAM[22674] = 8'b0;
    XRAM[22675] = 8'b0;
    XRAM[22676] = 8'b0;
    XRAM[22677] = 8'b0;
    XRAM[22678] = 8'b0;
    XRAM[22679] = 8'b0;
    XRAM[22680] = 8'b0;
    XRAM[22681] = 8'b0;
    XRAM[22682] = 8'b0;
    XRAM[22683] = 8'b0;
    XRAM[22684] = 8'b0;
    XRAM[22685] = 8'b0;
    XRAM[22686] = 8'b0;
    XRAM[22687] = 8'b0;
    XRAM[22688] = 8'b0;
    XRAM[22689] = 8'b0;
    XRAM[22690] = 8'b0;
    XRAM[22691] = 8'b0;
    XRAM[22692] = 8'b0;
    XRAM[22693] = 8'b0;
    XRAM[22694] = 8'b0;
    XRAM[22695] = 8'b0;
    XRAM[22696] = 8'b0;
    XRAM[22697] = 8'b0;
    XRAM[22698] = 8'b0;
    XRAM[22699] = 8'b0;
    XRAM[22700] = 8'b0;
    XRAM[22701] = 8'b0;
    XRAM[22702] = 8'b0;
    XRAM[22703] = 8'b0;
    XRAM[22704] = 8'b0;
    XRAM[22705] = 8'b0;
    XRAM[22706] = 8'b0;
    XRAM[22707] = 8'b0;
    XRAM[22708] = 8'b0;
    XRAM[22709] = 8'b0;
    XRAM[22710] = 8'b0;
    XRAM[22711] = 8'b0;
    XRAM[22712] = 8'b0;
    XRAM[22713] = 8'b0;
    XRAM[22714] = 8'b0;
    XRAM[22715] = 8'b0;
    XRAM[22716] = 8'b0;
    XRAM[22717] = 8'b0;
    XRAM[22718] = 8'b0;
    XRAM[22719] = 8'b0;
    XRAM[22720] = 8'b0;
    XRAM[22721] = 8'b0;
    XRAM[22722] = 8'b0;
    XRAM[22723] = 8'b0;
    XRAM[22724] = 8'b0;
    XRAM[22725] = 8'b0;
    XRAM[22726] = 8'b0;
    XRAM[22727] = 8'b0;
    XRAM[22728] = 8'b0;
    XRAM[22729] = 8'b0;
    XRAM[22730] = 8'b0;
    XRAM[22731] = 8'b0;
    XRAM[22732] = 8'b0;
    XRAM[22733] = 8'b0;
    XRAM[22734] = 8'b0;
    XRAM[22735] = 8'b0;
    XRAM[22736] = 8'b0;
    XRAM[22737] = 8'b0;
    XRAM[22738] = 8'b0;
    XRAM[22739] = 8'b0;
    XRAM[22740] = 8'b0;
    XRAM[22741] = 8'b0;
    XRAM[22742] = 8'b0;
    XRAM[22743] = 8'b0;
    XRAM[22744] = 8'b0;
    XRAM[22745] = 8'b0;
    XRAM[22746] = 8'b0;
    XRAM[22747] = 8'b0;
    XRAM[22748] = 8'b0;
    XRAM[22749] = 8'b0;
    XRAM[22750] = 8'b0;
    XRAM[22751] = 8'b0;
    XRAM[22752] = 8'b0;
    XRAM[22753] = 8'b0;
    XRAM[22754] = 8'b0;
    XRAM[22755] = 8'b0;
    XRAM[22756] = 8'b0;
    XRAM[22757] = 8'b0;
    XRAM[22758] = 8'b0;
    XRAM[22759] = 8'b0;
    XRAM[22760] = 8'b0;
    XRAM[22761] = 8'b0;
    XRAM[22762] = 8'b0;
    XRAM[22763] = 8'b0;
    XRAM[22764] = 8'b0;
    XRAM[22765] = 8'b0;
    XRAM[22766] = 8'b0;
    XRAM[22767] = 8'b0;
    XRAM[22768] = 8'b0;
    XRAM[22769] = 8'b0;
    XRAM[22770] = 8'b0;
    XRAM[22771] = 8'b0;
    XRAM[22772] = 8'b0;
    XRAM[22773] = 8'b0;
    XRAM[22774] = 8'b0;
    XRAM[22775] = 8'b0;
    XRAM[22776] = 8'b0;
    XRAM[22777] = 8'b0;
    XRAM[22778] = 8'b0;
    XRAM[22779] = 8'b0;
    XRAM[22780] = 8'b0;
    XRAM[22781] = 8'b0;
    XRAM[22782] = 8'b0;
    XRAM[22783] = 8'b0;
    XRAM[22784] = 8'b0;
    XRAM[22785] = 8'b0;
    XRAM[22786] = 8'b0;
    XRAM[22787] = 8'b0;
    XRAM[22788] = 8'b0;
    XRAM[22789] = 8'b0;
    XRAM[22790] = 8'b0;
    XRAM[22791] = 8'b0;
    XRAM[22792] = 8'b0;
    XRAM[22793] = 8'b0;
    XRAM[22794] = 8'b0;
    XRAM[22795] = 8'b0;
    XRAM[22796] = 8'b0;
    XRAM[22797] = 8'b0;
    XRAM[22798] = 8'b0;
    XRAM[22799] = 8'b0;
    XRAM[22800] = 8'b0;
    XRAM[22801] = 8'b0;
    XRAM[22802] = 8'b0;
    XRAM[22803] = 8'b0;
    XRAM[22804] = 8'b0;
    XRAM[22805] = 8'b0;
    XRAM[22806] = 8'b0;
    XRAM[22807] = 8'b0;
    XRAM[22808] = 8'b0;
    XRAM[22809] = 8'b0;
    XRAM[22810] = 8'b0;
    XRAM[22811] = 8'b0;
    XRAM[22812] = 8'b0;
    XRAM[22813] = 8'b0;
    XRAM[22814] = 8'b0;
    XRAM[22815] = 8'b0;
    XRAM[22816] = 8'b0;
    XRAM[22817] = 8'b0;
    XRAM[22818] = 8'b0;
    XRAM[22819] = 8'b0;
    XRAM[22820] = 8'b0;
    XRAM[22821] = 8'b0;
    XRAM[22822] = 8'b0;
    XRAM[22823] = 8'b0;
    XRAM[22824] = 8'b0;
    XRAM[22825] = 8'b0;
    XRAM[22826] = 8'b0;
    XRAM[22827] = 8'b0;
    XRAM[22828] = 8'b0;
    XRAM[22829] = 8'b0;
    XRAM[22830] = 8'b0;
    XRAM[22831] = 8'b0;
    XRAM[22832] = 8'b0;
    XRAM[22833] = 8'b0;
    XRAM[22834] = 8'b0;
    XRAM[22835] = 8'b0;
    XRAM[22836] = 8'b0;
    XRAM[22837] = 8'b0;
    XRAM[22838] = 8'b0;
    XRAM[22839] = 8'b0;
    XRAM[22840] = 8'b0;
    XRAM[22841] = 8'b0;
    XRAM[22842] = 8'b0;
    XRAM[22843] = 8'b0;
    XRAM[22844] = 8'b0;
    XRAM[22845] = 8'b0;
    XRAM[22846] = 8'b0;
    XRAM[22847] = 8'b0;
    XRAM[22848] = 8'b0;
    XRAM[22849] = 8'b0;
    XRAM[22850] = 8'b0;
    XRAM[22851] = 8'b0;
    XRAM[22852] = 8'b0;
    XRAM[22853] = 8'b0;
    XRAM[22854] = 8'b0;
    XRAM[22855] = 8'b0;
    XRAM[22856] = 8'b0;
    XRAM[22857] = 8'b0;
    XRAM[22858] = 8'b0;
    XRAM[22859] = 8'b0;
    XRAM[22860] = 8'b0;
    XRAM[22861] = 8'b0;
    XRAM[22862] = 8'b0;
    XRAM[22863] = 8'b0;
    XRAM[22864] = 8'b0;
    XRAM[22865] = 8'b0;
    XRAM[22866] = 8'b0;
    XRAM[22867] = 8'b0;
    XRAM[22868] = 8'b0;
    XRAM[22869] = 8'b0;
    XRAM[22870] = 8'b0;
    XRAM[22871] = 8'b0;
    XRAM[22872] = 8'b0;
    XRAM[22873] = 8'b0;
    XRAM[22874] = 8'b0;
    XRAM[22875] = 8'b0;
    XRAM[22876] = 8'b0;
    XRAM[22877] = 8'b0;
    XRAM[22878] = 8'b0;
    XRAM[22879] = 8'b0;
    XRAM[22880] = 8'b0;
    XRAM[22881] = 8'b0;
    XRAM[22882] = 8'b0;
    XRAM[22883] = 8'b0;
    XRAM[22884] = 8'b0;
    XRAM[22885] = 8'b0;
    XRAM[22886] = 8'b0;
    XRAM[22887] = 8'b0;
    XRAM[22888] = 8'b0;
    XRAM[22889] = 8'b0;
    XRAM[22890] = 8'b0;
    XRAM[22891] = 8'b0;
    XRAM[22892] = 8'b0;
    XRAM[22893] = 8'b0;
    XRAM[22894] = 8'b0;
    XRAM[22895] = 8'b0;
    XRAM[22896] = 8'b0;
    XRAM[22897] = 8'b0;
    XRAM[22898] = 8'b0;
    XRAM[22899] = 8'b0;
    XRAM[22900] = 8'b0;
    XRAM[22901] = 8'b0;
    XRAM[22902] = 8'b0;
    XRAM[22903] = 8'b0;
    XRAM[22904] = 8'b0;
    XRAM[22905] = 8'b0;
    XRAM[22906] = 8'b0;
    XRAM[22907] = 8'b0;
    XRAM[22908] = 8'b0;
    XRAM[22909] = 8'b0;
    XRAM[22910] = 8'b0;
    XRAM[22911] = 8'b0;
    XRAM[22912] = 8'b0;
    XRAM[22913] = 8'b0;
    XRAM[22914] = 8'b0;
    XRAM[22915] = 8'b0;
    XRAM[22916] = 8'b0;
    XRAM[22917] = 8'b0;
    XRAM[22918] = 8'b0;
    XRAM[22919] = 8'b0;
    XRAM[22920] = 8'b0;
    XRAM[22921] = 8'b0;
    XRAM[22922] = 8'b0;
    XRAM[22923] = 8'b0;
    XRAM[22924] = 8'b0;
    XRAM[22925] = 8'b0;
    XRAM[22926] = 8'b0;
    XRAM[22927] = 8'b0;
    XRAM[22928] = 8'b0;
    XRAM[22929] = 8'b0;
    XRAM[22930] = 8'b0;
    XRAM[22931] = 8'b0;
    XRAM[22932] = 8'b0;
    XRAM[22933] = 8'b0;
    XRAM[22934] = 8'b0;
    XRAM[22935] = 8'b0;
    XRAM[22936] = 8'b0;
    XRAM[22937] = 8'b0;
    XRAM[22938] = 8'b0;
    XRAM[22939] = 8'b0;
    XRAM[22940] = 8'b0;
    XRAM[22941] = 8'b0;
    XRAM[22942] = 8'b0;
    XRAM[22943] = 8'b0;
    XRAM[22944] = 8'b0;
    XRAM[22945] = 8'b0;
    XRAM[22946] = 8'b0;
    XRAM[22947] = 8'b0;
    XRAM[22948] = 8'b0;
    XRAM[22949] = 8'b0;
    XRAM[22950] = 8'b0;
    XRAM[22951] = 8'b0;
    XRAM[22952] = 8'b0;
    XRAM[22953] = 8'b0;
    XRAM[22954] = 8'b0;
    XRAM[22955] = 8'b0;
    XRAM[22956] = 8'b0;
    XRAM[22957] = 8'b0;
    XRAM[22958] = 8'b0;
    XRAM[22959] = 8'b0;
    XRAM[22960] = 8'b0;
    XRAM[22961] = 8'b0;
    XRAM[22962] = 8'b0;
    XRAM[22963] = 8'b0;
    XRAM[22964] = 8'b0;
    XRAM[22965] = 8'b0;
    XRAM[22966] = 8'b0;
    XRAM[22967] = 8'b0;
    XRAM[22968] = 8'b0;
    XRAM[22969] = 8'b0;
    XRAM[22970] = 8'b0;
    XRAM[22971] = 8'b0;
    XRAM[22972] = 8'b0;
    XRAM[22973] = 8'b0;
    XRAM[22974] = 8'b0;
    XRAM[22975] = 8'b0;
    XRAM[22976] = 8'b0;
    XRAM[22977] = 8'b0;
    XRAM[22978] = 8'b0;
    XRAM[22979] = 8'b0;
    XRAM[22980] = 8'b0;
    XRAM[22981] = 8'b0;
    XRAM[22982] = 8'b0;
    XRAM[22983] = 8'b0;
    XRAM[22984] = 8'b0;
    XRAM[22985] = 8'b0;
    XRAM[22986] = 8'b0;
    XRAM[22987] = 8'b0;
    XRAM[22988] = 8'b0;
    XRAM[22989] = 8'b0;
    XRAM[22990] = 8'b0;
    XRAM[22991] = 8'b0;
    XRAM[22992] = 8'b0;
    XRAM[22993] = 8'b0;
    XRAM[22994] = 8'b0;
    XRAM[22995] = 8'b0;
    XRAM[22996] = 8'b0;
    XRAM[22997] = 8'b0;
    XRAM[22998] = 8'b0;
    XRAM[22999] = 8'b0;
    XRAM[23000] = 8'b0;
    XRAM[23001] = 8'b0;
    XRAM[23002] = 8'b0;
    XRAM[23003] = 8'b0;
    XRAM[23004] = 8'b0;
    XRAM[23005] = 8'b0;
    XRAM[23006] = 8'b0;
    XRAM[23007] = 8'b0;
    XRAM[23008] = 8'b0;
    XRAM[23009] = 8'b0;
    XRAM[23010] = 8'b0;
    XRAM[23011] = 8'b0;
    XRAM[23012] = 8'b0;
    XRAM[23013] = 8'b0;
    XRAM[23014] = 8'b0;
    XRAM[23015] = 8'b0;
    XRAM[23016] = 8'b0;
    XRAM[23017] = 8'b0;
    XRAM[23018] = 8'b0;
    XRAM[23019] = 8'b0;
    XRAM[23020] = 8'b0;
    XRAM[23021] = 8'b0;
    XRAM[23022] = 8'b0;
    XRAM[23023] = 8'b0;
    XRAM[23024] = 8'b0;
    XRAM[23025] = 8'b0;
    XRAM[23026] = 8'b0;
    XRAM[23027] = 8'b0;
    XRAM[23028] = 8'b0;
    XRAM[23029] = 8'b0;
    XRAM[23030] = 8'b0;
    XRAM[23031] = 8'b0;
    XRAM[23032] = 8'b0;
    XRAM[23033] = 8'b0;
    XRAM[23034] = 8'b0;
    XRAM[23035] = 8'b0;
    XRAM[23036] = 8'b0;
    XRAM[23037] = 8'b0;
    XRAM[23038] = 8'b0;
    XRAM[23039] = 8'b0;
    XRAM[23040] = 8'b0;
    XRAM[23041] = 8'b0;
    XRAM[23042] = 8'b0;
    XRAM[23043] = 8'b0;
    XRAM[23044] = 8'b0;
    XRAM[23045] = 8'b0;
    XRAM[23046] = 8'b0;
    XRAM[23047] = 8'b0;
    XRAM[23048] = 8'b0;
    XRAM[23049] = 8'b0;
    XRAM[23050] = 8'b0;
    XRAM[23051] = 8'b0;
    XRAM[23052] = 8'b0;
    XRAM[23053] = 8'b0;
    XRAM[23054] = 8'b0;
    XRAM[23055] = 8'b0;
    XRAM[23056] = 8'b0;
    XRAM[23057] = 8'b0;
    XRAM[23058] = 8'b0;
    XRAM[23059] = 8'b0;
    XRAM[23060] = 8'b0;
    XRAM[23061] = 8'b0;
    XRAM[23062] = 8'b0;
    XRAM[23063] = 8'b0;
    XRAM[23064] = 8'b0;
    XRAM[23065] = 8'b0;
    XRAM[23066] = 8'b0;
    XRAM[23067] = 8'b0;
    XRAM[23068] = 8'b0;
    XRAM[23069] = 8'b0;
    XRAM[23070] = 8'b0;
    XRAM[23071] = 8'b0;
    XRAM[23072] = 8'b0;
    XRAM[23073] = 8'b0;
    XRAM[23074] = 8'b0;
    XRAM[23075] = 8'b0;
    XRAM[23076] = 8'b0;
    XRAM[23077] = 8'b0;
    XRAM[23078] = 8'b0;
    XRAM[23079] = 8'b0;
    XRAM[23080] = 8'b0;
    XRAM[23081] = 8'b0;
    XRAM[23082] = 8'b0;
    XRAM[23083] = 8'b0;
    XRAM[23084] = 8'b0;
    XRAM[23085] = 8'b0;
    XRAM[23086] = 8'b0;
    XRAM[23087] = 8'b0;
    XRAM[23088] = 8'b0;
    XRAM[23089] = 8'b0;
    XRAM[23090] = 8'b0;
    XRAM[23091] = 8'b0;
    XRAM[23092] = 8'b0;
    XRAM[23093] = 8'b0;
    XRAM[23094] = 8'b0;
    XRAM[23095] = 8'b0;
    XRAM[23096] = 8'b0;
    XRAM[23097] = 8'b0;
    XRAM[23098] = 8'b0;
    XRAM[23099] = 8'b0;
    XRAM[23100] = 8'b0;
    XRAM[23101] = 8'b0;
    XRAM[23102] = 8'b0;
    XRAM[23103] = 8'b0;
    XRAM[23104] = 8'b0;
    XRAM[23105] = 8'b0;
    XRAM[23106] = 8'b0;
    XRAM[23107] = 8'b0;
    XRAM[23108] = 8'b0;
    XRAM[23109] = 8'b0;
    XRAM[23110] = 8'b0;
    XRAM[23111] = 8'b0;
    XRAM[23112] = 8'b0;
    XRAM[23113] = 8'b0;
    XRAM[23114] = 8'b0;
    XRAM[23115] = 8'b0;
    XRAM[23116] = 8'b0;
    XRAM[23117] = 8'b0;
    XRAM[23118] = 8'b0;
    XRAM[23119] = 8'b0;
    XRAM[23120] = 8'b0;
    XRAM[23121] = 8'b0;
    XRAM[23122] = 8'b0;
    XRAM[23123] = 8'b0;
    XRAM[23124] = 8'b0;
    XRAM[23125] = 8'b0;
    XRAM[23126] = 8'b0;
    XRAM[23127] = 8'b0;
    XRAM[23128] = 8'b0;
    XRAM[23129] = 8'b0;
    XRAM[23130] = 8'b0;
    XRAM[23131] = 8'b0;
    XRAM[23132] = 8'b0;
    XRAM[23133] = 8'b0;
    XRAM[23134] = 8'b0;
    XRAM[23135] = 8'b0;
    XRAM[23136] = 8'b0;
    XRAM[23137] = 8'b0;
    XRAM[23138] = 8'b0;
    XRAM[23139] = 8'b0;
    XRAM[23140] = 8'b0;
    XRAM[23141] = 8'b0;
    XRAM[23142] = 8'b0;
    XRAM[23143] = 8'b0;
    XRAM[23144] = 8'b0;
    XRAM[23145] = 8'b0;
    XRAM[23146] = 8'b0;
    XRAM[23147] = 8'b0;
    XRAM[23148] = 8'b0;
    XRAM[23149] = 8'b0;
    XRAM[23150] = 8'b0;
    XRAM[23151] = 8'b0;
    XRAM[23152] = 8'b0;
    XRAM[23153] = 8'b0;
    XRAM[23154] = 8'b0;
    XRAM[23155] = 8'b0;
    XRAM[23156] = 8'b0;
    XRAM[23157] = 8'b0;
    XRAM[23158] = 8'b0;
    XRAM[23159] = 8'b0;
    XRAM[23160] = 8'b0;
    XRAM[23161] = 8'b0;
    XRAM[23162] = 8'b0;
    XRAM[23163] = 8'b0;
    XRAM[23164] = 8'b0;
    XRAM[23165] = 8'b0;
    XRAM[23166] = 8'b0;
    XRAM[23167] = 8'b0;
    XRAM[23168] = 8'b0;
    XRAM[23169] = 8'b0;
    XRAM[23170] = 8'b0;
    XRAM[23171] = 8'b0;
    XRAM[23172] = 8'b0;
    XRAM[23173] = 8'b0;
    XRAM[23174] = 8'b0;
    XRAM[23175] = 8'b0;
    XRAM[23176] = 8'b0;
    XRAM[23177] = 8'b0;
    XRAM[23178] = 8'b0;
    XRAM[23179] = 8'b0;
    XRAM[23180] = 8'b0;
    XRAM[23181] = 8'b0;
    XRAM[23182] = 8'b0;
    XRAM[23183] = 8'b0;
    XRAM[23184] = 8'b0;
    XRAM[23185] = 8'b0;
    XRAM[23186] = 8'b0;
    XRAM[23187] = 8'b0;
    XRAM[23188] = 8'b0;
    XRAM[23189] = 8'b0;
    XRAM[23190] = 8'b0;
    XRAM[23191] = 8'b0;
    XRAM[23192] = 8'b0;
    XRAM[23193] = 8'b0;
    XRAM[23194] = 8'b0;
    XRAM[23195] = 8'b0;
    XRAM[23196] = 8'b0;
    XRAM[23197] = 8'b0;
    XRAM[23198] = 8'b0;
    XRAM[23199] = 8'b0;
    XRAM[23200] = 8'b0;
    XRAM[23201] = 8'b0;
    XRAM[23202] = 8'b0;
    XRAM[23203] = 8'b0;
    XRAM[23204] = 8'b0;
    XRAM[23205] = 8'b0;
    XRAM[23206] = 8'b0;
    XRAM[23207] = 8'b0;
    XRAM[23208] = 8'b0;
    XRAM[23209] = 8'b0;
    XRAM[23210] = 8'b0;
    XRAM[23211] = 8'b0;
    XRAM[23212] = 8'b0;
    XRAM[23213] = 8'b0;
    XRAM[23214] = 8'b0;
    XRAM[23215] = 8'b0;
    XRAM[23216] = 8'b0;
    XRAM[23217] = 8'b0;
    XRAM[23218] = 8'b0;
    XRAM[23219] = 8'b0;
    XRAM[23220] = 8'b0;
    XRAM[23221] = 8'b0;
    XRAM[23222] = 8'b0;
    XRAM[23223] = 8'b0;
    XRAM[23224] = 8'b0;
    XRAM[23225] = 8'b0;
    XRAM[23226] = 8'b0;
    XRAM[23227] = 8'b0;
    XRAM[23228] = 8'b0;
    XRAM[23229] = 8'b0;
    XRAM[23230] = 8'b0;
    XRAM[23231] = 8'b0;
    XRAM[23232] = 8'b0;
    XRAM[23233] = 8'b0;
    XRAM[23234] = 8'b0;
    XRAM[23235] = 8'b0;
    XRAM[23236] = 8'b0;
    XRAM[23237] = 8'b0;
    XRAM[23238] = 8'b0;
    XRAM[23239] = 8'b0;
    XRAM[23240] = 8'b0;
    XRAM[23241] = 8'b0;
    XRAM[23242] = 8'b0;
    XRAM[23243] = 8'b0;
    XRAM[23244] = 8'b0;
    XRAM[23245] = 8'b0;
    XRAM[23246] = 8'b0;
    XRAM[23247] = 8'b0;
    XRAM[23248] = 8'b0;
    XRAM[23249] = 8'b0;
    XRAM[23250] = 8'b0;
    XRAM[23251] = 8'b0;
    XRAM[23252] = 8'b0;
    XRAM[23253] = 8'b0;
    XRAM[23254] = 8'b0;
    XRAM[23255] = 8'b0;
    XRAM[23256] = 8'b0;
    XRAM[23257] = 8'b0;
    XRAM[23258] = 8'b0;
    XRAM[23259] = 8'b0;
    XRAM[23260] = 8'b0;
    XRAM[23261] = 8'b0;
    XRAM[23262] = 8'b0;
    XRAM[23263] = 8'b0;
    XRAM[23264] = 8'b0;
    XRAM[23265] = 8'b0;
    XRAM[23266] = 8'b0;
    XRAM[23267] = 8'b0;
    XRAM[23268] = 8'b0;
    XRAM[23269] = 8'b0;
    XRAM[23270] = 8'b0;
    XRAM[23271] = 8'b0;
    XRAM[23272] = 8'b0;
    XRAM[23273] = 8'b0;
    XRAM[23274] = 8'b0;
    XRAM[23275] = 8'b0;
    XRAM[23276] = 8'b0;
    XRAM[23277] = 8'b0;
    XRAM[23278] = 8'b0;
    XRAM[23279] = 8'b0;
    XRAM[23280] = 8'b0;
    XRAM[23281] = 8'b0;
    XRAM[23282] = 8'b0;
    XRAM[23283] = 8'b0;
    XRAM[23284] = 8'b0;
    XRAM[23285] = 8'b0;
    XRAM[23286] = 8'b0;
    XRAM[23287] = 8'b0;
    XRAM[23288] = 8'b0;
    XRAM[23289] = 8'b0;
    XRAM[23290] = 8'b0;
    XRAM[23291] = 8'b0;
    XRAM[23292] = 8'b0;
    XRAM[23293] = 8'b0;
    XRAM[23294] = 8'b0;
    XRAM[23295] = 8'b0;
    XRAM[23296] = 8'b0;
    XRAM[23297] = 8'b0;
    XRAM[23298] = 8'b0;
    XRAM[23299] = 8'b0;
    XRAM[23300] = 8'b0;
    XRAM[23301] = 8'b0;
    XRAM[23302] = 8'b0;
    XRAM[23303] = 8'b0;
    XRAM[23304] = 8'b0;
    XRAM[23305] = 8'b0;
    XRAM[23306] = 8'b0;
    XRAM[23307] = 8'b0;
    XRAM[23308] = 8'b0;
    XRAM[23309] = 8'b0;
    XRAM[23310] = 8'b0;
    XRAM[23311] = 8'b0;
    XRAM[23312] = 8'b0;
    XRAM[23313] = 8'b0;
    XRAM[23314] = 8'b0;
    XRAM[23315] = 8'b0;
    XRAM[23316] = 8'b0;
    XRAM[23317] = 8'b0;
    XRAM[23318] = 8'b0;
    XRAM[23319] = 8'b0;
    XRAM[23320] = 8'b0;
    XRAM[23321] = 8'b0;
    XRAM[23322] = 8'b0;
    XRAM[23323] = 8'b0;
    XRAM[23324] = 8'b0;
    XRAM[23325] = 8'b0;
    XRAM[23326] = 8'b0;
    XRAM[23327] = 8'b0;
    XRAM[23328] = 8'b0;
    XRAM[23329] = 8'b0;
    XRAM[23330] = 8'b0;
    XRAM[23331] = 8'b0;
    XRAM[23332] = 8'b0;
    XRAM[23333] = 8'b0;
    XRAM[23334] = 8'b0;
    XRAM[23335] = 8'b0;
    XRAM[23336] = 8'b0;
    XRAM[23337] = 8'b0;
    XRAM[23338] = 8'b0;
    XRAM[23339] = 8'b0;
    XRAM[23340] = 8'b0;
    XRAM[23341] = 8'b0;
    XRAM[23342] = 8'b0;
    XRAM[23343] = 8'b0;
    XRAM[23344] = 8'b0;
    XRAM[23345] = 8'b0;
    XRAM[23346] = 8'b0;
    XRAM[23347] = 8'b0;
    XRAM[23348] = 8'b0;
    XRAM[23349] = 8'b0;
    XRAM[23350] = 8'b0;
    XRAM[23351] = 8'b0;
    XRAM[23352] = 8'b0;
    XRAM[23353] = 8'b0;
    XRAM[23354] = 8'b0;
    XRAM[23355] = 8'b0;
    XRAM[23356] = 8'b0;
    XRAM[23357] = 8'b0;
    XRAM[23358] = 8'b0;
    XRAM[23359] = 8'b0;
    XRAM[23360] = 8'b0;
    XRAM[23361] = 8'b0;
    XRAM[23362] = 8'b0;
    XRAM[23363] = 8'b0;
    XRAM[23364] = 8'b0;
    XRAM[23365] = 8'b0;
    XRAM[23366] = 8'b0;
    XRAM[23367] = 8'b0;
    XRAM[23368] = 8'b0;
    XRAM[23369] = 8'b0;
    XRAM[23370] = 8'b0;
    XRAM[23371] = 8'b0;
    XRAM[23372] = 8'b0;
    XRAM[23373] = 8'b0;
    XRAM[23374] = 8'b0;
    XRAM[23375] = 8'b0;
    XRAM[23376] = 8'b0;
    XRAM[23377] = 8'b0;
    XRAM[23378] = 8'b0;
    XRAM[23379] = 8'b0;
    XRAM[23380] = 8'b0;
    XRAM[23381] = 8'b0;
    XRAM[23382] = 8'b0;
    XRAM[23383] = 8'b0;
    XRAM[23384] = 8'b0;
    XRAM[23385] = 8'b0;
    XRAM[23386] = 8'b0;
    XRAM[23387] = 8'b0;
    XRAM[23388] = 8'b0;
    XRAM[23389] = 8'b0;
    XRAM[23390] = 8'b0;
    XRAM[23391] = 8'b0;
    XRAM[23392] = 8'b0;
    XRAM[23393] = 8'b0;
    XRAM[23394] = 8'b0;
    XRAM[23395] = 8'b0;
    XRAM[23396] = 8'b0;
    XRAM[23397] = 8'b0;
    XRAM[23398] = 8'b0;
    XRAM[23399] = 8'b0;
    XRAM[23400] = 8'b0;
    XRAM[23401] = 8'b0;
    XRAM[23402] = 8'b0;
    XRAM[23403] = 8'b0;
    XRAM[23404] = 8'b0;
    XRAM[23405] = 8'b0;
    XRAM[23406] = 8'b0;
    XRAM[23407] = 8'b0;
    XRAM[23408] = 8'b0;
    XRAM[23409] = 8'b0;
    XRAM[23410] = 8'b0;
    XRAM[23411] = 8'b0;
    XRAM[23412] = 8'b0;
    XRAM[23413] = 8'b0;
    XRAM[23414] = 8'b0;
    XRAM[23415] = 8'b0;
    XRAM[23416] = 8'b0;
    XRAM[23417] = 8'b0;
    XRAM[23418] = 8'b0;
    XRAM[23419] = 8'b0;
    XRAM[23420] = 8'b0;
    XRAM[23421] = 8'b0;
    XRAM[23422] = 8'b0;
    XRAM[23423] = 8'b0;
    XRAM[23424] = 8'b0;
    XRAM[23425] = 8'b0;
    XRAM[23426] = 8'b0;
    XRAM[23427] = 8'b0;
    XRAM[23428] = 8'b0;
    XRAM[23429] = 8'b0;
    XRAM[23430] = 8'b0;
    XRAM[23431] = 8'b0;
    XRAM[23432] = 8'b0;
    XRAM[23433] = 8'b0;
    XRAM[23434] = 8'b0;
    XRAM[23435] = 8'b0;
    XRAM[23436] = 8'b0;
    XRAM[23437] = 8'b0;
    XRAM[23438] = 8'b0;
    XRAM[23439] = 8'b0;
    XRAM[23440] = 8'b0;
    XRAM[23441] = 8'b0;
    XRAM[23442] = 8'b0;
    XRAM[23443] = 8'b0;
    XRAM[23444] = 8'b0;
    XRAM[23445] = 8'b0;
    XRAM[23446] = 8'b0;
    XRAM[23447] = 8'b0;
    XRAM[23448] = 8'b0;
    XRAM[23449] = 8'b0;
    XRAM[23450] = 8'b0;
    XRAM[23451] = 8'b0;
    XRAM[23452] = 8'b0;
    XRAM[23453] = 8'b0;
    XRAM[23454] = 8'b0;
    XRAM[23455] = 8'b0;
    XRAM[23456] = 8'b0;
    XRAM[23457] = 8'b0;
    XRAM[23458] = 8'b0;
    XRAM[23459] = 8'b0;
    XRAM[23460] = 8'b0;
    XRAM[23461] = 8'b0;
    XRAM[23462] = 8'b0;
    XRAM[23463] = 8'b0;
    XRAM[23464] = 8'b0;
    XRAM[23465] = 8'b0;
    XRAM[23466] = 8'b0;
    XRAM[23467] = 8'b0;
    XRAM[23468] = 8'b0;
    XRAM[23469] = 8'b0;
    XRAM[23470] = 8'b0;
    XRAM[23471] = 8'b0;
    XRAM[23472] = 8'b0;
    XRAM[23473] = 8'b0;
    XRAM[23474] = 8'b0;
    XRAM[23475] = 8'b0;
    XRAM[23476] = 8'b0;
    XRAM[23477] = 8'b0;
    XRAM[23478] = 8'b0;
    XRAM[23479] = 8'b0;
    XRAM[23480] = 8'b0;
    XRAM[23481] = 8'b0;
    XRAM[23482] = 8'b0;
    XRAM[23483] = 8'b0;
    XRAM[23484] = 8'b0;
    XRAM[23485] = 8'b0;
    XRAM[23486] = 8'b0;
    XRAM[23487] = 8'b0;
    XRAM[23488] = 8'b0;
    XRAM[23489] = 8'b0;
    XRAM[23490] = 8'b0;
    XRAM[23491] = 8'b0;
    XRAM[23492] = 8'b0;
    XRAM[23493] = 8'b0;
    XRAM[23494] = 8'b0;
    XRAM[23495] = 8'b0;
    XRAM[23496] = 8'b0;
    XRAM[23497] = 8'b0;
    XRAM[23498] = 8'b0;
    XRAM[23499] = 8'b0;
    XRAM[23500] = 8'b0;
    XRAM[23501] = 8'b0;
    XRAM[23502] = 8'b0;
    XRAM[23503] = 8'b0;
    XRAM[23504] = 8'b0;
    XRAM[23505] = 8'b0;
    XRAM[23506] = 8'b0;
    XRAM[23507] = 8'b0;
    XRAM[23508] = 8'b0;
    XRAM[23509] = 8'b0;
    XRAM[23510] = 8'b0;
    XRAM[23511] = 8'b0;
    XRAM[23512] = 8'b0;
    XRAM[23513] = 8'b0;
    XRAM[23514] = 8'b0;
    XRAM[23515] = 8'b0;
    XRAM[23516] = 8'b0;
    XRAM[23517] = 8'b0;
    XRAM[23518] = 8'b0;
    XRAM[23519] = 8'b0;
    XRAM[23520] = 8'b0;
    XRAM[23521] = 8'b0;
    XRAM[23522] = 8'b0;
    XRAM[23523] = 8'b0;
    XRAM[23524] = 8'b0;
    XRAM[23525] = 8'b0;
    XRAM[23526] = 8'b0;
    XRAM[23527] = 8'b0;
    XRAM[23528] = 8'b0;
    XRAM[23529] = 8'b0;
    XRAM[23530] = 8'b0;
    XRAM[23531] = 8'b0;
    XRAM[23532] = 8'b0;
    XRAM[23533] = 8'b0;
    XRAM[23534] = 8'b0;
    XRAM[23535] = 8'b0;
    XRAM[23536] = 8'b0;
    XRAM[23537] = 8'b0;
    XRAM[23538] = 8'b0;
    XRAM[23539] = 8'b0;
    XRAM[23540] = 8'b0;
    XRAM[23541] = 8'b0;
    XRAM[23542] = 8'b0;
    XRAM[23543] = 8'b0;
    XRAM[23544] = 8'b0;
    XRAM[23545] = 8'b0;
    XRAM[23546] = 8'b0;
    XRAM[23547] = 8'b0;
    XRAM[23548] = 8'b0;
    XRAM[23549] = 8'b0;
    XRAM[23550] = 8'b0;
    XRAM[23551] = 8'b0;
    XRAM[23552] = 8'b0;
    XRAM[23553] = 8'b0;
    XRAM[23554] = 8'b0;
    XRAM[23555] = 8'b0;
    XRAM[23556] = 8'b0;
    XRAM[23557] = 8'b0;
    XRAM[23558] = 8'b0;
    XRAM[23559] = 8'b0;
    XRAM[23560] = 8'b0;
    XRAM[23561] = 8'b0;
    XRAM[23562] = 8'b0;
    XRAM[23563] = 8'b0;
    XRAM[23564] = 8'b0;
    XRAM[23565] = 8'b0;
    XRAM[23566] = 8'b0;
    XRAM[23567] = 8'b0;
    XRAM[23568] = 8'b0;
    XRAM[23569] = 8'b0;
    XRAM[23570] = 8'b0;
    XRAM[23571] = 8'b0;
    XRAM[23572] = 8'b0;
    XRAM[23573] = 8'b0;
    XRAM[23574] = 8'b0;
    XRAM[23575] = 8'b0;
    XRAM[23576] = 8'b0;
    XRAM[23577] = 8'b0;
    XRAM[23578] = 8'b0;
    XRAM[23579] = 8'b0;
    XRAM[23580] = 8'b0;
    XRAM[23581] = 8'b0;
    XRAM[23582] = 8'b0;
    XRAM[23583] = 8'b0;
    XRAM[23584] = 8'b0;
    XRAM[23585] = 8'b0;
    XRAM[23586] = 8'b0;
    XRAM[23587] = 8'b0;
    XRAM[23588] = 8'b0;
    XRAM[23589] = 8'b0;
    XRAM[23590] = 8'b0;
    XRAM[23591] = 8'b0;
    XRAM[23592] = 8'b0;
    XRAM[23593] = 8'b0;
    XRAM[23594] = 8'b0;
    XRAM[23595] = 8'b0;
    XRAM[23596] = 8'b0;
    XRAM[23597] = 8'b0;
    XRAM[23598] = 8'b0;
    XRAM[23599] = 8'b0;
    XRAM[23600] = 8'b0;
    XRAM[23601] = 8'b0;
    XRAM[23602] = 8'b0;
    XRAM[23603] = 8'b0;
    XRAM[23604] = 8'b0;
    XRAM[23605] = 8'b0;
    XRAM[23606] = 8'b0;
    XRAM[23607] = 8'b0;
    XRAM[23608] = 8'b0;
    XRAM[23609] = 8'b0;
    XRAM[23610] = 8'b0;
    XRAM[23611] = 8'b0;
    XRAM[23612] = 8'b0;
    XRAM[23613] = 8'b0;
    XRAM[23614] = 8'b0;
    XRAM[23615] = 8'b0;
    XRAM[23616] = 8'b0;
    XRAM[23617] = 8'b0;
    XRAM[23618] = 8'b0;
    XRAM[23619] = 8'b0;
    XRAM[23620] = 8'b0;
    XRAM[23621] = 8'b0;
    XRAM[23622] = 8'b0;
    XRAM[23623] = 8'b0;
    XRAM[23624] = 8'b0;
    XRAM[23625] = 8'b0;
    XRAM[23626] = 8'b0;
    XRAM[23627] = 8'b0;
    XRAM[23628] = 8'b0;
    XRAM[23629] = 8'b0;
    XRAM[23630] = 8'b0;
    XRAM[23631] = 8'b0;
    XRAM[23632] = 8'b0;
    XRAM[23633] = 8'b0;
    XRAM[23634] = 8'b0;
    XRAM[23635] = 8'b0;
    XRAM[23636] = 8'b0;
    XRAM[23637] = 8'b0;
    XRAM[23638] = 8'b0;
    XRAM[23639] = 8'b0;
    XRAM[23640] = 8'b0;
    XRAM[23641] = 8'b0;
    XRAM[23642] = 8'b0;
    XRAM[23643] = 8'b0;
    XRAM[23644] = 8'b0;
    XRAM[23645] = 8'b0;
    XRAM[23646] = 8'b0;
    XRAM[23647] = 8'b0;
    XRAM[23648] = 8'b0;
    XRAM[23649] = 8'b0;
    XRAM[23650] = 8'b0;
    XRAM[23651] = 8'b0;
    XRAM[23652] = 8'b0;
    XRAM[23653] = 8'b0;
    XRAM[23654] = 8'b0;
    XRAM[23655] = 8'b0;
    XRAM[23656] = 8'b0;
    XRAM[23657] = 8'b0;
    XRAM[23658] = 8'b0;
    XRAM[23659] = 8'b0;
    XRAM[23660] = 8'b0;
    XRAM[23661] = 8'b0;
    XRAM[23662] = 8'b0;
    XRAM[23663] = 8'b0;
    XRAM[23664] = 8'b0;
    XRAM[23665] = 8'b0;
    XRAM[23666] = 8'b0;
    XRAM[23667] = 8'b0;
    XRAM[23668] = 8'b0;
    XRAM[23669] = 8'b0;
    XRAM[23670] = 8'b0;
    XRAM[23671] = 8'b0;
    XRAM[23672] = 8'b0;
    XRAM[23673] = 8'b0;
    XRAM[23674] = 8'b0;
    XRAM[23675] = 8'b0;
    XRAM[23676] = 8'b0;
    XRAM[23677] = 8'b0;
    XRAM[23678] = 8'b0;
    XRAM[23679] = 8'b0;
    XRAM[23680] = 8'b0;
    XRAM[23681] = 8'b0;
    XRAM[23682] = 8'b0;
    XRAM[23683] = 8'b0;
    XRAM[23684] = 8'b0;
    XRAM[23685] = 8'b0;
    XRAM[23686] = 8'b0;
    XRAM[23687] = 8'b0;
    XRAM[23688] = 8'b0;
    XRAM[23689] = 8'b0;
    XRAM[23690] = 8'b0;
    XRAM[23691] = 8'b0;
    XRAM[23692] = 8'b0;
    XRAM[23693] = 8'b0;
    XRAM[23694] = 8'b0;
    XRAM[23695] = 8'b0;
    XRAM[23696] = 8'b0;
    XRAM[23697] = 8'b0;
    XRAM[23698] = 8'b0;
    XRAM[23699] = 8'b0;
    XRAM[23700] = 8'b0;
    XRAM[23701] = 8'b0;
    XRAM[23702] = 8'b0;
    XRAM[23703] = 8'b0;
    XRAM[23704] = 8'b0;
    XRAM[23705] = 8'b0;
    XRAM[23706] = 8'b0;
    XRAM[23707] = 8'b0;
    XRAM[23708] = 8'b0;
    XRAM[23709] = 8'b0;
    XRAM[23710] = 8'b0;
    XRAM[23711] = 8'b0;
    XRAM[23712] = 8'b0;
    XRAM[23713] = 8'b0;
    XRAM[23714] = 8'b0;
    XRAM[23715] = 8'b0;
    XRAM[23716] = 8'b0;
    XRAM[23717] = 8'b0;
    XRAM[23718] = 8'b0;
    XRAM[23719] = 8'b0;
    XRAM[23720] = 8'b0;
    XRAM[23721] = 8'b0;
    XRAM[23722] = 8'b0;
    XRAM[23723] = 8'b0;
    XRAM[23724] = 8'b0;
    XRAM[23725] = 8'b0;
    XRAM[23726] = 8'b0;
    XRAM[23727] = 8'b0;
    XRAM[23728] = 8'b0;
    XRAM[23729] = 8'b0;
    XRAM[23730] = 8'b0;
    XRAM[23731] = 8'b0;
    XRAM[23732] = 8'b0;
    XRAM[23733] = 8'b0;
    XRAM[23734] = 8'b0;
    XRAM[23735] = 8'b0;
    XRAM[23736] = 8'b0;
    XRAM[23737] = 8'b0;
    XRAM[23738] = 8'b0;
    XRAM[23739] = 8'b0;
    XRAM[23740] = 8'b0;
    XRAM[23741] = 8'b0;
    XRAM[23742] = 8'b0;
    XRAM[23743] = 8'b0;
    XRAM[23744] = 8'b0;
    XRAM[23745] = 8'b0;
    XRAM[23746] = 8'b0;
    XRAM[23747] = 8'b0;
    XRAM[23748] = 8'b0;
    XRAM[23749] = 8'b0;
    XRAM[23750] = 8'b0;
    XRAM[23751] = 8'b0;
    XRAM[23752] = 8'b0;
    XRAM[23753] = 8'b0;
    XRAM[23754] = 8'b0;
    XRAM[23755] = 8'b0;
    XRAM[23756] = 8'b0;
    XRAM[23757] = 8'b0;
    XRAM[23758] = 8'b0;
    XRAM[23759] = 8'b0;
    XRAM[23760] = 8'b0;
    XRAM[23761] = 8'b0;
    XRAM[23762] = 8'b0;
    XRAM[23763] = 8'b0;
    XRAM[23764] = 8'b0;
    XRAM[23765] = 8'b0;
    XRAM[23766] = 8'b0;
    XRAM[23767] = 8'b0;
    XRAM[23768] = 8'b0;
    XRAM[23769] = 8'b0;
    XRAM[23770] = 8'b0;
    XRAM[23771] = 8'b0;
    XRAM[23772] = 8'b0;
    XRAM[23773] = 8'b0;
    XRAM[23774] = 8'b0;
    XRAM[23775] = 8'b0;
    XRAM[23776] = 8'b0;
    XRAM[23777] = 8'b0;
    XRAM[23778] = 8'b0;
    XRAM[23779] = 8'b0;
    XRAM[23780] = 8'b0;
    XRAM[23781] = 8'b0;
    XRAM[23782] = 8'b0;
    XRAM[23783] = 8'b0;
    XRAM[23784] = 8'b0;
    XRAM[23785] = 8'b0;
    XRAM[23786] = 8'b0;
    XRAM[23787] = 8'b0;
    XRAM[23788] = 8'b0;
    XRAM[23789] = 8'b0;
    XRAM[23790] = 8'b0;
    XRAM[23791] = 8'b0;
    XRAM[23792] = 8'b0;
    XRAM[23793] = 8'b0;
    XRAM[23794] = 8'b0;
    XRAM[23795] = 8'b0;
    XRAM[23796] = 8'b0;
    XRAM[23797] = 8'b0;
    XRAM[23798] = 8'b0;
    XRAM[23799] = 8'b0;
    XRAM[23800] = 8'b0;
    XRAM[23801] = 8'b0;
    XRAM[23802] = 8'b0;
    XRAM[23803] = 8'b0;
    XRAM[23804] = 8'b0;
    XRAM[23805] = 8'b0;
    XRAM[23806] = 8'b0;
    XRAM[23807] = 8'b0;
    XRAM[23808] = 8'b0;
    XRAM[23809] = 8'b0;
    XRAM[23810] = 8'b0;
    XRAM[23811] = 8'b0;
    XRAM[23812] = 8'b0;
    XRAM[23813] = 8'b0;
    XRAM[23814] = 8'b0;
    XRAM[23815] = 8'b0;
    XRAM[23816] = 8'b0;
    XRAM[23817] = 8'b0;
    XRAM[23818] = 8'b0;
    XRAM[23819] = 8'b0;
    XRAM[23820] = 8'b0;
    XRAM[23821] = 8'b0;
    XRAM[23822] = 8'b0;
    XRAM[23823] = 8'b0;
    XRAM[23824] = 8'b0;
    XRAM[23825] = 8'b0;
    XRAM[23826] = 8'b0;
    XRAM[23827] = 8'b0;
    XRAM[23828] = 8'b0;
    XRAM[23829] = 8'b0;
    XRAM[23830] = 8'b0;
    XRAM[23831] = 8'b0;
    XRAM[23832] = 8'b0;
    XRAM[23833] = 8'b0;
    XRAM[23834] = 8'b0;
    XRAM[23835] = 8'b0;
    XRAM[23836] = 8'b0;
    XRAM[23837] = 8'b0;
    XRAM[23838] = 8'b0;
    XRAM[23839] = 8'b0;
    XRAM[23840] = 8'b0;
    XRAM[23841] = 8'b0;
    XRAM[23842] = 8'b0;
    XRAM[23843] = 8'b0;
    XRAM[23844] = 8'b0;
    XRAM[23845] = 8'b0;
    XRAM[23846] = 8'b0;
    XRAM[23847] = 8'b0;
    XRAM[23848] = 8'b0;
    XRAM[23849] = 8'b0;
    XRAM[23850] = 8'b0;
    XRAM[23851] = 8'b0;
    XRAM[23852] = 8'b0;
    XRAM[23853] = 8'b0;
    XRAM[23854] = 8'b0;
    XRAM[23855] = 8'b0;
    XRAM[23856] = 8'b0;
    XRAM[23857] = 8'b0;
    XRAM[23858] = 8'b0;
    XRAM[23859] = 8'b0;
    XRAM[23860] = 8'b0;
    XRAM[23861] = 8'b0;
    XRAM[23862] = 8'b0;
    XRAM[23863] = 8'b0;
    XRAM[23864] = 8'b0;
    XRAM[23865] = 8'b0;
    XRAM[23866] = 8'b0;
    XRAM[23867] = 8'b0;
    XRAM[23868] = 8'b0;
    XRAM[23869] = 8'b0;
    XRAM[23870] = 8'b0;
    XRAM[23871] = 8'b0;
    XRAM[23872] = 8'b0;
    XRAM[23873] = 8'b0;
    XRAM[23874] = 8'b0;
    XRAM[23875] = 8'b0;
    XRAM[23876] = 8'b0;
    XRAM[23877] = 8'b0;
    XRAM[23878] = 8'b0;
    XRAM[23879] = 8'b0;
    XRAM[23880] = 8'b0;
    XRAM[23881] = 8'b0;
    XRAM[23882] = 8'b0;
    XRAM[23883] = 8'b0;
    XRAM[23884] = 8'b0;
    XRAM[23885] = 8'b0;
    XRAM[23886] = 8'b0;
    XRAM[23887] = 8'b0;
    XRAM[23888] = 8'b0;
    XRAM[23889] = 8'b0;
    XRAM[23890] = 8'b0;
    XRAM[23891] = 8'b0;
    XRAM[23892] = 8'b0;
    XRAM[23893] = 8'b0;
    XRAM[23894] = 8'b0;
    XRAM[23895] = 8'b0;
    XRAM[23896] = 8'b0;
    XRAM[23897] = 8'b0;
    XRAM[23898] = 8'b0;
    XRAM[23899] = 8'b0;
    XRAM[23900] = 8'b0;
    XRAM[23901] = 8'b0;
    XRAM[23902] = 8'b0;
    XRAM[23903] = 8'b0;
    XRAM[23904] = 8'b0;
    XRAM[23905] = 8'b0;
    XRAM[23906] = 8'b0;
    XRAM[23907] = 8'b0;
    XRAM[23908] = 8'b0;
    XRAM[23909] = 8'b0;
    XRAM[23910] = 8'b0;
    XRAM[23911] = 8'b0;
    XRAM[23912] = 8'b0;
    XRAM[23913] = 8'b0;
    XRAM[23914] = 8'b0;
    XRAM[23915] = 8'b0;
    XRAM[23916] = 8'b0;
    XRAM[23917] = 8'b0;
    XRAM[23918] = 8'b0;
    XRAM[23919] = 8'b0;
    XRAM[23920] = 8'b0;
    XRAM[23921] = 8'b0;
    XRAM[23922] = 8'b0;
    XRAM[23923] = 8'b0;
    XRAM[23924] = 8'b0;
    XRAM[23925] = 8'b0;
    XRAM[23926] = 8'b0;
    XRAM[23927] = 8'b0;
    XRAM[23928] = 8'b0;
    XRAM[23929] = 8'b0;
    XRAM[23930] = 8'b0;
    XRAM[23931] = 8'b0;
    XRAM[23932] = 8'b0;
    XRAM[23933] = 8'b0;
    XRAM[23934] = 8'b0;
    XRAM[23935] = 8'b0;
    XRAM[23936] = 8'b0;
    XRAM[23937] = 8'b0;
    XRAM[23938] = 8'b0;
    XRAM[23939] = 8'b0;
    XRAM[23940] = 8'b0;
    XRAM[23941] = 8'b0;
    XRAM[23942] = 8'b0;
    XRAM[23943] = 8'b0;
    XRAM[23944] = 8'b0;
    XRAM[23945] = 8'b0;
    XRAM[23946] = 8'b0;
    XRAM[23947] = 8'b0;
    XRAM[23948] = 8'b0;
    XRAM[23949] = 8'b0;
    XRAM[23950] = 8'b0;
    XRAM[23951] = 8'b0;
    XRAM[23952] = 8'b0;
    XRAM[23953] = 8'b0;
    XRAM[23954] = 8'b0;
    XRAM[23955] = 8'b0;
    XRAM[23956] = 8'b0;
    XRAM[23957] = 8'b0;
    XRAM[23958] = 8'b0;
    XRAM[23959] = 8'b0;
    XRAM[23960] = 8'b0;
    XRAM[23961] = 8'b0;
    XRAM[23962] = 8'b0;
    XRAM[23963] = 8'b0;
    XRAM[23964] = 8'b0;
    XRAM[23965] = 8'b0;
    XRAM[23966] = 8'b0;
    XRAM[23967] = 8'b0;
    XRAM[23968] = 8'b0;
    XRAM[23969] = 8'b0;
    XRAM[23970] = 8'b0;
    XRAM[23971] = 8'b0;
    XRAM[23972] = 8'b0;
    XRAM[23973] = 8'b0;
    XRAM[23974] = 8'b0;
    XRAM[23975] = 8'b0;
    XRAM[23976] = 8'b0;
    XRAM[23977] = 8'b0;
    XRAM[23978] = 8'b0;
    XRAM[23979] = 8'b0;
    XRAM[23980] = 8'b0;
    XRAM[23981] = 8'b0;
    XRAM[23982] = 8'b0;
    XRAM[23983] = 8'b0;
    XRAM[23984] = 8'b0;
    XRAM[23985] = 8'b0;
    XRAM[23986] = 8'b0;
    XRAM[23987] = 8'b0;
    XRAM[23988] = 8'b0;
    XRAM[23989] = 8'b0;
    XRAM[23990] = 8'b0;
    XRAM[23991] = 8'b0;
    XRAM[23992] = 8'b0;
    XRAM[23993] = 8'b0;
    XRAM[23994] = 8'b0;
    XRAM[23995] = 8'b0;
    XRAM[23996] = 8'b0;
    XRAM[23997] = 8'b0;
    XRAM[23998] = 8'b0;
    XRAM[23999] = 8'b0;
    XRAM[24000] = 8'b0;
    XRAM[24001] = 8'b0;
    XRAM[24002] = 8'b0;
    XRAM[24003] = 8'b0;
    XRAM[24004] = 8'b0;
    XRAM[24005] = 8'b0;
    XRAM[24006] = 8'b0;
    XRAM[24007] = 8'b0;
    XRAM[24008] = 8'b0;
    XRAM[24009] = 8'b0;
    XRAM[24010] = 8'b0;
    XRAM[24011] = 8'b0;
    XRAM[24012] = 8'b0;
    XRAM[24013] = 8'b0;
    XRAM[24014] = 8'b0;
    XRAM[24015] = 8'b0;
    XRAM[24016] = 8'b0;
    XRAM[24017] = 8'b0;
    XRAM[24018] = 8'b0;
    XRAM[24019] = 8'b0;
    XRAM[24020] = 8'b0;
    XRAM[24021] = 8'b0;
    XRAM[24022] = 8'b0;
    XRAM[24023] = 8'b0;
    XRAM[24024] = 8'b0;
    XRAM[24025] = 8'b0;
    XRAM[24026] = 8'b0;
    XRAM[24027] = 8'b0;
    XRAM[24028] = 8'b0;
    XRAM[24029] = 8'b0;
    XRAM[24030] = 8'b0;
    XRAM[24031] = 8'b0;
    XRAM[24032] = 8'b0;
    XRAM[24033] = 8'b0;
    XRAM[24034] = 8'b0;
    XRAM[24035] = 8'b0;
    XRAM[24036] = 8'b0;
    XRAM[24037] = 8'b0;
    XRAM[24038] = 8'b0;
    XRAM[24039] = 8'b0;
    XRAM[24040] = 8'b0;
    XRAM[24041] = 8'b0;
    XRAM[24042] = 8'b0;
    XRAM[24043] = 8'b0;
    XRAM[24044] = 8'b0;
    XRAM[24045] = 8'b0;
    XRAM[24046] = 8'b0;
    XRAM[24047] = 8'b0;
    XRAM[24048] = 8'b0;
    XRAM[24049] = 8'b0;
    XRAM[24050] = 8'b0;
    XRAM[24051] = 8'b0;
    XRAM[24052] = 8'b0;
    XRAM[24053] = 8'b0;
    XRAM[24054] = 8'b0;
    XRAM[24055] = 8'b0;
    XRAM[24056] = 8'b0;
    XRAM[24057] = 8'b0;
    XRAM[24058] = 8'b0;
    XRAM[24059] = 8'b0;
    XRAM[24060] = 8'b0;
    XRAM[24061] = 8'b0;
    XRAM[24062] = 8'b0;
    XRAM[24063] = 8'b0;
    XRAM[24064] = 8'b0;
    XRAM[24065] = 8'b0;
    XRAM[24066] = 8'b0;
    XRAM[24067] = 8'b0;
    XRAM[24068] = 8'b0;
    XRAM[24069] = 8'b0;
    XRAM[24070] = 8'b0;
    XRAM[24071] = 8'b0;
    XRAM[24072] = 8'b0;
    XRAM[24073] = 8'b0;
    XRAM[24074] = 8'b0;
    XRAM[24075] = 8'b0;
    XRAM[24076] = 8'b0;
    XRAM[24077] = 8'b0;
    XRAM[24078] = 8'b0;
    XRAM[24079] = 8'b0;
    XRAM[24080] = 8'b0;
    XRAM[24081] = 8'b0;
    XRAM[24082] = 8'b0;
    XRAM[24083] = 8'b0;
    XRAM[24084] = 8'b0;
    XRAM[24085] = 8'b0;
    XRAM[24086] = 8'b0;
    XRAM[24087] = 8'b0;
    XRAM[24088] = 8'b0;
    XRAM[24089] = 8'b0;
    XRAM[24090] = 8'b0;
    XRAM[24091] = 8'b0;
    XRAM[24092] = 8'b0;
    XRAM[24093] = 8'b0;
    XRAM[24094] = 8'b0;
    XRAM[24095] = 8'b0;
    XRAM[24096] = 8'b0;
    XRAM[24097] = 8'b0;
    XRAM[24098] = 8'b0;
    XRAM[24099] = 8'b0;
    XRAM[24100] = 8'b0;
    XRAM[24101] = 8'b0;
    XRAM[24102] = 8'b0;
    XRAM[24103] = 8'b0;
    XRAM[24104] = 8'b0;
    XRAM[24105] = 8'b0;
    XRAM[24106] = 8'b0;
    XRAM[24107] = 8'b0;
    XRAM[24108] = 8'b0;
    XRAM[24109] = 8'b0;
    XRAM[24110] = 8'b0;
    XRAM[24111] = 8'b0;
    XRAM[24112] = 8'b0;
    XRAM[24113] = 8'b0;
    XRAM[24114] = 8'b0;
    XRAM[24115] = 8'b0;
    XRAM[24116] = 8'b0;
    XRAM[24117] = 8'b0;
    XRAM[24118] = 8'b0;
    XRAM[24119] = 8'b0;
    XRAM[24120] = 8'b0;
    XRAM[24121] = 8'b0;
    XRAM[24122] = 8'b0;
    XRAM[24123] = 8'b0;
    XRAM[24124] = 8'b0;
    XRAM[24125] = 8'b0;
    XRAM[24126] = 8'b0;
    XRAM[24127] = 8'b0;
    XRAM[24128] = 8'b0;
    XRAM[24129] = 8'b0;
    XRAM[24130] = 8'b0;
    XRAM[24131] = 8'b0;
    XRAM[24132] = 8'b0;
    XRAM[24133] = 8'b0;
    XRAM[24134] = 8'b0;
    XRAM[24135] = 8'b0;
    XRAM[24136] = 8'b0;
    XRAM[24137] = 8'b0;
    XRAM[24138] = 8'b0;
    XRAM[24139] = 8'b0;
    XRAM[24140] = 8'b0;
    XRAM[24141] = 8'b0;
    XRAM[24142] = 8'b0;
    XRAM[24143] = 8'b0;
    XRAM[24144] = 8'b0;
    XRAM[24145] = 8'b0;
    XRAM[24146] = 8'b0;
    XRAM[24147] = 8'b0;
    XRAM[24148] = 8'b0;
    XRAM[24149] = 8'b0;
    XRAM[24150] = 8'b0;
    XRAM[24151] = 8'b0;
    XRAM[24152] = 8'b0;
    XRAM[24153] = 8'b0;
    XRAM[24154] = 8'b0;
    XRAM[24155] = 8'b0;
    XRAM[24156] = 8'b0;
    XRAM[24157] = 8'b0;
    XRAM[24158] = 8'b0;
    XRAM[24159] = 8'b0;
    XRAM[24160] = 8'b0;
    XRAM[24161] = 8'b0;
    XRAM[24162] = 8'b0;
    XRAM[24163] = 8'b0;
    XRAM[24164] = 8'b0;
    XRAM[24165] = 8'b0;
    XRAM[24166] = 8'b0;
    XRAM[24167] = 8'b0;
    XRAM[24168] = 8'b0;
    XRAM[24169] = 8'b0;
    XRAM[24170] = 8'b0;
    XRAM[24171] = 8'b0;
    XRAM[24172] = 8'b0;
    XRAM[24173] = 8'b0;
    XRAM[24174] = 8'b0;
    XRAM[24175] = 8'b0;
    XRAM[24176] = 8'b0;
    XRAM[24177] = 8'b0;
    XRAM[24178] = 8'b0;
    XRAM[24179] = 8'b0;
    XRAM[24180] = 8'b0;
    XRAM[24181] = 8'b0;
    XRAM[24182] = 8'b0;
    XRAM[24183] = 8'b0;
    XRAM[24184] = 8'b0;
    XRAM[24185] = 8'b0;
    XRAM[24186] = 8'b0;
    XRAM[24187] = 8'b0;
    XRAM[24188] = 8'b0;
    XRAM[24189] = 8'b0;
    XRAM[24190] = 8'b0;
    XRAM[24191] = 8'b0;
    XRAM[24192] = 8'b0;
    XRAM[24193] = 8'b0;
    XRAM[24194] = 8'b0;
    XRAM[24195] = 8'b0;
    XRAM[24196] = 8'b0;
    XRAM[24197] = 8'b0;
    XRAM[24198] = 8'b0;
    XRAM[24199] = 8'b0;
    XRAM[24200] = 8'b0;
    XRAM[24201] = 8'b0;
    XRAM[24202] = 8'b0;
    XRAM[24203] = 8'b0;
    XRAM[24204] = 8'b0;
    XRAM[24205] = 8'b0;
    XRAM[24206] = 8'b0;
    XRAM[24207] = 8'b0;
    XRAM[24208] = 8'b0;
    XRAM[24209] = 8'b0;
    XRAM[24210] = 8'b0;
    XRAM[24211] = 8'b0;
    XRAM[24212] = 8'b0;
    XRAM[24213] = 8'b0;
    XRAM[24214] = 8'b0;
    XRAM[24215] = 8'b0;
    XRAM[24216] = 8'b0;
    XRAM[24217] = 8'b0;
    XRAM[24218] = 8'b0;
    XRAM[24219] = 8'b0;
    XRAM[24220] = 8'b0;
    XRAM[24221] = 8'b0;
    XRAM[24222] = 8'b0;
    XRAM[24223] = 8'b0;
    XRAM[24224] = 8'b0;
    XRAM[24225] = 8'b0;
    XRAM[24226] = 8'b0;
    XRAM[24227] = 8'b0;
    XRAM[24228] = 8'b0;
    XRAM[24229] = 8'b0;
    XRAM[24230] = 8'b0;
    XRAM[24231] = 8'b0;
    XRAM[24232] = 8'b0;
    XRAM[24233] = 8'b0;
    XRAM[24234] = 8'b0;
    XRAM[24235] = 8'b0;
    XRAM[24236] = 8'b0;
    XRAM[24237] = 8'b0;
    XRAM[24238] = 8'b0;
    XRAM[24239] = 8'b0;
    XRAM[24240] = 8'b0;
    XRAM[24241] = 8'b0;
    XRAM[24242] = 8'b0;
    XRAM[24243] = 8'b0;
    XRAM[24244] = 8'b0;
    XRAM[24245] = 8'b0;
    XRAM[24246] = 8'b0;
    XRAM[24247] = 8'b0;
    XRAM[24248] = 8'b0;
    XRAM[24249] = 8'b0;
    XRAM[24250] = 8'b0;
    XRAM[24251] = 8'b0;
    XRAM[24252] = 8'b0;
    XRAM[24253] = 8'b0;
    XRAM[24254] = 8'b0;
    XRAM[24255] = 8'b0;
    XRAM[24256] = 8'b0;
    XRAM[24257] = 8'b0;
    XRAM[24258] = 8'b0;
    XRAM[24259] = 8'b0;
    XRAM[24260] = 8'b0;
    XRAM[24261] = 8'b0;
    XRAM[24262] = 8'b0;
    XRAM[24263] = 8'b0;
    XRAM[24264] = 8'b0;
    XRAM[24265] = 8'b0;
    XRAM[24266] = 8'b0;
    XRAM[24267] = 8'b0;
    XRAM[24268] = 8'b0;
    XRAM[24269] = 8'b0;
    XRAM[24270] = 8'b0;
    XRAM[24271] = 8'b0;
    XRAM[24272] = 8'b0;
    XRAM[24273] = 8'b0;
    XRAM[24274] = 8'b0;
    XRAM[24275] = 8'b0;
    XRAM[24276] = 8'b0;
    XRAM[24277] = 8'b0;
    XRAM[24278] = 8'b0;
    XRAM[24279] = 8'b0;
    XRAM[24280] = 8'b0;
    XRAM[24281] = 8'b0;
    XRAM[24282] = 8'b0;
    XRAM[24283] = 8'b0;
    XRAM[24284] = 8'b0;
    XRAM[24285] = 8'b0;
    XRAM[24286] = 8'b0;
    XRAM[24287] = 8'b0;
    XRAM[24288] = 8'b0;
    XRAM[24289] = 8'b0;
    XRAM[24290] = 8'b0;
    XRAM[24291] = 8'b0;
    XRAM[24292] = 8'b0;
    XRAM[24293] = 8'b0;
    XRAM[24294] = 8'b0;
    XRAM[24295] = 8'b0;
    XRAM[24296] = 8'b0;
    XRAM[24297] = 8'b0;
    XRAM[24298] = 8'b0;
    XRAM[24299] = 8'b0;
    XRAM[24300] = 8'b0;
    XRAM[24301] = 8'b0;
    XRAM[24302] = 8'b0;
    XRAM[24303] = 8'b0;
    XRAM[24304] = 8'b0;
    XRAM[24305] = 8'b0;
    XRAM[24306] = 8'b0;
    XRAM[24307] = 8'b0;
    XRAM[24308] = 8'b0;
    XRAM[24309] = 8'b0;
    XRAM[24310] = 8'b0;
    XRAM[24311] = 8'b0;
    XRAM[24312] = 8'b0;
    XRAM[24313] = 8'b0;
    XRAM[24314] = 8'b0;
    XRAM[24315] = 8'b0;
    XRAM[24316] = 8'b0;
    XRAM[24317] = 8'b0;
    XRAM[24318] = 8'b0;
    XRAM[24319] = 8'b0;
    XRAM[24320] = 8'b0;
    XRAM[24321] = 8'b0;
    XRAM[24322] = 8'b0;
    XRAM[24323] = 8'b0;
    XRAM[24324] = 8'b0;
    XRAM[24325] = 8'b0;
    XRAM[24326] = 8'b0;
    XRAM[24327] = 8'b0;
    XRAM[24328] = 8'b0;
    XRAM[24329] = 8'b0;
    XRAM[24330] = 8'b0;
    XRAM[24331] = 8'b0;
    XRAM[24332] = 8'b0;
    XRAM[24333] = 8'b0;
    XRAM[24334] = 8'b0;
    XRAM[24335] = 8'b0;
    XRAM[24336] = 8'b0;
    XRAM[24337] = 8'b0;
    XRAM[24338] = 8'b0;
    XRAM[24339] = 8'b0;
    XRAM[24340] = 8'b0;
    XRAM[24341] = 8'b0;
    XRAM[24342] = 8'b0;
    XRAM[24343] = 8'b0;
    XRAM[24344] = 8'b0;
    XRAM[24345] = 8'b0;
    XRAM[24346] = 8'b0;
    XRAM[24347] = 8'b0;
    XRAM[24348] = 8'b0;
    XRAM[24349] = 8'b0;
    XRAM[24350] = 8'b0;
    XRAM[24351] = 8'b0;
    XRAM[24352] = 8'b0;
    XRAM[24353] = 8'b0;
    XRAM[24354] = 8'b0;
    XRAM[24355] = 8'b0;
    XRAM[24356] = 8'b0;
    XRAM[24357] = 8'b0;
    XRAM[24358] = 8'b0;
    XRAM[24359] = 8'b0;
    XRAM[24360] = 8'b0;
    XRAM[24361] = 8'b0;
    XRAM[24362] = 8'b0;
    XRAM[24363] = 8'b0;
    XRAM[24364] = 8'b0;
    XRAM[24365] = 8'b0;
    XRAM[24366] = 8'b0;
    XRAM[24367] = 8'b0;
    XRAM[24368] = 8'b0;
    XRAM[24369] = 8'b0;
    XRAM[24370] = 8'b0;
    XRAM[24371] = 8'b0;
    XRAM[24372] = 8'b0;
    XRAM[24373] = 8'b0;
    XRAM[24374] = 8'b0;
    XRAM[24375] = 8'b0;
    XRAM[24376] = 8'b0;
    XRAM[24377] = 8'b0;
    XRAM[24378] = 8'b0;
    XRAM[24379] = 8'b0;
    XRAM[24380] = 8'b0;
    XRAM[24381] = 8'b0;
    XRAM[24382] = 8'b0;
    XRAM[24383] = 8'b0;
    XRAM[24384] = 8'b0;
    XRAM[24385] = 8'b0;
    XRAM[24386] = 8'b0;
    XRAM[24387] = 8'b0;
    XRAM[24388] = 8'b0;
    XRAM[24389] = 8'b0;
    XRAM[24390] = 8'b0;
    XRAM[24391] = 8'b0;
    XRAM[24392] = 8'b0;
    XRAM[24393] = 8'b0;
    XRAM[24394] = 8'b0;
    XRAM[24395] = 8'b0;
    XRAM[24396] = 8'b0;
    XRAM[24397] = 8'b0;
    XRAM[24398] = 8'b0;
    XRAM[24399] = 8'b0;
    XRAM[24400] = 8'b0;
    XRAM[24401] = 8'b0;
    XRAM[24402] = 8'b0;
    XRAM[24403] = 8'b0;
    XRAM[24404] = 8'b0;
    XRAM[24405] = 8'b0;
    XRAM[24406] = 8'b0;
    XRAM[24407] = 8'b0;
    XRAM[24408] = 8'b0;
    XRAM[24409] = 8'b0;
    XRAM[24410] = 8'b0;
    XRAM[24411] = 8'b0;
    XRAM[24412] = 8'b0;
    XRAM[24413] = 8'b0;
    XRAM[24414] = 8'b0;
    XRAM[24415] = 8'b0;
    XRAM[24416] = 8'b0;
    XRAM[24417] = 8'b0;
    XRAM[24418] = 8'b0;
    XRAM[24419] = 8'b0;
    XRAM[24420] = 8'b0;
    XRAM[24421] = 8'b0;
    XRAM[24422] = 8'b0;
    XRAM[24423] = 8'b0;
    XRAM[24424] = 8'b0;
    XRAM[24425] = 8'b0;
    XRAM[24426] = 8'b0;
    XRAM[24427] = 8'b0;
    XRAM[24428] = 8'b0;
    XRAM[24429] = 8'b0;
    XRAM[24430] = 8'b0;
    XRAM[24431] = 8'b0;
    XRAM[24432] = 8'b0;
    XRAM[24433] = 8'b0;
    XRAM[24434] = 8'b0;
    XRAM[24435] = 8'b0;
    XRAM[24436] = 8'b0;
    XRAM[24437] = 8'b0;
    XRAM[24438] = 8'b0;
    XRAM[24439] = 8'b0;
    XRAM[24440] = 8'b0;
    XRAM[24441] = 8'b0;
    XRAM[24442] = 8'b0;
    XRAM[24443] = 8'b0;
    XRAM[24444] = 8'b0;
    XRAM[24445] = 8'b0;
    XRAM[24446] = 8'b0;
    XRAM[24447] = 8'b0;
    XRAM[24448] = 8'b0;
    XRAM[24449] = 8'b0;
    XRAM[24450] = 8'b0;
    XRAM[24451] = 8'b0;
    XRAM[24452] = 8'b0;
    XRAM[24453] = 8'b0;
    XRAM[24454] = 8'b0;
    XRAM[24455] = 8'b0;
    XRAM[24456] = 8'b0;
    XRAM[24457] = 8'b0;
    XRAM[24458] = 8'b0;
    XRAM[24459] = 8'b0;
    XRAM[24460] = 8'b0;
    XRAM[24461] = 8'b0;
    XRAM[24462] = 8'b0;
    XRAM[24463] = 8'b0;
    XRAM[24464] = 8'b0;
    XRAM[24465] = 8'b0;
    XRAM[24466] = 8'b0;
    XRAM[24467] = 8'b0;
    XRAM[24468] = 8'b0;
    XRAM[24469] = 8'b0;
    XRAM[24470] = 8'b0;
    XRAM[24471] = 8'b0;
    XRAM[24472] = 8'b0;
    XRAM[24473] = 8'b0;
    XRAM[24474] = 8'b0;
    XRAM[24475] = 8'b0;
    XRAM[24476] = 8'b0;
    XRAM[24477] = 8'b0;
    XRAM[24478] = 8'b0;
    XRAM[24479] = 8'b0;
    XRAM[24480] = 8'b0;
    XRAM[24481] = 8'b0;
    XRAM[24482] = 8'b0;
    XRAM[24483] = 8'b0;
    XRAM[24484] = 8'b0;
    XRAM[24485] = 8'b0;
    XRAM[24486] = 8'b0;
    XRAM[24487] = 8'b0;
    XRAM[24488] = 8'b0;
    XRAM[24489] = 8'b0;
    XRAM[24490] = 8'b0;
    XRAM[24491] = 8'b0;
    XRAM[24492] = 8'b0;
    XRAM[24493] = 8'b0;
    XRAM[24494] = 8'b0;
    XRAM[24495] = 8'b0;
    XRAM[24496] = 8'b0;
    XRAM[24497] = 8'b0;
    XRAM[24498] = 8'b0;
    XRAM[24499] = 8'b0;
    XRAM[24500] = 8'b0;
    XRAM[24501] = 8'b0;
    XRAM[24502] = 8'b0;
    XRAM[24503] = 8'b0;
    XRAM[24504] = 8'b0;
    XRAM[24505] = 8'b0;
    XRAM[24506] = 8'b0;
    XRAM[24507] = 8'b0;
    XRAM[24508] = 8'b0;
    XRAM[24509] = 8'b0;
    XRAM[24510] = 8'b0;
    XRAM[24511] = 8'b0;
    XRAM[24512] = 8'b0;
    XRAM[24513] = 8'b0;
    XRAM[24514] = 8'b0;
    XRAM[24515] = 8'b0;
    XRAM[24516] = 8'b0;
    XRAM[24517] = 8'b0;
    XRAM[24518] = 8'b0;
    XRAM[24519] = 8'b0;
    XRAM[24520] = 8'b0;
    XRAM[24521] = 8'b0;
    XRAM[24522] = 8'b0;
    XRAM[24523] = 8'b0;
    XRAM[24524] = 8'b0;
    XRAM[24525] = 8'b0;
    XRAM[24526] = 8'b0;
    XRAM[24527] = 8'b0;
    XRAM[24528] = 8'b0;
    XRAM[24529] = 8'b0;
    XRAM[24530] = 8'b0;
    XRAM[24531] = 8'b0;
    XRAM[24532] = 8'b0;
    XRAM[24533] = 8'b0;
    XRAM[24534] = 8'b0;
    XRAM[24535] = 8'b0;
    XRAM[24536] = 8'b0;
    XRAM[24537] = 8'b0;
    XRAM[24538] = 8'b0;
    XRAM[24539] = 8'b0;
    XRAM[24540] = 8'b0;
    XRAM[24541] = 8'b0;
    XRAM[24542] = 8'b0;
    XRAM[24543] = 8'b0;
    XRAM[24544] = 8'b0;
    XRAM[24545] = 8'b0;
    XRAM[24546] = 8'b0;
    XRAM[24547] = 8'b0;
    XRAM[24548] = 8'b0;
    XRAM[24549] = 8'b0;
    XRAM[24550] = 8'b0;
    XRAM[24551] = 8'b0;
    XRAM[24552] = 8'b0;
    XRAM[24553] = 8'b0;
    XRAM[24554] = 8'b0;
    XRAM[24555] = 8'b0;
    XRAM[24556] = 8'b0;
    XRAM[24557] = 8'b0;
    XRAM[24558] = 8'b0;
    XRAM[24559] = 8'b0;
    XRAM[24560] = 8'b0;
    XRAM[24561] = 8'b0;
    XRAM[24562] = 8'b0;
    XRAM[24563] = 8'b0;
    XRAM[24564] = 8'b0;
    XRAM[24565] = 8'b0;
    XRAM[24566] = 8'b0;
    XRAM[24567] = 8'b0;
    XRAM[24568] = 8'b0;
    XRAM[24569] = 8'b0;
    XRAM[24570] = 8'b0;
    XRAM[24571] = 8'b0;
    XRAM[24572] = 8'b0;
    XRAM[24573] = 8'b0;
    XRAM[24574] = 8'b0;
    XRAM[24575] = 8'b0;
    XRAM[24576] = 8'b0;
    XRAM[24577] = 8'b0;
    XRAM[24578] = 8'b0;
    XRAM[24579] = 8'b0;
    XRAM[24580] = 8'b0;
    XRAM[24581] = 8'b0;
    XRAM[24582] = 8'b0;
    XRAM[24583] = 8'b0;
    XRAM[24584] = 8'b0;
    XRAM[24585] = 8'b0;
    XRAM[24586] = 8'b0;
    XRAM[24587] = 8'b0;
    XRAM[24588] = 8'b0;
    XRAM[24589] = 8'b0;
    XRAM[24590] = 8'b0;
    XRAM[24591] = 8'b0;
    XRAM[24592] = 8'b0;
    XRAM[24593] = 8'b0;
    XRAM[24594] = 8'b0;
    XRAM[24595] = 8'b0;
    XRAM[24596] = 8'b0;
    XRAM[24597] = 8'b0;
    XRAM[24598] = 8'b0;
    XRAM[24599] = 8'b0;
    XRAM[24600] = 8'b0;
    XRAM[24601] = 8'b0;
    XRAM[24602] = 8'b0;
    XRAM[24603] = 8'b0;
    XRAM[24604] = 8'b0;
    XRAM[24605] = 8'b0;
    XRAM[24606] = 8'b0;
    XRAM[24607] = 8'b0;
    XRAM[24608] = 8'b0;
    XRAM[24609] = 8'b0;
    XRAM[24610] = 8'b0;
    XRAM[24611] = 8'b0;
    XRAM[24612] = 8'b0;
    XRAM[24613] = 8'b0;
    XRAM[24614] = 8'b0;
    XRAM[24615] = 8'b0;
    XRAM[24616] = 8'b0;
    XRAM[24617] = 8'b0;
    XRAM[24618] = 8'b0;
    XRAM[24619] = 8'b0;
    XRAM[24620] = 8'b0;
    XRAM[24621] = 8'b0;
    XRAM[24622] = 8'b0;
    XRAM[24623] = 8'b0;
    XRAM[24624] = 8'b0;
    XRAM[24625] = 8'b0;
    XRAM[24626] = 8'b0;
    XRAM[24627] = 8'b0;
    XRAM[24628] = 8'b0;
    XRAM[24629] = 8'b0;
    XRAM[24630] = 8'b0;
    XRAM[24631] = 8'b0;
    XRAM[24632] = 8'b0;
    XRAM[24633] = 8'b0;
    XRAM[24634] = 8'b0;
    XRAM[24635] = 8'b0;
    XRAM[24636] = 8'b0;
    XRAM[24637] = 8'b0;
    XRAM[24638] = 8'b0;
    XRAM[24639] = 8'b0;
    XRAM[24640] = 8'b0;
    XRAM[24641] = 8'b0;
    XRAM[24642] = 8'b0;
    XRAM[24643] = 8'b0;
    XRAM[24644] = 8'b0;
    XRAM[24645] = 8'b0;
    XRAM[24646] = 8'b0;
    XRAM[24647] = 8'b0;
    XRAM[24648] = 8'b0;
    XRAM[24649] = 8'b0;
    XRAM[24650] = 8'b0;
    XRAM[24651] = 8'b0;
    XRAM[24652] = 8'b0;
    XRAM[24653] = 8'b0;
    XRAM[24654] = 8'b0;
    XRAM[24655] = 8'b0;
    XRAM[24656] = 8'b0;
    XRAM[24657] = 8'b0;
    XRAM[24658] = 8'b0;
    XRAM[24659] = 8'b0;
    XRAM[24660] = 8'b0;
    XRAM[24661] = 8'b0;
    XRAM[24662] = 8'b0;
    XRAM[24663] = 8'b0;
    XRAM[24664] = 8'b0;
    XRAM[24665] = 8'b0;
    XRAM[24666] = 8'b0;
    XRAM[24667] = 8'b0;
    XRAM[24668] = 8'b0;
    XRAM[24669] = 8'b0;
    XRAM[24670] = 8'b0;
    XRAM[24671] = 8'b0;
    XRAM[24672] = 8'b0;
    XRAM[24673] = 8'b0;
    XRAM[24674] = 8'b0;
    XRAM[24675] = 8'b0;
    XRAM[24676] = 8'b0;
    XRAM[24677] = 8'b0;
    XRAM[24678] = 8'b0;
    XRAM[24679] = 8'b0;
    XRAM[24680] = 8'b0;
    XRAM[24681] = 8'b0;
    XRAM[24682] = 8'b0;
    XRAM[24683] = 8'b0;
    XRAM[24684] = 8'b0;
    XRAM[24685] = 8'b0;
    XRAM[24686] = 8'b0;
    XRAM[24687] = 8'b0;
    XRAM[24688] = 8'b0;
    XRAM[24689] = 8'b0;
    XRAM[24690] = 8'b0;
    XRAM[24691] = 8'b0;
    XRAM[24692] = 8'b0;
    XRAM[24693] = 8'b0;
    XRAM[24694] = 8'b0;
    XRAM[24695] = 8'b0;
    XRAM[24696] = 8'b0;
    XRAM[24697] = 8'b0;
    XRAM[24698] = 8'b0;
    XRAM[24699] = 8'b0;
    XRAM[24700] = 8'b0;
    XRAM[24701] = 8'b0;
    XRAM[24702] = 8'b0;
    XRAM[24703] = 8'b0;
    XRAM[24704] = 8'b0;
    XRAM[24705] = 8'b0;
    XRAM[24706] = 8'b0;
    XRAM[24707] = 8'b0;
    XRAM[24708] = 8'b0;
    XRAM[24709] = 8'b0;
    XRAM[24710] = 8'b0;
    XRAM[24711] = 8'b0;
    XRAM[24712] = 8'b0;
    XRAM[24713] = 8'b0;
    XRAM[24714] = 8'b0;
    XRAM[24715] = 8'b0;
    XRAM[24716] = 8'b0;
    XRAM[24717] = 8'b0;
    XRAM[24718] = 8'b0;
    XRAM[24719] = 8'b0;
    XRAM[24720] = 8'b0;
    XRAM[24721] = 8'b0;
    XRAM[24722] = 8'b0;
    XRAM[24723] = 8'b0;
    XRAM[24724] = 8'b0;
    XRAM[24725] = 8'b0;
    XRAM[24726] = 8'b0;
    XRAM[24727] = 8'b0;
    XRAM[24728] = 8'b0;
    XRAM[24729] = 8'b0;
    XRAM[24730] = 8'b0;
    XRAM[24731] = 8'b0;
    XRAM[24732] = 8'b0;
    XRAM[24733] = 8'b0;
    XRAM[24734] = 8'b0;
    XRAM[24735] = 8'b0;
    XRAM[24736] = 8'b0;
    XRAM[24737] = 8'b0;
    XRAM[24738] = 8'b0;
    XRAM[24739] = 8'b0;
    XRAM[24740] = 8'b0;
    XRAM[24741] = 8'b0;
    XRAM[24742] = 8'b0;
    XRAM[24743] = 8'b0;
    XRAM[24744] = 8'b0;
    XRAM[24745] = 8'b0;
    XRAM[24746] = 8'b0;
    XRAM[24747] = 8'b0;
    XRAM[24748] = 8'b0;
    XRAM[24749] = 8'b0;
    XRAM[24750] = 8'b0;
    XRAM[24751] = 8'b0;
    XRAM[24752] = 8'b0;
    XRAM[24753] = 8'b0;
    XRAM[24754] = 8'b0;
    XRAM[24755] = 8'b0;
    XRAM[24756] = 8'b0;
    XRAM[24757] = 8'b0;
    XRAM[24758] = 8'b0;
    XRAM[24759] = 8'b0;
    XRAM[24760] = 8'b0;
    XRAM[24761] = 8'b0;
    XRAM[24762] = 8'b0;
    XRAM[24763] = 8'b0;
    XRAM[24764] = 8'b0;
    XRAM[24765] = 8'b0;
    XRAM[24766] = 8'b0;
    XRAM[24767] = 8'b0;
    XRAM[24768] = 8'b0;
    XRAM[24769] = 8'b0;
    XRAM[24770] = 8'b0;
    XRAM[24771] = 8'b0;
    XRAM[24772] = 8'b0;
    XRAM[24773] = 8'b0;
    XRAM[24774] = 8'b0;
    XRAM[24775] = 8'b0;
    XRAM[24776] = 8'b0;
    XRAM[24777] = 8'b0;
    XRAM[24778] = 8'b0;
    XRAM[24779] = 8'b0;
    XRAM[24780] = 8'b0;
    XRAM[24781] = 8'b0;
    XRAM[24782] = 8'b0;
    XRAM[24783] = 8'b0;
    XRAM[24784] = 8'b0;
    XRAM[24785] = 8'b0;
    XRAM[24786] = 8'b0;
    XRAM[24787] = 8'b0;
    XRAM[24788] = 8'b0;
    XRAM[24789] = 8'b0;
    XRAM[24790] = 8'b0;
    XRAM[24791] = 8'b0;
    XRAM[24792] = 8'b0;
    XRAM[24793] = 8'b0;
    XRAM[24794] = 8'b0;
    XRAM[24795] = 8'b0;
    XRAM[24796] = 8'b0;
    XRAM[24797] = 8'b0;
    XRAM[24798] = 8'b0;
    XRAM[24799] = 8'b0;
    XRAM[24800] = 8'b0;
    XRAM[24801] = 8'b0;
    XRAM[24802] = 8'b0;
    XRAM[24803] = 8'b0;
    XRAM[24804] = 8'b0;
    XRAM[24805] = 8'b0;
    XRAM[24806] = 8'b0;
    XRAM[24807] = 8'b0;
    XRAM[24808] = 8'b0;
    XRAM[24809] = 8'b0;
    XRAM[24810] = 8'b0;
    XRAM[24811] = 8'b0;
    XRAM[24812] = 8'b0;
    XRAM[24813] = 8'b0;
    XRAM[24814] = 8'b0;
    XRAM[24815] = 8'b0;
    XRAM[24816] = 8'b0;
    XRAM[24817] = 8'b0;
    XRAM[24818] = 8'b0;
    XRAM[24819] = 8'b0;
    XRAM[24820] = 8'b0;
    XRAM[24821] = 8'b0;
    XRAM[24822] = 8'b0;
    XRAM[24823] = 8'b0;
    XRAM[24824] = 8'b0;
    XRAM[24825] = 8'b0;
    XRAM[24826] = 8'b0;
    XRAM[24827] = 8'b0;
    XRAM[24828] = 8'b0;
    XRAM[24829] = 8'b0;
    XRAM[24830] = 8'b0;
    XRAM[24831] = 8'b0;
    XRAM[24832] = 8'b0;
    XRAM[24833] = 8'b0;
    XRAM[24834] = 8'b0;
    XRAM[24835] = 8'b0;
    XRAM[24836] = 8'b0;
    XRAM[24837] = 8'b0;
    XRAM[24838] = 8'b0;
    XRAM[24839] = 8'b0;
    XRAM[24840] = 8'b0;
    XRAM[24841] = 8'b0;
    XRAM[24842] = 8'b0;
    XRAM[24843] = 8'b0;
    XRAM[24844] = 8'b0;
    XRAM[24845] = 8'b0;
    XRAM[24846] = 8'b0;
    XRAM[24847] = 8'b0;
    XRAM[24848] = 8'b0;
    XRAM[24849] = 8'b0;
    XRAM[24850] = 8'b0;
    XRAM[24851] = 8'b0;
    XRAM[24852] = 8'b0;
    XRAM[24853] = 8'b0;
    XRAM[24854] = 8'b0;
    XRAM[24855] = 8'b0;
    XRAM[24856] = 8'b0;
    XRAM[24857] = 8'b0;
    XRAM[24858] = 8'b0;
    XRAM[24859] = 8'b0;
    XRAM[24860] = 8'b0;
    XRAM[24861] = 8'b0;
    XRAM[24862] = 8'b0;
    XRAM[24863] = 8'b0;
    XRAM[24864] = 8'b0;
    XRAM[24865] = 8'b0;
    XRAM[24866] = 8'b0;
    XRAM[24867] = 8'b0;
    XRAM[24868] = 8'b0;
    XRAM[24869] = 8'b0;
    XRAM[24870] = 8'b0;
    XRAM[24871] = 8'b0;
    XRAM[24872] = 8'b0;
    XRAM[24873] = 8'b0;
    XRAM[24874] = 8'b0;
    XRAM[24875] = 8'b0;
    XRAM[24876] = 8'b0;
    XRAM[24877] = 8'b0;
    XRAM[24878] = 8'b0;
    XRAM[24879] = 8'b0;
    XRAM[24880] = 8'b0;
    XRAM[24881] = 8'b0;
    XRAM[24882] = 8'b0;
    XRAM[24883] = 8'b0;
    XRAM[24884] = 8'b0;
    XRAM[24885] = 8'b0;
    XRAM[24886] = 8'b0;
    XRAM[24887] = 8'b0;
    XRAM[24888] = 8'b0;
    XRAM[24889] = 8'b0;
    XRAM[24890] = 8'b0;
    XRAM[24891] = 8'b0;
    XRAM[24892] = 8'b0;
    XRAM[24893] = 8'b0;
    XRAM[24894] = 8'b0;
    XRAM[24895] = 8'b0;
    XRAM[24896] = 8'b0;
    XRAM[24897] = 8'b0;
    XRAM[24898] = 8'b0;
    XRAM[24899] = 8'b0;
    XRAM[24900] = 8'b0;
    XRAM[24901] = 8'b0;
    XRAM[24902] = 8'b0;
    XRAM[24903] = 8'b0;
    XRAM[24904] = 8'b0;
    XRAM[24905] = 8'b0;
    XRAM[24906] = 8'b0;
    XRAM[24907] = 8'b0;
    XRAM[24908] = 8'b0;
    XRAM[24909] = 8'b0;
    XRAM[24910] = 8'b0;
    XRAM[24911] = 8'b0;
    XRAM[24912] = 8'b0;
    XRAM[24913] = 8'b0;
    XRAM[24914] = 8'b0;
    XRAM[24915] = 8'b0;
    XRAM[24916] = 8'b0;
    XRAM[24917] = 8'b0;
    XRAM[24918] = 8'b0;
    XRAM[24919] = 8'b0;
    XRAM[24920] = 8'b0;
    XRAM[24921] = 8'b0;
    XRAM[24922] = 8'b0;
    XRAM[24923] = 8'b0;
    XRAM[24924] = 8'b0;
    XRAM[24925] = 8'b0;
    XRAM[24926] = 8'b0;
    XRAM[24927] = 8'b0;
    XRAM[24928] = 8'b0;
    XRAM[24929] = 8'b0;
    XRAM[24930] = 8'b0;
    XRAM[24931] = 8'b0;
    XRAM[24932] = 8'b0;
    XRAM[24933] = 8'b0;
    XRAM[24934] = 8'b0;
    XRAM[24935] = 8'b0;
    XRAM[24936] = 8'b0;
    XRAM[24937] = 8'b0;
    XRAM[24938] = 8'b0;
    XRAM[24939] = 8'b0;
    XRAM[24940] = 8'b0;
    XRAM[24941] = 8'b0;
    XRAM[24942] = 8'b0;
    XRAM[24943] = 8'b0;
    XRAM[24944] = 8'b0;
    XRAM[24945] = 8'b0;
    XRAM[24946] = 8'b0;
    XRAM[24947] = 8'b0;
    XRAM[24948] = 8'b0;
    XRAM[24949] = 8'b0;
    XRAM[24950] = 8'b0;
    XRAM[24951] = 8'b0;
    XRAM[24952] = 8'b0;
    XRAM[24953] = 8'b0;
    XRAM[24954] = 8'b0;
    XRAM[24955] = 8'b0;
    XRAM[24956] = 8'b0;
    XRAM[24957] = 8'b0;
    XRAM[24958] = 8'b0;
    XRAM[24959] = 8'b0;
    XRAM[24960] = 8'b0;
    XRAM[24961] = 8'b0;
    XRAM[24962] = 8'b0;
    XRAM[24963] = 8'b0;
    XRAM[24964] = 8'b0;
    XRAM[24965] = 8'b0;
    XRAM[24966] = 8'b0;
    XRAM[24967] = 8'b0;
    XRAM[24968] = 8'b0;
    XRAM[24969] = 8'b0;
    XRAM[24970] = 8'b0;
    XRAM[24971] = 8'b0;
    XRAM[24972] = 8'b0;
    XRAM[24973] = 8'b0;
    XRAM[24974] = 8'b0;
    XRAM[24975] = 8'b0;
    XRAM[24976] = 8'b0;
    XRAM[24977] = 8'b0;
    XRAM[24978] = 8'b0;
    XRAM[24979] = 8'b0;
    XRAM[24980] = 8'b0;
    XRAM[24981] = 8'b0;
    XRAM[24982] = 8'b0;
    XRAM[24983] = 8'b0;
    XRAM[24984] = 8'b0;
    XRAM[24985] = 8'b0;
    XRAM[24986] = 8'b0;
    XRAM[24987] = 8'b0;
    XRAM[24988] = 8'b0;
    XRAM[24989] = 8'b0;
    XRAM[24990] = 8'b0;
    XRAM[24991] = 8'b0;
    XRAM[24992] = 8'b0;
    XRAM[24993] = 8'b0;
    XRAM[24994] = 8'b0;
    XRAM[24995] = 8'b0;
    XRAM[24996] = 8'b0;
    XRAM[24997] = 8'b0;
    XRAM[24998] = 8'b0;
    XRAM[24999] = 8'b0;
    XRAM[25000] = 8'b0;
    XRAM[25001] = 8'b0;
    XRAM[25002] = 8'b0;
    XRAM[25003] = 8'b0;
    XRAM[25004] = 8'b0;
    XRAM[25005] = 8'b0;
    XRAM[25006] = 8'b0;
    XRAM[25007] = 8'b0;
    XRAM[25008] = 8'b0;
    XRAM[25009] = 8'b0;
    XRAM[25010] = 8'b0;
    XRAM[25011] = 8'b0;
    XRAM[25012] = 8'b0;
    XRAM[25013] = 8'b0;
    XRAM[25014] = 8'b0;
    XRAM[25015] = 8'b0;
    XRAM[25016] = 8'b0;
    XRAM[25017] = 8'b0;
    XRAM[25018] = 8'b0;
    XRAM[25019] = 8'b0;
    XRAM[25020] = 8'b0;
    XRAM[25021] = 8'b0;
    XRAM[25022] = 8'b0;
    XRAM[25023] = 8'b0;
    XRAM[25024] = 8'b0;
    XRAM[25025] = 8'b0;
    XRAM[25026] = 8'b0;
    XRAM[25027] = 8'b0;
    XRAM[25028] = 8'b0;
    XRAM[25029] = 8'b0;
    XRAM[25030] = 8'b0;
    XRAM[25031] = 8'b0;
    XRAM[25032] = 8'b0;
    XRAM[25033] = 8'b0;
    XRAM[25034] = 8'b0;
    XRAM[25035] = 8'b0;
    XRAM[25036] = 8'b0;
    XRAM[25037] = 8'b0;
    XRAM[25038] = 8'b0;
    XRAM[25039] = 8'b0;
    XRAM[25040] = 8'b0;
    XRAM[25041] = 8'b0;
    XRAM[25042] = 8'b0;
    XRAM[25043] = 8'b0;
    XRAM[25044] = 8'b0;
    XRAM[25045] = 8'b0;
    XRAM[25046] = 8'b0;
    XRAM[25047] = 8'b0;
    XRAM[25048] = 8'b0;
    XRAM[25049] = 8'b0;
    XRAM[25050] = 8'b0;
    XRAM[25051] = 8'b0;
    XRAM[25052] = 8'b0;
    XRAM[25053] = 8'b0;
    XRAM[25054] = 8'b0;
    XRAM[25055] = 8'b0;
    XRAM[25056] = 8'b0;
    XRAM[25057] = 8'b0;
    XRAM[25058] = 8'b0;
    XRAM[25059] = 8'b0;
    XRAM[25060] = 8'b0;
    XRAM[25061] = 8'b0;
    XRAM[25062] = 8'b0;
    XRAM[25063] = 8'b0;
    XRAM[25064] = 8'b0;
    XRAM[25065] = 8'b0;
    XRAM[25066] = 8'b0;
    XRAM[25067] = 8'b0;
    XRAM[25068] = 8'b0;
    XRAM[25069] = 8'b0;
    XRAM[25070] = 8'b0;
    XRAM[25071] = 8'b0;
    XRAM[25072] = 8'b0;
    XRAM[25073] = 8'b0;
    XRAM[25074] = 8'b0;
    XRAM[25075] = 8'b0;
    XRAM[25076] = 8'b0;
    XRAM[25077] = 8'b0;
    XRAM[25078] = 8'b0;
    XRAM[25079] = 8'b0;
    XRAM[25080] = 8'b0;
    XRAM[25081] = 8'b0;
    XRAM[25082] = 8'b0;
    XRAM[25083] = 8'b0;
    XRAM[25084] = 8'b0;
    XRAM[25085] = 8'b0;
    XRAM[25086] = 8'b0;
    XRAM[25087] = 8'b0;
    XRAM[25088] = 8'b0;
    XRAM[25089] = 8'b0;
    XRAM[25090] = 8'b0;
    XRAM[25091] = 8'b0;
    XRAM[25092] = 8'b0;
    XRAM[25093] = 8'b0;
    XRAM[25094] = 8'b0;
    XRAM[25095] = 8'b0;
    XRAM[25096] = 8'b0;
    XRAM[25097] = 8'b0;
    XRAM[25098] = 8'b0;
    XRAM[25099] = 8'b0;
    XRAM[25100] = 8'b0;
    XRAM[25101] = 8'b0;
    XRAM[25102] = 8'b0;
    XRAM[25103] = 8'b0;
    XRAM[25104] = 8'b0;
    XRAM[25105] = 8'b0;
    XRAM[25106] = 8'b0;
    XRAM[25107] = 8'b0;
    XRAM[25108] = 8'b0;
    XRAM[25109] = 8'b0;
    XRAM[25110] = 8'b0;
    XRAM[25111] = 8'b0;
    XRAM[25112] = 8'b0;
    XRAM[25113] = 8'b0;
    XRAM[25114] = 8'b0;
    XRAM[25115] = 8'b0;
    XRAM[25116] = 8'b0;
    XRAM[25117] = 8'b0;
    XRAM[25118] = 8'b0;
    XRAM[25119] = 8'b0;
    XRAM[25120] = 8'b0;
    XRAM[25121] = 8'b0;
    XRAM[25122] = 8'b0;
    XRAM[25123] = 8'b0;
    XRAM[25124] = 8'b0;
    XRAM[25125] = 8'b0;
    XRAM[25126] = 8'b0;
    XRAM[25127] = 8'b0;
    XRAM[25128] = 8'b0;
    XRAM[25129] = 8'b0;
    XRAM[25130] = 8'b0;
    XRAM[25131] = 8'b0;
    XRAM[25132] = 8'b0;
    XRAM[25133] = 8'b0;
    XRAM[25134] = 8'b0;
    XRAM[25135] = 8'b0;
    XRAM[25136] = 8'b0;
    XRAM[25137] = 8'b0;
    XRAM[25138] = 8'b0;
    XRAM[25139] = 8'b0;
    XRAM[25140] = 8'b0;
    XRAM[25141] = 8'b0;
    XRAM[25142] = 8'b0;
    XRAM[25143] = 8'b0;
    XRAM[25144] = 8'b0;
    XRAM[25145] = 8'b0;
    XRAM[25146] = 8'b0;
    XRAM[25147] = 8'b0;
    XRAM[25148] = 8'b0;
    XRAM[25149] = 8'b0;
    XRAM[25150] = 8'b0;
    XRAM[25151] = 8'b0;
    XRAM[25152] = 8'b0;
    XRAM[25153] = 8'b0;
    XRAM[25154] = 8'b0;
    XRAM[25155] = 8'b0;
    XRAM[25156] = 8'b0;
    XRAM[25157] = 8'b0;
    XRAM[25158] = 8'b0;
    XRAM[25159] = 8'b0;
    XRAM[25160] = 8'b0;
    XRAM[25161] = 8'b0;
    XRAM[25162] = 8'b0;
    XRAM[25163] = 8'b0;
    XRAM[25164] = 8'b0;
    XRAM[25165] = 8'b0;
    XRAM[25166] = 8'b0;
    XRAM[25167] = 8'b0;
    XRAM[25168] = 8'b0;
    XRAM[25169] = 8'b0;
    XRAM[25170] = 8'b0;
    XRAM[25171] = 8'b0;
    XRAM[25172] = 8'b0;
    XRAM[25173] = 8'b0;
    XRAM[25174] = 8'b0;
    XRAM[25175] = 8'b0;
    XRAM[25176] = 8'b0;
    XRAM[25177] = 8'b0;
    XRAM[25178] = 8'b0;
    XRAM[25179] = 8'b0;
    XRAM[25180] = 8'b0;
    XRAM[25181] = 8'b0;
    XRAM[25182] = 8'b0;
    XRAM[25183] = 8'b0;
    XRAM[25184] = 8'b0;
    XRAM[25185] = 8'b0;
    XRAM[25186] = 8'b0;
    XRAM[25187] = 8'b0;
    XRAM[25188] = 8'b0;
    XRAM[25189] = 8'b0;
    XRAM[25190] = 8'b0;
    XRAM[25191] = 8'b0;
    XRAM[25192] = 8'b0;
    XRAM[25193] = 8'b0;
    XRAM[25194] = 8'b0;
    XRAM[25195] = 8'b0;
    XRAM[25196] = 8'b0;
    XRAM[25197] = 8'b0;
    XRAM[25198] = 8'b0;
    XRAM[25199] = 8'b0;
    XRAM[25200] = 8'b0;
    XRAM[25201] = 8'b0;
    XRAM[25202] = 8'b0;
    XRAM[25203] = 8'b0;
    XRAM[25204] = 8'b0;
    XRAM[25205] = 8'b0;
    XRAM[25206] = 8'b0;
    XRAM[25207] = 8'b0;
    XRAM[25208] = 8'b0;
    XRAM[25209] = 8'b0;
    XRAM[25210] = 8'b0;
    XRAM[25211] = 8'b0;
    XRAM[25212] = 8'b0;
    XRAM[25213] = 8'b0;
    XRAM[25214] = 8'b0;
    XRAM[25215] = 8'b0;
    XRAM[25216] = 8'b0;
    XRAM[25217] = 8'b0;
    XRAM[25218] = 8'b0;
    XRAM[25219] = 8'b0;
    XRAM[25220] = 8'b0;
    XRAM[25221] = 8'b0;
    XRAM[25222] = 8'b0;
    XRAM[25223] = 8'b0;
    XRAM[25224] = 8'b0;
    XRAM[25225] = 8'b0;
    XRAM[25226] = 8'b0;
    XRAM[25227] = 8'b0;
    XRAM[25228] = 8'b0;
    XRAM[25229] = 8'b0;
    XRAM[25230] = 8'b0;
    XRAM[25231] = 8'b0;
    XRAM[25232] = 8'b0;
    XRAM[25233] = 8'b0;
    XRAM[25234] = 8'b0;
    XRAM[25235] = 8'b0;
    XRAM[25236] = 8'b0;
    XRAM[25237] = 8'b0;
    XRAM[25238] = 8'b0;
    XRAM[25239] = 8'b0;
    XRAM[25240] = 8'b0;
    XRAM[25241] = 8'b0;
    XRAM[25242] = 8'b0;
    XRAM[25243] = 8'b0;
    XRAM[25244] = 8'b0;
    XRAM[25245] = 8'b0;
    XRAM[25246] = 8'b0;
    XRAM[25247] = 8'b0;
    XRAM[25248] = 8'b0;
    XRAM[25249] = 8'b0;
    XRAM[25250] = 8'b0;
    XRAM[25251] = 8'b0;
    XRAM[25252] = 8'b0;
    XRAM[25253] = 8'b0;
    XRAM[25254] = 8'b0;
    XRAM[25255] = 8'b0;
    XRAM[25256] = 8'b0;
    XRAM[25257] = 8'b0;
    XRAM[25258] = 8'b0;
    XRAM[25259] = 8'b0;
    XRAM[25260] = 8'b0;
    XRAM[25261] = 8'b0;
    XRAM[25262] = 8'b0;
    XRAM[25263] = 8'b0;
    XRAM[25264] = 8'b0;
    XRAM[25265] = 8'b0;
    XRAM[25266] = 8'b0;
    XRAM[25267] = 8'b0;
    XRAM[25268] = 8'b0;
    XRAM[25269] = 8'b0;
    XRAM[25270] = 8'b0;
    XRAM[25271] = 8'b0;
    XRAM[25272] = 8'b0;
    XRAM[25273] = 8'b0;
    XRAM[25274] = 8'b0;
    XRAM[25275] = 8'b0;
    XRAM[25276] = 8'b0;
    XRAM[25277] = 8'b0;
    XRAM[25278] = 8'b0;
    XRAM[25279] = 8'b0;
    XRAM[25280] = 8'b0;
    XRAM[25281] = 8'b0;
    XRAM[25282] = 8'b0;
    XRAM[25283] = 8'b0;
    XRAM[25284] = 8'b0;
    XRAM[25285] = 8'b0;
    XRAM[25286] = 8'b0;
    XRAM[25287] = 8'b0;
    XRAM[25288] = 8'b0;
    XRAM[25289] = 8'b0;
    XRAM[25290] = 8'b0;
    XRAM[25291] = 8'b0;
    XRAM[25292] = 8'b0;
    XRAM[25293] = 8'b0;
    XRAM[25294] = 8'b0;
    XRAM[25295] = 8'b0;
    XRAM[25296] = 8'b0;
    XRAM[25297] = 8'b0;
    XRAM[25298] = 8'b0;
    XRAM[25299] = 8'b0;
    XRAM[25300] = 8'b0;
    XRAM[25301] = 8'b0;
    XRAM[25302] = 8'b0;
    XRAM[25303] = 8'b0;
    XRAM[25304] = 8'b0;
    XRAM[25305] = 8'b0;
    XRAM[25306] = 8'b0;
    XRAM[25307] = 8'b0;
    XRAM[25308] = 8'b0;
    XRAM[25309] = 8'b0;
    XRAM[25310] = 8'b0;
    XRAM[25311] = 8'b0;
    XRAM[25312] = 8'b0;
    XRAM[25313] = 8'b0;
    XRAM[25314] = 8'b0;
    XRAM[25315] = 8'b0;
    XRAM[25316] = 8'b0;
    XRAM[25317] = 8'b0;
    XRAM[25318] = 8'b0;
    XRAM[25319] = 8'b0;
    XRAM[25320] = 8'b0;
    XRAM[25321] = 8'b0;
    XRAM[25322] = 8'b0;
    XRAM[25323] = 8'b0;
    XRAM[25324] = 8'b0;
    XRAM[25325] = 8'b0;
    XRAM[25326] = 8'b0;
    XRAM[25327] = 8'b0;
    XRAM[25328] = 8'b0;
    XRAM[25329] = 8'b0;
    XRAM[25330] = 8'b0;
    XRAM[25331] = 8'b0;
    XRAM[25332] = 8'b0;
    XRAM[25333] = 8'b0;
    XRAM[25334] = 8'b0;
    XRAM[25335] = 8'b0;
    XRAM[25336] = 8'b0;
    XRAM[25337] = 8'b0;
    XRAM[25338] = 8'b0;
    XRAM[25339] = 8'b0;
    XRAM[25340] = 8'b0;
    XRAM[25341] = 8'b0;
    XRAM[25342] = 8'b0;
    XRAM[25343] = 8'b0;
    XRAM[25344] = 8'b0;
    XRAM[25345] = 8'b0;
    XRAM[25346] = 8'b0;
    XRAM[25347] = 8'b0;
    XRAM[25348] = 8'b0;
    XRAM[25349] = 8'b0;
    XRAM[25350] = 8'b0;
    XRAM[25351] = 8'b0;
    XRAM[25352] = 8'b0;
    XRAM[25353] = 8'b0;
    XRAM[25354] = 8'b0;
    XRAM[25355] = 8'b0;
    XRAM[25356] = 8'b0;
    XRAM[25357] = 8'b0;
    XRAM[25358] = 8'b0;
    XRAM[25359] = 8'b0;
    XRAM[25360] = 8'b0;
    XRAM[25361] = 8'b0;
    XRAM[25362] = 8'b0;
    XRAM[25363] = 8'b0;
    XRAM[25364] = 8'b0;
    XRAM[25365] = 8'b0;
    XRAM[25366] = 8'b0;
    XRAM[25367] = 8'b0;
    XRAM[25368] = 8'b0;
    XRAM[25369] = 8'b0;
    XRAM[25370] = 8'b0;
    XRAM[25371] = 8'b0;
    XRAM[25372] = 8'b0;
    XRAM[25373] = 8'b0;
    XRAM[25374] = 8'b0;
    XRAM[25375] = 8'b0;
    XRAM[25376] = 8'b0;
    XRAM[25377] = 8'b0;
    XRAM[25378] = 8'b0;
    XRAM[25379] = 8'b0;
    XRAM[25380] = 8'b0;
    XRAM[25381] = 8'b0;
    XRAM[25382] = 8'b0;
    XRAM[25383] = 8'b0;
    XRAM[25384] = 8'b0;
    XRAM[25385] = 8'b0;
    XRAM[25386] = 8'b0;
    XRAM[25387] = 8'b0;
    XRAM[25388] = 8'b0;
    XRAM[25389] = 8'b0;
    XRAM[25390] = 8'b0;
    XRAM[25391] = 8'b0;
    XRAM[25392] = 8'b0;
    XRAM[25393] = 8'b0;
    XRAM[25394] = 8'b0;
    XRAM[25395] = 8'b0;
    XRAM[25396] = 8'b0;
    XRAM[25397] = 8'b0;
    XRAM[25398] = 8'b0;
    XRAM[25399] = 8'b0;
    XRAM[25400] = 8'b0;
    XRAM[25401] = 8'b0;
    XRAM[25402] = 8'b0;
    XRAM[25403] = 8'b0;
    XRAM[25404] = 8'b0;
    XRAM[25405] = 8'b0;
    XRAM[25406] = 8'b0;
    XRAM[25407] = 8'b0;
    XRAM[25408] = 8'b0;
    XRAM[25409] = 8'b0;
    XRAM[25410] = 8'b0;
    XRAM[25411] = 8'b0;
    XRAM[25412] = 8'b0;
    XRAM[25413] = 8'b0;
    XRAM[25414] = 8'b0;
    XRAM[25415] = 8'b0;
    XRAM[25416] = 8'b0;
    XRAM[25417] = 8'b0;
    XRAM[25418] = 8'b0;
    XRAM[25419] = 8'b0;
    XRAM[25420] = 8'b0;
    XRAM[25421] = 8'b0;
    XRAM[25422] = 8'b0;
    XRAM[25423] = 8'b0;
    XRAM[25424] = 8'b0;
    XRAM[25425] = 8'b0;
    XRAM[25426] = 8'b0;
    XRAM[25427] = 8'b0;
    XRAM[25428] = 8'b0;
    XRAM[25429] = 8'b0;
    XRAM[25430] = 8'b0;
    XRAM[25431] = 8'b0;
    XRAM[25432] = 8'b0;
    XRAM[25433] = 8'b0;
    XRAM[25434] = 8'b0;
    XRAM[25435] = 8'b0;
    XRAM[25436] = 8'b0;
    XRAM[25437] = 8'b0;
    XRAM[25438] = 8'b0;
    XRAM[25439] = 8'b0;
    XRAM[25440] = 8'b0;
    XRAM[25441] = 8'b0;
    XRAM[25442] = 8'b0;
    XRAM[25443] = 8'b0;
    XRAM[25444] = 8'b0;
    XRAM[25445] = 8'b0;
    XRAM[25446] = 8'b0;
    XRAM[25447] = 8'b0;
    XRAM[25448] = 8'b0;
    XRAM[25449] = 8'b0;
    XRAM[25450] = 8'b0;
    XRAM[25451] = 8'b0;
    XRAM[25452] = 8'b0;
    XRAM[25453] = 8'b0;
    XRAM[25454] = 8'b0;
    XRAM[25455] = 8'b0;
    XRAM[25456] = 8'b0;
    XRAM[25457] = 8'b0;
    XRAM[25458] = 8'b0;
    XRAM[25459] = 8'b0;
    XRAM[25460] = 8'b0;
    XRAM[25461] = 8'b0;
    XRAM[25462] = 8'b0;
    XRAM[25463] = 8'b0;
    XRAM[25464] = 8'b0;
    XRAM[25465] = 8'b0;
    XRAM[25466] = 8'b0;
    XRAM[25467] = 8'b0;
    XRAM[25468] = 8'b0;
    XRAM[25469] = 8'b0;
    XRAM[25470] = 8'b0;
    XRAM[25471] = 8'b0;
    XRAM[25472] = 8'b0;
    XRAM[25473] = 8'b0;
    XRAM[25474] = 8'b0;
    XRAM[25475] = 8'b0;
    XRAM[25476] = 8'b0;
    XRAM[25477] = 8'b0;
    XRAM[25478] = 8'b0;
    XRAM[25479] = 8'b0;
    XRAM[25480] = 8'b0;
    XRAM[25481] = 8'b0;
    XRAM[25482] = 8'b0;
    XRAM[25483] = 8'b0;
    XRAM[25484] = 8'b0;
    XRAM[25485] = 8'b0;
    XRAM[25486] = 8'b0;
    XRAM[25487] = 8'b0;
    XRAM[25488] = 8'b0;
    XRAM[25489] = 8'b0;
    XRAM[25490] = 8'b0;
    XRAM[25491] = 8'b0;
    XRAM[25492] = 8'b0;
    XRAM[25493] = 8'b0;
    XRAM[25494] = 8'b0;
    XRAM[25495] = 8'b0;
    XRAM[25496] = 8'b0;
    XRAM[25497] = 8'b0;
    XRAM[25498] = 8'b0;
    XRAM[25499] = 8'b0;
    XRAM[25500] = 8'b0;
    XRAM[25501] = 8'b0;
    XRAM[25502] = 8'b0;
    XRAM[25503] = 8'b0;
    XRAM[25504] = 8'b0;
    XRAM[25505] = 8'b0;
    XRAM[25506] = 8'b0;
    XRAM[25507] = 8'b0;
    XRAM[25508] = 8'b0;
    XRAM[25509] = 8'b0;
    XRAM[25510] = 8'b0;
    XRAM[25511] = 8'b0;
    XRAM[25512] = 8'b0;
    XRAM[25513] = 8'b0;
    XRAM[25514] = 8'b0;
    XRAM[25515] = 8'b0;
    XRAM[25516] = 8'b0;
    XRAM[25517] = 8'b0;
    XRAM[25518] = 8'b0;
    XRAM[25519] = 8'b0;
    XRAM[25520] = 8'b0;
    XRAM[25521] = 8'b0;
    XRAM[25522] = 8'b0;
    XRAM[25523] = 8'b0;
    XRAM[25524] = 8'b0;
    XRAM[25525] = 8'b0;
    XRAM[25526] = 8'b0;
    XRAM[25527] = 8'b0;
    XRAM[25528] = 8'b0;
    XRAM[25529] = 8'b0;
    XRAM[25530] = 8'b0;
    XRAM[25531] = 8'b0;
    XRAM[25532] = 8'b0;
    XRAM[25533] = 8'b0;
    XRAM[25534] = 8'b0;
    XRAM[25535] = 8'b0;
    XRAM[25536] = 8'b0;
    XRAM[25537] = 8'b0;
    XRAM[25538] = 8'b0;
    XRAM[25539] = 8'b0;
    XRAM[25540] = 8'b0;
    XRAM[25541] = 8'b0;
    XRAM[25542] = 8'b0;
    XRAM[25543] = 8'b0;
    XRAM[25544] = 8'b0;
    XRAM[25545] = 8'b0;
    XRAM[25546] = 8'b0;
    XRAM[25547] = 8'b0;
    XRAM[25548] = 8'b0;
    XRAM[25549] = 8'b0;
    XRAM[25550] = 8'b0;
    XRAM[25551] = 8'b0;
    XRAM[25552] = 8'b0;
    XRAM[25553] = 8'b0;
    XRAM[25554] = 8'b0;
    XRAM[25555] = 8'b0;
    XRAM[25556] = 8'b0;
    XRAM[25557] = 8'b0;
    XRAM[25558] = 8'b0;
    XRAM[25559] = 8'b0;
    XRAM[25560] = 8'b0;
    XRAM[25561] = 8'b0;
    XRAM[25562] = 8'b0;
    XRAM[25563] = 8'b0;
    XRAM[25564] = 8'b0;
    XRAM[25565] = 8'b0;
    XRAM[25566] = 8'b0;
    XRAM[25567] = 8'b0;
    XRAM[25568] = 8'b0;
    XRAM[25569] = 8'b0;
    XRAM[25570] = 8'b0;
    XRAM[25571] = 8'b0;
    XRAM[25572] = 8'b0;
    XRAM[25573] = 8'b0;
    XRAM[25574] = 8'b0;
    XRAM[25575] = 8'b0;
    XRAM[25576] = 8'b0;
    XRAM[25577] = 8'b0;
    XRAM[25578] = 8'b0;
    XRAM[25579] = 8'b0;
    XRAM[25580] = 8'b0;
    XRAM[25581] = 8'b0;
    XRAM[25582] = 8'b0;
    XRAM[25583] = 8'b0;
    XRAM[25584] = 8'b0;
    XRAM[25585] = 8'b0;
    XRAM[25586] = 8'b0;
    XRAM[25587] = 8'b0;
    XRAM[25588] = 8'b0;
    XRAM[25589] = 8'b0;
    XRAM[25590] = 8'b0;
    XRAM[25591] = 8'b0;
    XRAM[25592] = 8'b0;
    XRAM[25593] = 8'b0;
    XRAM[25594] = 8'b0;
    XRAM[25595] = 8'b0;
    XRAM[25596] = 8'b0;
    XRAM[25597] = 8'b0;
    XRAM[25598] = 8'b0;
    XRAM[25599] = 8'b0;
    XRAM[25600] = 8'b0;
    XRAM[25601] = 8'b0;
    XRAM[25602] = 8'b0;
    XRAM[25603] = 8'b0;
    XRAM[25604] = 8'b0;
    XRAM[25605] = 8'b0;
    XRAM[25606] = 8'b0;
    XRAM[25607] = 8'b0;
    XRAM[25608] = 8'b0;
    XRAM[25609] = 8'b0;
    XRAM[25610] = 8'b0;
    XRAM[25611] = 8'b0;
    XRAM[25612] = 8'b0;
    XRAM[25613] = 8'b0;
    XRAM[25614] = 8'b0;
    XRAM[25615] = 8'b0;
    XRAM[25616] = 8'b0;
    XRAM[25617] = 8'b0;
    XRAM[25618] = 8'b0;
    XRAM[25619] = 8'b0;
    XRAM[25620] = 8'b0;
    XRAM[25621] = 8'b0;
    XRAM[25622] = 8'b0;
    XRAM[25623] = 8'b0;
    XRAM[25624] = 8'b0;
    XRAM[25625] = 8'b0;
    XRAM[25626] = 8'b0;
    XRAM[25627] = 8'b0;
    XRAM[25628] = 8'b0;
    XRAM[25629] = 8'b0;
    XRAM[25630] = 8'b0;
    XRAM[25631] = 8'b0;
    XRAM[25632] = 8'b0;
    XRAM[25633] = 8'b0;
    XRAM[25634] = 8'b0;
    XRAM[25635] = 8'b0;
    XRAM[25636] = 8'b0;
    XRAM[25637] = 8'b0;
    XRAM[25638] = 8'b0;
    XRAM[25639] = 8'b0;
    XRAM[25640] = 8'b0;
    XRAM[25641] = 8'b0;
    XRAM[25642] = 8'b0;
    XRAM[25643] = 8'b0;
    XRAM[25644] = 8'b0;
    XRAM[25645] = 8'b0;
    XRAM[25646] = 8'b0;
    XRAM[25647] = 8'b0;
    XRAM[25648] = 8'b0;
    XRAM[25649] = 8'b0;
    XRAM[25650] = 8'b0;
    XRAM[25651] = 8'b0;
    XRAM[25652] = 8'b0;
    XRAM[25653] = 8'b0;
    XRAM[25654] = 8'b0;
    XRAM[25655] = 8'b0;
    XRAM[25656] = 8'b0;
    XRAM[25657] = 8'b0;
    XRAM[25658] = 8'b0;
    XRAM[25659] = 8'b0;
    XRAM[25660] = 8'b0;
    XRAM[25661] = 8'b0;
    XRAM[25662] = 8'b0;
    XRAM[25663] = 8'b0;
    XRAM[25664] = 8'b0;
    XRAM[25665] = 8'b0;
    XRAM[25666] = 8'b0;
    XRAM[25667] = 8'b0;
    XRAM[25668] = 8'b0;
    XRAM[25669] = 8'b0;
    XRAM[25670] = 8'b0;
    XRAM[25671] = 8'b0;
    XRAM[25672] = 8'b0;
    XRAM[25673] = 8'b0;
    XRAM[25674] = 8'b0;
    XRAM[25675] = 8'b0;
    XRAM[25676] = 8'b0;
    XRAM[25677] = 8'b0;
    XRAM[25678] = 8'b0;
    XRAM[25679] = 8'b0;
    XRAM[25680] = 8'b0;
    XRAM[25681] = 8'b0;
    XRAM[25682] = 8'b0;
    XRAM[25683] = 8'b0;
    XRAM[25684] = 8'b0;
    XRAM[25685] = 8'b0;
    XRAM[25686] = 8'b0;
    XRAM[25687] = 8'b0;
    XRAM[25688] = 8'b0;
    XRAM[25689] = 8'b0;
    XRAM[25690] = 8'b0;
    XRAM[25691] = 8'b0;
    XRAM[25692] = 8'b0;
    XRAM[25693] = 8'b0;
    XRAM[25694] = 8'b0;
    XRAM[25695] = 8'b0;
    XRAM[25696] = 8'b0;
    XRAM[25697] = 8'b0;
    XRAM[25698] = 8'b0;
    XRAM[25699] = 8'b0;
    XRAM[25700] = 8'b0;
    XRAM[25701] = 8'b0;
    XRAM[25702] = 8'b0;
    XRAM[25703] = 8'b0;
    XRAM[25704] = 8'b0;
    XRAM[25705] = 8'b0;
    XRAM[25706] = 8'b0;
    XRAM[25707] = 8'b0;
    XRAM[25708] = 8'b0;
    XRAM[25709] = 8'b0;
    XRAM[25710] = 8'b0;
    XRAM[25711] = 8'b0;
    XRAM[25712] = 8'b0;
    XRAM[25713] = 8'b0;
    XRAM[25714] = 8'b0;
    XRAM[25715] = 8'b0;
    XRAM[25716] = 8'b0;
    XRAM[25717] = 8'b0;
    XRAM[25718] = 8'b0;
    XRAM[25719] = 8'b0;
    XRAM[25720] = 8'b0;
    XRAM[25721] = 8'b0;
    XRAM[25722] = 8'b0;
    XRAM[25723] = 8'b0;
    XRAM[25724] = 8'b0;
    XRAM[25725] = 8'b0;
    XRAM[25726] = 8'b0;
    XRAM[25727] = 8'b0;
    XRAM[25728] = 8'b0;
    XRAM[25729] = 8'b0;
    XRAM[25730] = 8'b0;
    XRAM[25731] = 8'b0;
    XRAM[25732] = 8'b0;
    XRAM[25733] = 8'b0;
    XRAM[25734] = 8'b0;
    XRAM[25735] = 8'b0;
    XRAM[25736] = 8'b0;
    XRAM[25737] = 8'b0;
    XRAM[25738] = 8'b0;
    XRAM[25739] = 8'b0;
    XRAM[25740] = 8'b0;
    XRAM[25741] = 8'b0;
    XRAM[25742] = 8'b0;
    XRAM[25743] = 8'b0;
    XRAM[25744] = 8'b0;
    XRAM[25745] = 8'b0;
    XRAM[25746] = 8'b0;
    XRAM[25747] = 8'b0;
    XRAM[25748] = 8'b0;
    XRAM[25749] = 8'b0;
    XRAM[25750] = 8'b0;
    XRAM[25751] = 8'b0;
    XRAM[25752] = 8'b0;
    XRAM[25753] = 8'b0;
    XRAM[25754] = 8'b0;
    XRAM[25755] = 8'b0;
    XRAM[25756] = 8'b0;
    XRAM[25757] = 8'b0;
    XRAM[25758] = 8'b0;
    XRAM[25759] = 8'b0;
    XRAM[25760] = 8'b0;
    XRAM[25761] = 8'b0;
    XRAM[25762] = 8'b0;
    XRAM[25763] = 8'b0;
    XRAM[25764] = 8'b0;
    XRAM[25765] = 8'b0;
    XRAM[25766] = 8'b0;
    XRAM[25767] = 8'b0;
    XRAM[25768] = 8'b0;
    XRAM[25769] = 8'b0;
    XRAM[25770] = 8'b0;
    XRAM[25771] = 8'b0;
    XRAM[25772] = 8'b0;
    XRAM[25773] = 8'b0;
    XRAM[25774] = 8'b0;
    XRAM[25775] = 8'b0;
    XRAM[25776] = 8'b0;
    XRAM[25777] = 8'b0;
    XRAM[25778] = 8'b0;
    XRAM[25779] = 8'b0;
    XRAM[25780] = 8'b0;
    XRAM[25781] = 8'b0;
    XRAM[25782] = 8'b0;
    XRAM[25783] = 8'b0;
    XRAM[25784] = 8'b0;
    XRAM[25785] = 8'b0;
    XRAM[25786] = 8'b0;
    XRAM[25787] = 8'b0;
    XRAM[25788] = 8'b0;
    XRAM[25789] = 8'b0;
    XRAM[25790] = 8'b0;
    XRAM[25791] = 8'b0;
    XRAM[25792] = 8'b0;
    XRAM[25793] = 8'b0;
    XRAM[25794] = 8'b0;
    XRAM[25795] = 8'b0;
    XRAM[25796] = 8'b0;
    XRAM[25797] = 8'b0;
    XRAM[25798] = 8'b0;
    XRAM[25799] = 8'b0;
    XRAM[25800] = 8'b0;
    XRAM[25801] = 8'b0;
    XRAM[25802] = 8'b0;
    XRAM[25803] = 8'b0;
    XRAM[25804] = 8'b0;
    XRAM[25805] = 8'b0;
    XRAM[25806] = 8'b0;
    XRAM[25807] = 8'b0;
    XRAM[25808] = 8'b0;
    XRAM[25809] = 8'b0;
    XRAM[25810] = 8'b0;
    XRAM[25811] = 8'b0;
    XRAM[25812] = 8'b0;
    XRAM[25813] = 8'b0;
    XRAM[25814] = 8'b0;
    XRAM[25815] = 8'b0;
    XRAM[25816] = 8'b0;
    XRAM[25817] = 8'b0;
    XRAM[25818] = 8'b0;
    XRAM[25819] = 8'b0;
    XRAM[25820] = 8'b0;
    XRAM[25821] = 8'b0;
    XRAM[25822] = 8'b0;
    XRAM[25823] = 8'b0;
    XRAM[25824] = 8'b0;
    XRAM[25825] = 8'b0;
    XRAM[25826] = 8'b0;
    XRAM[25827] = 8'b0;
    XRAM[25828] = 8'b0;
    XRAM[25829] = 8'b0;
    XRAM[25830] = 8'b0;
    XRAM[25831] = 8'b0;
    XRAM[25832] = 8'b0;
    XRAM[25833] = 8'b0;
    XRAM[25834] = 8'b0;
    XRAM[25835] = 8'b0;
    XRAM[25836] = 8'b0;
    XRAM[25837] = 8'b0;
    XRAM[25838] = 8'b0;
    XRAM[25839] = 8'b0;
    XRAM[25840] = 8'b0;
    XRAM[25841] = 8'b0;
    XRAM[25842] = 8'b0;
    XRAM[25843] = 8'b0;
    XRAM[25844] = 8'b0;
    XRAM[25845] = 8'b0;
    XRAM[25846] = 8'b0;
    XRAM[25847] = 8'b0;
    XRAM[25848] = 8'b0;
    XRAM[25849] = 8'b0;
    XRAM[25850] = 8'b0;
    XRAM[25851] = 8'b0;
    XRAM[25852] = 8'b0;
    XRAM[25853] = 8'b0;
    XRAM[25854] = 8'b0;
    XRAM[25855] = 8'b0;
    XRAM[25856] = 8'b0;
    XRAM[25857] = 8'b0;
    XRAM[25858] = 8'b0;
    XRAM[25859] = 8'b0;
    XRAM[25860] = 8'b0;
    XRAM[25861] = 8'b0;
    XRAM[25862] = 8'b0;
    XRAM[25863] = 8'b0;
    XRAM[25864] = 8'b0;
    XRAM[25865] = 8'b0;
    XRAM[25866] = 8'b0;
    XRAM[25867] = 8'b0;
    XRAM[25868] = 8'b0;
    XRAM[25869] = 8'b0;
    XRAM[25870] = 8'b0;
    XRAM[25871] = 8'b0;
    XRAM[25872] = 8'b0;
    XRAM[25873] = 8'b0;
    XRAM[25874] = 8'b0;
    XRAM[25875] = 8'b0;
    XRAM[25876] = 8'b0;
    XRAM[25877] = 8'b0;
    XRAM[25878] = 8'b0;
    XRAM[25879] = 8'b0;
    XRAM[25880] = 8'b0;
    XRAM[25881] = 8'b0;
    XRAM[25882] = 8'b0;
    XRAM[25883] = 8'b0;
    XRAM[25884] = 8'b0;
    XRAM[25885] = 8'b0;
    XRAM[25886] = 8'b0;
    XRAM[25887] = 8'b0;
    XRAM[25888] = 8'b0;
    XRAM[25889] = 8'b0;
    XRAM[25890] = 8'b0;
    XRAM[25891] = 8'b0;
    XRAM[25892] = 8'b0;
    XRAM[25893] = 8'b0;
    XRAM[25894] = 8'b0;
    XRAM[25895] = 8'b0;
    XRAM[25896] = 8'b0;
    XRAM[25897] = 8'b0;
    XRAM[25898] = 8'b0;
    XRAM[25899] = 8'b0;
    XRAM[25900] = 8'b0;
    XRAM[25901] = 8'b0;
    XRAM[25902] = 8'b0;
    XRAM[25903] = 8'b0;
    XRAM[25904] = 8'b0;
    XRAM[25905] = 8'b0;
    XRAM[25906] = 8'b0;
    XRAM[25907] = 8'b0;
    XRAM[25908] = 8'b0;
    XRAM[25909] = 8'b0;
    XRAM[25910] = 8'b0;
    XRAM[25911] = 8'b0;
    XRAM[25912] = 8'b0;
    XRAM[25913] = 8'b0;
    XRAM[25914] = 8'b0;
    XRAM[25915] = 8'b0;
    XRAM[25916] = 8'b0;
    XRAM[25917] = 8'b0;
    XRAM[25918] = 8'b0;
    XRAM[25919] = 8'b0;
    XRAM[25920] = 8'b0;
    XRAM[25921] = 8'b0;
    XRAM[25922] = 8'b0;
    XRAM[25923] = 8'b0;
    XRAM[25924] = 8'b0;
    XRAM[25925] = 8'b0;
    XRAM[25926] = 8'b0;
    XRAM[25927] = 8'b0;
    XRAM[25928] = 8'b0;
    XRAM[25929] = 8'b0;
    XRAM[25930] = 8'b0;
    XRAM[25931] = 8'b0;
    XRAM[25932] = 8'b0;
    XRAM[25933] = 8'b0;
    XRAM[25934] = 8'b0;
    XRAM[25935] = 8'b0;
    XRAM[25936] = 8'b0;
    XRAM[25937] = 8'b0;
    XRAM[25938] = 8'b0;
    XRAM[25939] = 8'b0;
    XRAM[25940] = 8'b0;
    XRAM[25941] = 8'b0;
    XRAM[25942] = 8'b0;
    XRAM[25943] = 8'b0;
    XRAM[25944] = 8'b0;
    XRAM[25945] = 8'b0;
    XRAM[25946] = 8'b0;
    XRAM[25947] = 8'b0;
    XRAM[25948] = 8'b0;
    XRAM[25949] = 8'b0;
    XRAM[25950] = 8'b0;
    XRAM[25951] = 8'b0;
    XRAM[25952] = 8'b0;
    XRAM[25953] = 8'b0;
    XRAM[25954] = 8'b0;
    XRAM[25955] = 8'b0;
    XRAM[25956] = 8'b0;
    XRAM[25957] = 8'b0;
    XRAM[25958] = 8'b0;
    XRAM[25959] = 8'b0;
    XRAM[25960] = 8'b0;
    XRAM[25961] = 8'b0;
    XRAM[25962] = 8'b0;
    XRAM[25963] = 8'b0;
    XRAM[25964] = 8'b0;
    XRAM[25965] = 8'b0;
    XRAM[25966] = 8'b0;
    XRAM[25967] = 8'b0;
    XRAM[25968] = 8'b0;
    XRAM[25969] = 8'b0;
    XRAM[25970] = 8'b0;
    XRAM[25971] = 8'b0;
    XRAM[25972] = 8'b0;
    XRAM[25973] = 8'b0;
    XRAM[25974] = 8'b0;
    XRAM[25975] = 8'b0;
    XRAM[25976] = 8'b0;
    XRAM[25977] = 8'b0;
    XRAM[25978] = 8'b0;
    XRAM[25979] = 8'b0;
    XRAM[25980] = 8'b0;
    XRAM[25981] = 8'b0;
    XRAM[25982] = 8'b0;
    XRAM[25983] = 8'b0;
    XRAM[25984] = 8'b0;
    XRAM[25985] = 8'b0;
    XRAM[25986] = 8'b0;
    XRAM[25987] = 8'b0;
    XRAM[25988] = 8'b0;
    XRAM[25989] = 8'b0;
    XRAM[25990] = 8'b0;
    XRAM[25991] = 8'b0;
    XRAM[25992] = 8'b0;
    XRAM[25993] = 8'b0;
    XRAM[25994] = 8'b0;
    XRAM[25995] = 8'b0;
    XRAM[25996] = 8'b0;
    XRAM[25997] = 8'b0;
    XRAM[25998] = 8'b0;
    XRAM[25999] = 8'b0;
    XRAM[26000] = 8'b0;
    XRAM[26001] = 8'b0;
    XRAM[26002] = 8'b0;
    XRAM[26003] = 8'b0;
    XRAM[26004] = 8'b0;
    XRAM[26005] = 8'b0;
    XRAM[26006] = 8'b0;
    XRAM[26007] = 8'b0;
    XRAM[26008] = 8'b0;
    XRAM[26009] = 8'b0;
    XRAM[26010] = 8'b0;
    XRAM[26011] = 8'b0;
    XRAM[26012] = 8'b0;
    XRAM[26013] = 8'b0;
    XRAM[26014] = 8'b0;
    XRAM[26015] = 8'b0;
    XRAM[26016] = 8'b0;
    XRAM[26017] = 8'b0;
    XRAM[26018] = 8'b0;
    XRAM[26019] = 8'b0;
    XRAM[26020] = 8'b0;
    XRAM[26021] = 8'b0;
    XRAM[26022] = 8'b0;
    XRAM[26023] = 8'b0;
    XRAM[26024] = 8'b0;
    XRAM[26025] = 8'b0;
    XRAM[26026] = 8'b0;
    XRAM[26027] = 8'b0;
    XRAM[26028] = 8'b0;
    XRAM[26029] = 8'b0;
    XRAM[26030] = 8'b0;
    XRAM[26031] = 8'b0;
    XRAM[26032] = 8'b0;
    XRAM[26033] = 8'b0;
    XRAM[26034] = 8'b0;
    XRAM[26035] = 8'b0;
    XRAM[26036] = 8'b0;
    XRAM[26037] = 8'b0;
    XRAM[26038] = 8'b0;
    XRAM[26039] = 8'b0;
    XRAM[26040] = 8'b0;
    XRAM[26041] = 8'b0;
    XRAM[26042] = 8'b0;
    XRAM[26043] = 8'b0;
    XRAM[26044] = 8'b0;
    XRAM[26045] = 8'b0;
    XRAM[26046] = 8'b0;
    XRAM[26047] = 8'b0;
    XRAM[26048] = 8'b0;
    XRAM[26049] = 8'b0;
    XRAM[26050] = 8'b0;
    XRAM[26051] = 8'b0;
    XRAM[26052] = 8'b0;
    XRAM[26053] = 8'b0;
    XRAM[26054] = 8'b0;
    XRAM[26055] = 8'b0;
    XRAM[26056] = 8'b0;
    XRAM[26057] = 8'b0;
    XRAM[26058] = 8'b0;
    XRAM[26059] = 8'b0;
    XRAM[26060] = 8'b0;
    XRAM[26061] = 8'b0;
    XRAM[26062] = 8'b0;
    XRAM[26063] = 8'b0;
    XRAM[26064] = 8'b0;
    XRAM[26065] = 8'b0;
    XRAM[26066] = 8'b0;
    XRAM[26067] = 8'b0;
    XRAM[26068] = 8'b0;
    XRAM[26069] = 8'b0;
    XRAM[26070] = 8'b0;
    XRAM[26071] = 8'b0;
    XRAM[26072] = 8'b0;
    XRAM[26073] = 8'b0;
    XRAM[26074] = 8'b0;
    XRAM[26075] = 8'b0;
    XRAM[26076] = 8'b0;
    XRAM[26077] = 8'b0;
    XRAM[26078] = 8'b0;
    XRAM[26079] = 8'b0;
    XRAM[26080] = 8'b0;
    XRAM[26081] = 8'b0;
    XRAM[26082] = 8'b0;
    XRAM[26083] = 8'b0;
    XRAM[26084] = 8'b0;
    XRAM[26085] = 8'b0;
    XRAM[26086] = 8'b0;
    XRAM[26087] = 8'b0;
    XRAM[26088] = 8'b0;
    XRAM[26089] = 8'b0;
    XRAM[26090] = 8'b0;
    XRAM[26091] = 8'b0;
    XRAM[26092] = 8'b0;
    XRAM[26093] = 8'b0;
    XRAM[26094] = 8'b0;
    XRAM[26095] = 8'b0;
    XRAM[26096] = 8'b0;
    XRAM[26097] = 8'b0;
    XRAM[26098] = 8'b0;
    XRAM[26099] = 8'b0;
    XRAM[26100] = 8'b0;
    XRAM[26101] = 8'b0;
    XRAM[26102] = 8'b0;
    XRAM[26103] = 8'b0;
    XRAM[26104] = 8'b0;
    XRAM[26105] = 8'b0;
    XRAM[26106] = 8'b0;
    XRAM[26107] = 8'b0;
    XRAM[26108] = 8'b0;
    XRAM[26109] = 8'b0;
    XRAM[26110] = 8'b0;
    XRAM[26111] = 8'b0;
    XRAM[26112] = 8'b0;
    XRAM[26113] = 8'b0;
    XRAM[26114] = 8'b0;
    XRAM[26115] = 8'b0;
    XRAM[26116] = 8'b0;
    XRAM[26117] = 8'b0;
    XRAM[26118] = 8'b0;
    XRAM[26119] = 8'b0;
    XRAM[26120] = 8'b0;
    XRAM[26121] = 8'b0;
    XRAM[26122] = 8'b0;
    XRAM[26123] = 8'b0;
    XRAM[26124] = 8'b0;
    XRAM[26125] = 8'b0;
    XRAM[26126] = 8'b0;
    XRAM[26127] = 8'b0;
    XRAM[26128] = 8'b0;
    XRAM[26129] = 8'b0;
    XRAM[26130] = 8'b0;
    XRAM[26131] = 8'b0;
    XRAM[26132] = 8'b0;
    XRAM[26133] = 8'b0;
    XRAM[26134] = 8'b0;
    XRAM[26135] = 8'b0;
    XRAM[26136] = 8'b0;
    XRAM[26137] = 8'b0;
    XRAM[26138] = 8'b0;
    XRAM[26139] = 8'b0;
    XRAM[26140] = 8'b0;
    XRAM[26141] = 8'b0;
    XRAM[26142] = 8'b0;
    XRAM[26143] = 8'b0;
    XRAM[26144] = 8'b0;
    XRAM[26145] = 8'b0;
    XRAM[26146] = 8'b0;
    XRAM[26147] = 8'b0;
    XRAM[26148] = 8'b0;
    XRAM[26149] = 8'b0;
    XRAM[26150] = 8'b0;
    XRAM[26151] = 8'b0;
    XRAM[26152] = 8'b0;
    XRAM[26153] = 8'b0;
    XRAM[26154] = 8'b0;
    XRAM[26155] = 8'b0;
    XRAM[26156] = 8'b0;
    XRAM[26157] = 8'b0;
    XRAM[26158] = 8'b0;
    XRAM[26159] = 8'b0;
    XRAM[26160] = 8'b0;
    XRAM[26161] = 8'b0;
    XRAM[26162] = 8'b0;
    XRAM[26163] = 8'b0;
    XRAM[26164] = 8'b0;
    XRAM[26165] = 8'b0;
    XRAM[26166] = 8'b0;
    XRAM[26167] = 8'b0;
    XRAM[26168] = 8'b0;
    XRAM[26169] = 8'b0;
    XRAM[26170] = 8'b0;
    XRAM[26171] = 8'b0;
    XRAM[26172] = 8'b0;
    XRAM[26173] = 8'b0;
    XRAM[26174] = 8'b0;
    XRAM[26175] = 8'b0;
    XRAM[26176] = 8'b0;
    XRAM[26177] = 8'b0;
    XRAM[26178] = 8'b0;
    XRAM[26179] = 8'b0;
    XRAM[26180] = 8'b0;
    XRAM[26181] = 8'b0;
    XRAM[26182] = 8'b0;
    XRAM[26183] = 8'b0;
    XRAM[26184] = 8'b0;
    XRAM[26185] = 8'b0;
    XRAM[26186] = 8'b0;
    XRAM[26187] = 8'b0;
    XRAM[26188] = 8'b0;
    XRAM[26189] = 8'b0;
    XRAM[26190] = 8'b0;
    XRAM[26191] = 8'b0;
    XRAM[26192] = 8'b0;
    XRAM[26193] = 8'b0;
    XRAM[26194] = 8'b0;
    XRAM[26195] = 8'b0;
    XRAM[26196] = 8'b0;
    XRAM[26197] = 8'b0;
    XRAM[26198] = 8'b0;
    XRAM[26199] = 8'b0;
    XRAM[26200] = 8'b0;
    XRAM[26201] = 8'b0;
    XRAM[26202] = 8'b0;
    XRAM[26203] = 8'b0;
    XRAM[26204] = 8'b0;
    XRAM[26205] = 8'b0;
    XRAM[26206] = 8'b0;
    XRAM[26207] = 8'b0;
    XRAM[26208] = 8'b0;
    XRAM[26209] = 8'b0;
    XRAM[26210] = 8'b0;
    XRAM[26211] = 8'b0;
    XRAM[26212] = 8'b0;
    XRAM[26213] = 8'b0;
    XRAM[26214] = 8'b0;
    XRAM[26215] = 8'b0;
    XRAM[26216] = 8'b0;
    XRAM[26217] = 8'b0;
    XRAM[26218] = 8'b0;
    XRAM[26219] = 8'b0;
    XRAM[26220] = 8'b0;
    XRAM[26221] = 8'b0;
    XRAM[26222] = 8'b0;
    XRAM[26223] = 8'b0;
    XRAM[26224] = 8'b0;
    XRAM[26225] = 8'b0;
    XRAM[26226] = 8'b0;
    XRAM[26227] = 8'b0;
    XRAM[26228] = 8'b0;
    XRAM[26229] = 8'b0;
    XRAM[26230] = 8'b0;
    XRAM[26231] = 8'b0;
    XRAM[26232] = 8'b0;
    XRAM[26233] = 8'b0;
    XRAM[26234] = 8'b0;
    XRAM[26235] = 8'b0;
    XRAM[26236] = 8'b0;
    XRAM[26237] = 8'b0;
    XRAM[26238] = 8'b0;
    XRAM[26239] = 8'b0;
    XRAM[26240] = 8'b0;
    XRAM[26241] = 8'b0;
    XRAM[26242] = 8'b0;
    XRAM[26243] = 8'b0;
    XRAM[26244] = 8'b0;
    XRAM[26245] = 8'b0;
    XRAM[26246] = 8'b0;
    XRAM[26247] = 8'b0;
    XRAM[26248] = 8'b0;
    XRAM[26249] = 8'b0;
    XRAM[26250] = 8'b0;
    XRAM[26251] = 8'b0;
    XRAM[26252] = 8'b0;
    XRAM[26253] = 8'b0;
    XRAM[26254] = 8'b0;
    XRAM[26255] = 8'b0;
    XRAM[26256] = 8'b0;
    XRAM[26257] = 8'b0;
    XRAM[26258] = 8'b0;
    XRAM[26259] = 8'b0;
    XRAM[26260] = 8'b0;
    XRAM[26261] = 8'b0;
    XRAM[26262] = 8'b0;
    XRAM[26263] = 8'b0;
    XRAM[26264] = 8'b0;
    XRAM[26265] = 8'b0;
    XRAM[26266] = 8'b0;
    XRAM[26267] = 8'b0;
    XRAM[26268] = 8'b0;
    XRAM[26269] = 8'b0;
    XRAM[26270] = 8'b0;
    XRAM[26271] = 8'b0;
    XRAM[26272] = 8'b0;
    XRAM[26273] = 8'b0;
    XRAM[26274] = 8'b0;
    XRAM[26275] = 8'b0;
    XRAM[26276] = 8'b0;
    XRAM[26277] = 8'b0;
    XRAM[26278] = 8'b0;
    XRAM[26279] = 8'b0;
    XRAM[26280] = 8'b0;
    XRAM[26281] = 8'b0;
    XRAM[26282] = 8'b0;
    XRAM[26283] = 8'b0;
    XRAM[26284] = 8'b0;
    XRAM[26285] = 8'b0;
    XRAM[26286] = 8'b0;
    XRAM[26287] = 8'b0;
    XRAM[26288] = 8'b0;
    XRAM[26289] = 8'b0;
    XRAM[26290] = 8'b0;
    XRAM[26291] = 8'b0;
    XRAM[26292] = 8'b0;
    XRAM[26293] = 8'b0;
    XRAM[26294] = 8'b0;
    XRAM[26295] = 8'b0;
    XRAM[26296] = 8'b0;
    XRAM[26297] = 8'b0;
    XRAM[26298] = 8'b0;
    XRAM[26299] = 8'b0;
    XRAM[26300] = 8'b0;
    XRAM[26301] = 8'b0;
    XRAM[26302] = 8'b0;
    XRAM[26303] = 8'b0;
    XRAM[26304] = 8'b0;
    XRAM[26305] = 8'b0;
    XRAM[26306] = 8'b0;
    XRAM[26307] = 8'b0;
    XRAM[26308] = 8'b0;
    XRAM[26309] = 8'b0;
    XRAM[26310] = 8'b0;
    XRAM[26311] = 8'b0;
    XRAM[26312] = 8'b0;
    XRAM[26313] = 8'b0;
    XRAM[26314] = 8'b0;
    XRAM[26315] = 8'b0;
    XRAM[26316] = 8'b0;
    XRAM[26317] = 8'b0;
    XRAM[26318] = 8'b0;
    XRAM[26319] = 8'b0;
    XRAM[26320] = 8'b0;
    XRAM[26321] = 8'b0;
    XRAM[26322] = 8'b0;
    XRAM[26323] = 8'b0;
    XRAM[26324] = 8'b0;
    XRAM[26325] = 8'b0;
    XRAM[26326] = 8'b0;
    XRAM[26327] = 8'b0;
    XRAM[26328] = 8'b0;
    XRAM[26329] = 8'b0;
    XRAM[26330] = 8'b0;
    XRAM[26331] = 8'b0;
    XRAM[26332] = 8'b0;
    XRAM[26333] = 8'b0;
    XRAM[26334] = 8'b0;
    XRAM[26335] = 8'b0;
    XRAM[26336] = 8'b0;
    XRAM[26337] = 8'b0;
    XRAM[26338] = 8'b0;
    XRAM[26339] = 8'b0;
    XRAM[26340] = 8'b0;
    XRAM[26341] = 8'b0;
    XRAM[26342] = 8'b0;
    XRAM[26343] = 8'b0;
    XRAM[26344] = 8'b0;
    XRAM[26345] = 8'b0;
    XRAM[26346] = 8'b0;
    XRAM[26347] = 8'b0;
    XRAM[26348] = 8'b0;
    XRAM[26349] = 8'b0;
    XRAM[26350] = 8'b0;
    XRAM[26351] = 8'b0;
    XRAM[26352] = 8'b0;
    XRAM[26353] = 8'b0;
    XRAM[26354] = 8'b0;
    XRAM[26355] = 8'b0;
    XRAM[26356] = 8'b0;
    XRAM[26357] = 8'b0;
    XRAM[26358] = 8'b0;
    XRAM[26359] = 8'b0;
    XRAM[26360] = 8'b0;
    XRAM[26361] = 8'b0;
    XRAM[26362] = 8'b0;
    XRAM[26363] = 8'b0;
    XRAM[26364] = 8'b0;
    XRAM[26365] = 8'b0;
    XRAM[26366] = 8'b0;
    XRAM[26367] = 8'b0;
    XRAM[26368] = 8'b0;
    XRAM[26369] = 8'b0;
    XRAM[26370] = 8'b0;
    XRAM[26371] = 8'b0;
    XRAM[26372] = 8'b0;
    XRAM[26373] = 8'b0;
    XRAM[26374] = 8'b0;
    XRAM[26375] = 8'b0;
    XRAM[26376] = 8'b0;
    XRAM[26377] = 8'b0;
    XRAM[26378] = 8'b0;
    XRAM[26379] = 8'b0;
    XRAM[26380] = 8'b0;
    XRAM[26381] = 8'b0;
    XRAM[26382] = 8'b0;
    XRAM[26383] = 8'b0;
    XRAM[26384] = 8'b0;
    XRAM[26385] = 8'b0;
    XRAM[26386] = 8'b0;
    XRAM[26387] = 8'b0;
    XRAM[26388] = 8'b0;
    XRAM[26389] = 8'b0;
    XRAM[26390] = 8'b0;
    XRAM[26391] = 8'b0;
    XRAM[26392] = 8'b0;
    XRAM[26393] = 8'b0;
    XRAM[26394] = 8'b0;
    XRAM[26395] = 8'b0;
    XRAM[26396] = 8'b0;
    XRAM[26397] = 8'b0;
    XRAM[26398] = 8'b0;
    XRAM[26399] = 8'b0;
    XRAM[26400] = 8'b0;
    XRAM[26401] = 8'b0;
    XRAM[26402] = 8'b0;
    XRAM[26403] = 8'b0;
    XRAM[26404] = 8'b0;
    XRAM[26405] = 8'b0;
    XRAM[26406] = 8'b0;
    XRAM[26407] = 8'b0;
    XRAM[26408] = 8'b0;
    XRAM[26409] = 8'b0;
    XRAM[26410] = 8'b0;
    XRAM[26411] = 8'b0;
    XRAM[26412] = 8'b0;
    XRAM[26413] = 8'b0;
    XRAM[26414] = 8'b0;
    XRAM[26415] = 8'b0;
    XRAM[26416] = 8'b0;
    XRAM[26417] = 8'b0;
    XRAM[26418] = 8'b0;
    XRAM[26419] = 8'b0;
    XRAM[26420] = 8'b0;
    XRAM[26421] = 8'b0;
    XRAM[26422] = 8'b0;
    XRAM[26423] = 8'b0;
    XRAM[26424] = 8'b0;
    XRAM[26425] = 8'b0;
    XRAM[26426] = 8'b0;
    XRAM[26427] = 8'b0;
    XRAM[26428] = 8'b0;
    XRAM[26429] = 8'b0;
    XRAM[26430] = 8'b0;
    XRAM[26431] = 8'b0;
    XRAM[26432] = 8'b0;
    XRAM[26433] = 8'b0;
    XRAM[26434] = 8'b0;
    XRAM[26435] = 8'b0;
    XRAM[26436] = 8'b0;
    XRAM[26437] = 8'b0;
    XRAM[26438] = 8'b0;
    XRAM[26439] = 8'b0;
    XRAM[26440] = 8'b0;
    XRAM[26441] = 8'b0;
    XRAM[26442] = 8'b0;
    XRAM[26443] = 8'b0;
    XRAM[26444] = 8'b0;
    XRAM[26445] = 8'b0;
    XRAM[26446] = 8'b0;
    XRAM[26447] = 8'b0;
    XRAM[26448] = 8'b0;
    XRAM[26449] = 8'b0;
    XRAM[26450] = 8'b0;
    XRAM[26451] = 8'b0;
    XRAM[26452] = 8'b0;
    XRAM[26453] = 8'b0;
    XRAM[26454] = 8'b0;
    XRAM[26455] = 8'b0;
    XRAM[26456] = 8'b0;
    XRAM[26457] = 8'b0;
    XRAM[26458] = 8'b0;
    XRAM[26459] = 8'b0;
    XRAM[26460] = 8'b0;
    XRAM[26461] = 8'b0;
    XRAM[26462] = 8'b0;
    XRAM[26463] = 8'b0;
    XRAM[26464] = 8'b0;
    XRAM[26465] = 8'b0;
    XRAM[26466] = 8'b0;
    XRAM[26467] = 8'b0;
    XRAM[26468] = 8'b0;
    XRAM[26469] = 8'b0;
    XRAM[26470] = 8'b0;
    XRAM[26471] = 8'b0;
    XRAM[26472] = 8'b0;
    XRAM[26473] = 8'b0;
    XRAM[26474] = 8'b0;
    XRAM[26475] = 8'b0;
    XRAM[26476] = 8'b0;
    XRAM[26477] = 8'b0;
    XRAM[26478] = 8'b0;
    XRAM[26479] = 8'b0;
    XRAM[26480] = 8'b0;
    XRAM[26481] = 8'b0;
    XRAM[26482] = 8'b0;
    XRAM[26483] = 8'b0;
    XRAM[26484] = 8'b0;
    XRAM[26485] = 8'b0;
    XRAM[26486] = 8'b0;
    XRAM[26487] = 8'b0;
    XRAM[26488] = 8'b0;
    XRAM[26489] = 8'b0;
    XRAM[26490] = 8'b0;
    XRAM[26491] = 8'b0;
    XRAM[26492] = 8'b0;
    XRAM[26493] = 8'b0;
    XRAM[26494] = 8'b0;
    XRAM[26495] = 8'b0;
    XRAM[26496] = 8'b0;
    XRAM[26497] = 8'b0;
    XRAM[26498] = 8'b0;
    XRAM[26499] = 8'b0;
    XRAM[26500] = 8'b0;
    XRAM[26501] = 8'b0;
    XRAM[26502] = 8'b0;
    XRAM[26503] = 8'b0;
    XRAM[26504] = 8'b0;
    XRAM[26505] = 8'b0;
    XRAM[26506] = 8'b0;
    XRAM[26507] = 8'b0;
    XRAM[26508] = 8'b0;
    XRAM[26509] = 8'b0;
    XRAM[26510] = 8'b0;
    XRAM[26511] = 8'b0;
    XRAM[26512] = 8'b0;
    XRAM[26513] = 8'b0;
    XRAM[26514] = 8'b0;
    XRAM[26515] = 8'b0;
    XRAM[26516] = 8'b0;
    XRAM[26517] = 8'b0;
    XRAM[26518] = 8'b0;
    XRAM[26519] = 8'b0;
    XRAM[26520] = 8'b0;
    XRAM[26521] = 8'b0;
    XRAM[26522] = 8'b0;
    XRAM[26523] = 8'b0;
    XRAM[26524] = 8'b0;
    XRAM[26525] = 8'b0;
    XRAM[26526] = 8'b0;
    XRAM[26527] = 8'b0;
    XRAM[26528] = 8'b0;
    XRAM[26529] = 8'b0;
    XRAM[26530] = 8'b0;
    XRAM[26531] = 8'b0;
    XRAM[26532] = 8'b0;
    XRAM[26533] = 8'b0;
    XRAM[26534] = 8'b0;
    XRAM[26535] = 8'b0;
    XRAM[26536] = 8'b0;
    XRAM[26537] = 8'b0;
    XRAM[26538] = 8'b0;
    XRAM[26539] = 8'b0;
    XRAM[26540] = 8'b0;
    XRAM[26541] = 8'b0;
    XRAM[26542] = 8'b0;
    XRAM[26543] = 8'b0;
    XRAM[26544] = 8'b0;
    XRAM[26545] = 8'b0;
    XRAM[26546] = 8'b0;
    XRAM[26547] = 8'b0;
    XRAM[26548] = 8'b0;
    XRAM[26549] = 8'b0;
    XRAM[26550] = 8'b0;
    XRAM[26551] = 8'b0;
    XRAM[26552] = 8'b0;
    XRAM[26553] = 8'b0;
    XRAM[26554] = 8'b0;
    XRAM[26555] = 8'b0;
    XRAM[26556] = 8'b0;
    XRAM[26557] = 8'b0;
    XRAM[26558] = 8'b0;
    XRAM[26559] = 8'b0;
    XRAM[26560] = 8'b0;
    XRAM[26561] = 8'b0;
    XRAM[26562] = 8'b0;
    XRAM[26563] = 8'b0;
    XRAM[26564] = 8'b0;
    XRAM[26565] = 8'b0;
    XRAM[26566] = 8'b0;
    XRAM[26567] = 8'b0;
    XRAM[26568] = 8'b0;
    XRAM[26569] = 8'b0;
    XRAM[26570] = 8'b0;
    XRAM[26571] = 8'b0;
    XRAM[26572] = 8'b0;
    XRAM[26573] = 8'b0;
    XRAM[26574] = 8'b0;
    XRAM[26575] = 8'b0;
    XRAM[26576] = 8'b0;
    XRAM[26577] = 8'b0;
    XRAM[26578] = 8'b0;
    XRAM[26579] = 8'b0;
    XRAM[26580] = 8'b0;
    XRAM[26581] = 8'b0;
    XRAM[26582] = 8'b0;
    XRAM[26583] = 8'b0;
    XRAM[26584] = 8'b0;
    XRAM[26585] = 8'b0;
    XRAM[26586] = 8'b0;
    XRAM[26587] = 8'b0;
    XRAM[26588] = 8'b0;
    XRAM[26589] = 8'b0;
    XRAM[26590] = 8'b0;
    XRAM[26591] = 8'b0;
    XRAM[26592] = 8'b0;
    XRAM[26593] = 8'b0;
    XRAM[26594] = 8'b0;
    XRAM[26595] = 8'b0;
    XRAM[26596] = 8'b0;
    XRAM[26597] = 8'b0;
    XRAM[26598] = 8'b0;
    XRAM[26599] = 8'b0;
    XRAM[26600] = 8'b0;
    XRAM[26601] = 8'b0;
    XRAM[26602] = 8'b0;
    XRAM[26603] = 8'b0;
    XRAM[26604] = 8'b0;
    XRAM[26605] = 8'b0;
    XRAM[26606] = 8'b0;
    XRAM[26607] = 8'b0;
    XRAM[26608] = 8'b0;
    XRAM[26609] = 8'b0;
    XRAM[26610] = 8'b0;
    XRAM[26611] = 8'b0;
    XRAM[26612] = 8'b0;
    XRAM[26613] = 8'b0;
    XRAM[26614] = 8'b0;
    XRAM[26615] = 8'b0;
    XRAM[26616] = 8'b0;
    XRAM[26617] = 8'b0;
    XRAM[26618] = 8'b0;
    XRAM[26619] = 8'b0;
    XRAM[26620] = 8'b0;
    XRAM[26621] = 8'b0;
    XRAM[26622] = 8'b0;
    XRAM[26623] = 8'b0;
    XRAM[26624] = 8'b0;
    XRAM[26625] = 8'b0;
    XRAM[26626] = 8'b0;
    XRAM[26627] = 8'b0;
    XRAM[26628] = 8'b0;
    XRAM[26629] = 8'b0;
    XRAM[26630] = 8'b0;
    XRAM[26631] = 8'b0;
    XRAM[26632] = 8'b0;
    XRAM[26633] = 8'b0;
    XRAM[26634] = 8'b0;
    XRAM[26635] = 8'b0;
    XRAM[26636] = 8'b0;
    XRAM[26637] = 8'b0;
    XRAM[26638] = 8'b0;
    XRAM[26639] = 8'b0;
    XRAM[26640] = 8'b0;
    XRAM[26641] = 8'b0;
    XRAM[26642] = 8'b0;
    XRAM[26643] = 8'b0;
    XRAM[26644] = 8'b0;
    XRAM[26645] = 8'b0;
    XRAM[26646] = 8'b0;
    XRAM[26647] = 8'b0;
    XRAM[26648] = 8'b0;
    XRAM[26649] = 8'b0;
    XRAM[26650] = 8'b0;
    XRAM[26651] = 8'b0;
    XRAM[26652] = 8'b0;
    XRAM[26653] = 8'b0;
    XRAM[26654] = 8'b0;
    XRAM[26655] = 8'b0;
    XRAM[26656] = 8'b0;
    XRAM[26657] = 8'b0;
    XRAM[26658] = 8'b0;
    XRAM[26659] = 8'b0;
    XRAM[26660] = 8'b0;
    XRAM[26661] = 8'b0;
    XRAM[26662] = 8'b0;
    XRAM[26663] = 8'b0;
    XRAM[26664] = 8'b0;
    XRAM[26665] = 8'b0;
    XRAM[26666] = 8'b0;
    XRAM[26667] = 8'b0;
    XRAM[26668] = 8'b0;
    XRAM[26669] = 8'b0;
    XRAM[26670] = 8'b0;
    XRAM[26671] = 8'b0;
    XRAM[26672] = 8'b0;
    XRAM[26673] = 8'b0;
    XRAM[26674] = 8'b0;
    XRAM[26675] = 8'b0;
    XRAM[26676] = 8'b0;
    XRAM[26677] = 8'b0;
    XRAM[26678] = 8'b0;
    XRAM[26679] = 8'b0;
    XRAM[26680] = 8'b0;
    XRAM[26681] = 8'b0;
    XRAM[26682] = 8'b0;
    XRAM[26683] = 8'b0;
    XRAM[26684] = 8'b0;
    XRAM[26685] = 8'b0;
    XRAM[26686] = 8'b0;
    XRAM[26687] = 8'b0;
    XRAM[26688] = 8'b0;
    XRAM[26689] = 8'b0;
    XRAM[26690] = 8'b0;
    XRAM[26691] = 8'b0;
    XRAM[26692] = 8'b0;
    XRAM[26693] = 8'b0;
    XRAM[26694] = 8'b0;
    XRAM[26695] = 8'b0;
    XRAM[26696] = 8'b0;
    XRAM[26697] = 8'b0;
    XRAM[26698] = 8'b0;
    XRAM[26699] = 8'b0;
    XRAM[26700] = 8'b0;
    XRAM[26701] = 8'b0;
    XRAM[26702] = 8'b0;
    XRAM[26703] = 8'b0;
    XRAM[26704] = 8'b0;
    XRAM[26705] = 8'b0;
    XRAM[26706] = 8'b0;
    XRAM[26707] = 8'b0;
    XRAM[26708] = 8'b0;
    XRAM[26709] = 8'b0;
    XRAM[26710] = 8'b0;
    XRAM[26711] = 8'b0;
    XRAM[26712] = 8'b0;
    XRAM[26713] = 8'b0;
    XRAM[26714] = 8'b0;
    XRAM[26715] = 8'b0;
    XRAM[26716] = 8'b0;
    XRAM[26717] = 8'b0;
    XRAM[26718] = 8'b0;
    XRAM[26719] = 8'b0;
    XRAM[26720] = 8'b0;
    XRAM[26721] = 8'b0;
    XRAM[26722] = 8'b0;
    XRAM[26723] = 8'b0;
    XRAM[26724] = 8'b0;
    XRAM[26725] = 8'b0;
    XRAM[26726] = 8'b0;
    XRAM[26727] = 8'b0;
    XRAM[26728] = 8'b0;
    XRAM[26729] = 8'b0;
    XRAM[26730] = 8'b0;
    XRAM[26731] = 8'b0;
    XRAM[26732] = 8'b0;
    XRAM[26733] = 8'b0;
    XRAM[26734] = 8'b0;
    XRAM[26735] = 8'b0;
    XRAM[26736] = 8'b0;
    XRAM[26737] = 8'b0;
    XRAM[26738] = 8'b0;
    XRAM[26739] = 8'b0;
    XRAM[26740] = 8'b0;
    XRAM[26741] = 8'b0;
    XRAM[26742] = 8'b0;
    XRAM[26743] = 8'b0;
    XRAM[26744] = 8'b0;
    XRAM[26745] = 8'b0;
    XRAM[26746] = 8'b0;
    XRAM[26747] = 8'b0;
    XRAM[26748] = 8'b0;
    XRAM[26749] = 8'b0;
    XRAM[26750] = 8'b0;
    XRAM[26751] = 8'b0;
    XRAM[26752] = 8'b0;
    XRAM[26753] = 8'b0;
    XRAM[26754] = 8'b0;
    XRAM[26755] = 8'b0;
    XRAM[26756] = 8'b0;
    XRAM[26757] = 8'b0;
    XRAM[26758] = 8'b0;
    XRAM[26759] = 8'b0;
    XRAM[26760] = 8'b0;
    XRAM[26761] = 8'b0;
    XRAM[26762] = 8'b0;
    XRAM[26763] = 8'b0;
    XRAM[26764] = 8'b0;
    XRAM[26765] = 8'b0;
    XRAM[26766] = 8'b0;
    XRAM[26767] = 8'b0;
    XRAM[26768] = 8'b0;
    XRAM[26769] = 8'b0;
    XRAM[26770] = 8'b0;
    XRAM[26771] = 8'b0;
    XRAM[26772] = 8'b0;
    XRAM[26773] = 8'b0;
    XRAM[26774] = 8'b0;
    XRAM[26775] = 8'b0;
    XRAM[26776] = 8'b0;
    XRAM[26777] = 8'b0;
    XRAM[26778] = 8'b0;
    XRAM[26779] = 8'b0;
    XRAM[26780] = 8'b0;
    XRAM[26781] = 8'b0;
    XRAM[26782] = 8'b0;
    XRAM[26783] = 8'b0;
    XRAM[26784] = 8'b0;
    XRAM[26785] = 8'b0;
    XRAM[26786] = 8'b0;
    XRAM[26787] = 8'b0;
    XRAM[26788] = 8'b0;
    XRAM[26789] = 8'b0;
    XRAM[26790] = 8'b0;
    XRAM[26791] = 8'b0;
    XRAM[26792] = 8'b0;
    XRAM[26793] = 8'b0;
    XRAM[26794] = 8'b0;
    XRAM[26795] = 8'b0;
    XRAM[26796] = 8'b0;
    XRAM[26797] = 8'b0;
    XRAM[26798] = 8'b0;
    XRAM[26799] = 8'b0;
    XRAM[26800] = 8'b0;
    XRAM[26801] = 8'b0;
    XRAM[26802] = 8'b0;
    XRAM[26803] = 8'b0;
    XRAM[26804] = 8'b0;
    XRAM[26805] = 8'b0;
    XRAM[26806] = 8'b0;
    XRAM[26807] = 8'b0;
    XRAM[26808] = 8'b0;
    XRAM[26809] = 8'b0;
    XRAM[26810] = 8'b0;
    XRAM[26811] = 8'b0;
    XRAM[26812] = 8'b0;
    XRAM[26813] = 8'b0;
    XRAM[26814] = 8'b0;
    XRAM[26815] = 8'b0;
    XRAM[26816] = 8'b0;
    XRAM[26817] = 8'b0;
    XRAM[26818] = 8'b0;
    XRAM[26819] = 8'b0;
    XRAM[26820] = 8'b0;
    XRAM[26821] = 8'b0;
    XRAM[26822] = 8'b0;
    XRAM[26823] = 8'b0;
    XRAM[26824] = 8'b0;
    XRAM[26825] = 8'b0;
    XRAM[26826] = 8'b0;
    XRAM[26827] = 8'b0;
    XRAM[26828] = 8'b0;
    XRAM[26829] = 8'b0;
    XRAM[26830] = 8'b0;
    XRAM[26831] = 8'b0;
    XRAM[26832] = 8'b0;
    XRAM[26833] = 8'b0;
    XRAM[26834] = 8'b0;
    XRAM[26835] = 8'b0;
    XRAM[26836] = 8'b0;
    XRAM[26837] = 8'b0;
    XRAM[26838] = 8'b0;
    XRAM[26839] = 8'b0;
    XRAM[26840] = 8'b0;
    XRAM[26841] = 8'b0;
    XRAM[26842] = 8'b0;
    XRAM[26843] = 8'b0;
    XRAM[26844] = 8'b0;
    XRAM[26845] = 8'b0;
    XRAM[26846] = 8'b0;
    XRAM[26847] = 8'b0;
    XRAM[26848] = 8'b0;
    XRAM[26849] = 8'b0;
    XRAM[26850] = 8'b0;
    XRAM[26851] = 8'b0;
    XRAM[26852] = 8'b0;
    XRAM[26853] = 8'b0;
    XRAM[26854] = 8'b0;
    XRAM[26855] = 8'b0;
    XRAM[26856] = 8'b0;
    XRAM[26857] = 8'b0;
    XRAM[26858] = 8'b0;
    XRAM[26859] = 8'b0;
    XRAM[26860] = 8'b0;
    XRAM[26861] = 8'b0;
    XRAM[26862] = 8'b0;
    XRAM[26863] = 8'b0;
    XRAM[26864] = 8'b0;
    XRAM[26865] = 8'b0;
    XRAM[26866] = 8'b0;
    XRAM[26867] = 8'b0;
    XRAM[26868] = 8'b0;
    XRAM[26869] = 8'b0;
    XRAM[26870] = 8'b0;
    XRAM[26871] = 8'b0;
    XRAM[26872] = 8'b0;
    XRAM[26873] = 8'b0;
    XRAM[26874] = 8'b0;
    XRAM[26875] = 8'b0;
    XRAM[26876] = 8'b0;
    XRAM[26877] = 8'b0;
    XRAM[26878] = 8'b0;
    XRAM[26879] = 8'b0;
    XRAM[26880] = 8'b0;
    XRAM[26881] = 8'b0;
    XRAM[26882] = 8'b0;
    XRAM[26883] = 8'b0;
    XRAM[26884] = 8'b0;
    XRAM[26885] = 8'b0;
    XRAM[26886] = 8'b0;
    XRAM[26887] = 8'b0;
    XRAM[26888] = 8'b0;
    XRAM[26889] = 8'b0;
    XRAM[26890] = 8'b0;
    XRAM[26891] = 8'b0;
    XRAM[26892] = 8'b0;
    XRAM[26893] = 8'b0;
    XRAM[26894] = 8'b0;
    XRAM[26895] = 8'b0;
    XRAM[26896] = 8'b0;
    XRAM[26897] = 8'b0;
    XRAM[26898] = 8'b0;
    XRAM[26899] = 8'b0;
    XRAM[26900] = 8'b0;
    XRAM[26901] = 8'b0;
    XRAM[26902] = 8'b0;
    XRAM[26903] = 8'b0;
    XRAM[26904] = 8'b0;
    XRAM[26905] = 8'b0;
    XRAM[26906] = 8'b0;
    XRAM[26907] = 8'b0;
    XRAM[26908] = 8'b0;
    XRAM[26909] = 8'b0;
    XRAM[26910] = 8'b0;
    XRAM[26911] = 8'b0;
    XRAM[26912] = 8'b0;
    XRAM[26913] = 8'b0;
    XRAM[26914] = 8'b0;
    XRAM[26915] = 8'b0;
    XRAM[26916] = 8'b0;
    XRAM[26917] = 8'b0;
    XRAM[26918] = 8'b0;
    XRAM[26919] = 8'b0;
    XRAM[26920] = 8'b0;
    XRAM[26921] = 8'b0;
    XRAM[26922] = 8'b0;
    XRAM[26923] = 8'b0;
    XRAM[26924] = 8'b0;
    XRAM[26925] = 8'b0;
    XRAM[26926] = 8'b0;
    XRAM[26927] = 8'b0;
    XRAM[26928] = 8'b0;
    XRAM[26929] = 8'b0;
    XRAM[26930] = 8'b0;
    XRAM[26931] = 8'b0;
    XRAM[26932] = 8'b0;
    XRAM[26933] = 8'b0;
    XRAM[26934] = 8'b0;
    XRAM[26935] = 8'b0;
    XRAM[26936] = 8'b0;
    XRAM[26937] = 8'b0;
    XRAM[26938] = 8'b0;
    XRAM[26939] = 8'b0;
    XRAM[26940] = 8'b0;
    XRAM[26941] = 8'b0;
    XRAM[26942] = 8'b0;
    XRAM[26943] = 8'b0;
    XRAM[26944] = 8'b0;
    XRAM[26945] = 8'b0;
    XRAM[26946] = 8'b0;
    XRAM[26947] = 8'b0;
    XRAM[26948] = 8'b0;
    XRAM[26949] = 8'b0;
    XRAM[26950] = 8'b0;
    XRAM[26951] = 8'b0;
    XRAM[26952] = 8'b0;
    XRAM[26953] = 8'b0;
    XRAM[26954] = 8'b0;
    XRAM[26955] = 8'b0;
    XRAM[26956] = 8'b0;
    XRAM[26957] = 8'b0;
    XRAM[26958] = 8'b0;
    XRAM[26959] = 8'b0;
    XRAM[26960] = 8'b0;
    XRAM[26961] = 8'b0;
    XRAM[26962] = 8'b0;
    XRAM[26963] = 8'b0;
    XRAM[26964] = 8'b0;
    XRAM[26965] = 8'b0;
    XRAM[26966] = 8'b0;
    XRAM[26967] = 8'b0;
    XRAM[26968] = 8'b0;
    XRAM[26969] = 8'b0;
    XRAM[26970] = 8'b0;
    XRAM[26971] = 8'b0;
    XRAM[26972] = 8'b0;
    XRAM[26973] = 8'b0;
    XRAM[26974] = 8'b0;
    XRAM[26975] = 8'b0;
    XRAM[26976] = 8'b0;
    XRAM[26977] = 8'b0;
    XRAM[26978] = 8'b0;
    XRAM[26979] = 8'b0;
    XRAM[26980] = 8'b0;
    XRAM[26981] = 8'b0;
    XRAM[26982] = 8'b0;
    XRAM[26983] = 8'b0;
    XRAM[26984] = 8'b0;
    XRAM[26985] = 8'b0;
    XRAM[26986] = 8'b0;
    XRAM[26987] = 8'b0;
    XRAM[26988] = 8'b0;
    XRAM[26989] = 8'b0;
    XRAM[26990] = 8'b0;
    XRAM[26991] = 8'b0;
    XRAM[26992] = 8'b0;
    XRAM[26993] = 8'b0;
    XRAM[26994] = 8'b0;
    XRAM[26995] = 8'b0;
    XRAM[26996] = 8'b0;
    XRAM[26997] = 8'b0;
    XRAM[26998] = 8'b0;
    XRAM[26999] = 8'b0;
    XRAM[27000] = 8'b0;
    XRAM[27001] = 8'b0;
    XRAM[27002] = 8'b0;
    XRAM[27003] = 8'b0;
    XRAM[27004] = 8'b0;
    XRAM[27005] = 8'b0;
    XRAM[27006] = 8'b0;
    XRAM[27007] = 8'b0;
    XRAM[27008] = 8'b0;
    XRAM[27009] = 8'b0;
    XRAM[27010] = 8'b0;
    XRAM[27011] = 8'b0;
    XRAM[27012] = 8'b0;
    XRAM[27013] = 8'b0;
    XRAM[27014] = 8'b0;
    XRAM[27015] = 8'b0;
    XRAM[27016] = 8'b0;
    XRAM[27017] = 8'b0;
    XRAM[27018] = 8'b0;
    XRAM[27019] = 8'b0;
    XRAM[27020] = 8'b0;
    XRAM[27021] = 8'b0;
    XRAM[27022] = 8'b0;
    XRAM[27023] = 8'b0;
    XRAM[27024] = 8'b0;
    XRAM[27025] = 8'b0;
    XRAM[27026] = 8'b0;
    XRAM[27027] = 8'b0;
    XRAM[27028] = 8'b0;
    XRAM[27029] = 8'b0;
    XRAM[27030] = 8'b0;
    XRAM[27031] = 8'b0;
    XRAM[27032] = 8'b0;
    XRAM[27033] = 8'b0;
    XRAM[27034] = 8'b0;
    XRAM[27035] = 8'b0;
    XRAM[27036] = 8'b0;
    XRAM[27037] = 8'b0;
    XRAM[27038] = 8'b0;
    XRAM[27039] = 8'b0;
    XRAM[27040] = 8'b0;
    XRAM[27041] = 8'b0;
    XRAM[27042] = 8'b0;
    XRAM[27043] = 8'b0;
    XRAM[27044] = 8'b0;
    XRAM[27045] = 8'b0;
    XRAM[27046] = 8'b0;
    XRAM[27047] = 8'b0;
    XRAM[27048] = 8'b0;
    XRAM[27049] = 8'b0;
    XRAM[27050] = 8'b0;
    XRAM[27051] = 8'b0;
    XRAM[27052] = 8'b0;
    XRAM[27053] = 8'b0;
    XRAM[27054] = 8'b0;
    XRAM[27055] = 8'b0;
    XRAM[27056] = 8'b0;
    XRAM[27057] = 8'b0;
    XRAM[27058] = 8'b0;
    XRAM[27059] = 8'b0;
    XRAM[27060] = 8'b0;
    XRAM[27061] = 8'b0;
    XRAM[27062] = 8'b0;
    XRAM[27063] = 8'b0;
    XRAM[27064] = 8'b0;
    XRAM[27065] = 8'b0;
    XRAM[27066] = 8'b0;
    XRAM[27067] = 8'b0;
    XRAM[27068] = 8'b0;
    XRAM[27069] = 8'b0;
    XRAM[27070] = 8'b0;
    XRAM[27071] = 8'b0;
    XRAM[27072] = 8'b0;
    XRAM[27073] = 8'b0;
    XRAM[27074] = 8'b0;
    XRAM[27075] = 8'b0;
    XRAM[27076] = 8'b0;
    XRAM[27077] = 8'b0;
    XRAM[27078] = 8'b0;
    XRAM[27079] = 8'b0;
    XRAM[27080] = 8'b0;
    XRAM[27081] = 8'b0;
    XRAM[27082] = 8'b0;
    XRAM[27083] = 8'b0;
    XRAM[27084] = 8'b0;
    XRAM[27085] = 8'b0;
    XRAM[27086] = 8'b0;
    XRAM[27087] = 8'b0;
    XRAM[27088] = 8'b0;
    XRAM[27089] = 8'b0;
    XRAM[27090] = 8'b0;
    XRAM[27091] = 8'b0;
    XRAM[27092] = 8'b0;
    XRAM[27093] = 8'b0;
    XRAM[27094] = 8'b0;
    XRAM[27095] = 8'b0;
    XRAM[27096] = 8'b0;
    XRAM[27097] = 8'b0;
    XRAM[27098] = 8'b0;
    XRAM[27099] = 8'b0;
    XRAM[27100] = 8'b0;
    XRAM[27101] = 8'b0;
    XRAM[27102] = 8'b0;
    XRAM[27103] = 8'b0;
    XRAM[27104] = 8'b0;
    XRAM[27105] = 8'b0;
    XRAM[27106] = 8'b0;
    XRAM[27107] = 8'b0;
    XRAM[27108] = 8'b0;
    XRAM[27109] = 8'b0;
    XRAM[27110] = 8'b0;
    XRAM[27111] = 8'b0;
    XRAM[27112] = 8'b0;
    XRAM[27113] = 8'b0;
    XRAM[27114] = 8'b0;
    XRAM[27115] = 8'b0;
    XRAM[27116] = 8'b0;
    XRAM[27117] = 8'b0;
    XRAM[27118] = 8'b0;
    XRAM[27119] = 8'b0;
    XRAM[27120] = 8'b0;
    XRAM[27121] = 8'b0;
    XRAM[27122] = 8'b0;
    XRAM[27123] = 8'b0;
    XRAM[27124] = 8'b0;
    XRAM[27125] = 8'b0;
    XRAM[27126] = 8'b0;
    XRAM[27127] = 8'b0;
    XRAM[27128] = 8'b0;
    XRAM[27129] = 8'b0;
    XRAM[27130] = 8'b0;
    XRAM[27131] = 8'b0;
    XRAM[27132] = 8'b0;
    XRAM[27133] = 8'b0;
    XRAM[27134] = 8'b0;
    XRAM[27135] = 8'b0;
    XRAM[27136] = 8'b0;
    XRAM[27137] = 8'b0;
    XRAM[27138] = 8'b0;
    XRAM[27139] = 8'b0;
    XRAM[27140] = 8'b0;
    XRAM[27141] = 8'b0;
    XRAM[27142] = 8'b0;
    XRAM[27143] = 8'b0;
    XRAM[27144] = 8'b0;
    XRAM[27145] = 8'b0;
    XRAM[27146] = 8'b0;
    XRAM[27147] = 8'b0;
    XRAM[27148] = 8'b0;
    XRAM[27149] = 8'b0;
    XRAM[27150] = 8'b0;
    XRAM[27151] = 8'b0;
    XRAM[27152] = 8'b0;
    XRAM[27153] = 8'b0;
    XRAM[27154] = 8'b0;
    XRAM[27155] = 8'b0;
    XRAM[27156] = 8'b0;
    XRAM[27157] = 8'b0;
    XRAM[27158] = 8'b0;
    XRAM[27159] = 8'b0;
    XRAM[27160] = 8'b0;
    XRAM[27161] = 8'b0;
    XRAM[27162] = 8'b0;
    XRAM[27163] = 8'b0;
    XRAM[27164] = 8'b0;
    XRAM[27165] = 8'b0;
    XRAM[27166] = 8'b0;
    XRAM[27167] = 8'b0;
    XRAM[27168] = 8'b0;
    XRAM[27169] = 8'b0;
    XRAM[27170] = 8'b0;
    XRAM[27171] = 8'b0;
    XRAM[27172] = 8'b0;
    XRAM[27173] = 8'b0;
    XRAM[27174] = 8'b0;
    XRAM[27175] = 8'b0;
    XRAM[27176] = 8'b0;
    XRAM[27177] = 8'b0;
    XRAM[27178] = 8'b0;
    XRAM[27179] = 8'b0;
    XRAM[27180] = 8'b0;
    XRAM[27181] = 8'b0;
    XRAM[27182] = 8'b0;
    XRAM[27183] = 8'b0;
    XRAM[27184] = 8'b0;
    XRAM[27185] = 8'b0;
    XRAM[27186] = 8'b0;
    XRAM[27187] = 8'b0;
    XRAM[27188] = 8'b0;
    XRAM[27189] = 8'b0;
    XRAM[27190] = 8'b0;
    XRAM[27191] = 8'b0;
    XRAM[27192] = 8'b0;
    XRAM[27193] = 8'b0;
    XRAM[27194] = 8'b0;
    XRAM[27195] = 8'b0;
    XRAM[27196] = 8'b0;
    XRAM[27197] = 8'b0;
    XRAM[27198] = 8'b0;
    XRAM[27199] = 8'b0;
    XRAM[27200] = 8'b0;
    XRAM[27201] = 8'b0;
    XRAM[27202] = 8'b0;
    XRAM[27203] = 8'b0;
    XRAM[27204] = 8'b0;
    XRAM[27205] = 8'b0;
    XRAM[27206] = 8'b0;
    XRAM[27207] = 8'b0;
    XRAM[27208] = 8'b0;
    XRAM[27209] = 8'b0;
    XRAM[27210] = 8'b0;
    XRAM[27211] = 8'b0;
    XRAM[27212] = 8'b0;
    XRAM[27213] = 8'b0;
    XRAM[27214] = 8'b0;
    XRAM[27215] = 8'b0;
    XRAM[27216] = 8'b0;
    XRAM[27217] = 8'b0;
    XRAM[27218] = 8'b0;
    XRAM[27219] = 8'b0;
    XRAM[27220] = 8'b0;
    XRAM[27221] = 8'b0;
    XRAM[27222] = 8'b0;
    XRAM[27223] = 8'b0;
    XRAM[27224] = 8'b0;
    XRAM[27225] = 8'b0;
    XRAM[27226] = 8'b0;
    XRAM[27227] = 8'b0;
    XRAM[27228] = 8'b0;
    XRAM[27229] = 8'b0;
    XRAM[27230] = 8'b0;
    XRAM[27231] = 8'b0;
    XRAM[27232] = 8'b0;
    XRAM[27233] = 8'b0;
    XRAM[27234] = 8'b0;
    XRAM[27235] = 8'b0;
    XRAM[27236] = 8'b0;
    XRAM[27237] = 8'b0;
    XRAM[27238] = 8'b0;
    XRAM[27239] = 8'b0;
    XRAM[27240] = 8'b0;
    XRAM[27241] = 8'b0;
    XRAM[27242] = 8'b0;
    XRAM[27243] = 8'b0;
    XRAM[27244] = 8'b0;
    XRAM[27245] = 8'b0;
    XRAM[27246] = 8'b0;
    XRAM[27247] = 8'b0;
    XRAM[27248] = 8'b0;
    XRAM[27249] = 8'b0;
    XRAM[27250] = 8'b0;
    XRAM[27251] = 8'b0;
    XRAM[27252] = 8'b0;
    XRAM[27253] = 8'b0;
    XRAM[27254] = 8'b0;
    XRAM[27255] = 8'b0;
    XRAM[27256] = 8'b0;
    XRAM[27257] = 8'b0;
    XRAM[27258] = 8'b0;
    XRAM[27259] = 8'b0;
    XRAM[27260] = 8'b0;
    XRAM[27261] = 8'b0;
    XRAM[27262] = 8'b0;
    XRAM[27263] = 8'b0;
    XRAM[27264] = 8'b0;
    XRAM[27265] = 8'b0;
    XRAM[27266] = 8'b0;
    XRAM[27267] = 8'b0;
    XRAM[27268] = 8'b0;
    XRAM[27269] = 8'b0;
    XRAM[27270] = 8'b0;
    XRAM[27271] = 8'b0;
    XRAM[27272] = 8'b0;
    XRAM[27273] = 8'b0;
    XRAM[27274] = 8'b0;
    XRAM[27275] = 8'b0;
    XRAM[27276] = 8'b0;
    XRAM[27277] = 8'b0;
    XRAM[27278] = 8'b0;
    XRAM[27279] = 8'b0;
    XRAM[27280] = 8'b0;
    XRAM[27281] = 8'b0;
    XRAM[27282] = 8'b0;
    XRAM[27283] = 8'b0;
    XRAM[27284] = 8'b0;
    XRAM[27285] = 8'b0;
    XRAM[27286] = 8'b0;
    XRAM[27287] = 8'b0;
    XRAM[27288] = 8'b0;
    XRAM[27289] = 8'b0;
    XRAM[27290] = 8'b0;
    XRAM[27291] = 8'b0;
    XRAM[27292] = 8'b0;
    XRAM[27293] = 8'b0;
    XRAM[27294] = 8'b0;
    XRAM[27295] = 8'b0;
    XRAM[27296] = 8'b0;
    XRAM[27297] = 8'b0;
    XRAM[27298] = 8'b0;
    XRAM[27299] = 8'b0;
    XRAM[27300] = 8'b0;
    XRAM[27301] = 8'b0;
    XRAM[27302] = 8'b0;
    XRAM[27303] = 8'b0;
    XRAM[27304] = 8'b0;
    XRAM[27305] = 8'b0;
    XRAM[27306] = 8'b0;
    XRAM[27307] = 8'b0;
    XRAM[27308] = 8'b0;
    XRAM[27309] = 8'b0;
    XRAM[27310] = 8'b0;
    XRAM[27311] = 8'b0;
    XRAM[27312] = 8'b0;
    XRAM[27313] = 8'b0;
    XRAM[27314] = 8'b0;
    XRAM[27315] = 8'b0;
    XRAM[27316] = 8'b0;
    XRAM[27317] = 8'b0;
    XRAM[27318] = 8'b0;
    XRAM[27319] = 8'b0;
    XRAM[27320] = 8'b0;
    XRAM[27321] = 8'b0;
    XRAM[27322] = 8'b0;
    XRAM[27323] = 8'b0;
    XRAM[27324] = 8'b0;
    XRAM[27325] = 8'b0;
    XRAM[27326] = 8'b0;
    XRAM[27327] = 8'b0;
    XRAM[27328] = 8'b0;
    XRAM[27329] = 8'b0;
    XRAM[27330] = 8'b0;
    XRAM[27331] = 8'b0;
    XRAM[27332] = 8'b0;
    XRAM[27333] = 8'b0;
    XRAM[27334] = 8'b0;
    XRAM[27335] = 8'b0;
    XRAM[27336] = 8'b0;
    XRAM[27337] = 8'b0;
    XRAM[27338] = 8'b0;
    XRAM[27339] = 8'b0;
    XRAM[27340] = 8'b0;
    XRAM[27341] = 8'b0;
    XRAM[27342] = 8'b0;
    XRAM[27343] = 8'b0;
    XRAM[27344] = 8'b0;
    XRAM[27345] = 8'b0;
    XRAM[27346] = 8'b0;
    XRAM[27347] = 8'b0;
    XRAM[27348] = 8'b0;
    XRAM[27349] = 8'b0;
    XRAM[27350] = 8'b0;
    XRAM[27351] = 8'b0;
    XRAM[27352] = 8'b0;
    XRAM[27353] = 8'b0;
    XRAM[27354] = 8'b0;
    XRAM[27355] = 8'b0;
    XRAM[27356] = 8'b0;
    XRAM[27357] = 8'b0;
    XRAM[27358] = 8'b0;
    XRAM[27359] = 8'b0;
    XRAM[27360] = 8'b0;
    XRAM[27361] = 8'b0;
    XRAM[27362] = 8'b0;
    XRAM[27363] = 8'b0;
    XRAM[27364] = 8'b0;
    XRAM[27365] = 8'b0;
    XRAM[27366] = 8'b0;
    XRAM[27367] = 8'b0;
    XRAM[27368] = 8'b0;
    XRAM[27369] = 8'b0;
    XRAM[27370] = 8'b0;
    XRAM[27371] = 8'b0;
    XRAM[27372] = 8'b0;
    XRAM[27373] = 8'b0;
    XRAM[27374] = 8'b0;
    XRAM[27375] = 8'b0;
    XRAM[27376] = 8'b0;
    XRAM[27377] = 8'b0;
    XRAM[27378] = 8'b0;
    XRAM[27379] = 8'b0;
    XRAM[27380] = 8'b0;
    XRAM[27381] = 8'b0;
    XRAM[27382] = 8'b0;
    XRAM[27383] = 8'b0;
    XRAM[27384] = 8'b0;
    XRAM[27385] = 8'b0;
    XRAM[27386] = 8'b0;
    XRAM[27387] = 8'b0;
    XRAM[27388] = 8'b0;
    XRAM[27389] = 8'b0;
    XRAM[27390] = 8'b0;
    XRAM[27391] = 8'b0;
    XRAM[27392] = 8'b0;
    XRAM[27393] = 8'b0;
    XRAM[27394] = 8'b0;
    XRAM[27395] = 8'b0;
    XRAM[27396] = 8'b0;
    XRAM[27397] = 8'b0;
    XRAM[27398] = 8'b0;
    XRAM[27399] = 8'b0;
    XRAM[27400] = 8'b0;
    XRAM[27401] = 8'b0;
    XRAM[27402] = 8'b0;
    XRAM[27403] = 8'b0;
    XRAM[27404] = 8'b0;
    XRAM[27405] = 8'b0;
    XRAM[27406] = 8'b0;
    XRAM[27407] = 8'b0;
    XRAM[27408] = 8'b0;
    XRAM[27409] = 8'b0;
    XRAM[27410] = 8'b0;
    XRAM[27411] = 8'b0;
    XRAM[27412] = 8'b0;
    XRAM[27413] = 8'b0;
    XRAM[27414] = 8'b0;
    XRAM[27415] = 8'b0;
    XRAM[27416] = 8'b0;
    XRAM[27417] = 8'b0;
    XRAM[27418] = 8'b0;
    XRAM[27419] = 8'b0;
    XRAM[27420] = 8'b0;
    XRAM[27421] = 8'b0;
    XRAM[27422] = 8'b0;
    XRAM[27423] = 8'b0;
    XRAM[27424] = 8'b0;
    XRAM[27425] = 8'b0;
    XRAM[27426] = 8'b0;
    XRAM[27427] = 8'b0;
    XRAM[27428] = 8'b0;
    XRAM[27429] = 8'b0;
    XRAM[27430] = 8'b0;
    XRAM[27431] = 8'b0;
    XRAM[27432] = 8'b0;
    XRAM[27433] = 8'b0;
    XRAM[27434] = 8'b0;
    XRAM[27435] = 8'b0;
    XRAM[27436] = 8'b0;
    XRAM[27437] = 8'b0;
    XRAM[27438] = 8'b0;
    XRAM[27439] = 8'b0;
    XRAM[27440] = 8'b0;
    XRAM[27441] = 8'b0;
    XRAM[27442] = 8'b0;
    XRAM[27443] = 8'b0;
    XRAM[27444] = 8'b0;
    XRAM[27445] = 8'b0;
    XRAM[27446] = 8'b0;
    XRAM[27447] = 8'b0;
    XRAM[27448] = 8'b0;
    XRAM[27449] = 8'b0;
    XRAM[27450] = 8'b0;
    XRAM[27451] = 8'b0;
    XRAM[27452] = 8'b0;
    XRAM[27453] = 8'b0;
    XRAM[27454] = 8'b0;
    XRAM[27455] = 8'b0;
    XRAM[27456] = 8'b0;
    XRAM[27457] = 8'b0;
    XRAM[27458] = 8'b0;
    XRAM[27459] = 8'b0;
    XRAM[27460] = 8'b0;
    XRAM[27461] = 8'b0;
    XRAM[27462] = 8'b0;
    XRAM[27463] = 8'b0;
    XRAM[27464] = 8'b0;
    XRAM[27465] = 8'b0;
    XRAM[27466] = 8'b0;
    XRAM[27467] = 8'b0;
    XRAM[27468] = 8'b0;
    XRAM[27469] = 8'b0;
    XRAM[27470] = 8'b0;
    XRAM[27471] = 8'b0;
    XRAM[27472] = 8'b0;
    XRAM[27473] = 8'b0;
    XRAM[27474] = 8'b0;
    XRAM[27475] = 8'b0;
    XRAM[27476] = 8'b0;
    XRAM[27477] = 8'b0;
    XRAM[27478] = 8'b0;
    XRAM[27479] = 8'b0;
    XRAM[27480] = 8'b0;
    XRAM[27481] = 8'b0;
    XRAM[27482] = 8'b0;
    XRAM[27483] = 8'b0;
    XRAM[27484] = 8'b0;
    XRAM[27485] = 8'b0;
    XRAM[27486] = 8'b0;
    XRAM[27487] = 8'b0;
    XRAM[27488] = 8'b0;
    XRAM[27489] = 8'b0;
    XRAM[27490] = 8'b0;
    XRAM[27491] = 8'b0;
    XRAM[27492] = 8'b0;
    XRAM[27493] = 8'b0;
    XRAM[27494] = 8'b0;
    XRAM[27495] = 8'b0;
    XRAM[27496] = 8'b0;
    XRAM[27497] = 8'b0;
    XRAM[27498] = 8'b0;
    XRAM[27499] = 8'b0;
    XRAM[27500] = 8'b0;
    XRAM[27501] = 8'b0;
    XRAM[27502] = 8'b0;
    XRAM[27503] = 8'b0;
    XRAM[27504] = 8'b0;
    XRAM[27505] = 8'b0;
    XRAM[27506] = 8'b0;
    XRAM[27507] = 8'b0;
    XRAM[27508] = 8'b0;
    XRAM[27509] = 8'b0;
    XRAM[27510] = 8'b0;
    XRAM[27511] = 8'b0;
    XRAM[27512] = 8'b0;
    XRAM[27513] = 8'b0;
    XRAM[27514] = 8'b0;
    XRAM[27515] = 8'b0;
    XRAM[27516] = 8'b0;
    XRAM[27517] = 8'b0;
    XRAM[27518] = 8'b0;
    XRAM[27519] = 8'b0;
    XRAM[27520] = 8'b0;
    XRAM[27521] = 8'b0;
    XRAM[27522] = 8'b0;
    XRAM[27523] = 8'b0;
    XRAM[27524] = 8'b0;
    XRAM[27525] = 8'b0;
    XRAM[27526] = 8'b0;
    XRAM[27527] = 8'b0;
    XRAM[27528] = 8'b0;
    XRAM[27529] = 8'b0;
    XRAM[27530] = 8'b0;
    XRAM[27531] = 8'b0;
    XRAM[27532] = 8'b0;
    XRAM[27533] = 8'b0;
    XRAM[27534] = 8'b0;
    XRAM[27535] = 8'b0;
    XRAM[27536] = 8'b0;
    XRAM[27537] = 8'b0;
    XRAM[27538] = 8'b0;
    XRAM[27539] = 8'b0;
    XRAM[27540] = 8'b0;
    XRAM[27541] = 8'b0;
    XRAM[27542] = 8'b0;
    XRAM[27543] = 8'b0;
    XRAM[27544] = 8'b0;
    XRAM[27545] = 8'b0;
    XRAM[27546] = 8'b0;
    XRAM[27547] = 8'b0;
    XRAM[27548] = 8'b0;
    XRAM[27549] = 8'b0;
    XRAM[27550] = 8'b0;
    XRAM[27551] = 8'b0;
    XRAM[27552] = 8'b0;
    XRAM[27553] = 8'b0;
    XRAM[27554] = 8'b0;
    XRAM[27555] = 8'b0;
    XRAM[27556] = 8'b0;
    XRAM[27557] = 8'b0;
    XRAM[27558] = 8'b0;
    XRAM[27559] = 8'b0;
    XRAM[27560] = 8'b0;
    XRAM[27561] = 8'b0;
    XRAM[27562] = 8'b0;
    XRAM[27563] = 8'b0;
    XRAM[27564] = 8'b0;
    XRAM[27565] = 8'b0;
    XRAM[27566] = 8'b0;
    XRAM[27567] = 8'b0;
    XRAM[27568] = 8'b0;
    XRAM[27569] = 8'b0;
    XRAM[27570] = 8'b0;
    XRAM[27571] = 8'b0;
    XRAM[27572] = 8'b0;
    XRAM[27573] = 8'b0;
    XRAM[27574] = 8'b0;
    XRAM[27575] = 8'b0;
    XRAM[27576] = 8'b0;
    XRAM[27577] = 8'b0;
    XRAM[27578] = 8'b0;
    XRAM[27579] = 8'b0;
    XRAM[27580] = 8'b0;
    XRAM[27581] = 8'b0;
    XRAM[27582] = 8'b0;
    XRAM[27583] = 8'b0;
    XRAM[27584] = 8'b0;
    XRAM[27585] = 8'b0;
    XRAM[27586] = 8'b0;
    XRAM[27587] = 8'b0;
    XRAM[27588] = 8'b0;
    XRAM[27589] = 8'b0;
    XRAM[27590] = 8'b0;
    XRAM[27591] = 8'b0;
    XRAM[27592] = 8'b0;
    XRAM[27593] = 8'b0;
    XRAM[27594] = 8'b0;
    XRAM[27595] = 8'b0;
    XRAM[27596] = 8'b0;
    XRAM[27597] = 8'b0;
    XRAM[27598] = 8'b0;
    XRAM[27599] = 8'b0;
    XRAM[27600] = 8'b0;
    XRAM[27601] = 8'b0;
    XRAM[27602] = 8'b0;
    XRAM[27603] = 8'b0;
    XRAM[27604] = 8'b0;
    XRAM[27605] = 8'b0;
    XRAM[27606] = 8'b0;
    XRAM[27607] = 8'b0;
    XRAM[27608] = 8'b0;
    XRAM[27609] = 8'b0;
    XRAM[27610] = 8'b0;
    XRAM[27611] = 8'b0;
    XRAM[27612] = 8'b0;
    XRAM[27613] = 8'b0;
    XRAM[27614] = 8'b0;
    XRAM[27615] = 8'b0;
    XRAM[27616] = 8'b0;
    XRAM[27617] = 8'b0;
    XRAM[27618] = 8'b0;
    XRAM[27619] = 8'b0;
    XRAM[27620] = 8'b0;
    XRAM[27621] = 8'b0;
    XRAM[27622] = 8'b0;
    XRAM[27623] = 8'b0;
    XRAM[27624] = 8'b0;
    XRAM[27625] = 8'b0;
    XRAM[27626] = 8'b0;
    XRAM[27627] = 8'b0;
    XRAM[27628] = 8'b0;
    XRAM[27629] = 8'b0;
    XRAM[27630] = 8'b0;
    XRAM[27631] = 8'b0;
    XRAM[27632] = 8'b0;
    XRAM[27633] = 8'b0;
    XRAM[27634] = 8'b0;
    XRAM[27635] = 8'b0;
    XRAM[27636] = 8'b0;
    XRAM[27637] = 8'b0;
    XRAM[27638] = 8'b0;
    XRAM[27639] = 8'b0;
    XRAM[27640] = 8'b0;
    XRAM[27641] = 8'b0;
    XRAM[27642] = 8'b0;
    XRAM[27643] = 8'b0;
    XRAM[27644] = 8'b0;
    XRAM[27645] = 8'b0;
    XRAM[27646] = 8'b0;
    XRAM[27647] = 8'b0;
    XRAM[27648] = 8'b0;
    XRAM[27649] = 8'b0;
    XRAM[27650] = 8'b0;
    XRAM[27651] = 8'b0;
    XRAM[27652] = 8'b0;
    XRAM[27653] = 8'b0;
    XRAM[27654] = 8'b0;
    XRAM[27655] = 8'b0;
    XRAM[27656] = 8'b0;
    XRAM[27657] = 8'b0;
    XRAM[27658] = 8'b0;
    XRAM[27659] = 8'b0;
    XRAM[27660] = 8'b0;
    XRAM[27661] = 8'b0;
    XRAM[27662] = 8'b0;
    XRAM[27663] = 8'b0;
    XRAM[27664] = 8'b0;
    XRAM[27665] = 8'b0;
    XRAM[27666] = 8'b0;
    XRAM[27667] = 8'b0;
    XRAM[27668] = 8'b0;
    XRAM[27669] = 8'b0;
    XRAM[27670] = 8'b0;
    XRAM[27671] = 8'b0;
    XRAM[27672] = 8'b0;
    XRAM[27673] = 8'b0;
    XRAM[27674] = 8'b0;
    XRAM[27675] = 8'b0;
    XRAM[27676] = 8'b0;
    XRAM[27677] = 8'b0;
    XRAM[27678] = 8'b0;
    XRAM[27679] = 8'b0;
    XRAM[27680] = 8'b0;
    XRAM[27681] = 8'b0;
    XRAM[27682] = 8'b0;
    XRAM[27683] = 8'b0;
    XRAM[27684] = 8'b0;
    XRAM[27685] = 8'b0;
    XRAM[27686] = 8'b0;
    XRAM[27687] = 8'b0;
    XRAM[27688] = 8'b0;
    XRAM[27689] = 8'b0;
    XRAM[27690] = 8'b0;
    XRAM[27691] = 8'b0;
    XRAM[27692] = 8'b0;
    XRAM[27693] = 8'b0;
    XRAM[27694] = 8'b0;
    XRAM[27695] = 8'b0;
    XRAM[27696] = 8'b0;
    XRAM[27697] = 8'b0;
    XRAM[27698] = 8'b0;
    XRAM[27699] = 8'b0;
    XRAM[27700] = 8'b0;
    XRAM[27701] = 8'b0;
    XRAM[27702] = 8'b0;
    XRAM[27703] = 8'b0;
    XRAM[27704] = 8'b0;
    XRAM[27705] = 8'b0;
    XRAM[27706] = 8'b0;
    XRAM[27707] = 8'b0;
    XRAM[27708] = 8'b0;
    XRAM[27709] = 8'b0;
    XRAM[27710] = 8'b0;
    XRAM[27711] = 8'b0;
    XRAM[27712] = 8'b0;
    XRAM[27713] = 8'b0;
    XRAM[27714] = 8'b0;
    XRAM[27715] = 8'b0;
    XRAM[27716] = 8'b0;
    XRAM[27717] = 8'b0;
    XRAM[27718] = 8'b0;
    XRAM[27719] = 8'b0;
    XRAM[27720] = 8'b0;
    XRAM[27721] = 8'b0;
    XRAM[27722] = 8'b0;
    XRAM[27723] = 8'b0;
    XRAM[27724] = 8'b0;
    XRAM[27725] = 8'b0;
    XRAM[27726] = 8'b0;
    XRAM[27727] = 8'b0;
    XRAM[27728] = 8'b0;
    XRAM[27729] = 8'b0;
    XRAM[27730] = 8'b0;
    XRAM[27731] = 8'b0;
    XRAM[27732] = 8'b0;
    XRAM[27733] = 8'b0;
    XRAM[27734] = 8'b0;
    XRAM[27735] = 8'b0;
    XRAM[27736] = 8'b0;
    XRAM[27737] = 8'b0;
    XRAM[27738] = 8'b0;
    XRAM[27739] = 8'b0;
    XRAM[27740] = 8'b0;
    XRAM[27741] = 8'b0;
    XRAM[27742] = 8'b0;
    XRAM[27743] = 8'b0;
    XRAM[27744] = 8'b0;
    XRAM[27745] = 8'b0;
    XRAM[27746] = 8'b0;
    XRAM[27747] = 8'b0;
    XRAM[27748] = 8'b0;
    XRAM[27749] = 8'b0;
    XRAM[27750] = 8'b0;
    XRAM[27751] = 8'b0;
    XRAM[27752] = 8'b0;
    XRAM[27753] = 8'b0;
    XRAM[27754] = 8'b0;
    XRAM[27755] = 8'b0;
    XRAM[27756] = 8'b0;
    XRAM[27757] = 8'b0;
    XRAM[27758] = 8'b0;
    XRAM[27759] = 8'b0;
    XRAM[27760] = 8'b0;
    XRAM[27761] = 8'b0;
    XRAM[27762] = 8'b0;
    XRAM[27763] = 8'b0;
    XRAM[27764] = 8'b0;
    XRAM[27765] = 8'b0;
    XRAM[27766] = 8'b0;
    XRAM[27767] = 8'b0;
    XRAM[27768] = 8'b0;
    XRAM[27769] = 8'b0;
    XRAM[27770] = 8'b0;
    XRAM[27771] = 8'b0;
    XRAM[27772] = 8'b0;
    XRAM[27773] = 8'b0;
    XRAM[27774] = 8'b0;
    XRAM[27775] = 8'b0;
    XRAM[27776] = 8'b0;
    XRAM[27777] = 8'b0;
    XRAM[27778] = 8'b0;
    XRAM[27779] = 8'b0;
    XRAM[27780] = 8'b0;
    XRAM[27781] = 8'b0;
    XRAM[27782] = 8'b0;
    XRAM[27783] = 8'b0;
    XRAM[27784] = 8'b0;
    XRAM[27785] = 8'b0;
    XRAM[27786] = 8'b0;
    XRAM[27787] = 8'b0;
    XRAM[27788] = 8'b0;
    XRAM[27789] = 8'b0;
    XRAM[27790] = 8'b0;
    XRAM[27791] = 8'b0;
    XRAM[27792] = 8'b0;
    XRAM[27793] = 8'b0;
    XRAM[27794] = 8'b0;
    XRAM[27795] = 8'b0;
    XRAM[27796] = 8'b0;
    XRAM[27797] = 8'b0;
    XRAM[27798] = 8'b0;
    XRAM[27799] = 8'b0;
    XRAM[27800] = 8'b0;
    XRAM[27801] = 8'b0;
    XRAM[27802] = 8'b0;
    XRAM[27803] = 8'b0;
    XRAM[27804] = 8'b0;
    XRAM[27805] = 8'b0;
    XRAM[27806] = 8'b0;
    XRAM[27807] = 8'b0;
    XRAM[27808] = 8'b0;
    XRAM[27809] = 8'b0;
    XRAM[27810] = 8'b0;
    XRAM[27811] = 8'b0;
    XRAM[27812] = 8'b0;
    XRAM[27813] = 8'b0;
    XRAM[27814] = 8'b0;
    XRAM[27815] = 8'b0;
    XRAM[27816] = 8'b0;
    XRAM[27817] = 8'b0;
    XRAM[27818] = 8'b0;
    XRAM[27819] = 8'b0;
    XRAM[27820] = 8'b0;
    XRAM[27821] = 8'b0;
    XRAM[27822] = 8'b0;
    XRAM[27823] = 8'b0;
    XRAM[27824] = 8'b0;
    XRAM[27825] = 8'b0;
    XRAM[27826] = 8'b0;
    XRAM[27827] = 8'b0;
    XRAM[27828] = 8'b0;
    XRAM[27829] = 8'b0;
    XRAM[27830] = 8'b0;
    XRAM[27831] = 8'b0;
    XRAM[27832] = 8'b0;
    XRAM[27833] = 8'b0;
    XRAM[27834] = 8'b0;
    XRAM[27835] = 8'b0;
    XRAM[27836] = 8'b0;
    XRAM[27837] = 8'b0;
    XRAM[27838] = 8'b0;
    XRAM[27839] = 8'b0;
    XRAM[27840] = 8'b0;
    XRAM[27841] = 8'b0;
    XRAM[27842] = 8'b0;
    XRAM[27843] = 8'b0;
    XRAM[27844] = 8'b0;
    XRAM[27845] = 8'b0;
    XRAM[27846] = 8'b0;
    XRAM[27847] = 8'b0;
    XRAM[27848] = 8'b0;
    XRAM[27849] = 8'b0;
    XRAM[27850] = 8'b0;
    XRAM[27851] = 8'b0;
    XRAM[27852] = 8'b0;
    XRAM[27853] = 8'b0;
    XRAM[27854] = 8'b0;
    XRAM[27855] = 8'b0;
    XRAM[27856] = 8'b0;
    XRAM[27857] = 8'b0;
    XRAM[27858] = 8'b0;
    XRAM[27859] = 8'b0;
    XRAM[27860] = 8'b0;
    XRAM[27861] = 8'b0;
    XRAM[27862] = 8'b0;
    XRAM[27863] = 8'b0;
    XRAM[27864] = 8'b0;
    XRAM[27865] = 8'b0;
    XRAM[27866] = 8'b0;
    XRAM[27867] = 8'b0;
    XRAM[27868] = 8'b0;
    XRAM[27869] = 8'b0;
    XRAM[27870] = 8'b0;
    XRAM[27871] = 8'b0;
    XRAM[27872] = 8'b0;
    XRAM[27873] = 8'b0;
    XRAM[27874] = 8'b0;
    XRAM[27875] = 8'b0;
    XRAM[27876] = 8'b0;
    XRAM[27877] = 8'b0;
    XRAM[27878] = 8'b0;
    XRAM[27879] = 8'b0;
    XRAM[27880] = 8'b0;
    XRAM[27881] = 8'b0;
    XRAM[27882] = 8'b0;
    XRAM[27883] = 8'b0;
    XRAM[27884] = 8'b0;
    XRAM[27885] = 8'b0;
    XRAM[27886] = 8'b0;
    XRAM[27887] = 8'b0;
    XRAM[27888] = 8'b0;
    XRAM[27889] = 8'b0;
    XRAM[27890] = 8'b0;
    XRAM[27891] = 8'b0;
    XRAM[27892] = 8'b0;
    XRAM[27893] = 8'b0;
    XRAM[27894] = 8'b0;
    XRAM[27895] = 8'b0;
    XRAM[27896] = 8'b0;
    XRAM[27897] = 8'b0;
    XRAM[27898] = 8'b0;
    XRAM[27899] = 8'b0;
    XRAM[27900] = 8'b0;
    XRAM[27901] = 8'b0;
    XRAM[27902] = 8'b0;
    XRAM[27903] = 8'b0;
    XRAM[27904] = 8'b0;
    XRAM[27905] = 8'b0;
    XRAM[27906] = 8'b0;
    XRAM[27907] = 8'b0;
    XRAM[27908] = 8'b0;
    XRAM[27909] = 8'b0;
    XRAM[27910] = 8'b0;
    XRAM[27911] = 8'b0;
    XRAM[27912] = 8'b0;
    XRAM[27913] = 8'b0;
    XRAM[27914] = 8'b0;
    XRAM[27915] = 8'b0;
    XRAM[27916] = 8'b0;
    XRAM[27917] = 8'b0;
    XRAM[27918] = 8'b0;
    XRAM[27919] = 8'b0;
    XRAM[27920] = 8'b0;
    XRAM[27921] = 8'b0;
    XRAM[27922] = 8'b0;
    XRAM[27923] = 8'b0;
    XRAM[27924] = 8'b0;
    XRAM[27925] = 8'b0;
    XRAM[27926] = 8'b0;
    XRAM[27927] = 8'b0;
    XRAM[27928] = 8'b0;
    XRAM[27929] = 8'b0;
    XRAM[27930] = 8'b0;
    XRAM[27931] = 8'b0;
    XRAM[27932] = 8'b0;
    XRAM[27933] = 8'b0;
    XRAM[27934] = 8'b0;
    XRAM[27935] = 8'b0;
    XRAM[27936] = 8'b0;
    XRAM[27937] = 8'b0;
    XRAM[27938] = 8'b0;
    XRAM[27939] = 8'b0;
    XRAM[27940] = 8'b0;
    XRAM[27941] = 8'b0;
    XRAM[27942] = 8'b0;
    XRAM[27943] = 8'b0;
    XRAM[27944] = 8'b0;
    XRAM[27945] = 8'b0;
    XRAM[27946] = 8'b0;
    XRAM[27947] = 8'b0;
    XRAM[27948] = 8'b0;
    XRAM[27949] = 8'b0;
    XRAM[27950] = 8'b0;
    XRAM[27951] = 8'b0;
    XRAM[27952] = 8'b0;
    XRAM[27953] = 8'b0;
    XRAM[27954] = 8'b0;
    XRAM[27955] = 8'b0;
    XRAM[27956] = 8'b0;
    XRAM[27957] = 8'b0;
    XRAM[27958] = 8'b0;
    XRAM[27959] = 8'b0;
    XRAM[27960] = 8'b0;
    XRAM[27961] = 8'b0;
    XRAM[27962] = 8'b0;
    XRAM[27963] = 8'b0;
    XRAM[27964] = 8'b0;
    XRAM[27965] = 8'b0;
    XRAM[27966] = 8'b0;
    XRAM[27967] = 8'b0;
    XRAM[27968] = 8'b0;
    XRAM[27969] = 8'b0;
    XRAM[27970] = 8'b0;
    XRAM[27971] = 8'b0;
    XRAM[27972] = 8'b0;
    XRAM[27973] = 8'b0;
    XRAM[27974] = 8'b0;
    XRAM[27975] = 8'b0;
    XRAM[27976] = 8'b0;
    XRAM[27977] = 8'b0;
    XRAM[27978] = 8'b0;
    XRAM[27979] = 8'b0;
    XRAM[27980] = 8'b0;
    XRAM[27981] = 8'b0;
    XRAM[27982] = 8'b0;
    XRAM[27983] = 8'b0;
    XRAM[27984] = 8'b0;
    XRAM[27985] = 8'b0;
    XRAM[27986] = 8'b0;
    XRAM[27987] = 8'b0;
    XRAM[27988] = 8'b0;
    XRAM[27989] = 8'b0;
    XRAM[27990] = 8'b0;
    XRAM[27991] = 8'b0;
    XRAM[27992] = 8'b0;
    XRAM[27993] = 8'b0;
    XRAM[27994] = 8'b0;
    XRAM[27995] = 8'b0;
    XRAM[27996] = 8'b0;
    XRAM[27997] = 8'b0;
    XRAM[27998] = 8'b0;
    XRAM[27999] = 8'b0;
    XRAM[28000] = 8'b0;
    XRAM[28001] = 8'b0;
    XRAM[28002] = 8'b0;
    XRAM[28003] = 8'b0;
    XRAM[28004] = 8'b0;
    XRAM[28005] = 8'b0;
    XRAM[28006] = 8'b0;
    XRAM[28007] = 8'b0;
    XRAM[28008] = 8'b0;
    XRAM[28009] = 8'b0;
    XRAM[28010] = 8'b0;
    XRAM[28011] = 8'b0;
    XRAM[28012] = 8'b0;
    XRAM[28013] = 8'b0;
    XRAM[28014] = 8'b0;
    XRAM[28015] = 8'b0;
    XRAM[28016] = 8'b0;
    XRAM[28017] = 8'b0;
    XRAM[28018] = 8'b0;
    XRAM[28019] = 8'b0;
    XRAM[28020] = 8'b0;
    XRAM[28021] = 8'b0;
    XRAM[28022] = 8'b0;
    XRAM[28023] = 8'b0;
    XRAM[28024] = 8'b0;
    XRAM[28025] = 8'b0;
    XRAM[28026] = 8'b0;
    XRAM[28027] = 8'b0;
    XRAM[28028] = 8'b0;
    XRAM[28029] = 8'b0;
    XRAM[28030] = 8'b0;
    XRAM[28031] = 8'b0;
    XRAM[28032] = 8'b0;
    XRAM[28033] = 8'b0;
    XRAM[28034] = 8'b0;
    XRAM[28035] = 8'b0;
    XRAM[28036] = 8'b0;
    XRAM[28037] = 8'b0;
    XRAM[28038] = 8'b0;
    XRAM[28039] = 8'b0;
    XRAM[28040] = 8'b0;
    XRAM[28041] = 8'b0;
    XRAM[28042] = 8'b0;
    XRAM[28043] = 8'b0;
    XRAM[28044] = 8'b0;
    XRAM[28045] = 8'b0;
    XRAM[28046] = 8'b0;
    XRAM[28047] = 8'b0;
    XRAM[28048] = 8'b0;
    XRAM[28049] = 8'b0;
    XRAM[28050] = 8'b0;
    XRAM[28051] = 8'b0;
    XRAM[28052] = 8'b0;
    XRAM[28053] = 8'b0;
    XRAM[28054] = 8'b0;
    XRAM[28055] = 8'b0;
    XRAM[28056] = 8'b0;
    XRAM[28057] = 8'b0;
    XRAM[28058] = 8'b0;
    XRAM[28059] = 8'b0;
    XRAM[28060] = 8'b0;
    XRAM[28061] = 8'b0;
    XRAM[28062] = 8'b0;
    XRAM[28063] = 8'b0;
    XRAM[28064] = 8'b0;
    XRAM[28065] = 8'b0;
    XRAM[28066] = 8'b0;
    XRAM[28067] = 8'b0;
    XRAM[28068] = 8'b0;
    XRAM[28069] = 8'b0;
    XRAM[28070] = 8'b0;
    XRAM[28071] = 8'b0;
    XRAM[28072] = 8'b0;
    XRAM[28073] = 8'b0;
    XRAM[28074] = 8'b0;
    XRAM[28075] = 8'b0;
    XRAM[28076] = 8'b0;
    XRAM[28077] = 8'b0;
    XRAM[28078] = 8'b0;
    XRAM[28079] = 8'b0;
    XRAM[28080] = 8'b0;
    XRAM[28081] = 8'b0;
    XRAM[28082] = 8'b0;
    XRAM[28083] = 8'b0;
    XRAM[28084] = 8'b0;
    XRAM[28085] = 8'b0;
    XRAM[28086] = 8'b0;
    XRAM[28087] = 8'b0;
    XRAM[28088] = 8'b0;
    XRAM[28089] = 8'b0;
    XRAM[28090] = 8'b0;
    XRAM[28091] = 8'b0;
    XRAM[28092] = 8'b0;
    XRAM[28093] = 8'b0;
    XRAM[28094] = 8'b0;
    XRAM[28095] = 8'b0;
    XRAM[28096] = 8'b0;
    XRAM[28097] = 8'b0;
    XRAM[28098] = 8'b0;
    XRAM[28099] = 8'b0;
    XRAM[28100] = 8'b0;
    XRAM[28101] = 8'b0;
    XRAM[28102] = 8'b0;
    XRAM[28103] = 8'b0;
    XRAM[28104] = 8'b0;
    XRAM[28105] = 8'b0;
    XRAM[28106] = 8'b0;
    XRAM[28107] = 8'b0;
    XRAM[28108] = 8'b0;
    XRAM[28109] = 8'b0;
    XRAM[28110] = 8'b0;
    XRAM[28111] = 8'b0;
    XRAM[28112] = 8'b0;
    XRAM[28113] = 8'b0;
    XRAM[28114] = 8'b0;
    XRAM[28115] = 8'b0;
    XRAM[28116] = 8'b0;
    XRAM[28117] = 8'b0;
    XRAM[28118] = 8'b0;
    XRAM[28119] = 8'b0;
    XRAM[28120] = 8'b0;
    XRAM[28121] = 8'b0;
    XRAM[28122] = 8'b0;
    XRAM[28123] = 8'b0;
    XRAM[28124] = 8'b0;
    XRAM[28125] = 8'b0;
    XRAM[28126] = 8'b0;
    XRAM[28127] = 8'b0;
    XRAM[28128] = 8'b0;
    XRAM[28129] = 8'b0;
    XRAM[28130] = 8'b0;
    XRAM[28131] = 8'b0;
    XRAM[28132] = 8'b0;
    XRAM[28133] = 8'b0;
    XRAM[28134] = 8'b0;
    XRAM[28135] = 8'b0;
    XRAM[28136] = 8'b0;
    XRAM[28137] = 8'b0;
    XRAM[28138] = 8'b0;
    XRAM[28139] = 8'b0;
    XRAM[28140] = 8'b0;
    XRAM[28141] = 8'b0;
    XRAM[28142] = 8'b0;
    XRAM[28143] = 8'b0;
    XRAM[28144] = 8'b0;
    XRAM[28145] = 8'b0;
    XRAM[28146] = 8'b0;
    XRAM[28147] = 8'b0;
    XRAM[28148] = 8'b0;
    XRAM[28149] = 8'b0;
    XRAM[28150] = 8'b0;
    XRAM[28151] = 8'b0;
    XRAM[28152] = 8'b0;
    XRAM[28153] = 8'b0;
    XRAM[28154] = 8'b0;
    XRAM[28155] = 8'b0;
    XRAM[28156] = 8'b0;
    XRAM[28157] = 8'b0;
    XRAM[28158] = 8'b0;
    XRAM[28159] = 8'b0;
    XRAM[28160] = 8'b0;
    XRAM[28161] = 8'b0;
    XRAM[28162] = 8'b0;
    XRAM[28163] = 8'b0;
    XRAM[28164] = 8'b0;
    XRAM[28165] = 8'b0;
    XRAM[28166] = 8'b0;
    XRAM[28167] = 8'b0;
    XRAM[28168] = 8'b0;
    XRAM[28169] = 8'b0;
    XRAM[28170] = 8'b0;
    XRAM[28171] = 8'b0;
    XRAM[28172] = 8'b0;
    XRAM[28173] = 8'b0;
    XRAM[28174] = 8'b0;
    XRAM[28175] = 8'b0;
    XRAM[28176] = 8'b0;
    XRAM[28177] = 8'b0;
    XRAM[28178] = 8'b0;
    XRAM[28179] = 8'b0;
    XRAM[28180] = 8'b0;
    XRAM[28181] = 8'b0;
    XRAM[28182] = 8'b0;
    XRAM[28183] = 8'b0;
    XRAM[28184] = 8'b0;
    XRAM[28185] = 8'b0;
    XRAM[28186] = 8'b0;
    XRAM[28187] = 8'b0;
    XRAM[28188] = 8'b0;
    XRAM[28189] = 8'b0;
    XRAM[28190] = 8'b0;
    XRAM[28191] = 8'b0;
    XRAM[28192] = 8'b0;
    XRAM[28193] = 8'b0;
    XRAM[28194] = 8'b0;
    XRAM[28195] = 8'b0;
    XRAM[28196] = 8'b0;
    XRAM[28197] = 8'b0;
    XRAM[28198] = 8'b0;
    XRAM[28199] = 8'b0;
    XRAM[28200] = 8'b0;
    XRAM[28201] = 8'b0;
    XRAM[28202] = 8'b0;
    XRAM[28203] = 8'b0;
    XRAM[28204] = 8'b0;
    XRAM[28205] = 8'b0;
    XRAM[28206] = 8'b0;
    XRAM[28207] = 8'b0;
    XRAM[28208] = 8'b0;
    XRAM[28209] = 8'b0;
    XRAM[28210] = 8'b0;
    XRAM[28211] = 8'b0;
    XRAM[28212] = 8'b0;
    XRAM[28213] = 8'b0;
    XRAM[28214] = 8'b0;
    XRAM[28215] = 8'b0;
    XRAM[28216] = 8'b0;
    XRAM[28217] = 8'b0;
    XRAM[28218] = 8'b0;
    XRAM[28219] = 8'b0;
    XRAM[28220] = 8'b0;
    XRAM[28221] = 8'b0;
    XRAM[28222] = 8'b0;
    XRAM[28223] = 8'b0;
    XRAM[28224] = 8'b0;
    XRAM[28225] = 8'b0;
    XRAM[28226] = 8'b0;
    XRAM[28227] = 8'b0;
    XRAM[28228] = 8'b0;
    XRAM[28229] = 8'b0;
    XRAM[28230] = 8'b0;
    XRAM[28231] = 8'b0;
    XRAM[28232] = 8'b0;
    XRAM[28233] = 8'b0;
    XRAM[28234] = 8'b0;
    XRAM[28235] = 8'b0;
    XRAM[28236] = 8'b0;
    XRAM[28237] = 8'b0;
    XRAM[28238] = 8'b0;
    XRAM[28239] = 8'b0;
    XRAM[28240] = 8'b0;
    XRAM[28241] = 8'b0;
    XRAM[28242] = 8'b0;
    XRAM[28243] = 8'b0;
    XRAM[28244] = 8'b0;
    XRAM[28245] = 8'b0;
    XRAM[28246] = 8'b0;
    XRAM[28247] = 8'b0;
    XRAM[28248] = 8'b0;
    XRAM[28249] = 8'b0;
    XRAM[28250] = 8'b0;
    XRAM[28251] = 8'b0;
    XRAM[28252] = 8'b0;
    XRAM[28253] = 8'b0;
    XRAM[28254] = 8'b0;
    XRAM[28255] = 8'b0;
    XRAM[28256] = 8'b0;
    XRAM[28257] = 8'b0;
    XRAM[28258] = 8'b0;
    XRAM[28259] = 8'b0;
    XRAM[28260] = 8'b0;
    XRAM[28261] = 8'b0;
    XRAM[28262] = 8'b0;
    XRAM[28263] = 8'b0;
    XRAM[28264] = 8'b0;
    XRAM[28265] = 8'b0;
    XRAM[28266] = 8'b0;
    XRAM[28267] = 8'b0;
    XRAM[28268] = 8'b0;
    XRAM[28269] = 8'b0;
    XRAM[28270] = 8'b0;
    XRAM[28271] = 8'b0;
    XRAM[28272] = 8'b0;
    XRAM[28273] = 8'b0;
    XRAM[28274] = 8'b0;
    XRAM[28275] = 8'b0;
    XRAM[28276] = 8'b0;
    XRAM[28277] = 8'b0;
    XRAM[28278] = 8'b0;
    XRAM[28279] = 8'b0;
    XRAM[28280] = 8'b0;
    XRAM[28281] = 8'b0;
    XRAM[28282] = 8'b0;
    XRAM[28283] = 8'b0;
    XRAM[28284] = 8'b0;
    XRAM[28285] = 8'b0;
    XRAM[28286] = 8'b0;
    XRAM[28287] = 8'b0;
    XRAM[28288] = 8'b0;
    XRAM[28289] = 8'b0;
    XRAM[28290] = 8'b0;
    XRAM[28291] = 8'b0;
    XRAM[28292] = 8'b0;
    XRAM[28293] = 8'b0;
    XRAM[28294] = 8'b0;
    XRAM[28295] = 8'b0;
    XRAM[28296] = 8'b0;
    XRAM[28297] = 8'b0;
    XRAM[28298] = 8'b0;
    XRAM[28299] = 8'b0;
    XRAM[28300] = 8'b0;
    XRAM[28301] = 8'b0;
    XRAM[28302] = 8'b0;
    XRAM[28303] = 8'b0;
    XRAM[28304] = 8'b0;
    XRAM[28305] = 8'b0;
    XRAM[28306] = 8'b0;
    XRAM[28307] = 8'b0;
    XRAM[28308] = 8'b0;
    XRAM[28309] = 8'b0;
    XRAM[28310] = 8'b0;
    XRAM[28311] = 8'b0;
    XRAM[28312] = 8'b0;
    XRAM[28313] = 8'b0;
    XRAM[28314] = 8'b0;
    XRAM[28315] = 8'b0;
    XRAM[28316] = 8'b0;
    XRAM[28317] = 8'b0;
    XRAM[28318] = 8'b0;
    XRAM[28319] = 8'b0;
    XRAM[28320] = 8'b0;
    XRAM[28321] = 8'b0;
    XRAM[28322] = 8'b0;
    XRAM[28323] = 8'b0;
    XRAM[28324] = 8'b0;
    XRAM[28325] = 8'b0;
    XRAM[28326] = 8'b0;
    XRAM[28327] = 8'b0;
    XRAM[28328] = 8'b0;
    XRAM[28329] = 8'b0;
    XRAM[28330] = 8'b0;
    XRAM[28331] = 8'b0;
    XRAM[28332] = 8'b0;
    XRAM[28333] = 8'b0;
    XRAM[28334] = 8'b0;
    XRAM[28335] = 8'b0;
    XRAM[28336] = 8'b0;
    XRAM[28337] = 8'b0;
    XRAM[28338] = 8'b0;
    XRAM[28339] = 8'b0;
    XRAM[28340] = 8'b0;
    XRAM[28341] = 8'b0;
    XRAM[28342] = 8'b0;
    XRAM[28343] = 8'b0;
    XRAM[28344] = 8'b0;
    XRAM[28345] = 8'b0;
    XRAM[28346] = 8'b0;
    XRAM[28347] = 8'b0;
    XRAM[28348] = 8'b0;
    XRAM[28349] = 8'b0;
    XRAM[28350] = 8'b0;
    XRAM[28351] = 8'b0;
    XRAM[28352] = 8'b0;
    XRAM[28353] = 8'b0;
    XRAM[28354] = 8'b0;
    XRAM[28355] = 8'b0;
    XRAM[28356] = 8'b0;
    XRAM[28357] = 8'b0;
    XRAM[28358] = 8'b0;
    XRAM[28359] = 8'b0;
    XRAM[28360] = 8'b0;
    XRAM[28361] = 8'b0;
    XRAM[28362] = 8'b0;
    XRAM[28363] = 8'b0;
    XRAM[28364] = 8'b0;
    XRAM[28365] = 8'b0;
    XRAM[28366] = 8'b0;
    XRAM[28367] = 8'b0;
    XRAM[28368] = 8'b0;
    XRAM[28369] = 8'b0;
    XRAM[28370] = 8'b0;
    XRAM[28371] = 8'b0;
    XRAM[28372] = 8'b0;
    XRAM[28373] = 8'b0;
    XRAM[28374] = 8'b0;
    XRAM[28375] = 8'b0;
    XRAM[28376] = 8'b0;
    XRAM[28377] = 8'b0;
    XRAM[28378] = 8'b0;
    XRAM[28379] = 8'b0;
    XRAM[28380] = 8'b0;
    XRAM[28381] = 8'b0;
    XRAM[28382] = 8'b0;
    XRAM[28383] = 8'b0;
    XRAM[28384] = 8'b0;
    XRAM[28385] = 8'b0;
    XRAM[28386] = 8'b0;
    XRAM[28387] = 8'b0;
    XRAM[28388] = 8'b0;
    XRAM[28389] = 8'b0;
    XRAM[28390] = 8'b0;
    XRAM[28391] = 8'b0;
    XRAM[28392] = 8'b0;
    XRAM[28393] = 8'b0;
    XRAM[28394] = 8'b0;
    XRAM[28395] = 8'b0;
    XRAM[28396] = 8'b0;
    XRAM[28397] = 8'b0;
    XRAM[28398] = 8'b0;
    XRAM[28399] = 8'b0;
    XRAM[28400] = 8'b0;
    XRAM[28401] = 8'b0;
    XRAM[28402] = 8'b0;
    XRAM[28403] = 8'b0;
    XRAM[28404] = 8'b0;
    XRAM[28405] = 8'b0;
    XRAM[28406] = 8'b0;
    XRAM[28407] = 8'b0;
    XRAM[28408] = 8'b0;
    XRAM[28409] = 8'b0;
    XRAM[28410] = 8'b0;
    XRAM[28411] = 8'b0;
    XRAM[28412] = 8'b0;
    XRAM[28413] = 8'b0;
    XRAM[28414] = 8'b0;
    XRAM[28415] = 8'b0;
    XRAM[28416] = 8'b0;
    XRAM[28417] = 8'b0;
    XRAM[28418] = 8'b0;
    XRAM[28419] = 8'b0;
    XRAM[28420] = 8'b0;
    XRAM[28421] = 8'b0;
    XRAM[28422] = 8'b0;
    XRAM[28423] = 8'b0;
    XRAM[28424] = 8'b0;
    XRAM[28425] = 8'b0;
    XRAM[28426] = 8'b0;
    XRAM[28427] = 8'b0;
    XRAM[28428] = 8'b0;
    XRAM[28429] = 8'b0;
    XRAM[28430] = 8'b0;
    XRAM[28431] = 8'b0;
    XRAM[28432] = 8'b0;
    XRAM[28433] = 8'b0;
    XRAM[28434] = 8'b0;
    XRAM[28435] = 8'b0;
    XRAM[28436] = 8'b0;
    XRAM[28437] = 8'b0;
    XRAM[28438] = 8'b0;
    XRAM[28439] = 8'b0;
    XRAM[28440] = 8'b0;
    XRAM[28441] = 8'b0;
    XRAM[28442] = 8'b0;
    XRAM[28443] = 8'b0;
    XRAM[28444] = 8'b0;
    XRAM[28445] = 8'b0;
    XRAM[28446] = 8'b0;
    XRAM[28447] = 8'b0;
    XRAM[28448] = 8'b0;
    XRAM[28449] = 8'b0;
    XRAM[28450] = 8'b0;
    XRAM[28451] = 8'b0;
    XRAM[28452] = 8'b0;
    XRAM[28453] = 8'b0;
    XRAM[28454] = 8'b0;
    XRAM[28455] = 8'b0;
    XRAM[28456] = 8'b0;
    XRAM[28457] = 8'b0;
    XRAM[28458] = 8'b0;
    XRAM[28459] = 8'b0;
    XRAM[28460] = 8'b0;
    XRAM[28461] = 8'b0;
    XRAM[28462] = 8'b0;
    XRAM[28463] = 8'b0;
    XRAM[28464] = 8'b0;
    XRAM[28465] = 8'b0;
    XRAM[28466] = 8'b0;
    XRAM[28467] = 8'b0;
    XRAM[28468] = 8'b0;
    XRAM[28469] = 8'b0;
    XRAM[28470] = 8'b0;
    XRAM[28471] = 8'b0;
    XRAM[28472] = 8'b0;
    XRAM[28473] = 8'b0;
    XRAM[28474] = 8'b0;
    XRAM[28475] = 8'b0;
    XRAM[28476] = 8'b0;
    XRAM[28477] = 8'b0;
    XRAM[28478] = 8'b0;
    XRAM[28479] = 8'b0;
    XRAM[28480] = 8'b0;
    XRAM[28481] = 8'b0;
    XRAM[28482] = 8'b0;
    XRAM[28483] = 8'b0;
    XRAM[28484] = 8'b0;
    XRAM[28485] = 8'b0;
    XRAM[28486] = 8'b0;
    XRAM[28487] = 8'b0;
    XRAM[28488] = 8'b0;
    XRAM[28489] = 8'b0;
    XRAM[28490] = 8'b0;
    XRAM[28491] = 8'b0;
    XRAM[28492] = 8'b0;
    XRAM[28493] = 8'b0;
    XRAM[28494] = 8'b0;
    XRAM[28495] = 8'b0;
    XRAM[28496] = 8'b0;
    XRAM[28497] = 8'b0;
    XRAM[28498] = 8'b0;
    XRAM[28499] = 8'b0;
    XRAM[28500] = 8'b0;
    XRAM[28501] = 8'b0;
    XRAM[28502] = 8'b0;
    XRAM[28503] = 8'b0;
    XRAM[28504] = 8'b0;
    XRAM[28505] = 8'b0;
    XRAM[28506] = 8'b0;
    XRAM[28507] = 8'b0;
    XRAM[28508] = 8'b0;
    XRAM[28509] = 8'b0;
    XRAM[28510] = 8'b0;
    XRAM[28511] = 8'b0;
    XRAM[28512] = 8'b0;
    XRAM[28513] = 8'b0;
    XRAM[28514] = 8'b0;
    XRAM[28515] = 8'b0;
    XRAM[28516] = 8'b0;
    XRAM[28517] = 8'b0;
    XRAM[28518] = 8'b0;
    XRAM[28519] = 8'b0;
    XRAM[28520] = 8'b0;
    XRAM[28521] = 8'b0;
    XRAM[28522] = 8'b0;
    XRAM[28523] = 8'b0;
    XRAM[28524] = 8'b0;
    XRAM[28525] = 8'b0;
    XRAM[28526] = 8'b0;
    XRAM[28527] = 8'b0;
    XRAM[28528] = 8'b0;
    XRAM[28529] = 8'b0;
    XRAM[28530] = 8'b0;
    XRAM[28531] = 8'b0;
    XRAM[28532] = 8'b0;
    XRAM[28533] = 8'b0;
    XRAM[28534] = 8'b0;
    XRAM[28535] = 8'b0;
    XRAM[28536] = 8'b0;
    XRAM[28537] = 8'b0;
    XRAM[28538] = 8'b0;
    XRAM[28539] = 8'b0;
    XRAM[28540] = 8'b0;
    XRAM[28541] = 8'b0;
    XRAM[28542] = 8'b0;
    XRAM[28543] = 8'b0;
    XRAM[28544] = 8'b0;
    XRAM[28545] = 8'b0;
    XRAM[28546] = 8'b0;
    XRAM[28547] = 8'b0;
    XRAM[28548] = 8'b0;
    XRAM[28549] = 8'b0;
    XRAM[28550] = 8'b0;
    XRAM[28551] = 8'b0;
    XRAM[28552] = 8'b0;
    XRAM[28553] = 8'b0;
    XRAM[28554] = 8'b0;
    XRAM[28555] = 8'b0;
    XRAM[28556] = 8'b0;
    XRAM[28557] = 8'b0;
    XRAM[28558] = 8'b0;
    XRAM[28559] = 8'b0;
    XRAM[28560] = 8'b0;
    XRAM[28561] = 8'b0;
    XRAM[28562] = 8'b0;
    XRAM[28563] = 8'b0;
    XRAM[28564] = 8'b0;
    XRAM[28565] = 8'b0;
    XRAM[28566] = 8'b0;
    XRAM[28567] = 8'b0;
    XRAM[28568] = 8'b0;
    XRAM[28569] = 8'b0;
    XRAM[28570] = 8'b0;
    XRAM[28571] = 8'b0;
    XRAM[28572] = 8'b0;
    XRAM[28573] = 8'b0;
    XRAM[28574] = 8'b0;
    XRAM[28575] = 8'b0;
    XRAM[28576] = 8'b0;
    XRAM[28577] = 8'b0;
    XRAM[28578] = 8'b0;
    XRAM[28579] = 8'b0;
    XRAM[28580] = 8'b0;
    XRAM[28581] = 8'b0;
    XRAM[28582] = 8'b0;
    XRAM[28583] = 8'b0;
    XRAM[28584] = 8'b0;
    XRAM[28585] = 8'b0;
    XRAM[28586] = 8'b0;
    XRAM[28587] = 8'b0;
    XRAM[28588] = 8'b0;
    XRAM[28589] = 8'b0;
    XRAM[28590] = 8'b0;
    XRAM[28591] = 8'b0;
    XRAM[28592] = 8'b0;
    XRAM[28593] = 8'b0;
    XRAM[28594] = 8'b0;
    XRAM[28595] = 8'b0;
    XRAM[28596] = 8'b0;
    XRAM[28597] = 8'b0;
    XRAM[28598] = 8'b0;
    XRAM[28599] = 8'b0;
    XRAM[28600] = 8'b0;
    XRAM[28601] = 8'b0;
    XRAM[28602] = 8'b0;
    XRAM[28603] = 8'b0;
    XRAM[28604] = 8'b0;
    XRAM[28605] = 8'b0;
    XRAM[28606] = 8'b0;
    XRAM[28607] = 8'b0;
    XRAM[28608] = 8'b0;
    XRAM[28609] = 8'b0;
    XRAM[28610] = 8'b0;
    XRAM[28611] = 8'b0;
    XRAM[28612] = 8'b0;
    XRAM[28613] = 8'b0;
    XRAM[28614] = 8'b0;
    XRAM[28615] = 8'b0;
    XRAM[28616] = 8'b0;
    XRAM[28617] = 8'b0;
    XRAM[28618] = 8'b0;
    XRAM[28619] = 8'b0;
    XRAM[28620] = 8'b0;
    XRAM[28621] = 8'b0;
    XRAM[28622] = 8'b0;
    XRAM[28623] = 8'b0;
    XRAM[28624] = 8'b0;
    XRAM[28625] = 8'b0;
    XRAM[28626] = 8'b0;
    XRAM[28627] = 8'b0;
    XRAM[28628] = 8'b0;
    XRAM[28629] = 8'b0;
    XRAM[28630] = 8'b0;
    XRAM[28631] = 8'b0;
    XRAM[28632] = 8'b0;
    XRAM[28633] = 8'b0;
    XRAM[28634] = 8'b0;
    XRAM[28635] = 8'b0;
    XRAM[28636] = 8'b0;
    XRAM[28637] = 8'b0;
    XRAM[28638] = 8'b0;
    XRAM[28639] = 8'b0;
    XRAM[28640] = 8'b0;
    XRAM[28641] = 8'b0;
    XRAM[28642] = 8'b0;
    XRAM[28643] = 8'b0;
    XRAM[28644] = 8'b0;
    XRAM[28645] = 8'b0;
    XRAM[28646] = 8'b0;
    XRAM[28647] = 8'b0;
    XRAM[28648] = 8'b0;
    XRAM[28649] = 8'b0;
    XRAM[28650] = 8'b0;
    XRAM[28651] = 8'b0;
    XRAM[28652] = 8'b0;
    XRAM[28653] = 8'b0;
    XRAM[28654] = 8'b0;
    XRAM[28655] = 8'b0;
    XRAM[28656] = 8'b0;
    XRAM[28657] = 8'b0;
    XRAM[28658] = 8'b0;
    XRAM[28659] = 8'b0;
    XRAM[28660] = 8'b0;
    XRAM[28661] = 8'b0;
    XRAM[28662] = 8'b0;
    XRAM[28663] = 8'b0;
    XRAM[28664] = 8'b0;
    XRAM[28665] = 8'b0;
    XRAM[28666] = 8'b0;
    XRAM[28667] = 8'b0;
    XRAM[28668] = 8'b0;
    XRAM[28669] = 8'b0;
    XRAM[28670] = 8'b0;
    XRAM[28671] = 8'b0;
    XRAM[28672] = 8'b0;
    XRAM[28673] = 8'b0;
    XRAM[28674] = 8'b0;
    XRAM[28675] = 8'b0;
    XRAM[28676] = 8'b0;
    XRAM[28677] = 8'b0;
    XRAM[28678] = 8'b0;
    XRAM[28679] = 8'b0;
    XRAM[28680] = 8'b0;
    XRAM[28681] = 8'b0;
    XRAM[28682] = 8'b0;
    XRAM[28683] = 8'b0;
    XRAM[28684] = 8'b0;
    XRAM[28685] = 8'b0;
    XRAM[28686] = 8'b0;
    XRAM[28687] = 8'b0;
    XRAM[28688] = 8'b0;
    XRAM[28689] = 8'b0;
    XRAM[28690] = 8'b0;
    XRAM[28691] = 8'b0;
    XRAM[28692] = 8'b0;
    XRAM[28693] = 8'b0;
    XRAM[28694] = 8'b0;
    XRAM[28695] = 8'b0;
    XRAM[28696] = 8'b0;
    XRAM[28697] = 8'b0;
    XRAM[28698] = 8'b0;
    XRAM[28699] = 8'b0;
    XRAM[28700] = 8'b0;
    XRAM[28701] = 8'b0;
    XRAM[28702] = 8'b0;
    XRAM[28703] = 8'b0;
    XRAM[28704] = 8'b0;
    XRAM[28705] = 8'b0;
    XRAM[28706] = 8'b0;
    XRAM[28707] = 8'b0;
    XRAM[28708] = 8'b0;
    XRAM[28709] = 8'b0;
    XRAM[28710] = 8'b0;
    XRAM[28711] = 8'b0;
    XRAM[28712] = 8'b0;
    XRAM[28713] = 8'b0;
    XRAM[28714] = 8'b0;
    XRAM[28715] = 8'b0;
    XRAM[28716] = 8'b0;
    XRAM[28717] = 8'b0;
    XRAM[28718] = 8'b0;
    XRAM[28719] = 8'b0;
    XRAM[28720] = 8'b0;
    XRAM[28721] = 8'b0;
    XRAM[28722] = 8'b0;
    XRAM[28723] = 8'b0;
    XRAM[28724] = 8'b0;
    XRAM[28725] = 8'b0;
    XRAM[28726] = 8'b0;
    XRAM[28727] = 8'b0;
    XRAM[28728] = 8'b0;
    XRAM[28729] = 8'b0;
    XRAM[28730] = 8'b0;
    XRAM[28731] = 8'b0;
    XRAM[28732] = 8'b0;
    XRAM[28733] = 8'b0;
    XRAM[28734] = 8'b0;
    XRAM[28735] = 8'b0;
    XRAM[28736] = 8'b0;
    XRAM[28737] = 8'b0;
    XRAM[28738] = 8'b0;
    XRAM[28739] = 8'b0;
    XRAM[28740] = 8'b0;
    XRAM[28741] = 8'b0;
    XRAM[28742] = 8'b0;
    XRAM[28743] = 8'b0;
    XRAM[28744] = 8'b0;
    XRAM[28745] = 8'b0;
    XRAM[28746] = 8'b0;
    XRAM[28747] = 8'b0;
    XRAM[28748] = 8'b0;
    XRAM[28749] = 8'b0;
    XRAM[28750] = 8'b0;
    XRAM[28751] = 8'b0;
    XRAM[28752] = 8'b0;
    XRAM[28753] = 8'b0;
    XRAM[28754] = 8'b0;
    XRAM[28755] = 8'b0;
    XRAM[28756] = 8'b0;
    XRAM[28757] = 8'b0;
    XRAM[28758] = 8'b0;
    XRAM[28759] = 8'b0;
    XRAM[28760] = 8'b0;
    XRAM[28761] = 8'b0;
    XRAM[28762] = 8'b0;
    XRAM[28763] = 8'b0;
    XRAM[28764] = 8'b0;
    XRAM[28765] = 8'b0;
    XRAM[28766] = 8'b0;
    XRAM[28767] = 8'b0;
    XRAM[28768] = 8'b0;
    XRAM[28769] = 8'b0;
    XRAM[28770] = 8'b0;
    XRAM[28771] = 8'b0;
    XRAM[28772] = 8'b0;
    XRAM[28773] = 8'b0;
    XRAM[28774] = 8'b0;
    XRAM[28775] = 8'b0;
    XRAM[28776] = 8'b0;
    XRAM[28777] = 8'b0;
    XRAM[28778] = 8'b0;
    XRAM[28779] = 8'b0;
    XRAM[28780] = 8'b0;
    XRAM[28781] = 8'b0;
    XRAM[28782] = 8'b0;
    XRAM[28783] = 8'b0;
    XRAM[28784] = 8'b0;
    XRAM[28785] = 8'b0;
    XRAM[28786] = 8'b0;
    XRAM[28787] = 8'b0;
    XRAM[28788] = 8'b0;
    XRAM[28789] = 8'b0;
    XRAM[28790] = 8'b0;
    XRAM[28791] = 8'b0;
    XRAM[28792] = 8'b0;
    XRAM[28793] = 8'b0;
    XRAM[28794] = 8'b0;
    XRAM[28795] = 8'b0;
    XRAM[28796] = 8'b0;
    XRAM[28797] = 8'b0;
    XRAM[28798] = 8'b0;
    XRAM[28799] = 8'b0;
    XRAM[28800] = 8'b0;
    XRAM[28801] = 8'b0;
    XRAM[28802] = 8'b0;
    XRAM[28803] = 8'b0;
    XRAM[28804] = 8'b0;
    XRAM[28805] = 8'b0;
    XRAM[28806] = 8'b0;
    XRAM[28807] = 8'b0;
    XRAM[28808] = 8'b0;
    XRAM[28809] = 8'b0;
    XRAM[28810] = 8'b0;
    XRAM[28811] = 8'b0;
    XRAM[28812] = 8'b0;
    XRAM[28813] = 8'b0;
    XRAM[28814] = 8'b0;
    XRAM[28815] = 8'b0;
    XRAM[28816] = 8'b0;
    XRAM[28817] = 8'b0;
    XRAM[28818] = 8'b0;
    XRAM[28819] = 8'b0;
    XRAM[28820] = 8'b0;
    XRAM[28821] = 8'b0;
    XRAM[28822] = 8'b0;
    XRAM[28823] = 8'b0;
    XRAM[28824] = 8'b0;
    XRAM[28825] = 8'b0;
    XRAM[28826] = 8'b0;
    XRAM[28827] = 8'b0;
    XRAM[28828] = 8'b0;
    XRAM[28829] = 8'b0;
    XRAM[28830] = 8'b0;
    XRAM[28831] = 8'b0;
    XRAM[28832] = 8'b0;
    XRAM[28833] = 8'b0;
    XRAM[28834] = 8'b0;
    XRAM[28835] = 8'b0;
    XRAM[28836] = 8'b0;
    XRAM[28837] = 8'b0;
    XRAM[28838] = 8'b0;
    XRAM[28839] = 8'b0;
    XRAM[28840] = 8'b0;
    XRAM[28841] = 8'b0;
    XRAM[28842] = 8'b0;
    XRAM[28843] = 8'b0;
    XRAM[28844] = 8'b0;
    XRAM[28845] = 8'b0;
    XRAM[28846] = 8'b0;
    XRAM[28847] = 8'b0;
    XRAM[28848] = 8'b0;
    XRAM[28849] = 8'b0;
    XRAM[28850] = 8'b0;
    XRAM[28851] = 8'b0;
    XRAM[28852] = 8'b0;
    XRAM[28853] = 8'b0;
    XRAM[28854] = 8'b0;
    XRAM[28855] = 8'b0;
    XRAM[28856] = 8'b0;
    XRAM[28857] = 8'b0;
    XRAM[28858] = 8'b0;
    XRAM[28859] = 8'b0;
    XRAM[28860] = 8'b0;
    XRAM[28861] = 8'b0;
    XRAM[28862] = 8'b0;
    XRAM[28863] = 8'b0;
    XRAM[28864] = 8'b0;
    XRAM[28865] = 8'b0;
    XRAM[28866] = 8'b0;
    XRAM[28867] = 8'b0;
    XRAM[28868] = 8'b0;
    XRAM[28869] = 8'b0;
    XRAM[28870] = 8'b0;
    XRAM[28871] = 8'b0;
    XRAM[28872] = 8'b0;
    XRAM[28873] = 8'b0;
    XRAM[28874] = 8'b0;
    XRAM[28875] = 8'b0;
    XRAM[28876] = 8'b0;
    XRAM[28877] = 8'b0;
    XRAM[28878] = 8'b0;
    XRAM[28879] = 8'b0;
    XRAM[28880] = 8'b0;
    XRAM[28881] = 8'b0;
    XRAM[28882] = 8'b0;
    XRAM[28883] = 8'b0;
    XRAM[28884] = 8'b0;
    XRAM[28885] = 8'b0;
    XRAM[28886] = 8'b0;
    XRAM[28887] = 8'b0;
    XRAM[28888] = 8'b0;
    XRAM[28889] = 8'b0;
    XRAM[28890] = 8'b0;
    XRAM[28891] = 8'b0;
    XRAM[28892] = 8'b0;
    XRAM[28893] = 8'b0;
    XRAM[28894] = 8'b0;
    XRAM[28895] = 8'b0;
    XRAM[28896] = 8'b0;
    XRAM[28897] = 8'b0;
    XRAM[28898] = 8'b0;
    XRAM[28899] = 8'b0;
    XRAM[28900] = 8'b0;
    XRAM[28901] = 8'b0;
    XRAM[28902] = 8'b0;
    XRAM[28903] = 8'b0;
    XRAM[28904] = 8'b0;
    XRAM[28905] = 8'b0;
    XRAM[28906] = 8'b0;
    XRAM[28907] = 8'b0;
    XRAM[28908] = 8'b0;
    XRAM[28909] = 8'b0;
    XRAM[28910] = 8'b0;
    XRAM[28911] = 8'b0;
    XRAM[28912] = 8'b0;
    XRAM[28913] = 8'b0;
    XRAM[28914] = 8'b0;
    XRAM[28915] = 8'b0;
    XRAM[28916] = 8'b0;
    XRAM[28917] = 8'b0;
    XRAM[28918] = 8'b0;
    XRAM[28919] = 8'b0;
    XRAM[28920] = 8'b0;
    XRAM[28921] = 8'b0;
    XRAM[28922] = 8'b0;
    XRAM[28923] = 8'b0;
    XRAM[28924] = 8'b0;
    XRAM[28925] = 8'b0;
    XRAM[28926] = 8'b0;
    XRAM[28927] = 8'b0;
    XRAM[28928] = 8'b0;
    XRAM[28929] = 8'b0;
    XRAM[28930] = 8'b0;
    XRAM[28931] = 8'b0;
    XRAM[28932] = 8'b0;
    XRAM[28933] = 8'b0;
    XRAM[28934] = 8'b0;
    XRAM[28935] = 8'b0;
    XRAM[28936] = 8'b0;
    XRAM[28937] = 8'b0;
    XRAM[28938] = 8'b0;
    XRAM[28939] = 8'b0;
    XRAM[28940] = 8'b0;
    XRAM[28941] = 8'b0;
    XRAM[28942] = 8'b0;
    XRAM[28943] = 8'b0;
    XRAM[28944] = 8'b0;
    XRAM[28945] = 8'b0;
    XRAM[28946] = 8'b0;
    XRAM[28947] = 8'b0;
    XRAM[28948] = 8'b0;
    XRAM[28949] = 8'b0;
    XRAM[28950] = 8'b0;
    XRAM[28951] = 8'b0;
    XRAM[28952] = 8'b0;
    XRAM[28953] = 8'b0;
    XRAM[28954] = 8'b0;
    XRAM[28955] = 8'b0;
    XRAM[28956] = 8'b0;
    XRAM[28957] = 8'b0;
    XRAM[28958] = 8'b0;
    XRAM[28959] = 8'b0;
    XRAM[28960] = 8'b0;
    XRAM[28961] = 8'b0;
    XRAM[28962] = 8'b0;
    XRAM[28963] = 8'b0;
    XRAM[28964] = 8'b0;
    XRAM[28965] = 8'b0;
    XRAM[28966] = 8'b0;
    XRAM[28967] = 8'b0;
    XRAM[28968] = 8'b0;
    XRAM[28969] = 8'b0;
    XRAM[28970] = 8'b0;
    XRAM[28971] = 8'b0;
    XRAM[28972] = 8'b0;
    XRAM[28973] = 8'b0;
    XRAM[28974] = 8'b0;
    XRAM[28975] = 8'b0;
    XRAM[28976] = 8'b0;
    XRAM[28977] = 8'b0;
    XRAM[28978] = 8'b0;
    XRAM[28979] = 8'b0;
    XRAM[28980] = 8'b0;
    XRAM[28981] = 8'b0;
    XRAM[28982] = 8'b0;
    XRAM[28983] = 8'b0;
    XRAM[28984] = 8'b0;
    XRAM[28985] = 8'b0;
    XRAM[28986] = 8'b0;
    XRAM[28987] = 8'b0;
    XRAM[28988] = 8'b0;
    XRAM[28989] = 8'b0;
    XRAM[28990] = 8'b0;
    XRAM[28991] = 8'b0;
    XRAM[28992] = 8'b0;
    XRAM[28993] = 8'b0;
    XRAM[28994] = 8'b0;
    XRAM[28995] = 8'b0;
    XRAM[28996] = 8'b0;
    XRAM[28997] = 8'b0;
    XRAM[28998] = 8'b0;
    XRAM[28999] = 8'b0;
    XRAM[29000] = 8'b0;
    XRAM[29001] = 8'b0;
    XRAM[29002] = 8'b0;
    XRAM[29003] = 8'b0;
    XRAM[29004] = 8'b0;
    XRAM[29005] = 8'b0;
    XRAM[29006] = 8'b0;
    XRAM[29007] = 8'b0;
    XRAM[29008] = 8'b0;
    XRAM[29009] = 8'b0;
    XRAM[29010] = 8'b0;
    XRAM[29011] = 8'b0;
    XRAM[29012] = 8'b0;
    XRAM[29013] = 8'b0;
    XRAM[29014] = 8'b0;
    XRAM[29015] = 8'b0;
    XRAM[29016] = 8'b0;
    XRAM[29017] = 8'b0;
    XRAM[29018] = 8'b0;
    XRAM[29019] = 8'b0;
    XRAM[29020] = 8'b0;
    XRAM[29021] = 8'b0;
    XRAM[29022] = 8'b0;
    XRAM[29023] = 8'b0;
    XRAM[29024] = 8'b0;
    XRAM[29025] = 8'b0;
    XRAM[29026] = 8'b0;
    XRAM[29027] = 8'b0;
    XRAM[29028] = 8'b0;
    XRAM[29029] = 8'b0;
    XRAM[29030] = 8'b0;
    XRAM[29031] = 8'b0;
    XRAM[29032] = 8'b0;
    XRAM[29033] = 8'b0;
    XRAM[29034] = 8'b0;
    XRAM[29035] = 8'b0;
    XRAM[29036] = 8'b0;
    XRAM[29037] = 8'b0;
    XRAM[29038] = 8'b0;
    XRAM[29039] = 8'b0;
    XRAM[29040] = 8'b0;
    XRAM[29041] = 8'b0;
    XRAM[29042] = 8'b0;
    XRAM[29043] = 8'b0;
    XRAM[29044] = 8'b0;
    XRAM[29045] = 8'b0;
    XRAM[29046] = 8'b0;
    XRAM[29047] = 8'b0;
    XRAM[29048] = 8'b0;
    XRAM[29049] = 8'b0;
    XRAM[29050] = 8'b0;
    XRAM[29051] = 8'b0;
    XRAM[29052] = 8'b0;
    XRAM[29053] = 8'b0;
    XRAM[29054] = 8'b0;
    XRAM[29055] = 8'b0;
    XRAM[29056] = 8'b0;
    XRAM[29057] = 8'b0;
    XRAM[29058] = 8'b0;
    XRAM[29059] = 8'b0;
    XRAM[29060] = 8'b0;
    XRAM[29061] = 8'b0;
    XRAM[29062] = 8'b0;
    XRAM[29063] = 8'b0;
    XRAM[29064] = 8'b0;
    XRAM[29065] = 8'b0;
    XRAM[29066] = 8'b0;
    XRAM[29067] = 8'b0;
    XRAM[29068] = 8'b0;
    XRAM[29069] = 8'b0;
    XRAM[29070] = 8'b0;
    XRAM[29071] = 8'b0;
    XRAM[29072] = 8'b0;
    XRAM[29073] = 8'b0;
    XRAM[29074] = 8'b0;
    XRAM[29075] = 8'b0;
    XRAM[29076] = 8'b0;
    XRAM[29077] = 8'b0;
    XRAM[29078] = 8'b0;
    XRAM[29079] = 8'b0;
    XRAM[29080] = 8'b0;
    XRAM[29081] = 8'b0;
    XRAM[29082] = 8'b0;
    XRAM[29083] = 8'b0;
    XRAM[29084] = 8'b0;
    XRAM[29085] = 8'b0;
    XRAM[29086] = 8'b0;
    XRAM[29087] = 8'b0;
    XRAM[29088] = 8'b0;
    XRAM[29089] = 8'b0;
    XRAM[29090] = 8'b0;
    XRAM[29091] = 8'b0;
    XRAM[29092] = 8'b0;
    XRAM[29093] = 8'b0;
    XRAM[29094] = 8'b0;
    XRAM[29095] = 8'b0;
    XRAM[29096] = 8'b0;
    XRAM[29097] = 8'b0;
    XRAM[29098] = 8'b0;
    XRAM[29099] = 8'b0;
    XRAM[29100] = 8'b0;
    XRAM[29101] = 8'b0;
    XRAM[29102] = 8'b0;
    XRAM[29103] = 8'b0;
    XRAM[29104] = 8'b0;
    XRAM[29105] = 8'b0;
    XRAM[29106] = 8'b0;
    XRAM[29107] = 8'b0;
    XRAM[29108] = 8'b0;
    XRAM[29109] = 8'b0;
    XRAM[29110] = 8'b0;
    XRAM[29111] = 8'b0;
    XRAM[29112] = 8'b0;
    XRAM[29113] = 8'b0;
    XRAM[29114] = 8'b0;
    XRAM[29115] = 8'b0;
    XRAM[29116] = 8'b0;
    XRAM[29117] = 8'b0;
    XRAM[29118] = 8'b0;
    XRAM[29119] = 8'b0;
    XRAM[29120] = 8'b0;
    XRAM[29121] = 8'b0;
    XRAM[29122] = 8'b0;
    XRAM[29123] = 8'b0;
    XRAM[29124] = 8'b0;
    XRAM[29125] = 8'b0;
    XRAM[29126] = 8'b0;
    XRAM[29127] = 8'b0;
    XRAM[29128] = 8'b0;
    XRAM[29129] = 8'b0;
    XRAM[29130] = 8'b0;
    XRAM[29131] = 8'b0;
    XRAM[29132] = 8'b0;
    XRAM[29133] = 8'b0;
    XRAM[29134] = 8'b0;
    XRAM[29135] = 8'b0;
    XRAM[29136] = 8'b0;
    XRAM[29137] = 8'b0;
    XRAM[29138] = 8'b0;
    XRAM[29139] = 8'b0;
    XRAM[29140] = 8'b0;
    XRAM[29141] = 8'b0;
    XRAM[29142] = 8'b0;
    XRAM[29143] = 8'b0;
    XRAM[29144] = 8'b0;
    XRAM[29145] = 8'b0;
    XRAM[29146] = 8'b0;
    XRAM[29147] = 8'b0;
    XRAM[29148] = 8'b0;
    XRAM[29149] = 8'b0;
    XRAM[29150] = 8'b0;
    XRAM[29151] = 8'b0;
    XRAM[29152] = 8'b0;
    XRAM[29153] = 8'b0;
    XRAM[29154] = 8'b0;
    XRAM[29155] = 8'b0;
    XRAM[29156] = 8'b0;
    XRAM[29157] = 8'b0;
    XRAM[29158] = 8'b0;
    XRAM[29159] = 8'b0;
    XRAM[29160] = 8'b0;
    XRAM[29161] = 8'b0;
    XRAM[29162] = 8'b0;
    XRAM[29163] = 8'b0;
    XRAM[29164] = 8'b0;
    XRAM[29165] = 8'b0;
    XRAM[29166] = 8'b0;
    XRAM[29167] = 8'b0;
    XRAM[29168] = 8'b0;
    XRAM[29169] = 8'b0;
    XRAM[29170] = 8'b0;
    XRAM[29171] = 8'b0;
    XRAM[29172] = 8'b0;
    XRAM[29173] = 8'b0;
    XRAM[29174] = 8'b0;
    XRAM[29175] = 8'b0;
    XRAM[29176] = 8'b0;
    XRAM[29177] = 8'b0;
    XRAM[29178] = 8'b0;
    XRAM[29179] = 8'b0;
    XRAM[29180] = 8'b0;
    XRAM[29181] = 8'b0;
    XRAM[29182] = 8'b0;
    XRAM[29183] = 8'b0;
    XRAM[29184] = 8'b0;
    XRAM[29185] = 8'b0;
    XRAM[29186] = 8'b0;
    XRAM[29187] = 8'b0;
    XRAM[29188] = 8'b0;
    XRAM[29189] = 8'b0;
    XRAM[29190] = 8'b0;
    XRAM[29191] = 8'b0;
    XRAM[29192] = 8'b0;
    XRAM[29193] = 8'b0;
    XRAM[29194] = 8'b0;
    XRAM[29195] = 8'b0;
    XRAM[29196] = 8'b0;
    XRAM[29197] = 8'b0;
    XRAM[29198] = 8'b0;
    XRAM[29199] = 8'b0;
    XRAM[29200] = 8'b0;
    XRAM[29201] = 8'b0;
    XRAM[29202] = 8'b0;
    XRAM[29203] = 8'b0;
    XRAM[29204] = 8'b0;
    XRAM[29205] = 8'b0;
    XRAM[29206] = 8'b0;
    XRAM[29207] = 8'b0;
    XRAM[29208] = 8'b0;
    XRAM[29209] = 8'b0;
    XRAM[29210] = 8'b0;
    XRAM[29211] = 8'b0;
    XRAM[29212] = 8'b0;
    XRAM[29213] = 8'b0;
    XRAM[29214] = 8'b0;
    XRAM[29215] = 8'b0;
    XRAM[29216] = 8'b0;
    XRAM[29217] = 8'b0;
    XRAM[29218] = 8'b0;
    XRAM[29219] = 8'b0;
    XRAM[29220] = 8'b0;
    XRAM[29221] = 8'b0;
    XRAM[29222] = 8'b0;
    XRAM[29223] = 8'b0;
    XRAM[29224] = 8'b0;
    XRAM[29225] = 8'b0;
    XRAM[29226] = 8'b0;
    XRAM[29227] = 8'b0;
    XRAM[29228] = 8'b0;
    XRAM[29229] = 8'b0;
    XRAM[29230] = 8'b0;
    XRAM[29231] = 8'b0;
    XRAM[29232] = 8'b0;
    XRAM[29233] = 8'b0;
    XRAM[29234] = 8'b0;
    XRAM[29235] = 8'b0;
    XRAM[29236] = 8'b0;
    XRAM[29237] = 8'b0;
    XRAM[29238] = 8'b0;
    XRAM[29239] = 8'b0;
    XRAM[29240] = 8'b0;
    XRAM[29241] = 8'b0;
    XRAM[29242] = 8'b0;
    XRAM[29243] = 8'b0;
    XRAM[29244] = 8'b0;
    XRAM[29245] = 8'b0;
    XRAM[29246] = 8'b0;
    XRAM[29247] = 8'b0;
    XRAM[29248] = 8'b0;
    XRAM[29249] = 8'b0;
    XRAM[29250] = 8'b0;
    XRAM[29251] = 8'b0;
    XRAM[29252] = 8'b0;
    XRAM[29253] = 8'b0;
    XRAM[29254] = 8'b0;
    XRAM[29255] = 8'b0;
    XRAM[29256] = 8'b0;
    XRAM[29257] = 8'b0;
    XRAM[29258] = 8'b0;
    XRAM[29259] = 8'b0;
    XRAM[29260] = 8'b0;
    XRAM[29261] = 8'b0;
    XRAM[29262] = 8'b0;
    XRAM[29263] = 8'b0;
    XRAM[29264] = 8'b0;
    XRAM[29265] = 8'b0;
    XRAM[29266] = 8'b0;
    XRAM[29267] = 8'b0;
    XRAM[29268] = 8'b0;
    XRAM[29269] = 8'b0;
    XRAM[29270] = 8'b0;
    XRAM[29271] = 8'b0;
    XRAM[29272] = 8'b0;
    XRAM[29273] = 8'b0;
    XRAM[29274] = 8'b0;
    XRAM[29275] = 8'b0;
    XRAM[29276] = 8'b0;
    XRAM[29277] = 8'b0;
    XRAM[29278] = 8'b0;
    XRAM[29279] = 8'b0;
    XRAM[29280] = 8'b0;
    XRAM[29281] = 8'b0;
    XRAM[29282] = 8'b0;
    XRAM[29283] = 8'b0;
    XRAM[29284] = 8'b0;
    XRAM[29285] = 8'b0;
    XRAM[29286] = 8'b0;
    XRAM[29287] = 8'b0;
    XRAM[29288] = 8'b0;
    XRAM[29289] = 8'b0;
    XRAM[29290] = 8'b0;
    XRAM[29291] = 8'b0;
    XRAM[29292] = 8'b0;
    XRAM[29293] = 8'b0;
    XRAM[29294] = 8'b0;
    XRAM[29295] = 8'b0;
    XRAM[29296] = 8'b0;
    XRAM[29297] = 8'b0;
    XRAM[29298] = 8'b0;
    XRAM[29299] = 8'b0;
    XRAM[29300] = 8'b0;
    XRAM[29301] = 8'b0;
    XRAM[29302] = 8'b0;
    XRAM[29303] = 8'b0;
    XRAM[29304] = 8'b0;
    XRAM[29305] = 8'b0;
    XRAM[29306] = 8'b0;
    XRAM[29307] = 8'b0;
    XRAM[29308] = 8'b0;
    XRAM[29309] = 8'b0;
    XRAM[29310] = 8'b0;
    XRAM[29311] = 8'b0;
    XRAM[29312] = 8'b0;
    XRAM[29313] = 8'b0;
    XRAM[29314] = 8'b0;
    XRAM[29315] = 8'b0;
    XRAM[29316] = 8'b0;
    XRAM[29317] = 8'b0;
    XRAM[29318] = 8'b0;
    XRAM[29319] = 8'b0;
    XRAM[29320] = 8'b0;
    XRAM[29321] = 8'b0;
    XRAM[29322] = 8'b0;
    XRAM[29323] = 8'b0;
    XRAM[29324] = 8'b0;
    XRAM[29325] = 8'b0;
    XRAM[29326] = 8'b0;
    XRAM[29327] = 8'b0;
    XRAM[29328] = 8'b0;
    XRAM[29329] = 8'b0;
    XRAM[29330] = 8'b0;
    XRAM[29331] = 8'b0;
    XRAM[29332] = 8'b0;
    XRAM[29333] = 8'b0;
    XRAM[29334] = 8'b0;
    XRAM[29335] = 8'b0;
    XRAM[29336] = 8'b0;
    XRAM[29337] = 8'b0;
    XRAM[29338] = 8'b0;
    XRAM[29339] = 8'b0;
    XRAM[29340] = 8'b0;
    XRAM[29341] = 8'b0;
    XRAM[29342] = 8'b0;
    XRAM[29343] = 8'b0;
    XRAM[29344] = 8'b0;
    XRAM[29345] = 8'b0;
    XRAM[29346] = 8'b0;
    XRAM[29347] = 8'b0;
    XRAM[29348] = 8'b0;
    XRAM[29349] = 8'b0;
    XRAM[29350] = 8'b0;
    XRAM[29351] = 8'b0;
    XRAM[29352] = 8'b0;
    XRAM[29353] = 8'b0;
    XRAM[29354] = 8'b0;
    XRAM[29355] = 8'b0;
    XRAM[29356] = 8'b0;
    XRAM[29357] = 8'b0;
    XRAM[29358] = 8'b0;
    XRAM[29359] = 8'b0;
    XRAM[29360] = 8'b0;
    XRAM[29361] = 8'b0;
    XRAM[29362] = 8'b0;
    XRAM[29363] = 8'b0;
    XRAM[29364] = 8'b0;
    XRAM[29365] = 8'b0;
    XRAM[29366] = 8'b0;
    XRAM[29367] = 8'b0;
    XRAM[29368] = 8'b0;
    XRAM[29369] = 8'b0;
    XRAM[29370] = 8'b0;
    XRAM[29371] = 8'b0;
    XRAM[29372] = 8'b0;
    XRAM[29373] = 8'b0;
    XRAM[29374] = 8'b0;
    XRAM[29375] = 8'b0;
    XRAM[29376] = 8'b0;
    XRAM[29377] = 8'b0;
    XRAM[29378] = 8'b0;
    XRAM[29379] = 8'b0;
    XRAM[29380] = 8'b0;
    XRAM[29381] = 8'b0;
    XRAM[29382] = 8'b0;
    XRAM[29383] = 8'b0;
    XRAM[29384] = 8'b0;
    XRAM[29385] = 8'b0;
    XRAM[29386] = 8'b0;
    XRAM[29387] = 8'b0;
    XRAM[29388] = 8'b0;
    XRAM[29389] = 8'b0;
    XRAM[29390] = 8'b0;
    XRAM[29391] = 8'b0;
    XRAM[29392] = 8'b0;
    XRAM[29393] = 8'b0;
    XRAM[29394] = 8'b0;
    XRAM[29395] = 8'b0;
    XRAM[29396] = 8'b0;
    XRAM[29397] = 8'b0;
    XRAM[29398] = 8'b0;
    XRAM[29399] = 8'b0;
    XRAM[29400] = 8'b0;
    XRAM[29401] = 8'b0;
    XRAM[29402] = 8'b0;
    XRAM[29403] = 8'b0;
    XRAM[29404] = 8'b0;
    XRAM[29405] = 8'b0;
    XRAM[29406] = 8'b0;
    XRAM[29407] = 8'b0;
    XRAM[29408] = 8'b0;
    XRAM[29409] = 8'b0;
    XRAM[29410] = 8'b0;
    XRAM[29411] = 8'b0;
    XRAM[29412] = 8'b0;
    XRAM[29413] = 8'b0;
    XRAM[29414] = 8'b0;
    XRAM[29415] = 8'b0;
    XRAM[29416] = 8'b0;
    XRAM[29417] = 8'b0;
    XRAM[29418] = 8'b0;
    XRAM[29419] = 8'b0;
    XRAM[29420] = 8'b0;
    XRAM[29421] = 8'b0;
    XRAM[29422] = 8'b0;
    XRAM[29423] = 8'b0;
    XRAM[29424] = 8'b0;
    XRAM[29425] = 8'b0;
    XRAM[29426] = 8'b0;
    XRAM[29427] = 8'b0;
    XRAM[29428] = 8'b0;
    XRAM[29429] = 8'b0;
    XRAM[29430] = 8'b0;
    XRAM[29431] = 8'b0;
    XRAM[29432] = 8'b0;
    XRAM[29433] = 8'b0;
    XRAM[29434] = 8'b0;
    XRAM[29435] = 8'b0;
    XRAM[29436] = 8'b0;
    XRAM[29437] = 8'b0;
    XRAM[29438] = 8'b0;
    XRAM[29439] = 8'b0;
    XRAM[29440] = 8'b0;
    XRAM[29441] = 8'b0;
    XRAM[29442] = 8'b0;
    XRAM[29443] = 8'b0;
    XRAM[29444] = 8'b0;
    XRAM[29445] = 8'b0;
    XRAM[29446] = 8'b0;
    XRAM[29447] = 8'b0;
    XRAM[29448] = 8'b0;
    XRAM[29449] = 8'b0;
    XRAM[29450] = 8'b0;
    XRAM[29451] = 8'b0;
    XRAM[29452] = 8'b0;
    XRAM[29453] = 8'b0;
    XRAM[29454] = 8'b0;
    XRAM[29455] = 8'b0;
    XRAM[29456] = 8'b0;
    XRAM[29457] = 8'b0;
    XRAM[29458] = 8'b0;
    XRAM[29459] = 8'b0;
    XRAM[29460] = 8'b0;
    XRAM[29461] = 8'b0;
    XRAM[29462] = 8'b0;
    XRAM[29463] = 8'b0;
    XRAM[29464] = 8'b0;
    XRAM[29465] = 8'b0;
    XRAM[29466] = 8'b0;
    XRAM[29467] = 8'b0;
    XRAM[29468] = 8'b0;
    XRAM[29469] = 8'b0;
    XRAM[29470] = 8'b0;
    XRAM[29471] = 8'b0;
    XRAM[29472] = 8'b0;
    XRAM[29473] = 8'b0;
    XRAM[29474] = 8'b0;
    XRAM[29475] = 8'b0;
    XRAM[29476] = 8'b0;
    XRAM[29477] = 8'b0;
    XRAM[29478] = 8'b0;
    XRAM[29479] = 8'b0;
    XRAM[29480] = 8'b0;
    XRAM[29481] = 8'b0;
    XRAM[29482] = 8'b0;
    XRAM[29483] = 8'b0;
    XRAM[29484] = 8'b0;
    XRAM[29485] = 8'b0;
    XRAM[29486] = 8'b0;
    XRAM[29487] = 8'b0;
    XRAM[29488] = 8'b0;
    XRAM[29489] = 8'b0;
    XRAM[29490] = 8'b0;
    XRAM[29491] = 8'b0;
    XRAM[29492] = 8'b0;
    XRAM[29493] = 8'b0;
    XRAM[29494] = 8'b0;
    XRAM[29495] = 8'b0;
    XRAM[29496] = 8'b0;
    XRAM[29497] = 8'b0;
    XRAM[29498] = 8'b0;
    XRAM[29499] = 8'b0;
    XRAM[29500] = 8'b0;
    XRAM[29501] = 8'b0;
    XRAM[29502] = 8'b0;
    XRAM[29503] = 8'b0;
    XRAM[29504] = 8'b0;
    XRAM[29505] = 8'b0;
    XRAM[29506] = 8'b0;
    XRAM[29507] = 8'b0;
    XRAM[29508] = 8'b0;
    XRAM[29509] = 8'b0;
    XRAM[29510] = 8'b0;
    XRAM[29511] = 8'b0;
    XRAM[29512] = 8'b0;
    XRAM[29513] = 8'b0;
    XRAM[29514] = 8'b0;
    XRAM[29515] = 8'b0;
    XRAM[29516] = 8'b0;
    XRAM[29517] = 8'b0;
    XRAM[29518] = 8'b0;
    XRAM[29519] = 8'b0;
    XRAM[29520] = 8'b0;
    XRAM[29521] = 8'b0;
    XRAM[29522] = 8'b0;
    XRAM[29523] = 8'b0;
    XRAM[29524] = 8'b0;
    XRAM[29525] = 8'b0;
    XRAM[29526] = 8'b0;
    XRAM[29527] = 8'b0;
    XRAM[29528] = 8'b0;
    XRAM[29529] = 8'b0;
    XRAM[29530] = 8'b0;
    XRAM[29531] = 8'b0;
    XRAM[29532] = 8'b0;
    XRAM[29533] = 8'b0;
    XRAM[29534] = 8'b0;
    XRAM[29535] = 8'b0;
    XRAM[29536] = 8'b0;
    XRAM[29537] = 8'b0;
    XRAM[29538] = 8'b0;
    XRAM[29539] = 8'b0;
    XRAM[29540] = 8'b0;
    XRAM[29541] = 8'b0;
    XRAM[29542] = 8'b0;
    XRAM[29543] = 8'b0;
    XRAM[29544] = 8'b0;
    XRAM[29545] = 8'b0;
    XRAM[29546] = 8'b0;
    XRAM[29547] = 8'b0;
    XRAM[29548] = 8'b0;
    XRAM[29549] = 8'b0;
    XRAM[29550] = 8'b0;
    XRAM[29551] = 8'b0;
    XRAM[29552] = 8'b0;
    XRAM[29553] = 8'b0;
    XRAM[29554] = 8'b0;
    XRAM[29555] = 8'b0;
    XRAM[29556] = 8'b0;
    XRAM[29557] = 8'b0;
    XRAM[29558] = 8'b0;
    XRAM[29559] = 8'b0;
    XRAM[29560] = 8'b0;
    XRAM[29561] = 8'b0;
    XRAM[29562] = 8'b0;
    XRAM[29563] = 8'b0;
    XRAM[29564] = 8'b0;
    XRAM[29565] = 8'b0;
    XRAM[29566] = 8'b0;
    XRAM[29567] = 8'b0;
    XRAM[29568] = 8'b0;
    XRAM[29569] = 8'b0;
    XRAM[29570] = 8'b0;
    XRAM[29571] = 8'b0;
    XRAM[29572] = 8'b0;
    XRAM[29573] = 8'b0;
    XRAM[29574] = 8'b0;
    XRAM[29575] = 8'b0;
    XRAM[29576] = 8'b0;
    XRAM[29577] = 8'b0;
    XRAM[29578] = 8'b0;
    XRAM[29579] = 8'b0;
    XRAM[29580] = 8'b0;
    XRAM[29581] = 8'b0;
    XRAM[29582] = 8'b0;
    XRAM[29583] = 8'b0;
    XRAM[29584] = 8'b0;
    XRAM[29585] = 8'b0;
    XRAM[29586] = 8'b0;
    XRAM[29587] = 8'b0;
    XRAM[29588] = 8'b0;
    XRAM[29589] = 8'b0;
    XRAM[29590] = 8'b0;
    XRAM[29591] = 8'b0;
    XRAM[29592] = 8'b0;
    XRAM[29593] = 8'b0;
    XRAM[29594] = 8'b0;
    XRAM[29595] = 8'b0;
    XRAM[29596] = 8'b0;
    XRAM[29597] = 8'b0;
    XRAM[29598] = 8'b0;
    XRAM[29599] = 8'b0;
    XRAM[29600] = 8'b0;
    XRAM[29601] = 8'b0;
    XRAM[29602] = 8'b0;
    XRAM[29603] = 8'b0;
    XRAM[29604] = 8'b0;
    XRAM[29605] = 8'b0;
    XRAM[29606] = 8'b0;
    XRAM[29607] = 8'b0;
    XRAM[29608] = 8'b0;
    XRAM[29609] = 8'b0;
    XRAM[29610] = 8'b0;
    XRAM[29611] = 8'b0;
    XRAM[29612] = 8'b0;
    XRAM[29613] = 8'b0;
    XRAM[29614] = 8'b0;
    XRAM[29615] = 8'b0;
    XRAM[29616] = 8'b0;
    XRAM[29617] = 8'b0;
    XRAM[29618] = 8'b0;
    XRAM[29619] = 8'b0;
    XRAM[29620] = 8'b0;
    XRAM[29621] = 8'b0;
    XRAM[29622] = 8'b0;
    XRAM[29623] = 8'b0;
    XRAM[29624] = 8'b0;
    XRAM[29625] = 8'b0;
    XRAM[29626] = 8'b0;
    XRAM[29627] = 8'b0;
    XRAM[29628] = 8'b0;
    XRAM[29629] = 8'b0;
    XRAM[29630] = 8'b0;
    XRAM[29631] = 8'b0;
    XRAM[29632] = 8'b0;
    XRAM[29633] = 8'b0;
    XRAM[29634] = 8'b0;
    XRAM[29635] = 8'b0;
    XRAM[29636] = 8'b0;
    XRAM[29637] = 8'b0;
    XRAM[29638] = 8'b0;
    XRAM[29639] = 8'b0;
    XRAM[29640] = 8'b0;
    XRAM[29641] = 8'b0;
    XRAM[29642] = 8'b0;
    XRAM[29643] = 8'b0;
    XRAM[29644] = 8'b0;
    XRAM[29645] = 8'b0;
    XRAM[29646] = 8'b0;
    XRAM[29647] = 8'b0;
    XRAM[29648] = 8'b0;
    XRAM[29649] = 8'b0;
    XRAM[29650] = 8'b0;
    XRAM[29651] = 8'b0;
    XRAM[29652] = 8'b0;
    XRAM[29653] = 8'b0;
    XRAM[29654] = 8'b0;
    XRAM[29655] = 8'b0;
    XRAM[29656] = 8'b0;
    XRAM[29657] = 8'b0;
    XRAM[29658] = 8'b0;
    XRAM[29659] = 8'b0;
    XRAM[29660] = 8'b0;
    XRAM[29661] = 8'b0;
    XRAM[29662] = 8'b0;
    XRAM[29663] = 8'b0;
    XRAM[29664] = 8'b0;
    XRAM[29665] = 8'b0;
    XRAM[29666] = 8'b0;
    XRAM[29667] = 8'b0;
    XRAM[29668] = 8'b0;
    XRAM[29669] = 8'b0;
    XRAM[29670] = 8'b0;
    XRAM[29671] = 8'b0;
    XRAM[29672] = 8'b0;
    XRAM[29673] = 8'b0;
    XRAM[29674] = 8'b0;
    XRAM[29675] = 8'b0;
    XRAM[29676] = 8'b0;
    XRAM[29677] = 8'b0;
    XRAM[29678] = 8'b0;
    XRAM[29679] = 8'b0;
    XRAM[29680] = 8'b0;
    XRAM[29681] = 8'b0;
    XRAM[29682] = 8'b0;
    XRAM[29683] = 8'b0;
    XRAM[29684] = 8'b0;
    XRAM[29685] = 8'b0;
    XRAM[29686] = 8'b0;
    XRAM[29687] = 8'b0;
    XRAM[29688] = 8'b0;
    XRAM[29689] = 8'b0;
    XRAM[29690] = 8'b0;
    XRAM[29691] = 8'b0;
    XRAM[29692] = 8'b0;
    XRAM[29693] = 8'b0;
    XRAM[29694] = 8'b0;
    XRAM[29695] = 8'b0;
    XRAM[29696] = 8'b0;
    XRAM[29697] = 8'b0;
    XRAM[29698] = 8'b0;
    XRAM[29699] = 8'b0;
    XRAM[29700] = 8'b0;
    XRAM[29701] = 8'b0;
    XRAM[29702] = 8'b0;
    XRAM[29703] = 8'b0;
    XRAM[29704] = 8'b0;
    XRAM[29705] = 8'b0;
    XRAM[29706] = 8'b0;
    XRAM[29707] = 8'b0;
    XRAM[29708] = 8'b0;
    XRAM[29709] = 8'b0;
    XRAM[29710] = 8'b0;
    XRAM[29711] = 8'b0;
    XRAM[29712] = 8'b0;
    XRAM[29713] = 8'b0;
    XRAM[29714] = 8'b0;
    XRAM[29715] = 8'b0;
    XRAM[29716] = 8'b0;
    XRAM[29717] = 8'b0;
    XRAM[29718] = 8'b0;
    XRAM[29719] = 8'b0;
    XRAM[29720] = 8'b0;
    XRAM[29721] = 8'b0;
    XRAM[29722] = 8'b0;
    XRAM[29723] = 8'b0;
    XRAM[29724] = 8'b0;
    XRAM[29725] = 8'b0;
    XRAM[29726] = 8'b0;
    XRAM[29727] = 8'b0;
    XRAM[29728] = 8'b0;
    XRAM[29729] = 8'b0;
    XRAM[29730] = 8'b0;
    XRAM[29731] = 8'b0;
    XRAM[29732] = 8'b0;
    XRAM[29733] = 8'b0;
    XRAM[29734] = 8'b0;
    XRAM[29735] = 8'b0;
    XRAM[29736] = 8'b0;
    XRAM[29737] = 8'b0;
    XRAM[29738] = 8'b0;
    XRAM[29739] = 8'b0;
    XRAM[29740] = 8'b0;
    XRAM[29741] = 8'b0;
    XRAM[29742] = 8'b0;
    XRAM[29743] = 8'b0;
    XRAM[29744] = 8'b0;
    XRAM[29745] = 8'b0;
    XRAM[29746] = 8'b0;
    XRAM[29747] = 8'b0;
    XRAM[29748] = 8'b0;
    XRAM[29749] = 8'b0;
    XRAM[29750] = 8'b0;
    XRAM[29751] = 8'b0;
    XRAM[29752] = 8'b0;
    XRAM[29753] = 8'b0;
    XRAM[29754] = 8'b0;
    XRAM[29755] = 8'b0;
    XRAM[29756] = 8'b0;
    XRAM[29757] = 8'b0;
    XRAM[29758] = 8'b0;
    XRAM[29759] = 8'b0;
    XRAM[29760] = 8'b0;
    XRAM[29761] = 8'b0;
    XRAM[29762] = 8'b0;
    XRAM[29763] = 8'b0;
    XRAM[29764] = 8'b0;
    XRAM[29765] = 8'b0;
    XRAM[29766] = 8'b0;
    XRAM[29767] = 8'b0;
    XRAM[29768] = 8'b0;
    XRAM[29769] = 8'b0;
    XRAM[29770] = 8'b0;
    XRAM[29771] = 8'b0;
    XRAM[29772] = 8'b0;
    XRAM[29773] = 8'b0;
    XRAM[29774] = 8'b0;
    XRAM[29775] = 8'b0;
    XRAM[29776] = 8'b0;
    XRAM[29777] = 8'b0;
    XRAM[29778] = 8'b0;
    XRAM[29779] = 8'b0;
    XRAM[29780] = 8'b0;
    XRAM[29781] = 8'b0;
    XRAM[29782] = 8'b0;
    XRAM[29783] = 8'b0;
    XRAM[29784] = 8'b0;
    XRAM[29785] = 8'b0;
    XRAM[29786] = 8'b0;
    XRAM[29787] = 8'b0;
    XRAM[29788] = 8'b0;
    XRAM[29789] = 8'b0;
    XRAM[29790] = 8'b0;
    XRAM[29791] = 8'b0;
    XRAM[29792] = 8'b0;
    XRAM[29793] = 8'b0;
    XRAM[29794] = 8'b0;
    XRAM[29795] = 8'b0;
    XRAM[29796] = 8'b0;
    XRAM[29797] = 8'b0;
    XRAM[29798] = 8'b0;
    XRAM[29799] = 8'b0;
    XRAM[29800] = 8'b0;
    XRAM[29801] = 8'b0;
    XRAM[29802] = 8'b0;
    XRAM[29803] = 8'b0;
    XRAM[29804] = 8'b0;
    XRAM[29805] = 8'b0;
    XRAM[29806] = 8'b0;
    XRAM[29807] = 8'b0;
    XRAM[29808] = 8'b0;
    XRAM[29809] = 8'b0;
    XRAM[29810] = 8'b0;
    XRAM[29811] = 8'b0;
    XRAM[29812] = 8'b0;
    XRAM[29813] = 8'b0;
    XRAM[29814] = 8'b0;
    XRAM[29815] = 8'b0;
    XRAM[29816] = 8'b0;
    XRAM[29817] = 8'b0;
    XRAM[29818] = 8'b0;
    XRAM[29819] = 8'b0;
    XRAM[29820] = 8'b0;
    XRAM[29821] = 8'b0;
    XRAM[29822] = 8'b0;
    XRAM[29823] = 8'b0;
    XRAM[29824] = 8'b0;
    XRAM[29825] = 8'b0;
    XRAM[29826] = 8'b0;
    XRAM[29827] = 8'b0;
    XRAM[29828] = 8'b0;
    XRAM[29829] = 8'b0;
    XRAM[29830] = 8'b0;
    XRAM[29831] = 8'b0;
    XRAM[29832] = 8'b0;
    XRAM[29833] = 8'b0;
    XRAM[29834] = 8'b0;
    XRAM[29835] = 8'b0;
    XRAM[29836] = 8'b0;
    XRAM[29837] = 8'b0;
    XRAM[29838] = 8'b0;
    XRAM[29839] = 8'b0;
    XRAM[29840] = 8'b0;
    XRAM[29841] = 8'b0;
    XRAM[29842] = 8'b0;
    XRAM[29843] = 8'b0;
    XRAM[29844] = 8'b0;
    XRAM[29845] = 8'b0;
    XRAM[29846] = 8'b0;
    XRAM[29847] = 8'b0;
    XRAM[29848] = 8'b0;
    XRAM[29849] = 8'b0;
    XRAM[29850] = 8'b0;
    XRAM[29851] = 8'b0;
    XRAM[29852] = 8'b0;
    XRAM[29853] = 8'b0;
    XRAM[29854] = 8'b0;
    XRAM[29855] = 8'b0;
    XRAM[29856] = 8'b0;
    XRAM[29857] = 8'b0;
    XRAM[29858] = 8'b0;
    XRAM[29859] = 8'b0;
    XRAM[29860] = 8'b0;
    XRAM[29861] = 8'b0;
    XRAM[29862] = 8'b0;
    XRAM[29863] = 8'b0;
    XRAM[29864] = 8'b0;
    XRAM[29865] = 8'b0;
    XRAM[29866] = 8'b0;
    XRAM[29867] = 8'b0;
    XRAM[29868] = 8'b0;
    XRAM[29869] = 8'b0;
    XRAM[29870] = 8'b0;
    XRAM[29871] = 8'b0;
    XRAM[29872] = 8'b0;
    XRAM[29873] = 8'b0;
    XRAM[29874] = 8'b0;
    XRAM[29875] = 8'b0;
    XRAM[29876] = 8'b0;
    XRAM[29877] = 8'b0;
    XRAM[29878] = 8'b0;
    XRAM[29879] = 8'b0;
    XRAM[29880] = 8'b0;
    XRAM[29881] = 8'b0;
    XRAM[29882] = 8'b0;
    XRAM[29883] = 8'b0;
    XRAM[29884] = 8'b0;
    XRAM[29885] = 8'b0;
    XRAM[29886] = 8'b0;
    XRAM[29887] = 8'b0;
    XRAM[29888] = 8'b0;
    XRAM[29889] = 8'b0;
    XRAM[29890] = 8'b0;
    XRAM[29891] = 8'b0;
    XRAM[29892] = 8'b0;
    XRAM[29893] = 8'b0;
    XRAM[29894] = 8'b0;
    XRAM[29895] = 8'b0;
    XRAM[29896] = 8'b0;
    XRAM[29897] = 8'b0;
    XRAM[29898] = 8'b0;
    XRAM[29899] = 8'b0;
    XRAM[29900] = 8'b0;
    XRAM[29901] = 8'b0;
    XRAM[29902] = 8'b0;
    XRAM[29903] = 8'b0;
    XRAM[29904] = 8'b0;
    XRAM[29905] = 8'b0;
    XRAM[29906] = 8'b0;
    XRAM[29907] = 8'b0;
    XRAM[29908] = 8'b0;
    XRAM[29909] = 8'b0;
    XRAM[29910] = 8'b0;
    XRAM[29911] = 8'b0;
    XRAM[29912] = 8'b0;
    XRAM[29913] = 8'b0;
    XRAM[29914] = 8'b0;
    XRAM[29915] = 8'b0;
    XRAM[29916] = 8'b0;
    XRAM[29917] = 8'b0;
    XRAM[29918] = 8'b0;
    XRAM[29919] = 8'b0;
    XRAM[29920] = 8'b0;
    XRAM[29921] = 8'b0;
    XRAM[29922] = 8'b0;
    XRAM[29923] = 8'b0;
    XRAM[29924] = 8'b0;
    XRAM[29925] = 8'b0;
    XRAM[29926] = 8'b0;
    XRAM[29927] = 8'b0;
    XRAM[29928] = 8'b0;
    XRAM[29929] = 8'b0;
    XRAM[29930] = 8'b0;
    XRAM[29931] = 8'b0;
    XRAM[29932] = 8'b0;
    XRAM[29933] = 8'b0;
    XRAM[29934] = 8'b0;
    XRAM[29935] = 8'b0;
    XRAM[29936] = 8'b0;
    XRAM[29937] = 8'b0;
    XRAM[29938] = 8'b0;
    XRAM[29939] = 8'b0;
    XRAM[29940] = 8'b0;
    XRAM[29941] = 8'b0;
    XRAM[29942] = 8'b0;
    XRAM[29943] = 8'b0;
    XRAM[29944] = 8'b0;
    XRAM[29945] = 8'b0;
    XRAM[29946] = 8'b0;
    XRAM[29947] = 8'b0;
    XRAM[29948] = 8'b0;
    XRAM[29949] = 8'b0;
    XRAM[29950] = 8'b0;
    XRAM[29951] = 8'b0;
    XRAM[29952] = 8'b0;
    XRAM[29953] = 8'b0;
    XRAM[29954] = 8'b0;
    XRAM[29955] = 8'b0;
    XRAM[29956] = 8'b0;
    XRAM[29957] = 8'b0;
    XRAM[29958] = 8'b0;
    XRAM[29959] = 8'b0;
    XRAM[29960] = 8'b0;
    XRAM[29961] = 8'b0;
    XRAM[29962] = 8'b0;
    XRAM[29963] = 8'b0;
    XRAM[29964] = 8'b0;
    XRAM[29965] = 8'b0;
    XRAM[29966] = 8'b0;
    XRAM[29967] = 8'b0;
    XRAM[29968] = 8'b0;
    XRAM[29969] = 8'b0;
    XRAM[29970] = 8'b0;
    XRAM[29971] = 8'b0;
    XRAM[29972] = 8'b0;
    XRAM[29973] = 8'b0;
    XRAM[29974] = 8'b0;
    XRAM[29975] = 8'b0;
    XRAM[29976] = 8'b0;
    XRAM[29977] = 8'b0;
    XRAM[29978] = 8'b0;
    XRAM[29979] = 8'b0;
    XRAM[29980] = 8'b0;
    XRAM[29981] = 8'b0;
    XRAM[29982] = 8'b0;
    XRAM[29983] = 8'b0;
    XRAM[29984] = 8'b0;
    XRAM[29985] = 8'b0;
    XRAM[29986] = 8'b0;
    XRAM[29987] = 8'b0;
    XRAM[29988] = 8'b0;
    XRAM[29989] = 8'b0;
    XRAM[29990] = 8'b0;
    XRAM[29991] = 8'b0;
    XRAM[29992] = 8'b0;
    XRAM[29993] = 8'b0;
    XRAM[29994] = 8'b0;
    XRAM[29995] = 8'b0;
    XRAM[29996] = 8'b0;
    XRAM[29997] = 8'b0;
    XRAM[29998] = 8'b0;
    XRAM[29999] = 8'b0;
    XRAM[30000] = 8'b0;
    XRAM[30001] = 8'b0;
    XRAM[30002] = 8'b0;
    XRAM[30003] = 8'b0;
    XRAM[30004] = 8'b0;
    XRAM[30005] = 8'b0;
    XRAM[30006] = 8'b0;
    XRAM[30007] = 8'b0;
    XRAM[30008] = 8'b0;
    XRAM[30009] = 8'b0;
    XRAM[30010] = 8'b0;
    XRAM[30011] = 8'b0;
    XRAM[30012] = 8'b0;
    XRAM[30013] = 8'b0;
    XRAM[30014] = 8'b0;
    XRAM[30015] = 8'b0;
    XRAM[30016] = 8'b0;
    XRAM[30017] = 8'b0;
    XRAM[30018] = 8'b0;
    XRAM[30019] = 8'b0;
    XRAM[30020] = 8'b0;
    XRAM[30021] = 8'b0;
    XRAM[30022] = 8'b0;
    XRAM[30023] = 8'b0;
    XRAM[30024] = 8'b0;
    XRAM[30025] = 8'b0;
    XRAM[30026] = 8'b0;
    XRAM[30027] = 8'b0;
    XRAM[30028] = 8'b0;
    XRAM[30029] = 8'b0;
    XRAM[30030] = 8'b0;
    XRAM[30031] = 8'b0;
    XRAM[30032] = 8'b0;
    XRAM[30033] = 8'b0;
    XRAM[30034] = 8'b0;
    XRAM[30035] = 8'b0;
    XRAM[30036] = 8'b0;
    XRAM[30037] = 8'b0;
    XRAM[30038] = 8'b0;
    XRAM[30039] = 8'b0;
    XRAM[30040] = 8'b0;
    XRAM[30041] = 8'b0;
    XRAM[30042] = 8'b0;
    XRAM[30043] = 8'b0;
    XRAM[30044] = 8'b0;
    XRAM[30045] = 8'b0;
    XRAM[30046] = 8'b0;
    XRAM[30047] = 8'b0;
    XRAM[30048] = 8'b0;
    XRAM[30049] = 8'b0;
    XRAM[30050] = 8'b0;
    XRAM[30051] = 8'b0;
    XRAM[30052] = 8'b0;
    XRAM[30053] = 8'b0;
    XRAM[30054] = 8'b0;
    XRAM[30055] = 8'b0;
    XRAM[30056] = 8'b0;
    XRAM[30057] = 8'b0;
    XRAM[30058] = 8'b0;
    XRAM[30059] = 8'b0;
    XRAM[30060] = 8'b0;
    XRAM[30061] = 8'b0;
    XRAM[30062] = 8'b0;
    XRAM[30063] = 8'b0;
    XRAM[30064] = 8'b0;
    XRAM[30065] = 8'b0;
    XRAM[30066] = 8'b0;
    XRAM[30067] = 8'b0;
    XRAM[30068] = 8'b0;
    XRAM[30069] = 8'b0;
    XRAM[30070] = 8'b0;
    XRAM[30071] = 8'b0;
    XRAM[30072] = 8'b0;
    XRAM[30073] = 8'b0;
    XRAM[30074] = 8'b0;
    XRAM[30075] = 8'b0;
    XRAM[30076] = 8'b0;
    XRAM[30077] = 8'b0;
    XRAM[30078] = 8'b0;
    XRAM[30079] = 8'b0;
    XRAM[30080] = 8'b0;
    XRAM[30081] = 8'b0;
    XRAM[30082] = 8'b0;
    XRAM[30083] = 8'b0;
    XRAM[30084] = 8'b0;
    XRAM[30085] = 8'b0;
    XRAM[30086] = 8'b0;
    XRAM[30087] = 8'b0;
    XRAM[30088] = 8'b0;
    XRAM[30089] = 8'b0;
    XRAM[30090] = 8'b0;
    XRAM[30091] = 8'b0;
    XRAM[30092] = 8'b0;
    XRAM[30093] = 8'b0;
    XRAM[30094] = 8'b0;
    XRAM[30095] = 8'b0;
    XRAM[30096] = 8'b0;
    XRAM[30097] = 8'b0;
    XRAM[30098] = 8'b0;
    XRAM[30099] = 8'b0;
    XRAM[30100] = 8'b0;
    XRAM[30101] = 8'b0;
    XRAM[30102] = 8'b0;
    XRAM[30103] = 8'b0;
    XRAM[30104] = 8'b0;
    XRAM[30105] = 8'b0;
    XRAM[30106] = 8'b0;
    XRAM[30107] = 8'b0;
    XRAM[30108] = 8'b0;
    XRAM[30109] = 8'b0;
    XRAM[30110] = 8'b0;
    XRAM[30111] = 8'b0;
    XRAM[30112] = 8'b0;
    XRAM[30113] = 8'b0;
    XRAM[30114] = 8'b0;
    XRAM[30115] = 8'b0;
    XRAM[30116] = 8'b0;
    XRAM[30117] = 8'b0;
    XRAM[30118] = 8'b0;
    XRAM[30119] = 8'b0;
    XRAM[30120] = 8'b0;
    XRAM[30121] = 8'b0;
    XRAM[30122] = 8'b0;
    XRAM[30123] = 8'b0;
    XRAM[30124] = 8'b0;
    XRAM[30125] = 8'b0;
    XRAM[30126] = 8'b0;
    XRAM[30127] = 8'b0;
    XRAM[30128] = 8'b0;
    XRAM[30129] = 8'b0;
    XRAM[30130] = 8'b0;
    XRAM[30131] = 8'b0;
    XRAM[30132] = 8'b0;
    XRAM[30133] = 8'b0;
    XRAM[30134] = 8'b0;
    XRAM[30135] = 8'b0;
    XRAM[30136] = 8'b0;
    XRAM[30137] = 8'b0;
    XRAM[30138] = 8'b0;
    XRAM[30139] = 8'b0;
    XRAM[30140] = 8'b0;
    XRAM[30141] = 8'b0;
    XRAM[30142] = 8'b0;
    XRAM[30143] = 8'b0;
    XRAM[30144] = 8'b0;
    XRAM[30145] = 8'b0;
    XRAM[30146] = 8'b0;
    XRAM[30147] = 8'b0;
    XRAM[30148] = 8'b0;
    XRAM[30149] = 8'b0;
    XRAM[30150] = 8'b0;
    XRAM[30151] = 8'b0;
    XRAM[30152] = 8'b0;
    XRAM[30153] = 8'b0;
    XRAM[30154] = 8'b0;
    XRAM[30155] = 8'b0;
    XRAM[30156] = 8'b0;
    XRAM[30157] = 8'b0;
    XRAM[30158] = 8'b0;
    XRAM[30159] = 8'b0;
    XRAM[30160] = 8'b0;
    XRAM[30161] = 8'b0;
    XRAM[30162] = 8'b0;
    XRAM[30163] = 8'b0;
    XRAM[30164] = 8'b0;
    XRAM[30165] = 8'b0;
    XRAM[30166] = 8'b0;
    XRAM[30167] = 8'b0;
    XRAM[30168] = 8'b0;
    XRAM[30169] = 8'b0;
    XRAM[30170] = 8'b0;
    XRAM[30171] = 8'b0;
    XRAM[30172] = 8'b0;
    XRAM[30173] = 8'b0;
    XRAM[30174] = 8'b0;
    XRAM[30175] = 8'b0;
    XRAM[30176] = 8'b0;
    XRAM[30177] = 8'b0;
    XRAM[30178] = 8'b0;
    XRAM[30179] = 8'b0;
    XRAM[30180] = 8'b0;
    XRAM[30181] = 8'b0;
    XRAM[30182] = 8'b0;
    XRAM[30183] = 8'b0;
    XRAM[30184] = 8'b0;
    XRAM[30185] = 8'b0;
    XRAM[30186] = 8'b0;
    XRAM[30187] = 8'b0;
    XRAM[30188] = 8'b0;
    XRAM[30189] = 8'b0;
    XRAM[30190] = 8'b0;
    XRAM[30191] = 8'b0;
    XRAM[30192] = 8'b0;
    XRAM[30193] = 8'b0;
    XRAM[30194] = 8'b0;
    XRAM[30195] = 8'b0;
    XRAM[30196] = 8'b0;
    XRAM[30197] = 8'b0;
    XRAM[30198] = 8'b0;
    XRAM[30199] = 8'b0;
    XRAM[30200] = 8'b0;
    XRAM[30201] = 8'b0;
    XRAM[30202] = 8'b0;
    XRAM[30203] = 8'b0;
    XRAM[30204] = 8'b0;
    XRAM[30205] = 8'b0;
    XRAM[30206] = 8'b0;
    XRAM[30207] = 8'b0;
    XRAM[30208] = 8'b0;
    XRAM[30209] = 8'b0;
    XRAM[30210] = 8'b0;
    XRAM[30211] = 8'b0;
    XRAM[30212] = 8'b0;
    XRAM[30213] = 8'b0;
    XRAM[30214] = 8'b0;
    XRAM[30215] = 8'b0;
    XRAM[30216] = 8'b0;
    XRAM[30217] = 8'b0;
    XRAM[30218] = 8'b0;
    XRAM[30219] = 8'b0;
    XRAM[30220] = 8'b0;
    XRAM[30221] = 8'b0;
    XRAM[30222] = 8'b0;
    XRAM[30223] = 8'b0;
    XRAM[30224] = 8'b0;
    XRAM[30225] = 8'b0;
    XRAM[30226] = 8'b0;
    XRAM[30227] = 8'b0;
    XRAM[30228] = 8'b0;
    XRAM[30229] = 8'b0;
    XRAM[30230] = 8'b0;
    XRAM[30231] = 8'b0;
    XRAM[30232] = 8'b0;
    XRAM[30233] = 8'b0;
    XRAM[30234] = 8'b0;
    XRAM[30235] = 8'b0;
    XRAM[30236] = 8'b0;
    XRAM[30237] = 8'b0;
    XRAM[30238] = 8'b0;
    XRAM[30239] = 8'b0;
    XRAM[30240] = 8'b0;
    XRAM[30241] = 8'b0;
    XRAM[30242] = 8'b0;
    XRAM[30243] = 8'b0;
    XRAM[30244] = 8'b0;
    XRAM[30245] = 8'b0;
    XRAM[30246] = 8'b0;
    XRAM[30247] = 8'b0;
    XRAM[30248] = 8'b0;
    XRAM[30249] = 8'b0;
    XRAM[30250] = 8'b0;
    XRAM[30251] = 8'b0;
    XRAM[30252] = 8'b0;
    XRAM[30253] = 8'b0;
    XRAM[30254] = 8'b0;
    XRAM[30255] = 8'b0;
    XRAM[30256] = 8'b0;
    XRAM[30257] = 8'b0;
    XRAM[30258] = 8'b0;
    XRAM[30259] = 8'b0;
    XRAM[30260] = 8'b0;
    XRAM[30261] = 8'b0;
    XRAM[30262] = 8'b0;
    XRAM[30263] = 8'b0;
    XRAM[30264] = 8'b0;
    XRAM[30265] = 8'b0;
    XRAM[30266] = 8'b0;
    XRAM[30267] = 8'b0;
    XRAM[30268] = 8'b0;
    XRAM[30269] = 8'b0;
    XRAM[30270] = 8'b0;
    XRAM[30271] = 8'b0;
    XRAM[30272] = 8'b0;
    XRAM[30273] = 8'b0;
    XRAM[30274] = 8'b0;
    XRAM[30275] = 8'b0;
    XRAM[30276] = 8'b0;
    XRAM[30277] = 8'b0;
    XRAM[30278] = 8'b0;
    XRAM[30279] = 8'b0;
    XRAM[30280] = 8'b0;
    XRAM[30281] = 8'b0;
    XRAM[30282] = 8'b0;
    XRAM[30283] = 8'b0;
    XRAM[30284] = 8'b0;
    XRAM[30285] = 8'b0;
    XRAM[30286] = 8'b0;
    XRAM[30287] = 8'b0;
    XRAM[30288] = 8'b0;
    XRAM[30289] = 8'b0;
    XRAM[30290] = 8'b0;
    XRAM[30291] = 8'b0;
    XRAM[30292] = 8'b0;
    XRAM[30293] = 8'b0;
    XRAM[30294] = 8'b0;
    XRAM[30295] = 8'b0;
    XRAM[30296] = 8'b0;
    XRAM[30297] = 8'b0;
    XRAM[30298] = 8'b0;
    XRAM[30299] = 8'b0;
    XRAM[30300] = 8'b0;
    XRAM[30301] = 8'b0;
    XRAM[30302] = 8'b0;
    XRAM[30303] = 8'b0;
    XRAM[30304] = 8'b0;
    XRAM[30305] = 8'b0;
    XRAM[30306] = 8'b0;
    XRAM[30307] = 8'b0;
    XRAM[30308] = 8'b0;
    XRAM[30309] = 8'b0;
    XRAM[30310] = 8'b0;
    XRAM[30311] = 8'b0;
    XRAM[30312] = 8'b0;
    XRAM[30313] = 8'b0;
    XRAM[30314] = 8'b0;
    XRAM[30315] = 8'b0;
    XRAM[30316] = 8'b0;
    XRAM[30317] = 8'b0;
    XRAM[30318] = 8'b0;
    XRAM[30319] = 8'b0;
    XRAM[30320] = 8'b0;
    XRAM[30321] = 8'b0;
    XRAM[30322] = 8'b0;
    XRAM[30323] = 8'b0;
    XRAM[30324] = 8'b0;
    XRAM[30325] = 8'b0;
    XRAM[30326] = 8'b0;
    XRAM[30327] = 8'b0;
    XRAM[30328] = 8'b0;
    XRAM[30329] = 8'b0;
    XRAM[30330] = 8'b0;
    XRAM[30331] = 8'b0;
    XRAM[30332] = 8'b0;
    XRAM[30333] = 8'b0;
    XRAM[30334] = 8'b0;
    XRAM[30335] = 8'b0;
    XRAM[30336] = 8'b0;
    XRAM[30337] = 8'b0;
    XRAM[30338] = 8'b0;
    XRAM[30339] = 8'b0;
    XRAM[30340] = 8'b0;
    XRAM[30341] = 8'b0;
    XRAM[30342] = 8'b0;
    XRAM[30343] = 8'b0;
    XRAM[30344] = 8'b0;
    XRAM[30345] = 8'b0;
    XRAM[30346] = 8'b0;
    XRAM[30347] = 8'b0;
    XRAM[30348] = 8'b0;
    XRAM[30349] = 8'b0;
    XRAM[30350] = 8'b0;
    XRAM[30351] = 8'b0;
    XRAM[30352] = 8'b0;
    XRAM[30353] = 8'b0;
    XRAM[30354] = 8'b0;
    XRAM[30355] = 8'b0;
    XRAM[30356] = 8'b0;
    XRAM[30357] = 8'b0;
    XRAM[30358] = 8'b0;
    XRAM[30359] = 8'b0;
    XRAM[30360] = 8'b0;
    XRAM[30361] = 8'b0;
    XRAM[30362] = 8'b0;
    XRAM[30363] = 8'b0;
    XRAM[30364] = 8'b0;
    XRAM[30365] = 8'b0;
    XRAM[30366] = 8'b0;
    XRAM[30367] = 8'b0;
    XRAM[30368] = 8'b0;
    XRAM[30369] = 8'b0;
    XRAM[30370] = 8'b0;
    XRAM[30371] = 8'b0;
    XRAM[30372] = 8'b0;
    XRAM[30373] = 8'b0;
    XRAM[30374] = 8'b0;
    XRAM[30375] = 8'b0;
    XRAM[30376] = 8'b0;
    XRAM[30377] = 8'b0;
    XRAM[30378] = 8'b0;
    XRAM[30379] = 8'b0;
    XRAM[30380] = 8'b0;
    XRAM[30381] = 8'b0;
    XRAM[30382] = 8'b0;
    XRAM[30383] = 8'b0;
    XRAM[30384] = 8'b0;
    XRAM[30385] = 8'b0;
    XRAM[30386] = 8'b0;
    XRAM[30387] = 8'b0;
    XRAM[30388] = 8'b0;
    XRAM[30389] = 8'b0;
    XRAM[30390] = 8'b0;
    XRAM[30391] = 8'b0;
    XRAM[30392] = 8'b0;
    XRAM[30393] = 8'b0;
    XRAM[30394] = 8'b0;
    XRAM[30395] = 8'b0;
    XRAM[30396] = 8'b0;
    XRAM[30397] = 8'b0;
    XRAM[30398] = 8'b0;
    XRAM[30399] = 8'b0;
    XRAM[30400] = 8'b0;
    XRAM[30401] = 8'b0;
    XRAM[30402] = 8'b0;
    XRAM[30403] = 8'b0;
    XRAM[30404] = 8'b0;
    XRAM[30405] = 8'b0;
    XRAM[30406] = 8'b0;
    XRAM[30407] = 8'b0;
    XRAM[30408] = 8'b0;
    XRAM[30409] = 8'b0;
    XRAM[30410] = 8'b0;
    XRAM[30411] = 8'b0;
    XRAM[30412] = 8'b0;
    XRAM[30413] = 8'b0;
    XRAM[30414] = 8'b0;
    XRAM[30415] = 8'b0;
    XRAM[30416] = 8'b0;
    XRAM[30417] = 8'b0;
    XRAM[30418] = 8'b0;
    XRAM[30419] = 8'b0;
    XRAM[30420] = 8'b0;
    XRAM[30421] = 8'b0;
    XRAM[30422] = 8'b0;
    XRAM[30423] = 8'b0;
    XRAM[30424] = 8'b0;
    XRAM[30425] = 8'b0;
    XRAM[30426] = 8'b0;
    XRAM[30427] = 8'b0;
    XRAM[30428] = 8'b0;
    XRAM[30429] = 8'b0;
    XRAM[30430] = 8'b0;
    XRAM[30431] = 8'b0;
    XRAM[30432] = 8'b0;
    XRAM[30433] = 8'b0;
    XRAM[30434] = 8'b0;
    XRAM[30435] = 8'b0;
    XRAM[30436] = 8'b0;
    XRAM[30437] = 8'b0;
    XRAM[30438] = 8'b0;
    XRAM[30439] = 8'b0;
    XRAM[30440] = 8'b0;
    XRAM[30441] = 8'b0;
    XRAM[30442] = 8'b0;
    XRAM[30443] = 8'b0;
    XRAM[30444] = 8'b0;
    XRAM[30445] = 8'b0;
    XRAM[30446] = 8'b0;
    XRAM[30447] = 8'b0;
    XRAM[30448] = 8'b0;
    XRAM[30449] = 8'b0;
    XRAM[30450] = 8'b0;
    XRAM[30451] = 8'b0;
    XRAM[30452] = 8'b0;
    XRAM[30453] = 8'b0;
    XRAM[30454] = 8'b0;
    XRAM[30455] = 8'b0;
    XRAM[30456] = 8'b0;
    XRAM[30457] = 8'b0;
    XRAM[30458] = 8'b0;
    XRAM[30459] = 8'b0;
    XRAM[30460] = 8'b0;
    XRAM[30461] = 8'b0;
    XRAM[30462] = 8'b0;
    XRAM[30463] = 8'b0;
    XRAM[30464] = 8'b0;
    XRAM[30465] = 8'b0;
    XRAM[30466] = 8'b0;
    XRAM[30467] = 8'b0;
    XRAM[30468] = 8'b0;
    XRAM[30469] = 8'b0;
    XRAM[30470] = 8'b0;
    XRAM[30471] = 8'b0;
    XRAM[30472] = 8'b0;
    XRAM[30473] = 8'b0;
    XRAM[30474] = 8'b0;
    XRAM[30475] = 8'b0;
    XRAM[30476] = 8'b0;
    XRAM[30477] = 8'b0;
    XRAM[30478] = 8'b0;
    XRAM[30479] = 8'b0;
    XRAM[30480] = 8'b0;
    XRAM[30481] = 8'b0;
    XRAM[30482] = 8'b0;
    XRAM[30483] = 8'b0;
    XRAM[30484] = 8'b0;
    XRAM[30485] = 8'b0;
    XRAM[30486] = 8'b0;
    XRAM[30487] = 8'b0;
    XRAM[30488] = 8'b0;
    XRAM[30489] = 8'b0;
    XRAM[30490] = 8'b0;
    XRAM[30491] = 8'b0;
    XRAM[30492] = 8'b0;
    XRAM[30493] = 8'b0;
    XRAM[30494] = 8'b0;
    XRAM[30495] = 8'b0;
    XRAM[30496] = 8'b0;
    XRAM[30497] = 8'b0;
    XRAM[30498] = 8'b0;
    XRAM[30499] = 8'b0;
    XRAM[30500] = 8'b0;
    XRAM[30501] = 8'b0;
    XRAM[30502] = 8'b0;
    XRAM[30503] = 8'b0;
    XRAM[30504] = 8'b0;
    XRAM[30505] = 8'b0;
    XRAM[30506] = 8'b0;
    XRAM[30507] = 8'b0;
    XRAM[30508] = 8'b0;
    XRAM[30509] = 8'b0;
    XRAM[30510] = 8'b0;
    XRAM[30511] = 8'b0;
    XRAM[30512] = 8'b0;
    XRAM[30513] = 8'b0;
    XRAM[30514] = 8'b0;
    XRAM[30515] = 8'b0;
    XRAM[30516] = 8'b0;
    XRAM[30517] = 8'b0;
    XRAM[30518] = 8'b0;
    XRAM[30519] = 8'b0;
    XRAM[30520] = 8'b0;
    XRAM[30521] = 8'b0;
    XRAM[30522] = 8'b0;
    XRAM[30523] = 8'b0;
    XRAM[30524] = 8'b0;
    XRAM[30525] = 8'b0;
    XRAM[30526] = 8'b0;
    XRAM[30527] = 8'b0;
    XRAM[30528] = 8'b0;
    XRAM[30529] = 8'b0;
    XRAM[30530] = 8'b0;
    XRAM[30531] = 8'b0;
    XRAM[30532] = 8'b0;
    XRAM[30533] = 8'b0;
    XRAM[30534] = 8'b0;
    XRAM[30535] = 8'b0;
    XRAM[30536] = 8'b0;
    XRAM[30537] = 8'b0;
    XRAM[30538] = 8'b0;
    XRAM[30539] = 8'b0;
    XRAM[30540] = 8'b0;
    XRAM[30541] = 8'b0;
    XRAM[30542] = 8'b0;
    XRAM[30543] = 8'b0;
    XRAM[30544] = 8'b0;
    XRAM[30545] = 8'b0;
    XRAM[30546] = 8'b0;
    XRAM[30547] = 8'b0;
    XRAM[30548] = 8'b0;
    XRAM[30549] = 8'b0;
    XRAM[30550] = 8'b0;
    XRAM[30551] = 8'b0;
    XRAM[30552] = 8'b0;
    XRAM[30553] = 8'b0;
    XRAM[30554] = 8'b0;
    XRAM[30555] = 8'b0;
    XRAM[30556] = 8'b0;
    XRAM[30557] = 8'b0;
    XRAM[30558] = 8'b0;
    XRAM[30559] = 8'b0;
    XRAM[30560] = 8'b0;
    XRAM[30561] = 8'b0;
    XRAM[30562] = 8'b0;
    XRAM[30563] = 8'b0;
    XRAM[30564] = 8'b0;
    XRAM[30565] = 8'b0;
    XRAM[30566] = 8'b0;
    XRAM[30567] = 8'b0;
    XRAM[30568] = 8'b0;
    XRAM[30569] = 8'b0;
    XRAM[30570] = 8'b0;
    XRAM[30571] = 8'b0;
    XRAM[30572] = 8'b0;
    XRAM[30573] = 8'b0;
    XRAM[30574] = 8'b0;
    XRAM[30575] = 8'b0;
    XRAM[30576] = 8'b0;
    XRAM[30577] = 8'b0;
    XRAM[30578] = 8'b0;
    XRAM[30579] = 8'b0;
    XRAM[30580] = 8'b0;
    XRAM[30581] = 8'b0;
    XRAM[30582] = 8'b0;
    XRAM[30583] = 8'b0;
    XRAM[30584] = 8'b0;
    XRAM[30585] = 8'b0;
    XRAM[30586] = 8'b0;
    XRAM[30587] = 8'b0;
    XRAM[30588] = 8'b0;
    XRAM[30589] = 8'b0;
    XRAM[30590] = 8'b0;
    XRAM[30591] = 8'b0;
    XRAM[30592] = 8'b0;
    XRAM[30593] = 8'b0;
    XRAM[30594] = 8'b0;
    XRAM[30595] = 8'b0;
    XRAM[30596] = 8'b0;
    XRAM[30597] = 8'b0;
    XRAM[30598] = 8'b0;
    XRAM[30599] = 8'b0;
    XRAM[30600] = 8'b0;
    XRAM[30601] = 8'b0;
    XRAM[30602] = 8'b0;
    XRAM[30603] = 8'b0;
    XRAM[30604] = 8'b0;
    XRAM[30605] = 8'b0;
    XRAM[30606] = 8'b0;
    XRAM[30607] = 8'b0;
    XRAM[30608] = 8'b0;
    XRAM[30609] = 8'b0;
    XRAM[30610] = 8'b0;
    XRAM[30611] = 8'b0;
    XRAM[30612] = 8'b0;
    XRAM[30613] = 8'b0;
    XRAM[30614] = 8'b0;
    XRAM[30615] = 8'b0;
    XRAM[30616] = 8'b0;
    XRAM[30617] = 8'b0;
    XRAM[30618] = 8'b0;
    XRAM[30619] = 8'b0;
    XRAM[30620] = 8'b0;
    XRAM[30621] = 8'b0;
    XRAM[30622] = 8'b0;
    XRAM[30623] = 8'b0;
    XRAM[30624] = 8'b0;
    XRAM[30625] = 8'b0;
    XRAM[30626] = 8'b0;
    XRAM[30627] = 8'b0;
    XRAM[30628] = 8'b0;
    XRAM[30629] = 8'b0;
    XRAM[30630] = 8'b0;
    XRAM[30631] = 8'b0;
    XRAM[30632] = 8'b0;
    XRAM[30633] = 8'b0;
    XRAM[30634] = 8'b0;
    XRAM[30635] = 8'b0;
    XRAM[30636] = 8'b0;
    XRAM[30637] = 8'b0;
    XRAM[30638] = 8'b0;
    XRAM[30639] = 8'b0;
    XRAM[30640] = 8'b0;
    XRAM[30641] = 8'b0;
    XRAM[30642] = 8'b0;
    XRAM[30643] = 8'b0;
    XRAM[30644] = 8'b0;
    XRAM[30645] = 8'b0;
    XRAM[30646] = 8'b0;
    XRAM[30647] = 8'b0;
    XRAM[30648] = 8'b0;
    XRAM[30649] = 8'b0;
    XRAM[30650] = 8'b0;
    XRAM[30651] = 8'b0;
    XRAM[30652] = 8'b0;
    XRAM[30653] = 8'b0;
    XRAM[30654] = 8'b0;
    XRAM[30655] = 8'b0;
    XRAM[30656] = 8'b0;
    XRAM[30657] = 8'b0;
    XRAM[30658] = 8'b0;
    XRAM[30659] = 8'b0;
    XRAM[30660] = 8'b0;
    XRAM[30661] = 8'b0;
    XRAM[30662] = 8'b0;
    XRAM[30663] = 8'b0;
    XRAM[30664] = 8'b0;
    XRAM[30665] = 8'b0;
    XRAM[30666] = 8'b0;
    XRAM[30667] = 8'b0;
    XRAM[30668] = 8'b0;
    XRAM[30669] = 8'b0;
    XRAM[30670] = 8'b0;
    XRAM[30671] = 8'b0;
    XRAM[30672] = 8'b0;
    XRAM[30673] = 8'b0;
    XRAM[30674] = 8'b0;
    XRAM[30675] = 8'b0;
    XRAM[30676] = 8'b0;
    XRAM[30677] = 8'b0;
    XRAM[30678] = 8'b0;
    XRAM[30679] = 8'b0;
    XRAM[30680] = 8'b0;
    XRAM[30681] = 8'b0;
    XRAM[30682] = 8'b0;
    XRAM[30683] = 8'b0;
    XRAM[30684] = 8'b0;
    XRAM[30685] = 8'b0;
    XRAM[30686] = 8'b0;
    XRAM[30687] = 8'b0;
    XRAM[30688] = 8'b0;
    XRAM[30689] = 8'b0;
    XRAM[30690] = 8'b0;
    XRAM[30691] = 8'b0;
    XRAM[30692] = 8'b0;
    XRAM[30693] = 8'b0;
    XRAM[30694] = 8'b0;
    XRAM[30695] = 8'b0;
    XRAM[30696] = 8'b0;
    XRAM[30697] = 8'b0;
    XRAM[30698] = 8'b0;
    XRAM[30699] = 8'b0;
    XRAM[30700] = 8'b0;
    XRAM[30701] = 8'b0;
    XRAM[30702] = 8'b0;
    XRAM[30703] = 8'b0;
    XRAM[30704] = 8'b0;
    XRAM[30705] = 8'b0;
    XRAM[30706] = 8'b0;
    XRAM[30707] = 8'b0;
    XRAM[30708] = 8'b0;
    XRAM[30709] = 8'b0;
    XRAM[30710] = 8'b0;
    XRAM[30711] = 8'b0;
    XRAM[30712] = 8'b0;
    XRAM[30713] = 8'b0;
    XRAM[30714] = 8'b0;
    XRAM[30715] = 8'b0;
    XRAM[30716] = 8'b0;
    XRAM[30717] = 8'b0;
    XRAM[30718] = 8'b0;
    XRAM[30719] = 8'b0;
    XRAM[30720] = 8'b0;
    XRAM[30721] = 8'b0;
    XRAM[30722] = 8'b0;
    XRAM[30723] = 8'b0;
    XRAM[30724] = 8'b0;
    XRAM[30725] = 8'b0;
    XRAM[30726] = 8'b0;
    XRAM[30727] = 8'b0;
    XRAM[30728] = 8'b0;
    XRAM[30729] = 8'b0;
    XRAM[30730] = 8'b0;
    XRAM[30731] = 8'b0;
    XRAM[30732] = 8'b0;
    XRAM[30733] = 8'b0;
    XRAM[30734] = 8'b0;
    XRAM[30735] = 8'b0;
    XRAM[30736] = 8'b0;
    XRAM[30737] = 8'b0;
    XRAM[30738] = 8'b0;
    XRAM[30739] = 8'b0;
    XRAM[30740] = 8'b0;
    XRAM[30741] = 8'b0;
    XRAM[30742] = 8'b0;
    XRAM[30743] = 8'b0;
    XRAM[30744] = 8'b0;
    XRAM[30745] = 8'b0;
    XRAM[30746] = 8'b0;
    XRAM[30747] = 8'b0;
    XRAM[30748] = 8'b0;
    XRAM[30749] = 8'b0;
    XRAM[30750] = 8'b0;
    XRAM[30751] = 8'b0;
    XRAM[30752] = 8'b0;
    XRAM[30753] = 8'b0;
    XRAM[30754] = 8'b0;
    XRAM[30755] = 8'b0;
    XRAM[30756] = 8'b0;
    XRAM[30757] = 8'b0;
    XRAM[30758] = 8'b0;
    XRAM[30759] = 8'b0;
    XRAM[30760] = 8'b0;
    XRAM[30761] = 8'b0;
    XRAM[30762] = 8'b0;
    XRAM[30763] = 8'b0;
    XRAM[30764] = 8'b0;
    XRAM[30765] = 8'b0;
    XRAM[30766] = 8'b0;
    XRAM[30767] = 8'b0;
    XRAM[30768] = 8'b0;
    XRAM[30769] = 8'b0;
    XRAM[30770] = 8'b0;
    XRAM[30771] = 8'b0;
    XRAM[30772] = 8'b0;
    XRAM[30773] = 8'b0;
    XRAM[30774] = 8'b0;
    XRAM[30775] = 8'b0;
    XRAM[30776] = 8'b0;
    XRAM[30777] = 8'b0;
    XRAM[30778] = 8'b0;
    XRAM[30779] = 8'b0;
    XRAM[30780] = 8'b0;
    XRAM[30781] = 8'b0;
    XRAM[30782] = 8'b0;
    XRAM[30783] = 8'b0;
    XRAM[30784] = 8'b0;
    XRAM[30785] = 8'b0;
    XRAM[30786] = 8'b0;
    XRAM[30787] = 8'b0;
    XRAM[30788] = 8'b0;
    XRAM[30789] = 8'b0;
    XRAM[30790] = 8'b0;
    XRAM[30791] = 8'b0;
    XRAM[30792] = 8'b0;
    XRAM[30793] = 8'b0;
    XRAM[30794] = 8'b0;
    XRAM[30795] = 8'b0;
    XRAM[30796] = 8'b0;
    XRAM[30797] = 8'b0;
    XRAM[30798] = 8'b0;
    XRAM[30799] = 8'b0;
    XRAM[30800] = 8'b0;
    XRAM[30801] = 8'b0;
    XRAM[30802] = 8'b0;
    XRAM[30803] = 8'b0;
    XRAM[30804] = 8'b0;
    XRAM[30805] = 8'b0;
    XRAM[30806] = 8'b0;
    XRAM[30807] = 8'b0;
    XRAM[30808] = 8'b0;
    XRAM[30809] = 8'b0;
    XRAM[30810] = 8'b0;
    XRAM[30811] = 8'b0;
    XRAM[30812] = 8'b0;
    XRAM[30813] = 8'b0;
    XRAM[30814] = 8'b0;
    XRAM[30815] = 8'b0;
    XRAM[30816] = 8'b0;
    XRAM[30817] = 8'b0;
    XRAM[30818] = 8'b0;
    XRAM[30819] = 8'b0;
    XRAM[30820] = 8'b0;
    XRAM[30821] = 8'b0;
    XRAM[30822] = 8'b0;
    XRAM[30823] = 8'b0;
    XRAM[30824] = 8'b0;
    XRAM[30825] = 8'b0;
    XRAM[30826] = 8'b0;
    XRAM[30827] = 8'b0;
    XRAM[30828] = 8'b0;
    XRAM[30829] = 8'b0;
    XRAM[30830] = 8'b0;
    XRAM[30831] = 8'b0;
    XRAM[30832] = 8'b0;
    XRAM[30833] = 8'b0;
    XRAM[30834] = 8'b0;
    XRAM[30835] = 8'b0;
    XRAM[30836] = 8'b0;
    XRAM[30837] = 8'b0;
    XRAM[30838] = 8'b0;
    XRAM[30839] = 8'b0;
    XRAM[30840] = 8'b0;
    XRAM[30841] = 8'b0;
    XRAM[30842] = 8'b0;
    XRAM[30843] = 8'b0;
    XRAM[30844] = 8'b0;
    XRAM[30845] = 8'b0;
    XRAM[30846] = 8'b0;
    XRAM[30847] = 8'b0;
    XRAM[30848] = 8'b0;
    XRAM[30849] = 8'b0;
    XRAM[30850] = 8'b0;
    XRAM[30851] = 8'b0;
    XRAM[30852] = 8'b0;
    XRAM[30853] = 8'b0;
    XRAM[30854] = 8'b0;
    XRAM[30855] = 8'b0;
    XRAM[30856] = 8'b0;
    XRAM[30857] = 8'b0;
    XRAM[30858] = 8'b0;
    XRAM[30859] = 8'b0;
    XRAM[30860] = 8'b0;
    XRAM[30861] = 8'b0;
    XRAM[30862] = 8'b0;
    XRAM[30863] = 8'b0;
    XRAM[30864] = 8'b0;
    XRAM[30865] = 8'b0;
    XRAM[30866] = 8'b0;
    XRAM[30867] = 8'b0;
    XRAM[30868] = 8'b0;
    XRAM[30869] = 8'b0;
    XRAM[30870] = 8'b0;
    XRAM[30871] = 8'b0;
    XRAM[30872] = 8'b0;
    XRAM[30873] = 8'b0;
    XRAM[30874] = 8'b0;
    XRAM[30875] = 8'b0;
    XRAM[30876] = 8'b0;
    XRAM[30877] = 8'b0;
    XRAM[30878] = 8'b0;
    XRAM[30879] = 8'b0;
    XRAM[30880] = 8'b0;
    XRAM[30881] = 8'b0;
    XRAM[30882] = 8'b0;
    XRAM[30883] = 8'b0;
    XRAM[30884] = 8'b0;
    XRAM[30885] = 8'b0;
    XRAM[30886] = 8'b0;
    XRAM[30887] = 8'b0;
    XRAM[30888] = 8'b0;
    XRAM[30889] = 8'b0;
    XRAM[30890] = 8'b0;
    XRAM[30891] = 8'b0;
    XRAM[30892] = 8'b0;
    XRAM[30893] = 8'b0;
    XRAM[30894] = 8'b0;
    XRAM[30895] = 8'b0;
    XRAM[30896] = 8'b0;
    XRAM[30897] = 8'b0;
    XRAM[30898] = 8'b0;
    XRAM[30899] = 8'b0;
    XRAM[30900] = 8'b0;
    XRAM[30901] = 8'b0;
    XRAM[30902] = 8'b0;
    XRAM[30903] = 8'b0;
    XRAM[30904] = 8'b0;
    XRAM[30905] = 8'b0;
    XRAM[30906] = 8'b0;
    XRAM[30907] = 8'b0;
    XRAM[30908] = 8'b0;
    XRAM[30909] = 8'b0;
    XRAM[30910] = 8'b0;
    XRAM[30911] = 8'b0;
    XRAM[30912] = 8'b0;
    XRAM[30913] = 8'b0;
    XRAM[30914] = 8'b0;
    XRAM[30915] = 8'b0;
    XRAM[30916] = 8'b0;
    XRAM[30917] = 8'b0;
    XRAM[30918] = 8'b0;
    XRAM[30919] = 8'b0;
    XRAM[30920] = 8'b0;
    XRAM[30921] = 8'b0;
    XRAM[30922] = 8'b0;
    XRAM[30923] = 8'b0;
    XRAM[30924] = 8'b0;
    XRAM[30925] = 8'b0;
    XRAM[30926] = 8'b0;
    XRAM[30927] = 8'b0;
    XRAM[30928] = 8'b0;
    XRAM[30929] = 8'b0;
    XRAM[30930] = 8'b0;
    XRAM[30931] = 8'b0;
    XRAM[30932] = 8'b0;
    XRAM[30933] = 8'b0;
    XRAM[30934] = 8'b0;
    XRAM[30935] = 8'b0;
    XRAM[30936] = 8'b0;
    XRAM[30937] = 8'b0;
    XRAM[30938] = 8'b0;
    XRAM[30939] = 8'b0;
    XRAM[30940] = 8'b0;
    XRAM[30941] = 8'b0;
    XRAM[30942] = 8'b0;
    XRAM[30943] = 8'b0;
    XRAM[30944] = 8'b0;
    XRAM[30945] = 8'b0;
    XRAM[30946] = 8'b0;
    XRAM[30947] = 8'b0;
    XRAM[30948] = 8'b0;
    XRAM[30949] = 8'b0;
    XRAM[30950] = 8'b0;
    XRAM[30951] = 8'b0;
    XRAM[30952] = 8'b0;
    XRAM[30953] = 8'b0;
    XRAM[30954] = 8'b0;
    XRAM[30955] = 8'b0;
    XRAM[30956] = 8'b0;
    XRAM[30957] = 8'b0;
    XRAM[30958] = 8'b0;
    XRAM[30959] = 8'b0;
    XRAM[30960] = 8'b0;
    XRAM[30961] = 8'b0;
    XRAM[30962] = 8'b0;
    XRAM[30963] = 8'b0;
    XRAM[30964] = 8'b0;
    XRAM[30965] = 8'b0;
    XRAM[30966] = 8'b0;
    XRAM[30967] = 8'b0;
    XRAM[30968] = 8'b0;
    XRAM[30969] = 8'b0;
    XRAM[30970] = 8'b0;
    XRAM[30971] = 8'b0;
    XRAM[30972] = 8'b0;
    XRAM[30973] = 8'b0;
    XRAM[30974] = 8'b0;
    XRAM[30975] = 8'b0;
    XRAM[30976] = 8'b0;
    XRAM[30977] = 8'b0;
    XRAM[30978] = 8'b0;
    XRAM[30979] = 8'b0;
    XRAM[30980] = 8'b0;
    XRAM[30981] = 8'b0;
    XRAM[30982] = 8'b0;
    XRAM[30983] = 8'b0;
    XRAM[30984] = 8'b0;
    XRAM[30985] = 8'b0;
    XRAM[30986] = 8'b0;
    XRAM[30987] = 8'b0;
    XRAM[30988] = 8'b0;
    XRAM[30989] = 8'b0;
    XRAM[30990] = 8'b0;
    XRAM[30991] = 8'b0;
    XRAM[30992] = 8'b0;
    XRAM[30993] = 8'b0;
    XRAM[30994] = 8'b0;
    XRAM[30995] = 8'b0;
    XRAM[30996] = 8'b0;
    XRAM[30997] = 8'b0;
    XRAM[30998] = 8'b0;
    XRAM[30999] = 8'b0;
    XRAM[31000] = 8'b0;
    XRAM[31001] = 8'b0;
    XRAM[31002] = 8'b0;
    XRAM[31003] = 8'b0;
    XRAM[31004] = 8'b0;
    XRAM[31005] = 8'b0;
    XRAM[31006] = 8'b0;
    XRAM[31007] = 8'b0;
    XRAM[31008] = 8'b0;
    XRAM[31009] = 8'b0;
    XRAM[31010] = 8'b0;
    XRAM[31011] = 8'b0;
    XRAM[31012] = 8'b0;
    XRAM[31013] = 8'b0;
    XRAM[31014] = 8'b0;
    XRAM[31015] = 8'b0;
    XRAM[31016] = 8'b0;
    XRAM[31017] = 8'b0;
    XRAM[31018] = 8'b0;
    XRAM[31019] = 8'b0;
    XRAM[31020] = 8'b0;
    XRAM[31021] = 8'b0;
    XRAM[31022] = 8'b0;
    XRAM[31023] = 8'b0;
    XRAM[31024] = 8'b0;
    XRAM[31025] = 8'b0;
    XRAM[31026] = 8'b0;
    XRAM[31027] = 8'b0;
    XRAM[31028] = 8'b0;
    XRAM[31029] = 8'b0;
    XRAM[31030] = 8'b0;
    XRAM[31031] = 8'b0;
    XRAM[31032] = 8'b0;
    XRAM[31033] = 8'b0;
    XRAM[31034] = 8'b0;
    XRAM[31035] = 8'b0;
    XRAM[31036] = 8'b0;
    XRAM[31037] = 8'b0;
    XRAM[31038] = 8'b0;
    XRAM[31039] = 8'b0;
    XRAM[31040] = 8'b0;
    XRAM[31041] = 8'b0;
    XRAM[31042] = 8'b0;
    XRAM[31043] = 8'b0;
    XRAM[31044] = 8'b0;
    XRAM[31045] = 8'b0;
    XRAM[31046] = 8'b0;
    XRAM[31047] = 8'b0;
    XRAM[31048] = 8'b0;
    XRAM[31049] = 8'b0;
    XRAM[31050] = 8'b0;
    XRAM[31051] = 8'b0;
    XRAM[31052] = 8'b0;
    XRAM[31053] = 8'b0;
    XRAM[31054] = 8'b0;
    XRAM[31055] = 8'b0;
    XRAM[31056] = 8'b0;
    XRAM[31057] = 8'b0;
    XRAM[31058] = 8'b0;
    XRAM[31059] = 8'b0;
    XRAM[31060] = 8'b0;
    XRAM[31061] = 8'b0;
    XRAM[31062] = 8'b0;
    XRAM[31063] = 8'b0;
    XRAM[31064] = 8'b0;
    XRAM[31065] = 8'b0;
    XRAM[31066] = 8'b0;
    XRAM[31067] = 8'b0;
    XRAM[31068] = 8'b0;
    XRAM[31069] = 8'b0;
    XRAM[31070] = 8'b0;
    XRAM[31071] = 8'b0;
    XRAM[31072] = 8'b0;
    XRAM[31073] = 8'b0;
    XRAM[31074] = 8'b0;
    XRAM[31075] = 8'b0;
    XRAM[31076] = 8'b0;
    XRAM[31077] = 8'b0;
    XRAM[31078] = 8'b0;
    XRAM[31079] = 8'b0;
    XRAM[31080] = 8'b0;
    XRAM[31081] = 8'b0;
    XRAM[31082] = 8'b0;
    XRAM[31083] = 8'b0;
    XRAM[31084] = 8'b0;
    XRAM[31085] = 8'b0;
    XRAM[31086] = 8'b0;
    XRAM[31087] = 8'b0;
    XRAM[31088] = 8'b0;
    XRAM[31089] = 8'b0;
    XRAM[31090] = 8'b0;
    XRAM[31091] = 8'b0;
    XRAM[31092] = 8'b0;
    XRAM[31093] = 8'b0;
    XRAM[31094] = 8'b0;
    XRAM[31095] = 8'b0;
    XRAM[31096] = 8'b0;
    XRAM[31097] = 8'b0;
    XRAM[31098] = 8'b0;
    XRAM[31099] = 8'b0;
    XRAM[31100] = 8'b0;
    XRAM[31101] = 8'b0;
    XRAM[31102] = 8'b0;
    XRAM[31103] = 8'b0;
    XRAM[31104] = 8'b0;
    XRAM[31105] = 8'b0;
    XRAM[31106] = 8'b0;
    XRAM[31107] = 8'b0;
    XRAM[31108] = 8'b0;
    XRAM[31109] = 8'b0;
    XRAM[31110] = 8'b0;
    XRAM[31111] = 8'b0;
    XRAM[31112] = 8'b0;
    XRAM[31113] = 8'b0;
    XRAM[31114] = 8'b0;
    XRAM[31115] = 8'b0;
    XRAM[31116] = 8'b0;
    XRAM[31117] = 8'b0;
    XRAM[31118] = 8'b0;
    XRAM[31119] = 8'b0;
    XRAM[31120] = 8'b0;
    XRAM[31121] = 8'b0;
    XRAM[31122] = 8'b0;
    XRAM[31123] = 8'b0;
    XRAM[31124] = 8'b0;
    XRAM[31125] = 8'b0;
    XRAM[31126] = 8'b0;
    XRAM[31127] = 8'b0;
    XRAM[31128] = 8'b0;
    XRAM[31129] = 8'b0;
    XRAM[31130] = 8'b0;
    XRAM[31131] = 8'b0;
    XRAM[31132] = 8'b0;
    XRAM[31133] = 8'b0;
    XRAM[31134] = 8'b0;
    XRAM[31135] = 8'b0;
    XRAM[31136] = 8'b0;
    XRAM[31137] = 8'b0;
    XRAM[31138] = 8'b0;
    XRAM[31139] = 8'b0;
    XRAM[31140] = 8'b0;
    XRAM[31141] = 8'b0;
    XRAM[31142] = 8'b0;
    XRAM[31143] = 8'b0;
    XRAM[31144] = 8'b0;
    XRAM[31145] = 8'b0;
    XRAM[31146] = 8'b0;
    XRAM[31147] = 8'b0;
    XRAM[31148] = 8'b0;
    XRAM[31149] = 8'b0;
    XRAM[31150] = 8'b0;
    XRAM[31151] = 8'b0;
    XRAM[31152] = 8'b0;
    XRAM[31153] = 8'b0;
    XRAM[31154] = 8'b0;
    XRAM[31155] = 8'b0;
    XRAM[31156] = 8'b0;
    XRAM[31157] = 8'b0;
    XRAM[31158] = 8'b0;
    XRAM[31159] = 8'b0;
    XRAM[31160] = 8'b0;
    XRAM[31161] = 8'b0;
    XRAM[31162] = 8'b0;
    XRAM[31163] = 8'b0;
    XRAM[31164] = 8'b0;
    XRAM[31165] = 8'b0;
    XRAM[31166] = 8'b0;
    XRAM[31167] = 8'b0;
    XRAM[31168] = 8'b0;
    XRAM[31169] = 8'b0;
    XRAM[31170] = 8'b0;
    XRAM[31171] = 8'b0;
    XRAM[31172] = 8'b0;
    XRAM[31173] = 8'b0;
    XRAM[31174] = 8'b0;
    XRAM[31175] = 8'b0;
    XRAM[31176] = 8'b0;
    XRAM[31177] = 8'b0;
    XRAM[31178] = 8'b0;
    XRAM[31179] = 8'b0;
    XRAM[31180] = 8'b0;
    XRAM[31181] = 8'b0;
    XRAM[31182] = 8'b0;
    XRAM[31183] = 8'b0;
    XRAM[31184] = 8'b0;
    XRAM[31185] = 8'b0;
    XRAM[31186] = 8'b0;
    XRAM[31187] = 8'b0;
    XRAM[31188] = 8'b0;
    XRAM[31189] = 8'b0;
    XRAM[31190] = 8'b0;
    XRAM[31191] = 8'b0;
    XRAM[31192] = 8'b0;
    XRAM[31193] = 8'b0;
    XRAM[31194] = 8'b0;
    XRAM[31195] = 8'b0;
    XRAM[31196] = 8'b0;
    XRAM[31197] = 8'b0;
    XRAM[31198] = 8'b0;
    XRAM[31199] = 8'b0;
    XRAM[31200] = 8'b0;
    XRAM[31201] = 8'b0;
    XRAM[31202] = 8'b0;
    XRAM[31203] = 8'b0;
    XRAM[31204] = 8'b0;
    XRAM[31205] = 8'b0;
    XRAM[31206] = 8'b0;
    XRAM[31207] = 8'b0;
    XRAM[31208] = 8'b0;
    XRAM[31209] = 8'b0;
    XRAM[31210] = 8'b0;
    XRAM[31211] = 8'b0;
    XRAM[31212] = 8'b0;
    XRAM[31213] = 8'b0;
    XRAM[31214] = 8'b0;
    XRAM[31215] = 8'b0;
    XRAM[31216] = 8'b0;
    XRAM[31217] = 8'b0;
    XRAM[31218] = 8'b0;
    XRAM[31219] = 8'b0;
    XRAM[31220] = 8'b0;
    XRAM[31221] = 8'b0;
    XRAM[31222] = 8'b0;
    XRAM[31223] = 8'b0;
    XRAM[31224] = 8'b0;
    XRAM[31225] = 8'b0;
    XRAM[31226] = 8'b0;
    XRAM[31227] = 8'b0;
    XRAM[31228] = 8'b0;
    XRAM[31229] = 8'b0;
    XRAM[31230] = 8'b0;
    XRAM[31231] = 8'b0;
    XRAM[31232] = 8'b0;
    XRAM[31233] = 8'b0;
    XRAM[31234] = 8'b0;
    XRAM[31235] = 8'b0;
    XRAM[31236] = 8'b0;
    XRAM[31237] = 8'b0;
    XRAM[31238] = 8'b0;
    XRAM[31239] = 8'b0;
    XRAM[31240] = 8'b0;
    XRAM[31241] = 8'b0;
    XRAM[31242] = 8'b0;
    XRAM[31243] = 8'b0;
    XRAM[31244] = 8'b0;
    XRAM[31245] = 8'b0;
    XRAM[31246] = 8'b0;
    XRAM[31247] = 8'b0;
    XRAM[31248] = 8'b0;
    XRAM[31249] = 8'b0;
    XRAM[31250] = 8'b0;
    XRAM[31251] = 8'b0;
    XRAM[31252] = 8'b0;
    XRAM[31253] = 8'b0;
    XRAM[31254] = 8'b0;
    XRAM[31255] = 8'b0;
    XRAM[31256] = 8'b0;
    XRAM[31257] = 8'b0;
    XRAM[31258] = 8'b0;
    XRAM[31259] = 8'b0;
    XRAM[31260] = 8'b0;
    XRAM[31261] = 8'b0;
    XRAM[31262] = 8'b0;
    XRAM[31263] = 8'b0;
    XRAM[31264] = 8'b0;
    XRAM[31265] = 8'b0;
    XRAM[31266] = 8'b0;
    XRAM[31267] = 8'b0;
    XRAM[31268] = 8'b0;
    XRAM[31269] = 8'b0;
    XRAM[31270] = 8'b0;
    XRAM[31271] = 8'b0;
    XRAM[31272] = 8'b0;
    XRAM[31273] = 8'b0;
    XRAM[31274] = 8'b0;
    XRAM[31275] = 8'b0;
    XRAM[31276] = 8'b0;
    XRAM[31277] = 8'b0;
    XRAM[31278] = 8'b0;
    XRAM[31279] = 8'b0;
    XRAM[31280] = 8'b0;
    XRAM[31281] = 8'b0;
    XRAM[31282] = 8'b0;
    XRAM[31283] = 8'b0;
    XRAM[31284] = 8'b0;
    XRAM[31285] = 8'b0;
    XRAM[31286] = 8'b0;
    XRAM[31287] = 8'b0;
    XRAM[31288] = 8'b0;
    XRAM[31289] = 8'b0;
    XRAM[31290] = 8'b0;
    XRAM[31291] = 8'b0;
    XRAM[31292] = 8'b0;
    XRAM[31293] = 8'b0;
    XRAM[31294] = 8'b0;
    XRAM[31295] = 8'b0;
    XRAM[31296] = 8'b0;
    XRAM[31297] = 8'b0;
    XRAM[31298] = 8'b0;
    XRAM[31299] = 8'b0;
    XRAM[31300] = 8'b0;
    XRAM[31301] = 8'b0;
    XRAM[31302] = 8'b0;
    XRAM[31303] = 8'b0;
    XRAM[31304] = 8'b0;
    XRAM[31305] = 8'b0;
    XRAM[31306] = 8'b0;
    XRAM[31307] = 8'b0;
    XRAM[31308] = 8'b0;
    XRAM[31309] = 8'b0;
    XRAM[31310] = 8'b0;
    XRAM[31311] = 8'b0;
    XRAM[31312] = 8'b0;
    XRAM[31313] = 8'b0;
    XRAM[31314] = 8'b0;
    XRAM[31315] = 8'b0;
    XRAM[31316] = 8'b0;
    XRAM[31317] = 8'b0;
    XRAM[31318] = 8'b0;
    XRAM[31319] = 8'b0;
    XRAM[31320] = 8'b0;
    XRAM[31321] = 8'b0;
    XRAM[31322] = 8'b0;
    XRAM[31323] = 8'b0;
    XRAM[31324] = 8'b0;
    XRAM[31325] = 8'b0;
    XRAM[31326] = 8'b0;
    XRAM[31327] = 8'b0;
    XRAM[31328] = 8'b0;
    XRAM[31329] = 8'b0;
    XRAM[31330] = 8'b0;
    XRAM[31331] = 8'b0;
    XRAM[31332] = 8'b0;
    XRAM[31333] = 8'b0;
    XRAM[31334] = 8'b0;
    XRAM[31335] = 8'b0;
    XRAM[31336] = 8'b0;
    XRAM[31337] = 8'b0;
    XRAM[31338] = 8'b0;
    XRAM[31339] = 8'b0;
    XRAM[31340] = 8'b0;
    XRAM[31341] = 8'b0;
    XRAM[31342] = 8'b0;
    XRAM[31343] = 8'b0;
    XRAM[31344] = 8'b0;
    XRAM[31345] = 8'b0;
    XRAM[31346] = 8'b0;
    XRAM[31347] = 8'b0;
    XRAM[31348] = 8'b0;
    XRAM[31349] = 8'b0;
    XRAM[31350] = 8'b0;
    XRAM[31351] = 8'b0;
    XRAM[31352] = 8'b0;
    XRAM[31353] = 8'b0;
    XRAM[31354] = 8'b0;
    XRAM[31355] = 8'b0;
    XRAM[31356] = 8'b0;
    XRAM[31357] = 8'b0;
    XRAM[31358] = 8'b0;
    XRAM[31359] = 8'b0;
    XRAM[31360] = 8'b0;
    XRAM[31361] = 8'b0;
    XRAM[31362] = 8'b0;
    XRAM[31363] = 8'b0;
    XRAM[31364] = 8'b0;
    XRAM[31365] = 8'b0;
    XRAM[31366] = 8'b0;
    XRAM[31367] = 8'b0;
    XRAM[31368] = 8'b0;
    XRAM[31369] = 8'b0;
    XRAM[31370] = 8'b0;
    XRAM[31371] = 8'b0;
    XRAM[31372] = 8'b0;
    XRAM[31373] = 8'b0;
    XRAM[31374] = 8'b0;
    XRAM[31375] = 8'b0;
    XRAM[31376] = 8'b0;
    XRAM[31377] = 8'b0;
    XRAM[31378] = 8'b0;
    XRAM[31379] = 8'b0;
    XRAM[31380] = 8'b0;
    XRAM[31381] = 8'b0;
    XRAM[31382] = 8'b0;
    XRAM[31383] = 8'b0;
    XRAM[31384] = 8'b0;
    XRAM[31385] = 8'b0;
    XRAM[31386] = 8'b0;
    XRAM[31387] = 8'b0;
    XRAM[31388] = 8'b0;
    XRAM[31389] = 8'b0;
    XRAM[31390] = 8'b0;
    XRAM[31391] = 8'b0;
    XRAM[31392] = 8'b0;
    XRAM[31393] = 8'b0;
    XRAM[31394] = 8'b0;
    XRAM[31395] = 8'b0;
    XRAM[31396] = 8'b0;
    XRAM[31397] = 8'b0;
    XRAM[31398] = 8'b0;
    XRAM[31399] = 8'b0;
    XRAM[31400] = 8'b0;
    XRAM[31401] = 8'b0;
    XRAM[31402] = 8'b0;
    XRAM[31403] = 8'b0;
    XRAM[31404] = 8'b0;
    XRAM[31405] = 8'b0;
    XRAM[31406] = 8'b0;
    XRAM[31407] = 8'b0;
    XRAM[31408] = 8'b0;
    XRAM[31409] = 8'b0;
    XRAM[31410] = 8'b0;
    XRAM[31411] = 8'b0;
    XRAM[31412] = 8'b0;
    XRAM[31413] = 8'b0;
    XRAM[31414] = 8'b0;
    XRAM[31415] = 8'b0;
    XRAM[31416] = 8'b0;
    XRAM[31417] = 8'b0;
    XRAM[31418] = 8'b0;
    XRAM[31419] = 8'b0;
    XRAM[31420] = 8'b0;
    XRAM[31421] = 8'b0;
    XRAM[31422] = 8'b0;
    XRAM[31423] = 8'b0;
    XRAM[31424] = 8'b0;
    XRAM[31425] = 8'b0;
    XRAM[31426] = 8'b0;
    XRAM[31427] = 8'b0;
    XRAM[31428] = 8'b0;
    XRAM[31429] = 8'b0;
    XRAM[31430] = 8'b0;
    XRAM[31431] = 8'b0;
    XRAM[31432] = 8'b0;
    XRAM[31433] = 8'b0;
    XRAM[31434] = 8'b0;
    XRAM[31435] = 8'b0;
    XRAM[31436] = 8'b0;
    XRAM[31437] = 8'b0;
    XRAM[31438] = 8'b0;
    XRAM[31439] = 8'b0;
    XRAM[31440] = 8'b0;
    XRAM[31441] = 8'b0;
    XRAM[31442] = 8'b0;
    XRAM[31443] = 8'b0;
    XRAM[31444] = 8'b0;
    XRAM[31445] = 8'b0;
    XRAM[31446] = 8'b0;
    XRAM[31447] = 8'b0;
    XRAM[31448] = 8'b0;
    XRAM[31449] = 8'b0;
    XRAM[31450] = 8'b0;
    XRAM[31451] = 8'b0;
    XRAM[31452] = 8'b0;
    XRAM[31453] = 8'b0;
    XRAM[31454] = 8'b0;
    XRAM[31455] = 8'b0;
    XRAM[31456] = 8'b0;
    XRAM[31457] = 8'b0;
    XRAM[31458] = 8'b0;
    XRAM[31459] = 8'b0;
    XRAM[31460] = 8'b0;
    XRAM[31461] = 8'b0;
    XRAM[31462] = 8'b0;
    XRAM[31463] = 8'b0;
    XRAM[31464] = 8'b0;
    XRAM[31465] = 8'b0;
    XRAM[31466] = 8'b0;
    XRAM[31467] = 8'b0;
    XRAM[31468] = 8'b0;
    XRAM[31469] = 8'b0;
    XRAM[31470] = 8'b0;
    XRAM[31471] = 8'b0;
    XRAM[31472] = 8'b0;
    XRAM[31473] = 8'b0;
    XRAM[31474] = 8'b0;
    XRAM[31475] = 8'b0;
    XRAM[31476] = 8'b0;
    XRAM[31477] = 8'b0;
    XRAM[31478] = 8'b0;
    XRAM[31479] = 8'b0;
    XRAM[31480] = 8'b0;
    XRAM[31481] = 8'b0;
    XRAM[31482] = 8'b0;
    XRAM[31483] = 8'b0;
    XRAM[31484] = 8'b0;
    XRAM[31485] = 8'b0;
    XRAM[31486] = 8'b0;
    XRAM[31487] = 8'b0;
    XRAM[31488] = 8'b0;
    XRAM[31489] = 8'b0;
    XRAM[31490] = 8'b0;
    XRAM[31491] = 8'b0;
    XRAM[31492] = 8'b0;
    XRAM[31493] = 8'b0;
    XRAM[31494] = 8'b0;
    XRAM[31495] = 8'b0;
    XRAM[31496] = 8'b0;
    XRAM[31497] = 8'b0;
    XRAM[31498] = 8'b0;
    XRAM[31499] = 8'b0;
    XRAM[31500] = 8'b0;
    XRAM[31501] = 8'b0;
    XRAM[31502] = 8'b0;
    XRAM[31503] = 8'b0;
    XRAM[31504] = 8'b0;
    XRAM[31505] = 8'b0;
    XRAM[31506] = 8'b0;
    XRAM[31507] = 8'b0;
    XRAM[31508] = 8'b0;
    XRAM[31509] = 8'b0;
    XRAM[31510] = 8'b0;
    XRAM[31511] = 8'b0;
    XRAM[31512] = 8'b0;
    XRAM[31513] = 8'b0;
    XRAM[31514] = 8'b0;
    XRAM[31515] = 8'b0;
    XRAM[31516] = 8'b0;
    XRAM[31517] = 8'b0;
    XRAM[31518] = 8'b0;
    XRAM[31519] = 8'b0;
    XRAM[31520] = 8'b0;
    XRAM[31521] = 8'b0;
    XRAM[31522] = 8'b0;
    XRAM[31523] = 8'b0;
    XRAM[31524] = 8'b0;
    XRAM[31525] = 8'b0;
    XRAM[31526] = 8'b0;
    XRAM[31527] = 8'b0;
    XRAM[31528] = 8'b0;
    XRAM[31529] = 8'b0;
    XRAM[31530] = 8'b0;
    XRAM[31531] = 8'b0;
    XRAM[31532] = 8'b0;
    XRAM[31533] = 8'b0;
    XRAM[31534] = 8'b0;
    XRAM[31535] = 8'b0;
    XRAM[31536] = 8'b0;
    XRAM[31537] = 8'b0;
    XRAM[31538] = 8'b0;
    XRAM[31539] = 8'b0;
    XRAM[31540] = 8'b0;
    XRAM[31541] = 8'b0;
    XRAM[31542] = 8'b0;
    XRAM[31543] = 8'b0;
    XRAM[31544] = 8'b0;
    XRAM[31545] = 8'b0;
    XRAM[31546] = 8'b0;
    XRAM[31547] = 8'b0;
    XRAM[31548] = 8'b0;
    XRAM[31549] = 8'b0;
    XRAM[31550] = 8'b0;
    XRAM[31551] = 8'b0;
    XRAM[31552] = 8'b0;
    XRAM[31553] = 8'b0;
    XRAM[31554] = 8'b0;
    XRAM[31555] = 8'b0;
    XRAM[31556] = 8'b0;
    XRAM[31557] = 8'b0;
    XRAM[31558] = 8'b0;
    XRAM[31559] = 8'b0;
    XRAM[31560] = 8'b0;
    XRAM[31561] = 8'b0;
    XRAM[31562] = 8'b0;
    XRAM[31563] = 8'b0;
    XRAM[31564] = 8'b0;
    XRAM[31565] = 8'b0;
    XRAM[31566] = 8'b0;
    XRAM[31567] = 8'b0;
    XRAM[31568] = 8'b0;
    XRAM[31569] = 8'b0;
    XRAM[31570] = 8'b0;
    XRAM[31571] = 8'b0;
    XRAM[31572] = 8'b0;
    XRAM[31573] = 8'b0;
    XRAM[31574] = 8'b0;
    XRAM[31575] = 8'b0;
    XRAM[31576] = 8'b0;
    XRAM[31577] = 8'b0;
    XRAM[31578] = 8'b0;
    XRAM[31579] = 8'b0;
    XRAM[31580] = 8'b0;
    XRAM[31581] = 8'b0;
    XRAM[31582] = 8'b0;
    XRAM[31583] = 8'b0;
    XRAM[31584] = 8'b0;
    XRAM[31585] = 8'b0;
    XRAM[31586] = 8'b0;
    XRAM[31587] = 8'b0;
    XRAM[31588] = 8'b0;
    XRAM[31589] = 8'b0;
    XRAM[31590] = 8'b0;
    XRAM[31591] = 8'b0;
    XRAM[31592] = 8'b0;
    XRAM[31593] = 8'b0;
    XRAM[31594] = 8'b0;
    XRAM[31595] = 8'b0;
    XRAM[31596] = 8'b0;
    XRAM[31597] = 8'b0;
    XRAM[31598] = 8'b0;
    XRAM[31599] = 8'b0;
    XRAM[31600] = 8'b0;
    XRAM[31601] = 8'b0;
    XRAM[31602] = 8'b0;
    XRAM[31603] = 8'b0;
    XRAM[31604] = 8'b0;
    XRAM[31605] = 8'b0;
    XRAM[31606] = 8'b0;
    XRAM[31607] = 8'b0;
    XRAM[31608] = 8'b0;
    XRAM[31609] = 8'b0;
    XRAM[31610] = 8'b0;
    XRAM[31611] = 8'b0;
    XRAM[31612] = 8'b0;
    XRAM[31613] = 8'b0;
    XRAM[31614] = 8'b0;
    XRAM[31615] = 8'b0;
    XRAM[31616] = 8'b0;
    XRAM[31617] = 8'b0;
    XRAM[31618] = 8'b0;
    XRAM[31619] = 8'b0;
    XRAM[31620] = 8'b0;
    XRAM[31621] = 8'b0;
    XRAM[31622] = 8'b0;
    XRAM[31623] = 8'b0;
    XRAM[31624] = 8'b0;
    XRAM[31625] = 8'b0;
    XRAM[31626] = 8'b0;
    XRAM[31627] = 8'b0;
    XRAM[31628] = 8'b0;
    XRAM[31629] = 8'b0;
    XRAM[31630] = 8'b0;
    XRAM[31631] = 8'b0;
    XRAM[31632] = 8'b0;
    XRAM[31633] = 8'b0;
    XRAM[31634] = 8'b0;
    XRAM[31635] = 8'b0;
    XRAM[31636] = 8'b0;
    XRAM[31637] = 8'b0;
    XRAM[31638] = 8'b0;
    XRAM[31639] = 8'b0;
    XRAM[31640] = 8'b0;
    XRAM[31641] = 8'b0;
    XRAM[31642] = 8'b0;
    XRAM[31643] = 8'b0;
    XRAM[31644] = 8'b0;
    XRAM[31645] = 8'b0;
    XRAM[31646] = 8'b0;
    XRAM[31647] = 8'b0;
    XRAM[31648] = 8'b0;
    XRAM[31649] = 8'b0;
    XRAM[31650] = 8'b0;
    XRAM[31651] = 8'b0;
    XRAM[31652] = 8'b0;
    XRAM[31653] = 8'b0;
    XRAM[31654] = 8'b0;
    XRAM[31655] = 8'b0;
    XRAM[31656] = 8'b0;
    XRAM[31657] = 8'b0;
    XRAM[31658] = 8'b0;
    XRAM[31659] = 8'b0;
    XRAM[31660] = 8'b0;
    XRAM[31661] = 8'b0;
    XRAM[31662] = 8'b0;
    XRAM[31663] = 8'b0;
    XRAM[31664] = 8'b0;
    XRAM[31665] = 8'b0;
    XRAM[31666] = 8'b0;
    XRAM[31667] = 8'b0;
    XRAM[31668] = 8'b0;
    XRAM[31669] = 8'b0;
    XRAM[31670] = 8'b0;
    XRAM[31671] = 8'b0;
    XRAM[31672] = 8'b0;
    XRAM[31673] = 8'b0;
    XRAM[31674] = 8'b0;
    XRAM[31675] = 8'b0;
    XRAM[31676] = 8'b0;
    XRAM[31677] = 8'b0;
    XRAM[31678] = 8'b0;
    XRAM[31679] = 8'b0;
    XRAM[31680] = 8'b0;
    XRAM[31681] = 8'b0;
    XRAM[31682] = 8'b0;
    XRAM[31683] = 8'b0;
    XRAM[31684] = 8'b0;
    XRAM[31685] = 8'b0;
    XRAM[31686] = 8'b0;
    XRAM[31687] = 8'b0;
    XRAM[31688] = 8'b0;
    XRAM[31689] = 8'b0;
    XRAM[31690] = 8'b0;
    XRAM[31691] = 8'b0;
    XRAM[31692] = 8'b0;
    XRAM[31693] = 8'b0;
    XRAM[31694] = 8'b0;
    XRAM[31695] = 8'b0;
    XRAM[31696] = 8'b0;
    XRAM[31697] = 8'b0;
    XRAM[31698] = 8'b0;
    XRAM[31699] = 8'b0;
    XRAM[31700] = 8'b0;
    XRAM[31701] = 8'b0;
    XRAM[31702] = 8'b0;
    XRAM[31703] = 8'b0;
    XRAM[31704] = 8'b0;
    XRAM[31705] = 8'b0;
    XRAM[31706] = 8'b0;
    XRAM[31707] = 8'b0;
    XRAM[31708] = 8'b0;
    XRAM[31709] = 8'b0;
    XRAM[31710] = 8'b0;
    XRAM[31711] = 8'b0;
    XRAM[31712] = 8'b0;
    XRAM[31713] = 8'b0;
    XRAM[31714] = 8'b0;
    XRAM[31715] = 8'b0;
    XRAM[31716] = 8'b0;
    XRAM[31717] = 8'b0;
    XRAM[31718] = 8'b0;
    XRAM[31719] = 8'b0;
    XRAM[31720] = 8'b0;
    XRAM[31721] = 8'b0;
    XRAM[31722] = 8'b0;
    XRAM[31723] = 8'b0;
    XRAM[31724] = 8'b0;
    XRAM[31725] = 8'b0;
    XRAM[31726] = 8'b0;
    XRAM[31727] = 8'b0;
    XRAM[31728] = 8'b0;
    XRAM[31729] = 8'b0;
    XRAM[31730] = 8'b0;
    XRAM[31731] = 8'b0;
    XRAM[31732] = 8'b0;
    XRAM[31733] = 8'b0;
    XRAM[31734] = 8'b0;
    XRAM[31735] = 8'b0;
    XRAM[31736] = 8'b0;
    XRAM[31737] = 8'b0;
    XRAM[31738] = 8'b0;
    XRAM[31739] = 8'b0;
    XRAM[31740] = 8'b0;
    XRAM[31741] = 8'b0;
    XRAM[31742] = 8'b0;
    XRAM[31743] = 8'b0;
    XRAM[31744] = 8'b0;
    XRAM[31745] = 8'b0;
    XRAM[31746] = 8'b0;
    XRAM[31747] = 8'b0;
    XRAM[31748] = 8'b0;
    XRAM[31749] = 8'b0;
    XRAM[31750] = 8'b0;
    XRAM[31751] = 8'b0;
    XRAM[31752] = 8'b0;
    XRAM[31753] = 8'b0;
    XRAM[31754] = 8'b0;
    XRAM[31755] = 8'b0;
    XRAM[31756] = 8'b0;
    XRAM[31757] = 8'b0;
    XRAM[31758] = 8'b0;
    XRAM[31759] = 8'b0;
    XRAM[31760] = 8'b0;
    XRAM[31761] = 8'b0;
    XRAM[31762] = 8'b0;
    XRAM[31763] = 8'b0;
    XRAM[31764] = 8'b0;
    XRAM[31765] = 8'b0;
    XRAM[31766] = 8'b0;
    XRAM[31767] = 8'b0;
    XRAM[31768] = 8'b0;
    XRAM[31769] = 8'b0;
    XRAM[31770] = 8'b0;
    XRAM[31771] = 8'b0;
    XRAM[31772] = 8'b0;
    XRAM[31773] = 8'b0;
    XRAM[31774] = 8'b0;
    XRAM[31775] = 8'b0;
    XRAM[31776] = 8'b0;
    XRAM[31777] = 8'b0;
    XRAM[31778] = 8'b0;
    XRAM[31779] = 8'b0;
    XRAM[31780] = 8'b0;
    XRAM[31781] = 8'b0;
    XRAM[31782] = 8'b0;
    XRAM[31783] = 8'b0;
    XRAM[31784] = 8'b0;
    XRAM[31785] = 8'b0;
    XRAM[31786] = 8'b0;
    XRAM[31787] = 8'b0;
    XRAM[31788] = 8'b0;
    XRAM[31789] = 8'b0;
    XRAM[31790] = 8'b0;
    XRAM[31791] = 8'b0;
    XRAM[31792] = 8'b0;
    XRAM[31793] = 8'b0;
    XRAM[31794] = 8'b0;
    XRAM[31795] = 8'b0;
    XRAM[31796] = 8'b0;
    XRAM[31797] = 8'b0;
    XRAM[31798] = 8'b0;
    XRAM[31799] = 8'b0;
    XRAM[31800] = 8'b0;
    XRAM[31801] = 8'b0;
    XRAM[31802] = 8'b0;
    XRAM[31803] = 8'b0;
    XRAM[31804] = 8'b0;
    XRAM[31805] = 8'b0;
    XRAM[31806] = 8'b0;
    XRAM[31807] = 8'b0;
    XRAM[31808] = 8'b0;
    XRAM[31809] = 8'b0;
    XRAM[31810] = 8'b0;
    XRAM[31811] = 8'b0;
    XRAM[31812] = 8'b0;
    XRAM[31813] = 8'b0;
    XRAM[31814] = 8'b0;
    XRAM[31815] = 8'b0;
    XRAM[31816] = 8'b0;
    XRAM[31817] = 8'b0;
    XRAM[31818] = 8'b0;
    XRAM[31819] = 8'b0;
    XRAM[31820] = 8'b0;
    XRAM[31821] = 8'b0;
    XRAM[31822] = 8'b0;
    XRAM[31823] = 8'b0;
    XRAM[31824] = 8'b0;
    XRAM[31825] = 8'b0;
    XRAM[31826] = 8'b0;
    XRAM[31827] = 8'b0;
    XRAM[31828] = 8'b0;
    XRAM[31829] = 8'b0;
    XRAM[31830] = 8'b0;
    XRAM[31831] = 8'b0;
    XRAM[31832] = 8'b0;
    XRAM[31833] = 8'b0;
    XRAM[31834] = 8'b0;
    XRAM[31835] = 8'b0;
    XRAM[31836] = 8'b0;
    XRAM[31837] = 8'b0;
    XRAM[31838] = 8'b0;
    XRAM[31839] = 8'b0;
    XRAM[31840] = 8'b0;
    XRAM[31841] = 8'b0;
    XRAM[31842] = 8'b0;
    XRAM[31843] = 8'b0;
    XRAM[31844] = 8'b0;
    XRAM[31845] = 8'b0;
    XRAM[31846] = 8'b0;
    XRAM[31847] = 8'b0;
    XRAM[31848] = 8'b0;
    XRAM[31849] = 8'b0;
    XRAM[31850] = 8'b0;
    XRAM[31851] = 8'b0;
    XRAM[31852] = 8'b0;
    XRAM[31853] = 8'b0;
    XRAM[31854] = 8'b0;
    XRAM[31855] = 8'b0;
    XRAM[31856] = 8'b0;
    XRAM[31857] = 8'b0;
    XRAM[31858] = 8'b0;
    XRAM[31859] = 8'b0;
    XRAM[31860] = 8'b0;
    XRAM[31861] = 8'b0;
    XRAM[31862] = 8'b0;
    XRAM[31863] = 8'b0;
    XRAM[31864] = 8'b0;
    XRAM[31865] = 8'b0;
    XRAM[31866] = 8'b0;
    XRAM[31867] = 8'b0;
    XRAM[31868] = 8'b0;
    XRAM[31869] = 8'b0;
    XRAM[31870] = 8'b0;
    XRAM[31871] = 8'b0;
    XRAM[31872] = 8'b0;
    XRAM[31873] = 8'b0;
    XRAM[31874] = 8'b0;
    XRAM[31875] = 8'b0;
    XRAM[31876] = 8'b0;
    XRAM[31877] = 8'b0;
    XRAM[31878] = 8'b0;
    XRAM[31879] = 8'b0;
    XRAM[31880] = 8'b0;
    XRAM[31881] = 8'b0;
    XRAM[31882] = 8'b0;
    XRAM[31883] = 8'b0;
    XRAM[31884] = 8'b0;
    XRAM[31885] = 8'b0;
    XRAM[31886] = 8'b0;
    XRAM[31887] = 8'b0;
    XRAM[31888] = 8'b0;
    XRAM[31889] = 8'b0;
    XRAM[31890] = 8'b0;
    XRAM[31891] = 8'b0;
    XRAM[31892] = 8'b0;
    XRAM[31893] = 8'b0;
    XRAM[31894] = 8'b0;
    XRAM[31895] = 8'b0;
    XRAM[31896] = 8'b0;
    XRAM[31897] = 8'b0;
    XRAM[31898] = 8'b0;
    XRAM[31899] = 8'b0;
    XRAM[31900] = 8'b0;
    XRAM[31901] = 8'b0;
    XRAM[31902] = 8'b0;
    XRAM[31903] = 8'b0;
    XRAM[31904] = 8'b0;
    XRAM[31905] = 8'b0;
    XRAM[31906] = 8'b0;
    XRAM[31907] = 8'b0;
    XRAM[31908] = 8'b0;
    XRAM[31909] = 8'b0;
    XRAM[31910] = 8'b0;
    XRAM[31911] = 8'b0;
    XRAM[31912] = 8'b0;
    XRAM[31913] = 8'b0;
    XRAM[31914] = 8'b0;
    XRAM[31915] = 8'b0;
    XRAM[31916] = 8'b0;
    XRAM[31917] = 8'b0;
    XRAM[31918] = 8'b0;
    XRAM[31919] = 8'b0;
    XRAM[31920] = 8'b0;
    XRAM[31921] = 8'b0;
    XRAM[31922] = 8'b0;
    XRAM[31923] = 8'b0;
    XRAM[31924] = 8'b0;
    XRAM[31925] = 8'b0;
    XRAM[31926] = 8'b0;
    XRAM[31927] = 8'b0;
    XRAM[31928] = 8'b0;
    XRAM[31929] = 8'b0;
    XRAM[31930] = 8'b0;
    XRAM[31931] = 8'b0;
    XRAM[31932] = 8'b0;
    XRAM[31933] = 8'b0;
    XRAM[31934] = 8'b0;
    XRAM[31935] = 8'b0;
    XRAM[31936] = 8'b0;
    XRAM[31937] = 8'b0;
    XRAM[31938] = 8'b0;
    XRAM[31939] = 8'b0;
    XRAM[31940] = 8'b0;
    XRAM[31941] = 8'b0;
    XRAM[31942] = 8'b0;
    XRAM[31943] = 8'b0;
    XRAM[31944] = 8'b0;
    XRAM[31945] = 8'b0;
    XRAM[31946] = 8'b0;
    XRAM[31947] = 8'b0;
    XRAM[31948] = 8'b0;
    XRAM[31949] = 8'b0;
    XRAM[31950] = 8'b0;
    XRAM[31951] = 8'b0;
    XRAM[31952] = 8'b0;
    XRAM[31953] = 8'b0;
    XRAM[31954] = 8'b0;
    XRAM[31955] = 8'b0;
    XRAM[31956] = 8'b0;
    XRAM[31957] = 8'b0;
    XRAM[31958] = 8'b0;
    XRAM[31959] = 8'b0;
    XRAM[31960] = 8'b0;
    XRAM[31961] = 8'b0;
    XRAM[31962] = 8'b0;
    XRAM[31963] = 8'b0;
    XRAM[31964] = 8'b0;
    XRAM[31965] = 8'b0;
    XRAM[31966] = 8'b0;
    XRAM[31967] = 8'b0;
    XRAM[31968] = 8'b0;
    XRAM[31969] = 8'b0;
    XRAM[31970] = 8'b0;
    XRAM[31971] = 8'b0;
    XRAM[31972] = 8'b0;
    XRAM[31973] = 8'b0;
    XRAM[31974] = 8'b0;
    XRAM[31975] = 8'b0;
    XRAM[31976] = 8'b0;
    XRAM[31977] = 8'b0;
    XRAM[31978] = 8'b0;
    XRAM[31979] = 8'b0;
    XRAM[31980] = 8'b0;
    XRAM[31981] = 8'b0;
    XRAM[31982] = 8'b0;
    XRAM[31983] = 8'b0;
    XRAM[31984] = 8'b0;
    XRAM[31985] = 8'b0;
    XRAM[31986] = 8'b0;
    XRAM[31987] = 8'b0;
    XRAM[31988] = 8'b0;
    XRAM[31989] = 8'b0;
    XRAM[31990] = 8'b0;
    XRAM[31991] = 8'b0;
    XRAM[31992] = 8'b0;
    XRAM[31993] = 8'b0;
    XRAM[31994] = 8'b0;
    XRAM[31995] = 8'b0;
    XRAM[31996] = 8'b0;
    XRAM[31997] = 8'b0;
    XRAM[31998] = 8'b0;
    XRAM[31999] = 8'b0;
    XRAM[32000] = 8'b0;
    XRAM[32001] = 8'b0;
    XRAM[32002] = 8'b0;
    XRAM[32003] = 8'b0;
    XRAM[32004] = 8'b0;
    XRAM[32005] = 8'b0;
    XRAM[32006] = 8'b0;
    XRAM[32007] = 8'b0;
    XRAM[32008] = 8'b0;
    XRAM[32009] = 8'b0;
    XRAM[32010] = 8'b0;
    XRAM[32011] = 8'b0;
    XRAM[32012] = 8'b0;
    XRAM[32013] = 8'b0;
    XRAM[32014] = 8'b0;
    XRAM[32015] = 8'b0;
    XRAM[32016] = 8'b0;
    XRAM[32017] = 8'b0;
    XRAM[32018] = 8'b0;
    XRAM[32019] = 8'b0;
    XRAM[32020] = 8'b0;
    XRAM[32021] = 8'b0;
    XRAM[32022] = 8'b0;
    XRAM[32023] = 8'b0;
    XRAM[32024] = 8'b0;
    XRAM[32025] = 8'b0;
    XRAM[32026] = 8'b0;
    XRAM[32027] = 8'b0;
    XRAM[32028] = 8'b0;
    XRAM[32029] = 8'b0;
    XRAM[32030] = 8'b0;
    XRAM[32031] = 8'b0;
    XRAM[32032] = 8'b0;
    XRAM[32033] = 8'b0;
    XRAM[32034] = 8'b0;
    XRAM[32035] = 8'b0;
    XRAM[32036] = 8'b0;
    XRAM[32037] = 8'b0;
    XRAM[32038] = 8'b0;
    XRAM[32039] = 8'b0;
    XRAM[32040] = 8'b0;
    XRAM[32041] = 8'b0;
    XRAM[32042] = 8'b0;
    XRAM[32043] = 8'b0;
    XRAM[32044] = 8'b0;
    XRAM[32045] = 8'b0;
    XRAM[32046] = 8'b0;
    XRAM[32047] = 8'b0;
    XRAM[32048] = 8'b0;
    XRAM[32049] = 8'b0;
    XRAM[32050] = 8'b0;
    XRAM[32051] = 8'b0;
    XRAM[32052] = 8'b0;
    XRAM[32053] = 8'b0;
    XRAM[32054] = 8'b0;
    XRAM[32055] = 8'b0;
    XRAM[32056] = 8'b0;
    XRAM[32057] = 8'b0;
    XRAM[32058] = 8'b0;
    XRAM[32059] = 8'b0;
    XRAM[32060] = 8'b0;
    XRAM[32061] = 8'b0;
    XRAM[32062] = 8'b0;
    XRAM[32063] = 8'b0;
    XRAM[32064] = 8'b0;
    XRAM[32065] = 8'b0;
    XRAM[32066] = 8'b0;
    XRAM[32067] = 8'b0;
    XRAM[32068] = 8'b0;
    XRAM[32069] = 8'b0;
    XRAM[32070] = 8'b0;
    XRAM[32071] = 8'b0;
    XRAM[32072] = 8'b0;
    XRAM[32073] = 8'b0;
    XRAM[32074] = 8'b0;
    XRAM[32075] = 8'b0;
    XRAM[32076] = 8'b0;
    XRAM[32077] = 8'b0;
    XRAM[32078] = 8'b0;
    XRAM[32079] = 8'b0;
    XRAM[32080] = 8'b0;
    XRAM[32081] = 8'b0;
    XRAM[32082] = 8'b0;
    XRAM[32083] = 8'b0;
    XRAM[32084] = 8'b0;
    XRAM[32085] = 8'b0;
    XRAM[32086] = 8'b0;
    XRAM[32087] = 8'b0;
    XRAM[32088] = 8'b0;
    XRAM[32089] = 8'b0;
    XRAM[32090] = 8'b0;
    XRAM[32091] = 8'b0;
    XRAM[32092] = 8'b0;
    XRAM[32093] = 8'b0;
    XRAM[32094] = 8'b0;
    XRAM[32095] = 8'b0;
    XRAM[32096] = 8'b0;
    XRAM[32097] = 8'b0;
    XRAM[32098] = 8'b0;
    XRAM[32099] = 8'b0;
    XRAM[32100] = 8'b0;
    XRAM[32101] = 8'b0;
    XRAM[32102] = 8'b0;
    XRAM[32103] = 8'b0;
    XRAM[32104] = 8'b0;
    XRAM[32105] = 8'b0;
    XRAM[32106] = 8'b0;
    XRAM[32107] = 8'b0;
    XRAM[32108] = 8'b0;
    XRAM[32109] = 8'b0;
    XRAM[32110] = 8'b0;
    XRAM[32111] = 8'b0;
    XRAM[32112] = 8'b0;
    XRAM[32113] = 8'b0;
    XRAM[32114] = 8'b0;
    XRAM[32115] = 8'b0;
    XRAM[32116] = 8'b0;
    XRAM[32117] = 8'b0;
    XRAM[32118] = 8'b0;
    XRAM[32119] = 8'b0;
    XRAM[32120] = 8'b0;
    XRAM[32121] = 8'b0;
    XRAM[32122] = 8'b0;
    XRAM[32123] = 8'b0;
    XRAM[32124] = 8'b0;
    XRAM[32125] = 8'b0;
    XRAM[32126] = 8'b0;
    XRAM[32127] = 8'b0;
    XRAM[32128] = 8'b0;
    XRAM[32129] = 8'b0;
    XRAM[32130] = 8'b0;
    XRAM[32131] = 8'b0;
    XRAM[32132] = 8'b0;
    XRAM[32133] = 8'b0;
    XRAM[32134] = 8'b0;
    XRAM[32135] = 8'b0;
    XRAM[32136] = 8'b0;
    XRAM[32137] = 8'b0;
    XRAM[32138] = 8'b0;
    XRAM[32139] = 8'b0;
    XRAM[32140] = 8'b0;
    XRAM[32141] = 8'b0;
    XRAM[32142] = 8'b0;
    XRAM[32143] = 8'b0;
    XRAM[32144] = 8'b0;
    XRAM[32145] = 8'b0;
    XRAM[32146] = 8'b0;
    XRAM[32147] = 8'b0;
    XRAM[32148] = 8'b0;
    XRAM[32149] = 8'b0;
    XRAM[32150] = 8'b0;
    XRAM[32151] = 8'b0;
    XRAM[32152] = 8'b0;
    XRAM[32153] = 8'b0;
    XRAM[32154] = 8'b0;
    XRAM[32155] = 8'b0;
    XRAM[32156] = 8'b0;
    XRAM[32157] = 8'b0;
    XRAM[32158] = 8'b0;
    XRAM[32159] = 8'b0;
    XRAM[32160] = 8'b0;
    XRAM[32161] = 8'b0;
    XRAM[32162] = 8'b0;
    XRAM[32163] = 8'b0;
    XRAM[32164] = 8'b0;
    XRAM[32165] = 8'b0;
    XRAM[32166] = 8'b0;
    XRAM[32167] = 8'b0;
    XRAM[32168] = 8'b0;
    XRAM[32169] = 8'b0;
    XRAM[32170] = 8'b0;
    XRAM[32171] = 8'b0;
    XRAM[32172] = 8'b0;
    XRAM[32173] = 8'b0;
    XRAM[32174] = 8'b0;
    XRAM[32175] = 8'b0;
    XRAM[32176] = 8'b0;
    XRAM[32177] = 8'b0;
    XRAM[32178] = 8'b0;
    XRAM[32179] = 8'b0;
    XRAM[32180] = 8'b0;
    XRAM[32181] = 8'b0;
    XRAM[32182] = 8'b0;
    XRAM[32183] = 8'b0;
    XRAM[32184] = 8'b0;
    XRAM[32185] = 8'b0;
    XRAM[32186] = 8'b0;
    XRAM[32187] = 8'b0;
    XRAM[32188] = 8'b0;
    XRAM[32189] = 8'b0;
    XRAM[32190] = 8'b0;
    XRAM[32191] = 8'b0;
    XRAM[32192] = 8'b0;
    XRAM[32193] = 8'b0;
    XRAM[32194] = 8'b0;
    XRAM[32195] = 8'b0;
    XRAM[32196] = 8'b0;
    XRAM[32197] = 8'b0;
    XRAM[32198] = 8'b0;
    XRAM[32199] = 8'b0;
    XRAM[32200] = 8'b0;
    XRAM[32201] = 8'b0;
    XRAM[32202] = 8'b0;
    XRAM[32203] = 8'b0;
    XRAM[32204] = 8'b0;
    XRAM[32205] = 8'b0;
    XRAM[32206] = 8'b0;
    XRAM[32207] = 8'b0;
    XRAM[32208] = 8'b0;
    XRAM[32209] = 8'b0;
    XRAM[32210] = 8'b0;
    XRAM[32211] = 8'b0;
    XRAM[32212] = 8'b0;
    XRAM[32213] = 8'b0;
    XRAM[32214] = 8'b0;
    XRAM[32215] = 8'b0;
    XRAM[32216] = 8'b0;
    XRAM[32217] = 8'b0;
    XRAM[32218] = 8'b0;
    XRAM[32219] = 8'b0;
    XRAM[32220] = 8'b0;
    XRAM[32221] = 8'b0;
    XRAM[32222] = 8'b0;
    XRAM[32223] = 8'b0;
    XRAM[32224] = 8'b0;
    XRAM[32225] = 8'b0;
    XRAM[32226] = 8'b0;
    XRAM[32227] = 8'b0;
    XRAM[32228] = 8'b0;
    XRAM[32229] = 8'b0;
    XRAM[32230] = 8'b0;
    XRAM[32231] = 8'b0;
    XRAM[32232] = 8'b0;
    XRAM[32233] = 8'b0;
    XRAM[32234] = 8'b0;
    XRAM[32235] = 8'b0;
    XRAM[32236] = 8'b0;
    XRAM[32237] = 8'b0;
    XRAM[32238] = 8'b0;
    XRAM[32239] = 8'b0;
    XRAM[32240] = 8'b0;
    XRAM[32241] = 8'b0;
    XRAM[32242] = 8'b0;
    XRAM[32243] = 8'b0;
    XRAM[32244] = 8'b0;
    XRAM[32245] = 8'b0;
    XRAM[32246] = 8'b0;
    XRAM[32247] = 8'b0;
    XRAM[32248] = 8'b0;
    XRAM[32249] = 8'b0;
    XRAM[32250] = 8'b0;
    XRAM[32251] = 8'b0;
    XRAM[32252] = 8'b0;
    XRAM[32253] = 8'b0;
    XRAM[32254] = 8'b0;
    XRAM[32255] = 8'b0;
    XRAM[32256] = 8'b0;
    XRAM[32257] = 8'b0;
    XRAM[32258] = 8'b0;
    XRAM[32259] = 8'b0;
    XRAM[32260] = 8'b0;
    XRAM[32261] = 8'b0;
    XRAM[32262] = 8'b0;
    XRAM[32263] = 8'b0;
    XRAM[32264] = 8'b0;
    XRAM[32265] = 8'b0;
    XRAM[32266] = 8'b0;
    XRAM[32267] = 8'b0;
    XRAM[32268] = 8'b0;
    XRAM[32269] = 8'b0;
    XRAM[32270] = 8'b0;
    XRAM[32271] = 8'b0;
    XRAM[32272] = 8'b0;
    XRAM[32273] = 8'b0;
    XRAM[32274] = 8'b0;
    XRAM[32275] = 8'b0;
    XRAM[32276] = 8'b0;
    XRAM[32277] = 8'b0;
    XRAM[32278] = 8'b0;
    XRAM[32279] = 8'b0;
    XRAM[32280] = 8'b0;
    XRAM[32281] = 8'b0;
    XRAM[32282] = 8'b0;
    XRAM[32283] = 8'b0;
    XRAM[32284] = 8'b0;
    XRAM[32285] = 8'b0;
    XRAM[32286] = 8'b0;
    XRAM[32287] = 8'b0;
    XRAM[32288] = 8'b0;
    XRAM[32289] = 8'b0;
    XRAM[32290] = 8'b0;
    XRAM[32291] = 8'b0;
    XRAM[32292] = 8'b0;
    XRAM[32293] = 8'b0;
    XRAM[32294] = 8'b0;
    XRAM[32295] = 8'b0;
    XRAM[32296] = 8'b0;
    XRAM[32297] = 8'b0;
    XRAM[32298] = 8'b0;
    XRAM[32299] = 8'b0;
    XRAM[32300] = 8'b0;
    XRAM[32301] = 8'b0;
    XRAM[32302] = 8'b0;
    XRAM[32303] = 8'b0;
    XRAM[32304] = 8'b0;
    XRAM[32305] = 8'b0;
    XRAM[32306] = 8'b0;
    XRAM[32307] = 8'b0;
    XRAM[32308] = 8'b0;
    XRAM[32309] = 8'b0;
    XRAM[32310] = 8'b0;
    XRAM[32311] = 8'b0;
    XRAM[32312] = 8'b0;
    XRAM[32313] = 8'b0;
    XRAM[32314] = 8'b0;
    XRAM[32315] = 8'b0;
    XRAM[32316] = 8'b0;
    XRAM[32317] = 8'b0;
    XRAM[32318] = 8'b0;
    XRAM[32319] = 8'b0;
    XRAM[32320] = 8'b0;
    XRAM[32321] = 8'b0;
    XRAM[32322] = 8'b0;
    XRAM[32323] = 8'b0;
    XRAM[32324] = 8'b0;
    XRAM[32325] = 8'b0;
    XRAM[32326] = 8'b0;
    XRAM[32327] = 8'b0;
    XRAM[32328] = 8'b0;
    XRAM[32329] = 8'b0;
    XRAM[32330] = 8'b0;
    XRAM[32331] = 8'b0;
    XRAM[32332] = 8'b0;
    XRAM[32333] = 8'b0;
    XRAM[32334] = 8'b0;
    XRAM[32335] = 8'b0;
    XRAM[32336] = 8'b0;
    XRAM[32337] = 8'b0;
    XRAM[32338] = 8'b0;
    XRAM[32339] = 8'b0;
    XRAM[32340] = 8'b0;
    XRAM[32341] = 8'b0;
    XRAM[32342] = 8'b0;
    XRAM[32343] = 8'b0;
    XRAM[32344] = 8'b0;
    XRAM[32345] = 8'b0;
    XRAM[32346] = 8'b0;
    XRAM[32347] = 8'b0;
    XRAM[32348] = 8'b0;
    XRAM[32349] = 8'b0;
    XRAM[32350] = 8'b0;
    XRAM[32351] = 8'b0;
    XRAM[32352] = 8'b0;
    XRAM[32353] = 8'b0;
    XRAM[32354] = 8'b0;
    XRAM[32355] = 8'b0;
    XRAM[32356] = 8'b0;
    XRAM[32357] = 8'b0;
    XRAM[32358] = 8'b0;
    XRAM[32359] = 8'b0;
    XRAM[32360] = 8'b0;
    XRAM[32361] = 8'b0;
    XRAM[32362] = 8'b0;
    XRAM[32363] = 8'b0;
    XRAM[32364] = 8'b0;
    XRAM[32365] = 8'b0;
    XRAM[32366] = 8'b0;
    XRAM[32367] = 8'b0;
    XRAM[32368] = 8'b0;
    XRAM[32369] = 8'b0;
    XRAM[32370] = 8'b0;
    XRAM[32371] = 8'b0;
    XRAM[32372] = 8'b0;
    XRAM[32373] = 8'b0;
    XRAM[32374] = 8'b0;
    XRAM[32375] = 8'b0;
    XRAM[32376] = 8'b0;
    XRAM[32377] = 8'b0;
    XRAM[32378] = 8'b0;
    XRAM[32379] = 8'b0;
    XRAM[32380] = 8'b0;
    XRAM[32381] = 8'b0;
    XRAM[32382] = 8'b0;
    XRAM[32383] = 8'b0;
    XRAM[32384] = 8'b0;
    XRAM[32385] = 8'b0;
    XRAM[32386] = 8'b0;
    XRAM[32387] = 8'b0;
    XRAM[32388] = 8'b0;
    XRAM[32389] = 8'b0;
    XRAM[32390] = 8'b0;
    XRAM[32391] = 8'b0;
    XRAM[32392] = 8'b0;
    XRAM[32393] = 8'b0;
    XRAM[32394] = 8'b0;
    XRAM[32395] = 8'b0;
    XRAM[32396] = 8'b0;
    XRAM[32397] = 8'b0;
    XRAM[32398] = 8'b0;
    XRAM[32399] = 8'b0;
    XRAM[32400] = 8'b0;
    XRAM[32401] = 8'b0;
    XRAM[32402] = 8'b0;
    XRAM[32403] = 8'b0;
    XRAM[32404] = 8'b0;
    XRAM[32405] = 8'b0;
    XRAM[32406] = 8'b0;
    XRAM[32407] = 8'b0;
    XRAM[32408] = 8'b0;
    XRAM[32409] = 8'b0;
    XRAM[32410] = 8'b0;
    XRAM[32411] = 8'b0;
    XRAM[32412] = 8'b0;
    XRAM[32413] = 8'b0;
    XRAM[32414] = 8'b0;
    XRAM[32415] = 8'b0;
    XRAM[32416] = 8'b0;
    XRAM[32417] = 8'b0;
    XRAM[32418] = 8'b0;
    XRAM[32419] = 8'b0;
    XRAM[32420] = 8'b0;
    XRAM[32421] = 8'b0;
    XRAM[32422] = 8'b0;
    XRAM[32423] = 8'b0;
    XRAM[32424] = 8'b0;
    XRAM[32425] = 8'b0;
    XRAM[32426] = 8'b0;
    XRAM[32427] = 8'b0;
    XRAM[32428] = 8'b0;
    XRAM[32429] = 8'b0;
    XRAM[32430] = 8'b0;
    XRAM[32431] = 8'b0;
    XRAM[32432] = 8'b0;
    XRAM[32433] = 8'b0;
    XRAM[32434] = 8'b0;
    XRAM[32435] = 8'b0;
    XRAM[32436] = 8'b0;
    XRAM[32437] = 8'b0;
    XRAM[32438] = 8'b0;
    XRAM[32439] = 8'b0;
    XRAM[32440] = 8'b0;
    XRAM[32441] = 8'b0;
    XRAM[32442] = 8'b0;
    XRAM[32443] = 8'b0;
    XRAM[32444] = 8'b0;
    XRAM[32445] = 8'b0;
    XRAM[32446] = 8'b0;
    XRAM[32447] = 8'b0;
    XRAM[32448] = 8'b0;
    XRAM[32449] = 8'b0;
    XRAM[32450] = 8'b0;
    XRAM[32451] = 8'b0;
    XRAM[32452] = 8'b0;
    XRAM[32453] = 8'b0;
    XRAM[32454] = 8'b0;
    XRAM[32455] = 8'b0;
    XRAM[32456] = 8'b0;
    XRAM[32457] = 8'b0;
    XRAM[32458] = 8'b0;
    XRAM[32459] = 8'b0;
    XRAM[32460] = 8'b0;
    XRAM[32461] = 8'b0;
    XRAM[32462] = 8'b0;
    XRAM[32463] = 8'b0;
    XRAM[32464] = 8'b0;
    XRAM[32465] = 8'b0;
    XRAM[32466] = 8'b0;
    XRAM[32467] = 8'b0;
    XRAM[32468] = 8'b0;
    XRAM[32469] = 8'b0;
    XRAM[32470] = 8'b0;
    XRAM[32471] = 8'b0;
    XRAM[32472] = 8'b0;
    XRAM[32473] = 8'b0;
    XRAM[32474] = 8'b0;
    XRAM[32475] = 8'b0;
    XRAM[32476] = 8'b0;
    XRAM[32477] = 8'b0;
    XRAM[32478] = 8'b0;
    XRAM[32479] = 8'b0;
    XRAM[32480] = 8'b0;
    XRAM[32481] = 8'b0;
    XRAM[32482] = 8'b0;
    XRAM[32483] = 8'b0;
    XRAM[32484] = 8'b0;
    XRAM[32485] = 8'b0;
    XRAM[32486] = 8'b0;
    XRAM[32487] = 8'b0;
    XRAM[32488] = 8'b0;
    XRAM[32489] = 8'b0;
    XRAM[32490] = 8'b0;
    XRAM[32491] = 8'b0;
    XRAM[32492] = 8'b0;
    XRAM[32493] = 8'b0;
    XRAM[32494] = 8'b0;
    XRAM[32495] = 8'b0;
    XRAM[32496] = 8'b0;
    XRAM[32497] = 8'b0;
    XRAM[32498] = 8'b0;
    XRAM[32499] = 8'b0;
    XRAM[32500] = 8'b0;
    XRAM[32501] = 8'b0;
    XRAM[32502] = 8'b0;
    XRAM[32503] = 8'b0;
    XRAM[32504] = 8'b0;
    XRAM[32505] = 8'b0;
    XRAM[32506] = 8'b0;
    XRAM[32507] = 8'b0;
    XRAM[32508] = 8'b0;
    XRAM[32509] = 8'b0;
    XRAM[32510] = 8'b0;
    XRAM[32511] = 8'b0;
    XRAM[32512] = 8'b0;
    XRAM[32513] = 8'b0;
    XRAM[32514] = 8'b0;
    XRAM[32515] = 8'b0;
    XRAM[32516] = 8'b0;
    XRAM[32517] = 8'b0;
    XRAM[32518] = 8'b0;
    XRAM[32519] = 8'b0;
    XRAM[32520] = 8'b0;
    XRAM[32521] = 8'b0;
    XRAM[32522] = 8'b0;
    XRAM[32523] = 8'b0;
    XRAM[32524] = 8'b0;
    XRAM[32525] = 8'b0;
    XRAM[32526] = 8'b0;
    XRAM[32527] = 8'b0;
    XRAM[32528] = 8'b0;
    XRAM[32529] = 8'b0;
    XRAM[32530] = 8'b0;
    XRAM[32531] = 8'b0;
    XRAM[32532] = 8'b0;
    XRAM[32533] = 8'b0;
    XRAM[32534] = 8'b0;
    XRAM[32535] = 8'b0;
    XRAM[32536] = 8'b0;
    XRAM[32537] = 8'b0;
    XRAM[32538] = 8'b0;
    XRAM[32539] = 8'b0;
    XRAM[32540] = 8'b0;
    XRAM[32541] = 8'b0;
    XRAM[32542] = 8'b0;
    XRAM[32543] = 8'b0;
    XRAM[32544] = 8'b0;
    XRAM[32545] = 8'b0;
    XRAM[32546] = 8'b0;
    XRAM[32547] = 8'b0;
    XRAM[32548] = 8'b0;
    XRAM[32549] = 8'b0;
    XRAM[32550] = 8'b0;
    XRAM[32551] = 8'b0;
    XRAM[32552] = 8'b0;
    XRAM[32553] = 8'b0;
    XRAM[32554] = 8'b0;
    XRAM[32555] = 8'b0;
    XRAM[32556] = 8'b0;
    XRAM[32557] = 8'b0;
    XRAM[32558] = 8'b0;
    XRAM[32559] = 8'b0;
    XRAM[32560] = 8'b0;
    XRAM[32561] = 8'b0;
    XRAM[32562] = 8'b0;
    XRAM[32563] = 8'b0;
    XRAM[32564] = 8'b0;
    XRAM[32565] = 8'b0;
    XRAM[32566] = 8'b0;
    XRAM[32567] = 8'b0;
    XRAM[32568] = 8'b0;
    XRAM[32569] = 8'b0;
    XRAM[32570] = 8'b0;
    XRAM[32571] = 8'b0;
    XRAM[32572] = 8'b0;
    XRAM[32573] = 8'b0;
    XRAM[32574] = 8'b0;
    XRAM[32575] = 8'b0;
    XRAM[32576] = 8'b0;
    XRAM[32577] = 8'b0;
    XRAM[32578] = 8'b0;
    XRAM[32579] = 8'b0;
    XRAM[32580] = 8'b0;
    XRAM[32581] = 8'b0;
    XRAM[32582] = 8'b0;
    XRAM[32583] = 8'b0;
    XRAM[32584] = 8'b0;
    XRAM[32585] = 8'b0;
    XRAM[32586] = 8'b0;
    XRAM[32587] = 8'b0;
    XRAM[32588] = 8'b0;
    XRAM[32589] = 8'b0;
    XRAM[32590] = 8'b0;
    XRAM[32591] = 8'b0;
    XRAM[32592] = 8'b0;
    XRAM[32593] = 8'b0;
    XRAM[32594] = 8'b0;
    XRAM[32595] = 8'b0;
    XRAM[32596] = 8'b0;
    XRAM[32597] = 8'b0;
    XRAM[32598] = 8'b0;
    XRAM[32599] = 8'b0;
    XRAM[32600] = 8'b0;
    XRAM[32601] = 8'b0;
    XRAM[32602] = 8'b0;
    XRAM[32603] = 8'b0;
    XRAM[32604] = 8'b0;
    XRAM[32605] = 8'b0;
    XRAM[32606] = 8'b0;
    XRAM[32607] = 8'b0;
    XRAM[32608] = 8'b0;
    XRAM[32609] = 8'b0;
    XRAM[32610] = 8'b0;
    XRAM[32611] = 8'b0;
    XRAM[32612] = 8'b0;
    XRAM[32613] = 8'b0;
    XRAM[32614] = 8'b0;
    XRAM[32615] = 8'b0;
    XRAM[32616] = 8'b0;
    XRAM[32617] = 8'b0;
    XRAM[32618] = 8'b0;
    XRAM[32619] = 8'b0;
    XRAM[32620] = 8'b0;
    XRAM[32621] = 8'b0;
    XRAM[32622] = 8'b0;
    XRAM[32623] = 8'b0;
    XRAM[32624] = 8'b0;
    XRAM[32625] = 8'b0;
    XRAM[32626] = 8'b0;
    XRAM[32627] = 8'b0;
    XRAM[32628] = 8'b0;
    XRAM[32629] = 8'b0;
    XRAM[32630] = 8'b0;
    XRAM[32631] = 8'b0;
    XRAM[32632] = 8'b0;
    XRAM[32633] = 8'b0;
    XRAM[32634] = 8'b0;
    XRAM[32635] = 8'b0;
    XRAM[32636] = 8'b0;
    XRAM[32637] = 8'b0;
    XRAM[32638] = 8'b0;
    XRAM[32639] = 8'b0;
    XRAM[32640] = 8'b0;
    XRAM[32641] = 8'b0;
    XRAM[32642] = 8'b0;
    XRAM[32643] = 8'b0;
    XRAM[32644] = 8'b0;
    XRAM[32645] = 8'b0;
    XRAM[32646] = 8'b0;
    XRAM[32647] = 8'b0;
    XRAM[32648] = 8'b0;
    XRAM[32649] = 8'b0;
    XRAM[32650] = 8'b0;
    XRAM[32651] = 8'b0;
    XRAM[32652] = 8'b0;
    XRAM[32653] = 8'b0;
    XRAM[32654] = 8'b0;
    XRAM[32655] = 8'b0;
    XRAM[32656] = 8'b0;
    XRAM[32657] = 8'b0;
    XRAM[32658] = 8'b0;
    XRAM[32659] = 8'b0;
    XRAM[32660] = 8'b0;
    XRAM[32661] = 8'b0;
    XRAM[32662] = 8'b0;
    XRAM[32663] = 8'b0;
    XRAM[32664] = 8'b0;
    XRAM[32665] = 8'b0;
    XRAM[32666] = 8'b0;
    XRAM[32667] = 8'b0;
    XRAM[32668] = 8'b0;
    XRAM[32669] = 8'b0;
    XRAM[32670] = 8'b0;
    XRAM[32671] = 8'b0;
    XRAM[32672] = 8'b0;
    XRAM[32673] = 8'b0;
    XRAM[32674] = 8'b0;
    XRAM[32675] = 8'b0;
    XRAM[32676] = 8'b0;
    XRAM[32677] = 8'b0;
    XRAM[32678] = 8'b0;
    XRAM[32679] = 8'b0;
    XRAM[32680] = 8'b0;
    XRAM[32681] = 8'b0;
    XRAM[32682] = 8'b0;
    XRAM[32683] = 8'b0;
    XRAM[32684] = 8'b0;
    XRAM[32685] = 8'b0;
    XRAM[32686] = 8'b0;
    XRAM[32687] = 8'b0;
    XRAM[32688] = 8'b0;
    XRAM[32689] = 8'b0;
    XRAM[32690] = 8'b0;
    XRAM[32691] = 8'b0;
    XRAM[32692] = 8'b0;
    XRAM[32693] = 8'b0;
    XRAM[32694] = 8'b0;
    XRAM[32695] = 8'b0;
    XRAM[32696] = 8'b0;
    XRAM[32697] = 8'b0;
    XRAM[32698] = 8'b0;
    XRAM[32699] = 8'b0;
    XRAM[32700] = 8'b0;
    XRAM[32701] = 8'b0;
    XRAM[32702] = 8'b0;
    XRAM[32703] = 8'b0;
    XRAM[32704] = 8'b0;
    XRAM[32705] = 8'b0;
    XRAM[32706] = 8'b0;
    XRAM[32707] = 8'b0;
    XRAM[32708] = 8'b0;
    XRAM[32709] = 8'b0;
    XRAM[32710] = 8'b0;
    XRAM[32711] = 8'b0;
    XRAM[32712] = 8'b0;
    XRAM[32713] = 8'b0;
    XRAM[32714] = 8'b0;
    XRAM[32715] = 8'b0;
    XRAM[32716] = 8'b0;
    XRAM[32717] = 8'b0;
    XRAM[32718] = 8'b0;
    XRAM[32719] = 8'b0;
    XRAM[32720] = 8'b0;
    XRAM[32721] = 8'b0;
    XRAM[32722] = 8'b0;
    XRAM[32723] = 8'b0;
    XRAM[32724] = 8'b0;
    XRAM[32725] = 8'b0;
    XRAM[32726] = 8'b0;
    XRAM[32727] = 8'b0;
    XRAM[32728] = 8'b0;
    XRAM[32729] = 8'b0;
    XRAM[32730] = 8'b0;
    XRAM[32731] = 8'b0;
    XRAM[32732] = 8'b0;
    XRAM[32733] = 8'b0;
    XRAM[32734] = 8'b0;
    XRAM[32735] = 8'b0;
    XRAM[32736] = 8'b0;
    XRAM[32737] = 8'b0;
    XRAM[32738] = 8'b0;
    XRAM[32739] = 8'b0;
    XRAM[32740] = 8'b0;
    XRAM[32741] = 8'b0;
    XRAM[32742] = 8'b0;
    XRAM[32743] = 8'b0;
    XRAM[32744] = 8'b0;
    XRAM[32745] = 8'b0;
    XRAM[32746] = 8'b0;
    XRAM[32747] = 8'b0;
    XRAM[32748] = 8'b0;
    XRAM[32749] = 8'b0;
    XRAM[32750] = 8'b0;
    XRAM[32751] = 8'b0;
    XRAM[32752] = 8'b0;
    XRAM[32753] = 8'b0;
    XRAM[32754] = 8'b0;
    XRAM[32755] = 8'b0;
    XRAM[32756] = 8'b0;
    XRAM[32757] = 8'b0;
    XRAM[32758] = 8'b0;
    XRAM[32759] = 8'b0;
    XRAM[32760] = 8'b0;
    XRAM[32761] = 8'b0;
    XRAM[32762] = 8'b0;
    XRAM[32763] = 8'b0;
    XRAM[32764] = 8'b0;
    XRAM[32765] = 8'b0;
    XRAM[32766] = 8'b0;
    XRAM[32767] = 8'b0;
    XRAM[32768] = 8'b0;
    XRAM[32769] = 8'b0;
    XRAM[32770] = 8'b0;
    XRAM[32771] = 8'b0;
    XRAM[32772] = 8'b0;
    XRAM[32773] = 8'b0;
    XRAM[32774] = 8'b0;
    XRAM[32775] = 8'b0;
    XRAM[32776] = 8'b0;
    XRAM[32777] = 8'b0;
    XRAM[32778] = 8'b0;
    XRAM[32779] = 8'b0;
    XRAM[32780] = 8'b0;
    XRAM[32781] = 8'b0;
    XRAM[32782] = 8'b0;
    XRAM[32783] = 8'b0;
    XRAM[32784] = 8'b0;
    XRAM[32785] = 8'b0;
    XRAM[32786] = 8'b0;
    XRAM[32787] = 8'b0;
    XRAM[32788] = 8'b0;
    XRAM[32789] = 8'b0;
    XRAM[32790] = 8'b0;
    XRAM[32791] = 8'b0;
    XRAM[32792] = 8'b0;
    XRAM[32793] = 8'b0;
    XRAM[32794] = 8'b0;
    XRAM[32795] = 8'b0;
    XRAM[32796] = 8'b0;
    XRAM[32797] = 8'b0;
    XRAM[32798] = 8'b0;
    XRAM[32799] = 8'b0;
    XRAM[32800] = 8'b0;
    XRAM[32801] = 8'b0;
    XRAM[32802] = 8'b0;
    XRAM[32803] = 8'b0;
    XRAM[32804] = 8'b0;
    XRAM[32805] = 8'b0;
    XRAM[32806] = 8'b0;
    XRAM[32807] = 8'b0;
    XRAM[32808] = 8'b0;
    XRAM[32809] = 8'b0;
    XRAM[32810] = 8'b0;
    XRAM[32811] = 8'b0;
    XRAM[32812] = 8'b0;
    XRAM[32813] = 8'b0;
    XRAM[32814] = 8'b0;
    XRAM[32815] = 8'b0;
    XRAM[32816] = 8'b0;
    XRAM[32817] = 8'b0;
    XRAM[32818] = 8'b0;
    XRAM[32819] = 8'b0;
    XRAM[32820] = 8'b0;
    XRAM[32821] = 8'b0;
    XRAM[32822] = 8'b0;
    XRAM[32823] = 8'b0;
    XRAM[32824] = 8'b0;
    XRAM[32825] = 8'b0;
    XRAM[32826] = 8'b0;
    XRAM[32827] = 8'b0;
    XRAM[32828] = 8'b0;
    XRAM[32829] = 8'b0;
    XRAM[32830] = 8'b0;
    XRAM[32831] = 8'b0;
    XRAM[32832] = 8'b0;
    XRAM[32833] = 8'b0;
    XRAM[32834] = 8'b0;
    XRAM[32835] = 8'b0;
    XRAM[32836] = 8'b0;
    XRAM[32837] = 8'b0;
    XRAM[32838] = 8'b0;
    XRAM[32839] = 8'b0;
    XRAM[32840] = 8'b0;
    XRAM[32841] = 8'b0;
    XRAM[32842] = 8'b0;
    XRAM[32843] = 8'b0;
    XRAM[32844] = 8'b0;
    XRAM[32845] = 8'b0;
    XRAM[32846] = 8'b0;
    XRAM[32847] = 8'b0;
    XRAM[32848] = 8'b0;
    XRAM[32849] = 8'b0;
    XRAM[32850] = 8'b0;
    XRAM[32851] = 8'b0;
    XRAM[32852] = 8'b0;
    XRAM[32853] = 8'b0;
    XRAM[32854] = 8'b0;
    XRAM[32855] = 8'b0;
    XRAM[32856] = 8'b0;
    XRAM[32857] = 8'b0;
    XRAM[32858] = 8'b0;
    XRAM[32859] = 8'b0;
    XRAM[32860] = 8'b0;
    XRAM[32861] = 8'b0;
    XRAM[32862] = 8'b0;
    XRAM[32863] = 8'b0;
    XRAM[32864] = 8'b0;
    XRAM[32865] = 8'b0;
    XRAM[32866] = 8'b0;
    XRAM[32867] = 8'b0;
    XRAM[32868] = 8'b0;
    XRAM[32869] = 8'b0;
    XRAM[32870] = 8'b0;
    XRAM[32871] = 8'b0;
    XRAM[32872] = 8'b0;
    XRAM[32873] = 8'b0;
    XRAM[32874] = 8'b0;
    XRAM[32875] = 8'b0;
    XRAM[32876] = 8'b0;
    XRAM[32877] = 8'b0;
    XRAM[32878] = 8'b0;
    XRAM[32879] = 8'b0;
    XRAM[32880] = 8'b0;
    XRAM[32881] = 8'b0;
    XRAM[32882] = 8'b0;
    XRAM[32883] = 8'b0;
    XRAM[32884] = 8'b0;
    XRAM[32885] = 8'b0;
    XRAM[32886] = 8'b0;
    XRAM[32887] = 8'b0;
    XRAM[32888] = 8'b0;
    XRAM[32889] = 8'b0;
    XRAM[32890] = 8'b0;
    XRAM[32891] = 8'b0;
    XRAM[32892] = 8'b0;
    XRAM[32893] = 8'b0;
    XRAM[32894] = 8'b0;
    XRAM[32895] = 8'b0;
    XRAM[32896] = 8'b0;
    XRAM[32897] = 8'b0;
    XRAM[32898] = 8'b0;
    XRAM[32899] = 8'b0;
    XRAM[32900] = 8'b0;
    XRAM[32901] = 8'b0;
    XRAM[32902] = 8'b0;
    XRAM[32903] = 8'b0;
    XRAM[32904] = 8'b0;
    XRAM[32905] = 8'b0;
    XRAM[32906] = 8'b0;
    XRAM[32907] = 8'b0;
    XRAM[32908] = 8'b0;
    XRAM[32909] = 8'b0;
    XRAM[32910] = 8'b0;
    XRAM[32911] = 8'b0;
    XRAM[32912] = 8'b0;
    XRAM[32913] = 8'b0;
    XRAM[32914] = 8'b0;
    XRAM[32915] = 8'b0;
    XRAM[32916] = 8'b0;
    XRAM[32917] = 8'b0;
    XRAM[32918] = 8'b0;
    XRAM[32919] = 8'b0;
    XRAM[32920] = 8'b0;
    XRAM[32921] = 8'b0;
    XRAM[32922] = 8'b0;
    XRAM[32923] = 8'b0;
    XRAM[32924] = 8'b0;
    XRAM[32925] = 8'b0;
    XRAM[32926] = 8'b0;
    XRAM[32927] = 8'b0;
    XRAM[32928] = 8'b0;
    XRAM[32929] = 8'b0;
    XRAM[32930] = 8'b0;
    XRAM[32931] = 8'b0;
    XRAM[32932] = 8'b0;
    XRAM[32933] = 8'b0;
    XRAM[32934] = 8'b0;
    XRAM[32935] = 8'b0;
    XRAM[32936] = 8'b0;
    XRAM[32937] = 8'b0;
    XRAM[32938] = 8'b0;
    XRAM[32939] = 8'b0;
    XRAM[32940] = 8'b0;
    XRAM[32941] = 8'b0;
    XRAM[32942] = 8'b0;
    XRAM[32943] = 8'b0;
    XRAM[32944] = 8'b0;
    XRAM[32945] = 8'b0;
    XRAM[32946] = 8'b0;
    XRAM[32947] = 8'b0;
    XRAM[32948] = 8'b0;
    XRAM[32949] = 8'b0;
    XRAM[32950] = 8'b0;
    XRAM[32951] = 8'b0;
    XRAM[32952] = 8'b0;
    XRAM[32953] = 8'b0;
    XRAM[32954] = 8'b0;
    XRAM[32955] = 8'b0;
    XRAM[32956] = 8'b0;
    XRAM[32957] = 8'b0;
    XRAM[32958] = 8'b0;
    XRAM[32959] = 8'b0;
    XRAM[32960] = 8'b0;
    XRAM[32961] = 8'b0;
    XRAM[32962] = 8'b0;
    XRAM[32963] = 8'b0;
    XRAM[32964] = 8'b0;
    XRAM[32965] = 8'b0;
    XRAM[32966] = 8'b0;
    XRAM[32967] = 8'b0;
    XRAM[32968] = 8'b0;
    XRAM[32969] = 8'b0;
    XRAM[32970] = 8'b0;
    XRAM[32971] = 8'b0;
    XRAM[32972] = 8'b0;
    XRAM[32973] = 8'b0;
    XRAM[32974] = 8'b0;
    XRAM[32975] = 8'b0;
    XRAM[32976] = 8'b0;
    XRAM[32977] = 8'b0;
    XRAM[32978] = 8'b0;
    XRAM[32979] = 8'b0;
    XRAM[32980] = 8'b0;
    XRAM[32981] = 8'b0;
    XRAM[32982] = 8'b0;
    XRAM[32983] = 8'b0;
    XRAM[32984] = 8'b0;
    XRAM[32985] = 8'b0;
    XRAM[32986] = 8'b0;
    XRAM[32987] = 8'b0;
    XRAM[32988] = 8'b0;
    XRAM[32989] = 8'b0;
    XRAM[32990] = 8'b0;
    XRAM[32991] = 8'b0;
    XRAM[32992] = 8'b0;
    XRAM[32993] = 8'b0;
    XRAM[32994] = 8'b0;
    XRAM[32995] = 8'b0;
    XRAM[32996] = 8'b0;
    XRAM[32997] = 8'b0;
    XRAM[32998] = 8'b0;
    XRAM[32999] = 8'b0;
    XRAM[33000] = 8'b0;
    XRAM[33001] = 8'b0;
    XRAM[33002] = 8'b0;
    XRAM[33003] = 8'b0;
    XRAM[33004] = 8'b0;
    XRAM[33005] = 8'b0;
    XRAM[33006] = 8'b0;
    XRAM[33007] = 8'b0;
    XRAM[33008] = 8'b0;
    XRAM[33009] = 8'b0;
    XRAM[33010] = 8'b0;
    XRAM[33011] = 8'b0;
    XRAM[33012] = 8'b0;
    XRAM[33013] = 8'b0;
    XRAM[33014] = 8'b0;
    XRAM[33015] = 8'b0;
    XRAM[33016] = 8'b0;
    XRAM[33017] = 8'b0;
    XRAM[33018] = 8'b0;
    XRAM[33019] = 8'b0;
    XRAM[33020] = 8'b0;
    XRAM[33021] = 8'b0;
    XRAM[33022] = 8'b0;
    XRAM[33023] = 8'b0;
    XRAM[33024] = 8'b0;
    XRAM[33025] = 8'b0;
    XRAM[33026] = 8'b0;
    XRAM[33027] = 8'b0;
    XRAM[33028] = 8'b0;
    XRAM[33029] = 8'b0;
    XRAM[33030] = 8'b0;
    XRAM[33031] = 8'b0;
    XRAM[33032] = 8'b0;
    XRAM[33033] = 8'b0;
    XRAM[33034] = 8'b0;
    XRAM[33035] = 8'b0;
    XRAM[33036] = 8'b0;
    XRAM[33037] = 8'b0;
    XRAM[33038] = 8'b0;
    XRAM[33039] = 8'b0;
    XRAM[33040] = 8'b0;
    XRAM[33041] = 8'b0;
    XRAM[33042] = 8'b0;
    XRAM[33043] = 8'b0;
    XRAM[33044] = 8'b0;
    XRAM[33045] = 8'b0;
    XRAM[33046] = 8'b0;
    XRAM[33047] = 8'b0;
    XRAM[33048] = 8'b0;
    XRAM[33049] = 8'b0;
    XRAM[33050] = 8'b0;
    XRAM[33051] = 8'b0;
    XRAM[33052] = 8'b0;
    XRAM[33053] = 8'b0;
    XRAM[33054] = 8'b0;
    XRAM[33055] = 8'b0;
    XRAM[33056] = 8'b0;
    XRAM[33057] = 8'b0;
    XRAM[33058] = 8'b0;
    XRAM[33059] = 8'b0;
    XRAM[33060] = 8'b0;
    XRAM[33061] = 8'b0;
    XRAM[33062] = 8'b0;
    XRAM[33063] = 8'b0;
    XRAM[33064] = 8'b0;
    XRAM[33065] = 8'b0;
    XRAM[33066] = 8'b0;
    XRAM[33067] = 8'b0;
    XRAM[33068] = 8'b0;
    XRAM[33069] = 8'b0;
    XRAM[33070] = 8'b0;
    XRAM[33071] = 8'b0;
    XRAM[33072] = 8'b0;
    XRAM[33073] = 8'b0;
    XRAM[33074] = 8'b0;
    XRAM[33075] = 8'b0;
    XRAM[33076] = 8'b0;
    XRAM[33077] = 8'b0;
    XRAM[33078] = 8'b0;
    XRAM[33079] = 8'b0;
    XRAM[33080] = 8'b0;
    XRAM[33081] = 8'b0;
    XRAM[33082] = 8'b0;
    XRAM[33083] = 8'b0;
    XRAM[33084] = 8'b0;
    XRAM[33085] = 8'b0;
    XRAM[33086] = 8'b0;
    XRAM[33087] = 8'b0;
    XRAM[33088] = 8'b0;
    XRAM[33089] = 8'b0;
    XRAM[33090] = 8'b0;
    XRAM[33091] = 8'b0;
    XRAM[33092] = 8'b0;
    XRAM[33093] = 8'b0;
    XRAM[33094] = 8'b0;
    XRAM[33095] = 8'b0;
    XRAM[33096] = 8'b0;
    XRAM[33097] = 8'b0;
    XRAM[33098] = 8'b0;
    XRAM[33099] = 8'b0;
    XRAM[33100] = 8'b0;
    XRAM[33101] = 8'b0;
    XRAM[33102] = 8'b0;
    XRAM[33103] = 8'b0;
    XRAM[33104] = 8'b0;
    XRAM[33105] = 8'b0;
    XRAM[33106] = 8'b0;
    XRAM[33107] = 8'b0;
    XRAM[33108] = 8'b0;
    XRAM[33109] = 8'b0;
    XRAM[33110] = 8'b0;
    XRAM[33111] = 8'b0;
    XRAM[33112] = 8'b0;
    XRAM[33113] = 8'b0;
    XRAM[33114] = 8'b0;
    XRAM[33115] = 8'b0;
    XRAM[33116] = 8'b0;
    XRAM[33117] = 8'b0;
    XRAM[33118] = 8'b0;
    XRAM[33119] = 8'b0;
    XRAM[33120] = 8'b0;
    XRAM[33121] = 8'b0;
    XRAM[33122] = 8'b0;
    XRAM[33123] = 8'b0;
    XRAM[33124] = 8'b0;
    XRAM[33125] = 8'b0;
    XRAM[33126] = 8'b0;
    XRAM[33127] = 8'b0;
    XRAM[33128] = 8'b0;
    XRAM[33129] = 8'b0;
    XRAM[33130] = 8'b0;
    XRAM[33131] = 8'b0;
    XRAM[33132] = 8'b0;
    XRAM[33133] = 8'b0;
    XRAM[33134] = 8'b0;
    XRAM[33135] = 8'b0;
    XRAM[33136] = 8'b0;
    XRAM[33137] = 8'b0;
    XRAM[33138] = 8'b0;
    XRAM[33139] = 8'b0;
    XRAM[33140] = 8'b0;
    XRAM[33141] = 8'b0;
    XRAM[33142] = 8'b0;
    XRAM[33143] = 8'b0;
    XRAM[33144] = 8'b0;
    XRAM[33145] = 8'b0;
    XRAM[33146] = 8'b0;
    XRAM[33147] = 8'b0;
    XRAM[33148] = 8'b0;
    XRAM[33149] = 8'b0;
    XRAM[33150] = 8'b0;
    XRAM[33151] = 8'b0;
    XRAM[33152] = 8'b0;
    XRAM[33153] = 8'b0;
    XRAM[33154] = 8'b0;
    XRAM[33155] = 8'b0;
    XRAM[33156] = 8'b0;
    XRAM[33157] = 8'b0;
    XRAM[33158] = 8'b0;
    XRAM[33159] = 8'b0;
    XRAM[33160] = 8'b0;
    XRAM[33161] = 8'b0;
    XRAM[33162] = 8'b0;
    XRAM[33163] = 8'b0;
    XRAM[33164] = 8'b0;
    XRAM[33165] = 8'b0;
    XRAM[33166] = 8'b0;
    XRAM[33167] = 8'b0;
    XRAM[33168] = 8'b0;
    XRAM[33169] = 8'b0;
    XRAM[33170] = 8'b0;
    XRAM[33171] = 8'b0;
    XRAM[33172] = 8'b0;
    XRAM[33173] = 8'b0;
    XRAM[33174] = 8'b0;
    XRAM[33175] = 8'b0;
    XRAM[33176] = 8'b0;
    XRAM[33177] = 8'b0;
    XRAM[33178] = 8'b0;
    XRAM[33179] = 8'b0;
    XRAM[33180] = 8'b0;
    XRAM[33181] = 8'b0;
    XRAM[33182] = 8'b0;
    XRAM[33183] = 8'b0;
    XRAM[33184] = 8'b0;
    XRAM[33185] = 8'b0;
    XRAM[33186] = 8'b0;
    XRAM[33187] = 8'b0;
    XRAM[33188] = 8'b0;
    XRAM[33189] = 8'b0;
    XRAM[33190] = 8'b0;
    XRAM[33191] = 8'b0;
    XRAM[33192] = 8'b0;
    XRAM[33193] = 8'b0;
    XRAM[33194] = 8'b0;
    XRAM[33195] = 8'b0;
    XRAM[33196] = 8'b0;
    XRAM[33197] = 8'b0;
    XRAM[33198] = 8'b0;
    XRAM[33199] = 8'b0;
    XRAM[33200] = 8'b0;
    XRAM[33201] = 8'b0;
    XRAM[33202] = 8'b0;
    XRAM[33203] = 8'b0;
    XRAM[33204] = 8'b0;
    XRAM[33205] = 8'b0;
    XRAM[33206] = 8'b0;
    XRAM[33207] = 8'b0;
    XRAM[33208] = 8'b0;
    XRAM[33209] = 8'b0;
    XRAM[33210] = 8'b0;
    XRAM[33211] = 8'b0;
    XRAM[33212] = 8'b0;
    XRAM[33213] = 8'b0;
    XRAM[33214] = 8'b0;
    XRAM[33215] = 8'b0;
    XRAM[33216] = 8'b0;
    XRAM[33217] = 8'b0;
    XRAM[33218] = 8'b0;
    XRAM[33219] = 8'b0;
    XRAM[33220] = 8'b0;
    XRAM[33221] = 8'b0;
    XRAM[33222] = 8'b0;
    XRAM[33223] = 8'b0;
    XRAM[33224] = 8'b0;
    XRAM[33225] = 8'b0;
    XRAM[33226] = 8'b0;
    XRAM[33227] = 8'b0;
    XRAM[33228] = 8'b0;
    XRAM[33229] = 8'b0;
    XRAM[33230] = 8'b0;
    XRAM[33231] = 8'b0;
    XRAM[33232] = 8'b0;
    XRAM[33233] = 8'b0;
    XRAM[33234] = 8'b0;
    XRAM[33235] = 8'b0;
    XRAM[33236] = 8'b0;
    XRAM[33237] = 8'b0;
    XRAM[33238] = 8'b0;
    XRAM[33239] = 8'b0;
    XRAM[33240] = 8'b0;
    XRAM[33241] = 8'b0;
    XRAM[33242] = 8'b0;
    XRAM[33243] = 8'b0;
    XRAM[33244] = 8'b0;
    XRAM[33245] = 8'b0;
    XRAM[33246] = 8'b0;
    XRAM[33247] = 8'b0;
    XRAM[33248] = 8'b0;
    XRAM[33249] = 8'b0;
    XRAM[33250] = 8'b0;
    XRAM[33251] = 8'b0;
    XRAM[33252] = 8'b0;
    XRAM[33253] = 8'b0;
    XRAM[33254] = 8'b0;
    XRAM[33255] = 8'b0;
    XRAM[33256] = 8'b0;
    XRAM[33257] = 8'b0;
    XRAM[33258] = 8'b0;
    XRAM[33259] = 8'b0;
    XRAM[33260] = 8'b0;
    XRAM[33261] = 8'b0;
    XRAM[33262] = 8'b0;
    XRAM[33263] = 8'b0;
    XRAM[33264] = 8'b0;
    XRAM[33265] = 8'b0;
    XRAM[33266] = 8'b0;
    XRAM[33267] = 8'b0;
    XRAM[33268] = 8'b0;
    XRAM[33269] = 8'b0;
    XRAM[33270] = 8'b0;
    XRAM[33271] = 8'b0;
    XRAM[33272] = 8'b0;
    XRAM[33273] = 8'b0;
    XRAM[33274] = 8'b0;
    XRAM[33275] = 8'b0;
    XRAM[33276] = 8'b0;
    XRAM[33277] = 8'b0;
    XRAM[33278] = 8'b0;
    XRAM[33279] = 8'b0;
    XRAM[33280] = 8'b0;
    XRAM[33281] = 8'b0;
    XRAM[33282] = 8'b0;
    XRAM[33283] = 8'b0;
    XRAM[33284] = 8'b0;
    XRAM[33285] = 8'b0;
    XRAM[33286] = 8'b0;
    XRAM[33287] = 8'b0;
    XRAM[33288] = 8'b0;
    XRAM[33289] = 8'b0;
    XRAM[33290] = 8'b0;
    XRAM[33291] = 8'b0;
    XRAM[33292] = 8'b0;
    XRAM[33293] = 8'b0;
    XRAM[33294] = 8'b0;
    XRAM[33295] = 8'b0;
    XRAM[33296] = 8'b0;
    XRAM[33297] = 8'b0;
    XRAM[33298] = 8'b0;
    XRAM[33299] = 8'b0;
    XRAM[33300] = 8'b0;
    XRAM[33301] = 8'b0;
    XRAM[33302] = 8'b0;
    XRAM[33303] = 8'b0;
    XRAM[33304] = 8'b0;
    XRAM[33305] = 8'b0;
    XRAM[33306] = 8'b0;
    XRAM[33307] = 8'b0;
    XRAM[33308] = 8'b0;
    XRAM[33309] = 8'b0;
    XRAM[33310] = 8'b0;
    XRAM[33311] = 8'b0;
    XRAM[33312] = 8'b0;
    XRAM[33313] = 8'b0;
    XRAM[33314] = 8'b0;
    XRAM[33315] = 8'b0;
    XRAM[33316] = 8'b0;
    XRAM[33317] = 8'b0;
    XRAM[33318] = 8'b0;
    XRAM[33319] = 8'b0;
    XRAM[33320] = 8'b0;
    XRAM[33321] = 8'b0;
    XRAM[33322] = 8'b0;
    XRAM[33323] = 8'b0;
    XRAM[33324] = 8'b0;
    XRAM[33325] = 8'b0;
    XRAM[33326] = 8'b0;
    XRAM[33327] = 8'b0;
    XRAM[33328] = 8'b0;
    XRAM[33329] = 8'b0;
    XRAM[33330] = 8'b0;
    XRAM[33331] = 8'b0;
    XRAM[33332] = 8'b0;
    XRAM[33333] = 8'b0;
    XRAM[33334] = 8'b0;
    XRAM[33335] = 8'b0;
    XRAM[33336] = 8'b0;
    XRAM[33337] = 8'b0;
    XRAM[33338] = 8'b0;
    XRAM[33339] = 8'b0;
    XRAM[33340] = 8'b0;
    XRAM[33341] = 8'b0;
    XRAM[33342] = 8'b0;
    XRAM[33343] = 8'b0;
    XRAM[33344] = 8'b0;
    XRAM[33345] = 8'b0;
    XRAM[33346] = 8'b0;
    XRAM[33347] = 8'b0;
    XRAM[33348] = 8'b0;
    XRAM[33349] = 8'b0;
    XRAM[33350] = 8'b0;
    XRAM[33351] = 8'b0;
    XRAM[33352] = 8'b0;
    XRAM[33353] = 8'b0;
    XRAM[33354] = 8'b0;
    XRAM[33355] = 8'b0;
    XRAM[33356] = 8'b0;
    XRAM[33357] = 8'b0;
    XRAM[33358] = 8'b0;
    XRAM[33359] = 8'b0;
    XRAM[33360] = 8'b0;
    XRAM[33361] = 8'b0;
    XRAM[33362] = 8'b0;
    XRAM[33363] = 8'b0;
    XRAM[33364] = 8'b0;
    XRAM[33365] = 8'b0;
    XRAM[33366] = 8'b0;
    XRAM[33367] = 8'b0;
    XRAM[33368] = 8'b0;
    XRAM[33369] = 8'b0;
    XRAM[33370] = 8'b0;
    XRAM[33371] = 8'b0;
    XRAM[33372] = 8'b0;
    XRAM[33373] = 8'b0;
    XRAM[33374] = 8'b0;
    XRAM[33375] = 8'b0;
    XRAM[33376] = 8'b0;
    XRAM[33377] = 8'b0;
    XRAM[33378] = 8'b0;
    XRAM[33379] = 8'b0;
    XRAM[33380] = 8'b0;
    XRAM[33381] = 8'b0;
    XRAM[33382] = 8'b0;
    XRAM[33383] = 8'b0;
    XRAM[33384] = 8'b0;
    XRAM[33385] = 8'b0;
    XRAM[33386] = 8'b0;
    XRAM[33387] = 8'b0;
    XRAM[33388] = 8'b0;
    XRAM[33389] = 8'b0;
    XRAM[33390] = 8'b0;
    XRAM[33391] = 8'b0;
    XRAM[33392] = 8'b0;
    XRAM[33393] = 8'b0;
    XRAM[33394] = 8'b0;
    XRAM[33395] = 8'b0;
    XRAM[33396] = 8'b0;
    XRAM[33397] = 8'b0;
    XRAM[33398] = 8'b0;
    XRAM[33399] = 8'b0;
    XRAM[33400] = 8'b0;
    XRAM[33401] = 8'b0;
    XRAM[33402] = 8'b0;
    XRAM[33403] = 8'b0;
    XRAM[33404] = 8'b0;
    XRAM[33405] = 8'b0;
    XRAM[33406] = 8'b0;
    XRAM[33407] = 8'b0;
    XRAM[33408] = 8'b0;
    XRAM[33409] = 8'b0;
    XRAM[33410] = 8'b0;
    XRAM[33411] = 8'b0;
    XRAM[33412] = 8'b0;
    XRAM[33413] = 8'b0;
    XRAM[33414] = 8'b0;
    XRAM[33415] = 8'b0;
    XRAM[33416] = 8'b0;
    XRAM[33417] = 8'b0;
    XRAM[33418] = 8'b0;
    XRAM[33419] = 8'b0;
    XRAM[33420] = 8'b0;
    XRAM[33421] = 8'b0;
    XRAM[33422] = 8'b0;
    XRAM[33423] = 8'b0;
    XRAM[33424] = 8'b0;
    XRAM[33425] = 8'b0;
    XRAM[33426] = 8'b0;
    XRAM[33427] = 8'b0;
    XRAM[33428] = 8'b0;
    XRAM[33429] = 8'b0;
    XRAM[33430] = 8'b0;
    XRAM[33431] = 8'b0;
    XRAM[33432] = 8'b0;
    XRAM[33433] = 8'b0;
    XRAM[33434] = 8'b0;
    XRAM[33435] = 8'b0;
    XRAM[33436] = 8'b0;
    XRAM[33437] = 8'b0;
    XRAM[33438] = 8'b0;
    XRAM[33439] = 8'b0;
    XRAM[33440] = 8'b0;
    XRAM[33441] = 8'b0;
    XRAM[33442] = 8'b0;
    XRAM[33443] = 8'b0;
    XRAM[33444] = 8'b0;
    XRAM[33445] = 8'b0;
    XRAM[33446] = 8'b0;
    XRAM[33447] = 8'b0;
    XRAM[33448] = 8'b0;
    XRAM[33449] = 8'b0;
    XRAM[33450] = 8'b0;
    XRAM[33451] = 8'b0;
    XRAM[33452] = 8'b0;
    XRAM[33453] = 8'b0;
    XRAM[33454] = 8'b0;
    XRAM[33455] = 8'b0;
    XRAM[33456] = 8'b0;
    XRAM[33457] = 8'b0;
    XRAM[33458] = 8'b0;
    XRAM[33459] = 8'b0;
    XRAM[33460] = 8'b0;
    XRAM[33461] = 8'b0;
    XRAM[33462] = 8'b0;
    XRAM[33463] = 8'b0;
    XRAM[33464] = 8'b0;
    XRAM[33465] = 8'b0;
    XRAM[33466] = 8'b0;
    XRAM[33467] = 8'b0;
    XRAM[33468] = 8'b0;
    XRAM[33469] = 8'b0;
    XRAM[33470] = 8'b0;
    XRAM[33471] = 8'b0;
    XRAM[33472] = 8'b0;
    XRAM[33473] = 8'b0;
    XRAM[33474] = 8'b0;
    XRAM[33475] = 8'b0;
    XRAM[33476] = 8'b0;
    XRAM[33477] = 8'b0;
    XRAM[33478] = 8'b0;
    XRAM[33479] = 8'b0;
    XRAM[33480] = 8'b0;
    XRAM[33481] = 8'b0;
    XRAM[33482] = 8'b0;
    XRAM[33483] = 8'b0;
    XRAM[33484] = 8'b0;
    XRAM[33485] = 8'b0;
    XRAM[33486] = 8'b0;
    XRAM[33487] = 8'b0;
    XRAM[33488] = 8'b0;
    XRAM[33489] = 8'b0;
    XRAM[33490] = 8'b0;
    XRAM[33491] = 8'b0;
    XRAM[33492] = 8'b0;
    XRAM[33493] = 8'b0;
    XRAM[33494] = 8'b0;
    XRAM[33495] = 8'b0;
    XRAM[33496] = 8'b0;
    XRAM[33497] = 8'b0;
    XRAM[33498] = 8'b0;
    XRAM[33499] = 8'b0;
    XRAM[33500] = 8'b0;
    XRAM[33501] = 8'b0;
    XRAM[33502] = 8'b0;
    XRAM[33503] = 8'b0;
    XRAM[33504] = 8'b0;
    XRAM[33505] = 8'b0;
    XRAM[33506] = 8'b0;
    XRAM[33507] = 8'b0;
    XRAM[33508] = 8'b0;
    XRAM[33509] = 8'b0;
    XRAM[33510] = 8'b0;
    XRAM[33511] = 8'b0;
    XRAM[33512] = 8'b0;
    XRAM[33513] = 8'b0;
    XRAM[33514] = 8'b0;
    XRAM[33515] = 8'b0;
    XRAM[33516] = 8'b0;
    XRAM[33517] = 8'b0;
    XRAM[33518] = 8'b0;
    XRAM[33519] = 8'b0;
    XRAM[33520] = 8'b0;
    XRAM[33521] = 8'b0;
    XRAM[33522] = 8'b0;
    XRAM[33523] = 8'b0;
    XRAM[33524] = 8'b0;
    XRAM[33525] = 8'b0;
    XRAM[33526] = 8'b0;
    XRAM[33527] = 8'b0;
    XRAM[33528] = 8'b0;
    XRAM[33529] = 8'b0;
    XRAM[33530] = 8'b0;
    XRAM[33531] = 8'b0;
    XRAM[33532] = 8'b0;
    XRAM[33533] = 8'b0;
    XRAM[33534] = 8'b0;
    XRAM[33535] = 8'b0;
    XRAM[33536] = 8'b0;
    XRAM[33537] = 8'b0;
    XRAM[33538] = 8'b0;
    XRAM[33539] = 8'b0;
    XRAM[33540] = 8'b0;
    XRAM[33541] = 8'b0;
    XRAM[33542] = 8'b0;
    XRAM[33543] = 8'b0;
    XRAM[33544] = 8'b0;
    XRAM[33545] = 8'b0;
    XRAM[33546] = 8'b0;
    XRAM[33547] = 8'b0;
    XRAM[33548] = 8'b0;
    XRAM[33549] = 8'b0;
    XRAM[33550] = 8'b0;
    XRAM[33551] = 8'b0;
    XRAM[33552] = 8'b0;
    XRAM[33553] = 8'b0;
    XRAM[33554] = 8'b0;
    XRAM[33555] = 8'b0;
    XRAM[33556] = 8'b0;
    XRAM[33557] = 8'b0;
    XRAM[33558] = 8'b0;
    XRAM[33559] = 8'b0;
    XRAM[33560] = 8'b0;
    XRAM[33561] = 8'b0;
    XRAM[33562] = 8'b0;
    XRAM[33563] = 8'b0;
    XRAM[33564] = 8'b0;
    XRAM[33565] = 8'b0;
    XRAM[33566] = 8'b0;
    XRAM[33567] = 8'b0;
    XRAM[33568] = 8'b0;
    XRAM[33569] = 8'b0;
    XRAM[33570] = 8'b0;
    XRAM[33571] = 8'b0;
    XRAM[33572] = 8'b0;
    XRAM[33573] = 8'b0;
    XRAM[33574] = 8'b0;
    XRAM[33575] = 8'b0;
    XRAM[33576] = 8'b0;
    XRAM[33577] = 8'b0;
    XRAM[33578] = 8'b0;
    XRAM[33579] = 8'b0;
    XRAM[33580] = 8'b0;
    XRAM[33581] = 8'b0;
    XRAM[33582] = 8'b0;
    XRAM[33583] = 8'b0;
    XRAM[33584] = 8'b0;
    XRAM[33585] = 8'b0;
    XRAM[33586] = 8'b0;
    XRAM[33587] = 8'b0;
    XRAM[33588] = 8'b0;
    XRAM[33589] = 8'b0;
    XRAM[33590] = 8'b0;
    XRAM[33591] = 8'b0;
    XRAM[33592] = 8'b0;
    XRAM[33593] = 8'b0;
    XRAM[33594] = 8'b0;
    XRAM[33595] = 8'b0;
    XRAM[33596] = 8'b0;
    XRAM[33597] = 8'b0;
    XRAM[33598] = 8'b0;
    XRAM[33599] = 8'b0;
    XRAM[33600] = 8'b0;
    XRAM[33601] = 8'b0;
    XRAM[33602] = 8'b0;
    XRAM[33603] = 8'b0;
    XRAM[33604] = 8'b0;
    XRAM[33605] = 8'b0;
    XRAM[33606] = 8'b0;
    XRAM[33607] = 8'b0;
    XRAM[33608] = 8'b0;
    XRAM[33609] = 8'b0;
    XRAM[33610] = 8'b0;
    XRAM[33611] = 8'b0;
    XRAM[33612] = 8'b0;
    XRAM[33613] = 8'b0;
    XRAM[33614] = 8'b0;
    XRAM[33615] = 8'b0;
    XRAM[33616] = 8'b0;
    XRAM[33617] = 8'b0;
    XRAM[33618] = 8'b0;
    XRAM[33619] = 8'b0;
    XRAM[33620] = 8'b0;
    XRAM[33621] = 8'b0;
    XRAM[33622] = 8'b0;
    XRAM[33623] = 8'b0;
    XRAM[33624] = 8'b0;
    XRAM[33625] = 8'b0;
    XRAM[33626] = 8'b0;
    XRAM[33627] = 8'b0;
    XRAM[33628] = 8'b0;
    XRAM[33629] = 8'b0;
    XRAM[33630] = 8'b0;
    XRAM[33631] = 8'b0;
    XRAM[33632] = 8'b0;
    XRAM[33633] = 8'b0;
    XRAM[33634] = 8'b0;
    XRAM[33635] = 8'b0;
    XRAM[33636] = 8'b0;
    XRAM[33637] = 8'b0;
    XRAM[33638] = 8'b0;
    XRAM[33639] = 8'b0;
    XRAM[33640] = 8'b0;
    XRAM[33641] = 8'b0;
    XRAM[33642] = 8'b0;
    XRAM[33643] = 8'b0;
    XRAM[33644] = 8'b0;
    XRAM[33645] = 8'b0;
    XRAM[33646] = 8'b0;
    XRAM[33647] = 8'b0;
    XRAM[33648] = 8'b0;
    XRAM[33649] = 8'b0;
    XRAM[33650] = 8'b0;
    XRAM[33651] = 8'b0;
    XRAM[33652] = 8'b0;
    XRAM[33653] = 8'b0;
    XRAM[33654] = 8'b0;
    XRAM[33655] = 8'b0;
    XRAM[33656] = 8'b0;
    XRAM[33657] = 8'b0;
    XRAM[33658] = 8'b0;
    XRAM[33659] = 8'b0;
    XRAM[33660] = 8'b0;
    XRAM[33661] = 8'b0;
    XRAM[33662] = 8'b0;
    XRAM[33663] = 8'b0;
    XRAM[33664] = 8'b0;
    XRAM[33665] = 8'b0;
    XRAM[33666] = 8'b0;
    XRAM[33667] = 8'b0;
    XRAM[33668] = 8'b0;
    XRAM[33669] = 8'b0;
    XRAM[33670] = 8'b0;
    XRAM[33671] = 8'b0;
    XRAM[33672] = 8'b0;
    XRAM[33673] = 8'b0;
    XRAM[33674] = 8'b0;
    XRAM[33675] = 8'b0;
    XRAM[33676] = 8'b0;
    XRAM[33677] = 8'b0;
    XRAM[33678] = 8'b0;
    XRAM[33679] = 8'b0;
    XRAM[33680] = 8'b0;
    XRAM[33681] = 8'b0;
    XRAM[33682] = 8'b0;
    XRAM[33683] = 8'b0;
    XRAM[33684] = 8'b0;
    XRAM[33685] = 8'b0;
    XRAM[33686] = 8'b0;
    XRAM[33687] = 8'b0;
    XRAM[33688] = 8'b0;
    XRAM[33689] = 8'b0;
    XRAM[33690] = 8'b0;
    XRAM[33691] = 8'b0;
    XRAM[33692] = 8'b0;
    XRAM[33693] = 8'b0;
    XRAM[33694] = 8'b0;
    XRAM[33695] = 8'b0;
    XRAM[33696] = 8'b0;
    XRAM[33697] = 8'b0;
    XRAM[33698] = 8'b0;
    XRAM[33699] = 8'b0;
    XRAM[33700] = 8'b0;
    XRAM[33701] = 8'b0;
    XRAM[33702] = 8'b0;
    XRAM[33703] = 8'b0;
    XRAM[33704] = 8'b0;
    XRAM[33705] = 8'b0;
    XRAM[33706] = 8'b0;
    XRAM[33707] = 8'b0;
    XRAM[33708] = 8'b0;
    XRAM[33709] = 8'b0;
    XRAM[33710] = 8'b0;
    XRAM[33711] = 8'b0;
    XRAM[33712] = 8'b0;
    XRAM[33713] = 8'b0;
    XRAM[33714] = 8'b0;
    XRAM[33715] = 8'b0;
    XRAM[33716] = 8'b0;
    XRAM[33717] = 8'b0;
    XRAM[33718] = 8'b0;
    XRAM[33719] = 8'b0;
    XRAM[33720] = 8'b0;
    XRAM[33721] = 8'b0;
    XRAM[33722] = 8'b0;
    XRAM[33723] = 8'b0;
    XRAM[33724] = 8'b0;
    XRAM[33725] = 8'b0;
    XRAM[33726] = 8'b0;
    XRAM[33727] = 8'b0;
    XRAM[33728] = 8'b0;
    XRAM[33729] = 8'b0;
    XRAM[33730] = 8'b0;
    XRAM[33731] = 8'b0;
    XRAM[33732] = 8'b0;
    XRAM[33733] = 8'b0;
    XRAM[33734] = 8'b0;
    XRAM[33735] = 8'b0;
    XRAM[33736] = 8'b0;
    XRAM[33737] = 8'b0;
    XRAM[33738] = 8'b0;
    XRAM[33739] = 8'b0;
    XRAM[33740] = 8'b0;
    XRAM[33741] = 8'b0;
    XRAM[33742] = 8'b0;
    XRAM[33743] = 8'b0;
    XRAM[33744] = 8'b0;
    XRAM[33745] = 8'b0;
    XRAM[33746] = 8'b0;
    XRAM[33747] = 8'b0;
    XRAM[33748] = 8'b0;
    XRAM[33749] = 8'b0;
    XRAM[33750] = 8'b0;
    XRAM[33751] = 8'b0;
    XRAM[33752] = 8'b0;
    XRAM[33753] = 8'b0;
    XRAM[33754] = 8'b0;
    XRAM[33755] = 8'b0;
    XRAM[33756] = 8'b0;
    XRAM[33757] = 8'b0;
    XRAM[33758] = 8'b0;
    XRAM[33759] = 8'b0;
    XRAM[33760] = 8'b0;
    XRAM[33761] = 8'b0;
    XRAM[33762] = 8'b0;
    XRAM[33763] = 8'b0;
    XRAM[33764] = 8'b0;
    XRAM[33765] = 8'b0;
    XRAM[33766] = 8'b0;
    XRAM[33767] = 8'b0;
    XRAM[33768] = 8'b0;
    XRAM[33769] = 8'b0;
    XRAM[33770] = 8'b0;
    XRAM[33771] = 8'b0;
    XRAM[33772] = 8'b0;
    XRAM[33773] = 8'b0;
    XRAM[33774] = 8'b0;
    XRAM[33775] = 8'b0;
    XRAM[33776] = 8'b0;
    XRAM[33777] = 8'b0;
    XRAM[33778] = 8'b0;
    XRAM[33779] = 8'b0;
    XRAM[33780] = 8'b0;
    XRAM[33781] = 8'b0;
    XRAM[33782] = 8'b0;
    XRAM[33783] = 8'b0;
    XRAM[33784] = 8'b0;
    XRAM[33785] = 8'b0;
    XRAM[33786] = 8'b0;
    XRAM[33787] = 8'b0;
    XRAM[33788] = 8'b0;
    XRAM[33789] = 8'b0;
    XRAM[33790] = 8'b0;
    XRAM[33791] = 8'b0;
    XRAM[33792] = 8'b0;
    XRAM[33793] = 8'b0;
    XRAM[33794] = 8'b0;
    XRAM[33795] = 8'b0;
    XRAM[33796] = 8'b0;
    XRAM[33797] = 8'b0;
    XRAM[33798] = 8'b0;
    XRAM[33799] = 8'b0;
    XRAM[33800] = 8'b0;
    XRAM[33801] = 8'b0;
    XRAM[33802] = 8'b0;
    XRAM[33803] = 8'b0;
    XRAM[33804] = 8'b0;
    XRAM[33805] = 8'b0;
    XRAM[33806] = 8'b0;
    XRAM[33807] = 8'b0;
    XRAM[33808] = 8'b0;
    XRAM[33809] = 8'b0;
    XRAM[33810] = 8'b0;
    XRAM[33811] = 8'b0;
    XRAM[33812] = 8'b0;
    XRAM[33813] = 8'b0;
    XRAM[33814] = 8'b0;
    XRAM[33815] = 8'b0;
    XRAM[33816] = 8'b0;
    XRAM[33817] = 8'b0;
    XRAM[33818] = 8'b0;
    XRAM[33819] = 8'b0;
    XRAM[33820] = 8'b0;
    XRAM[33821] = 8'b0;
    XRAM[33822] = 8'b0;
    XRAM[33823] = 8'b0;
    XRAM[33824] = 8'b0;
    XRAM[33825] = 8'b0;
    XRAM[33826] = 8'b0;
    XRAM[33827] = 8'b0;
    XRAM[33828] = 8'b0;
    XRAM[33829] = 8'b0;
    XRAM[33830] = 8'b0;
    XRAM[33831] = 8'b0;
    XRAM[33832] = 8'b0;
    XRAM[33833] = 8'b0;
    XRAM[33834] = 8'b0;
    XRAM[33835] = 8'b0;
    XRAM[33836] = 8'b0;
    XRAM[33837] = 8'b0;
    XRAM[33838] = 8'b0;
    XRAM[33839] = 8'b0;
    XRAM[33840] = 8'b0;
    XRAM[33841] = 8'b0;
    XRAM[33842] = 8'b0;
    XRAM[33843] = 8'b0;
    XRAM[33844] = 8'b0;
    XRAM[33845] = 8'b0;
    XRAM[33846] = 8'b0;
    XRAM[33847] = 8'b0;
    XRAM[33848] = 8'b0;
    XRAM[33849] = 8'b0;
    XRAM[33850] = 8'b0;
    XRAM[33851] = 8'b0;
    XRAM[33852] = 8'b0;
    XRAM[33853] = 8'b0;
    XRAM[33854] = 8'b0;
    XRAM[33855] = 8'b0;
    XRAM[33856] = 8'b0;
    XRAM[33857] = 8'b0;
    XRAM[33858] = 8'b0;
    XRAM[33859] = 8'b0;
    XRAM[33860] = 8'b0;
    XRAM[33861] = 8'b0;
    XRAM[33862] = 8'b0;
    XRAM[33863] = 8'b0;
    XRAM[33864] = 8'b0;
    XRAM[33865] = 8'b0;
    XRAM[33866] = 8'b0;
    XRAM[33867] = 8'b0;
    XRAM[33868] = 8'b0;
    XRAM[33869] = 8'b0;
    XRAM[33870] = 8'b0;
    XRAM[33871] = 8'b0;
    XRAM[33872] = 8'b0;
    XRAM[33873] = 8'b0;
    XRAM[33874] = 8'b0;
    XRAM[33875] = 8'b0;
    XRAM[33876] = 8'b0;
    XRAM[33877] = 8'b0;
    XRAM[33878] = 8'b0;
    XRAM[33879] = 8'b0;
    XRAM[33880] = 8'b0;
    XRAM[33881] = 8'b0;
    XRAM[33882] = 8'b0;
    XRAM[33883] = 8'b0;
    XRAM[33884] = 8'b0;
    XRAM[33885] = 8'b0;
    XRAM[33886] = 8'b0;
    XRAM[33887] = 8'b0;
    XRAM[33888] = 8'b0;
    XRAM[33889] = 8'b0;
    XRAM[33890] = 8'b0;
    XRAM[33891] = 8'b0;
    XRAM[33892] = 8'b0;
    XRAM[33893] = 8'b0;
    XRAM[33894] = 8'b0;
    XRAM[33895] = 8'b0;
    XRAM[33896] = 8'b0;
    XRAM[33897] = 8'b0;
    XRAM[33898] = 8'b0;
    XRAM[33899] = 8'b0;
    XRAM[33900] = 8'b0;
    XRAM[33901] = 8'b0;
    XRAM[33902] = 8'b0;
    XRAM[33903] = 8'b0;
    XRAM[33904] = 8'b0;
    XRAM[33905] = 8'b0;
    XRAM[33906] = 8'b0;
    XRAM[33907] = 8'b0;
    XRAM[33908] = 8'b0;
    XRAM[33909] = 8'b0;
    XRAM[33910] = 8'b0;
    XRAM[33911] = 8'b0;
    XRAM[33912] = 8'b0;
    XRAM[33913] = 8'b0;
    XRAM[33914] = 8'b0;
    XRAM[33915] = 8'b0;
    XRAM[33916] = 8'b0;
    XRAM[33917] = 8'b0;
    XRAM[33918] = 8'b0;
    XRAM[33919] = 8'b0;
    XRAM[33920] = 8'b0;
    XRAM[33921] = 8'b0;
    XRAM[33922] = 8'b0;
    XRAM[33923] = 8'b0;
    XRAM[33924] = 8'b0;
    XRAM[33925] = 8'b0;
    XRAM[33926] = 8'b0;
    XRAM[33927] = 8'b0;
    XRAM[33928] = 8'b0;
    XRAM[33929] = 8'b0;
    XRAM[33930] = 8'b0;
    XRAM[33931] = 8'b0;
    XRAM[33932] = 8'b0;
    XRAM[33933] = 8'b0;
    XRAM[33934] = 8'b0;
    XRAM[33935] = 8'b0;
    XRAM[33936] = 8'b0;
    XRAM[33937] = 8'b0;
    XRAM[33938] = 8'b0;
    XRAM[33939] = 8'b0;
    XRAM[33940] = 8'b0;
    XRAM[33941] = 8'b0;
    XRAM[33942] = 8'b0;
    XRAM[33943] = 8'b0;
    XRAM[33944] = 8'b0;
    XRAM[33945] = 8'b0;
    XRAM[33946] = 8'b0;
    XRAM[33947] = 8'b0;
    XRAM[33948] = 8'b0;
    XRAM[33949] = 8'b0;
    XRAM[33950] = 8'b0;
    XRAM[33951] = 8'b0;
    XRAM[33952] = 8'b0;
    XRAM[33953] = 8'b0;
    XRAM[33954] = 8'b0;
    XRAM[33955] = 8'b0;
    XRAM[33956] = 8'b0;
    XRAM[33957] = 8'b0;
    XRAM[33958] = 8'b0;
    XRAM[33959] = 8'b0;
    XRAM[33960] = 8'b0;
    XRAM[33961] = 8'b0;
    XRAM[33962] = 8'b0;
    XRAM[33963] = 8'b0;
    XRAM[33964] = 8'b0;
    XRAM[33965] = 8'b0;
    XRAM[33966] = 8'b0;
    XRAM[33967] = 8'b0;
    XRAM[33968] = 8'b0;
    XRAM[33969] = 8'b0;
    XRAM[33970] = 8'b0;
    XRAM[33971] = 8'b0;
    XRAM[33972] = 8'b0;
    XRAM[33973] = 8'b0;
    XRAM[33974] = 8'b0;
    XRAM[33975] = 8'b0;
    XRAM[33976] = 8'b0;
    XRAM[33977] = 8'b0;
    XRAM[33978] = 8'b0;
    XRAM[33979] = 8'b0;
    XRAM[33980] = 8'b0;
    XRAM[33981] = 8'b0;
    XRAM[33982] = 8'b0;
    XRAM[33983] = 8'b0;
    XRAM[33984] = 8'b0;
    XRAM[33985] = 8'b0;
    XRAM[33986] = 8'b0;
    XRAM[33987] = 8'b0;
    XRAM[33988] = 8'b0;
    XRAM[33989] = 8'b0;
    XRAM[33990] = 8'b0;
    XRAM[33991] = 8'b0;
    XRAM[33992] = 8'b0;
    XRAM[33993] = 8'b0;
    XRAM[33994] = 8'b0;
    XRAM[33995] = 8'b0;
    XRAM[33996] = 8'b0;
    XRAM[33997] = 8'b0;
    XRAM[33998] = 8'b0;
    XRAM[33999] = 8'b0;
    XRAM[34000] = 8'b0;
    XRAM[34001] = 8'b0;
    XRAM[34002] = 8'b0;
    XRAM[34003] = 8'b0;
    XRAM[34004] = 8'b0;
    XRAM[34005] = 8'b0;
    XRAM[34006] = 8'b0;
    XRAM[34007] = 8'b0;
    XRAM[34008] = 8'b0;
    XRAM[34009] = 8'b0;
    XRAM[34010] = 8'b0;
    XRAM[34011] = 8'b0;
    XRAM[34012] = 8'b0;
    XRAM[34013] = 8'b0;
    XRAM[34014] = 8'b0;
    XRAM[34015] = 8'b0;
    XRAM[34016] = 8'b0;
    XRAM[34017] = 8'b0;
    XRAM[34018] = 8'b0;
    XRAM[34019] = 8'b0;
    XRAM[34020] = 8'b0;
    XRAM[34021] = 8'b0;
    XRAM[34022] = 8'b0;
    XRAM[34023] = 8'b0;
    XRAM[34024] = 8'b0;
    XRAM[34025] = 8'b0;
    XRAM[34026] = 8'b0;
    XRAM[34027] = 8'b0;
    XRAM[34028] = 8'b0;
    XRAM[34029] = 8'b0;
    XRAM[34030] = 8'b0;
    XRAM[34031] = 8'b0;
    XRAM[34032] = 8'b0;
    XRAM[34033] = 8'b0;
    XRAM[34034] = 8'b0;
    XRAM[34035] = 8'b0;
    XRAM[34036] = 8'b0;
    XRAM[34037] = 8'b0;
    XRAM[34038] = 8'b0;
    XRAM[34039] = 8'b0;
    XRAM[34040] = 8'b0;
    XRAM[34041] = 8'b0;
    XRAM[34042] = 8'b0;
    XRAM[34043] = 8'b0;
    XRAM[34044] = 8'b0;
    XRAM[34045] = 8'b0;
    XRAM[34046] = 8'b0;
    XRAM[34047] = 8'b0;
    XRAM[34048] = 8'b0;
    XRAM[34049] = 8'b0;
    XRAM[34050] = 8'b0;
    XRAM[34051] = 8'b0;
    XRAM[34052] = 8'b0;
    XRAM[34053] = 8'b0;
    XRAM[34054] = 8'b0;
    XRAM[34055] = 8'b0;
    XRAM[34056] = 8'b0;
    XRAM[34057] = 8'b0;
    XRAM[34058] = 8'b0;
    XRAM[34059] = 8'b0;
    XRAM[34060] = 8'b0;
    XRAM[34061] = 8'b0;
    XRAM[34062] = 8'b0;
    XRAM[34063] = 8'b0;
    XRAM[34064] = 8'b0;
    XRAM[34065] = 8'b0;
    XRAM[34066] = 8'b0;
    XRAM[34067] = 8'b0;
    XRAM[34068] = 8'b0;
    XRAM[34069] = 8'b0;
    XRAM[34070] = 8'b0;
    XRAM[34071] = 8'b0;
    XRAM[34072] = 8'b0;
    XRAM[34073] = 8'b0;
    XRAM[34074] = 8'b0;
    XRAM[34075] = 8'b0;
    XRAM[34076] = 8'b0;
    XRAM[34077] = 8'b0;
    XRAM[34078] = 8'b0;
    XRAM[34079] = 8'b0;
    XRAM[34080] = 8'b0;
    XRAM[34081] = 8'b0;
    XRAM[34082] = 8'b0;
    XRAM[34083] = 8'b0;
    XRAM[34084] = 8'b0;
    XRAM[34085] = 8'b0;
    XRAM[34086] = 8'b0;
    XRAM[34087] = 8'b0;
    XRAM[34088] = 8'b0;
    XRAM[34089] = 8'b0;
    XRAM[34090] = 8'b0;
    XRAM[34091] = 8'b0;
    XRAM[34092] = 8'b0;
    XRAM[34093] = 8'b0;
    XRAM[34094] = 8'b0;
    XRAM[34095] = 8'b0;
    XRAM[34096] = 8'b0;
    XRAM[34097] = 8'b0;
    XRAM[34098] = 8'b0;
    XRAM[34099] = 8'b0;
    XRAM[34100] = 8'b0;
    XRAM[34101] = 8'b0;
    XRAM[34102] = 8'b0;
    XRAM[34103] = 8'b0;
    XRAM[34104] = 8'b0;
    XRAM[34105] = 8'b0;
    XRAM[34106] = 8'b0;
    XRAM[34107] = 8'b0;
    XRAM[34108] = 8'b0;
    XRAM[34109] = 8'b0;
    XRAM[34110] = 8'b0;
    XRAM[34111] = 8'b0;
    XRAM[34112] = 8'b0;
    XRAM[34113] = 8'b0;
    XRAM[34114] = 8'b0;
    XRAM[34115] = 8'b0;
    XRAM[34116] = 8'b0;
    XRAM[34117] = 8'b0;
    XRAM[34118] = 8'b0;
    XRAM[34119] = 8'b0;
    XRAM[34120] = 8'b0;
    XRAM[34121] = 8'b0;
    XRAM[34122] = 8'b0;
    XRAM[34123] = 8'b0;
    XRAM[34124] = 8'b0;
    XRAM[34125] = 8'b0;
    XRAM[34126] = 8'b0;
    XRAM[34127] = 8'b0;
    XRAM[34128] = 8'b0;
    XRAM[34129] = 8'b0;
    XRAM[34130] = 8'b0;
    XRAM[34131] = 8'b0;
    XRAM[34132] = 8'b0;
    XRAM[34133] = 8'b0;
    XRAM[34134] = 8'b0;
    XRAM[34135] = 8'b0;
    XRAM[34136] = 8'b0;
    XRAM[34137] = 8'b0;
    XRAM[34138] = 8'b0;
    XRAM[34139] = 8'b0;
    XRAM[34140] = 8'b0;
    XRAM[34141] = 8'b0;
    XRAM[34142] = 8'b0;
    XRAM[34143] = 8'b0;
    XRAM[34144] = 8'b0;
    XRAM[34145] = 8'b0;
    XRAM[34146] = 8'b0;
    XRAM[34147] = 8'b0;
    XRAM[34148] = 8'b0;
    XRAM[34149] = 8'b0;
    XRAM[34150] = 8'b0;
    XRAM[34151] = 8'b0;
    XRAM[34152] = 8'b0;
    XRAM[34153] = 8'b0;
    XRAM[34154] = 8'b0;
    XRAM[34155] = 8'b0;
    XRAM[34156] = 8'b0;
    XRAM[34157] = 8'b0;
    XRAM[34158] = 8'b0;
    XRAM[34159] = 8'b0;
    XRAM[34160] = 8'b0;
    XRAM[34161] = 8'b0;
    XRAM[34162] = 8'b0;
    XRAM[34163] = 8'b0;
    XRAM[34164] = 8'b0;
    XRAM[34165] = 8'b0;
    XRAM[34166] = 8'b0;
    XRAM[34167] = 8'b0;
    XRAM[34168] = 8'b0;
    XRAM[34169] = 8'b0;
    XRAM[34170] = 8'b0;
    XRAM[34171] = 8'b0;
    XRAM[34172] = 8'b0;
    XRAM[34173] = 8'b0;
    XRAM[34174] = 8'b0;
    XRAM[34175] = 8'b0;
    XRAM[34176] = 8'b0;
    XRAM[34177] = 8'b0;
    XRAM[34178] = 8'b0;
    XRAM[34179] = 8'b0;
    XRAM[34180] = 8'b0;
    XRAM[34181] = 8'b0;
    XRAM[34182] = 8'b0;
    XRAM[34183] = 8'b0;
    XRAM[34184] = 8'b0;
    XRAM[34185] = 8'b0;
    XRAM[34186] = 8'b0;
    XRAM[34187] = 8'b0;
    XRAM[34188] = 8'b0;
    XRAM[34189] = 8'b0;
    XRAM[34190] = 8'b0;
    XRAM[34191] = 8'b0;
    XRAM[34192] = 8'b0;
    XRAM[34193] = 8'b0;
    XRAM[34194] = 8'b0;
    XRAM[34195] = 8'b0;
    XRAM[34196] = 8'b0;
    XRAM[34197] = 8'b0;
    XRAM[34198] = 8'b0;
    XRAM[34199] = 8'b0;
    XRAM[34200] = 8'b0;
    XRAM[34201] = 8'b0;
    XRAM[34202] = 8'b0;
    XRAM[34203] = 8'b0;
    XRAM[34204] = 8'b0;
    XRAM[34205] = 8'b0;
    XRAM[34206] = 8'b0;
    XRAM[34207] = 8'b0;
    XRAM[34208] = 8'b0;
    XRAM[34209] = 8'b0;
    XRAM[34210] = 8'b0;
    XRAM[34211] = 8'b0;
    XRAM[34212] = 8'b0;
    XRAM[34213] = 8'b0;
    XRAM[34214] = 8'b0;
    XRAM[34215] = 8'b0;
    XRAM[34216] = 8'b0;
    XRAM[34217] = 8'b0;
    XRAM[34218] = 8'b0;
    XRAM[34219] = 8'b0;
    XRAM[34220] = 8'b0;
    XRAM[34221] = 8'b0;
    XRAM[34222] = 8'b0;
    XRAM[34223] = 8'b0;
    XRAM[34224] = 8'b0;
    XRAM[34225] = 8'b0;
    XRAM[34226] = 8'b0;
    XRAM[34227] = 8'b0;
    XRAM[34228] = 8'b0;
    XRAM[34229] = 8'b0;
    XRAM[34230] = 8'b0;
    XRAM[34231] = 8'b0;
    XRAM[34232] = 8'b0;
    XRAM[34233] = 8'b0;
    XRAM[34234] = 8'b0;
    XRAM[34235] = 8'b0;
    XRAM[34236] = 8'b0;
    XRAM[34237] = 8'b0;
    XRAM[34238] = 8'b0;
    XRAM[34239] = 8'b0;
    XRAM[34240] = 8'b0;
    XRAM[34241] = 8'b0;
    XRAM[34242] = 8'b0;
    XRAM[34243] = 8'b0;
    XRAM[34244] = 8'b0;
    XRAM[34245] = 8'b0;
    XRAM[34246] = 8'b0;
    XRAM[34247] = 8'b0;
    XRAM[34248] = 8'b0;
    XRAM[34249] = 8'b0;
    XRAM[34250] = 8'b0;
    XRAM[34251] = 8'b0;
    XRAM[34252] = 8'b0;
    XRAM[34253] = 8'b0;
    XRAM[34254] = 8'b0;
    XRAM[34255] = 8'b0;
    XRAM[34256] = 8'b0;
    XRAM[34257] = 8'b0;
    XRAM[34258] = 8'b0;
    XRAM[34259] = 8'b0;
    XRAM[34260] = 8'b0;
    XRAM[34261] = 8'b0;
    XRAM[34262] = 8'b0;
    XRAM[34263] = 8'b0;
    XRAM[34264] = 8'b0;
    XRAM[34265] = 8'b0;
    XRAM[34266] = 8'b0;
    XRAM[34267] = 8'b0;
    XRAM[34268] = 8'b0;
    XRAM[34269] = 8'b0;
    XRAM[34270] = 8'b0;
    XRAM[34271] = 8'b0;
    XRAM[34272] = 8'b0;
    XRAM[34273] = 8'b0;
    XRAM[34274] = 8'b0;
    XRAM[34275] = 8'b0;
    XRAM[34276] = 8'b0;
    XRAM[34277] = 8'b0;
    XRAM[34278] = 8'b0;
    XRAM[34279] = 8'b0;
    XRAM[34280] = 8'b0;
    XRAM[34281] = 8'b0;
    XRAM[34282] = 8'b0;
    XRAM[34283] = 8'b0;
    XRAM[34284] = 8'b0;
    XRAM[34285] = 8'b0;
    XRAM[34286] = 8'b0;
    XRAM[34287] = 8'b0;
    XRAM[34288] = 8'b0;
    XRAM[34289] = 8'b0;
    XRAM[34290] = 8'b0;
    XRAM[34291] = 8'b0;
    XRAM[34292] = 8'b0;
    XRAM[34293] = 8'b0;
    XRAM[34294] = 8'b0;
    XRAM[34295] = 8'b0;
    XRAM[34296] = 8'b0;
    XRAM[34297] = 8'b0;
    XRAM[34298] = 8'b0;
    XRAM[34299] = 8'b0;
    XRAM[34300] = 8'b0;
    XRAM[34301] = 8'b0;
    XRAM[34302] = 8'b0;
    XRAM[34303] = 8'b0;
    XRAM[34304] = 8'b0;
    XRAM[34305] = 8'b0;
    XRAM[34306] = 8'b0;
    XRAM[34307] = 8'b0;
    XRAM[34308] = 8'b0;
    XRAM[34309] = 8'b0;
    XRAM[34310] = 8'b0;
    XRAM[34311] = 8'b0;
    XRAM[34312] = 8'b0;
    XRAM[34313] = 8'b0;
    XRAM[34314] = 8'b0;
    XRAM[34315] = 8'b0;
    XRAM[34316] = 8'b0;
    XRAM[34317] = 8'b0;
    XRAM[34318] = 8'b0;
    XRAM[34319] = 8'b0;
    XRAM[34320] = 8'b0;
    XRAM[34321] = 8'b0;
    XRAM[34322] = 8'b0;
    XRAM[34323] = 8'b0;
    XRAM[34324] = 8'b0;
    XRAM[34325] = 8'b0;
    XRAM[34326] = 8'b0;
    XRAM[34327] = 8'b0;
    XRAM[34328] = 8'b0;
    XRAM[34329] = 8'b0;
    XRAM[34330] = 8'b0;
    XRAM[34331] = 8'b0;
    XRAM[34332] = 8'b0;
    XRAM[34333] = 8'b0;
    XRAM[34334] = 8'b0;
    XRAM[34335] = 8'b0;
    XRAM[34336] = 8'b0;
    XRAM[34337] = 8'b0;
    XRAM[34338] = 8'b0;
    XRAM[34339] = 8'b0;
    XRAM[34340] = 8'b0;
    XRAM[34341] = 8'b0;
    XRAM[34342] = 8'b0;
    XRAM[34343] = 8'b0;
    XRAM[34344] = 8'b0;
    XRAM[34345] = 8'b0;
    XRAM[34346] = 8'b0;
    XRAM[34347] = 8'b0;
    XRAM[34348] = 8'b0;
    XRAM[34349] = 8'b0;
    XRAM[34350] = 8'b0;
    XRAM[34351] = 8'b0;
    XRAM[34352] = 8'b0;
    XRAM[34353] = 8'b0;
    XRAM[34354] = 8'b0;
    XRAM[34355] = 8'b0;
    XRAM[34356] = 8'b0;
    XRAM[34357] = 8'b0;
    XRAM[34358] = 8'b0;
    XRAM[34359] = 8'b0;
    XRAM[34360] = 8'b0;
    XRAM[34361] = 8'b0;
    XRAM[34362] = 8'b0;
    XRAM[34363] = 8'b0;
    XRAM[34364] = 8'b0;
    XRAM[34365] = 8'b0;
    XRAM[34366] = 8'b0;
    XRAM[34367] = 8'b0;
    XRAM[34368] = 8'b0;
    XRAM[34369] = 8'b0;
    XRAM[34370] = 8'b0;
    XRAM[34371] = 8'b0;
    XRAM[34372] = 8'b0;
    XRAM[34373] = 8'b0;
    XRAM[34374] = 8'b0;
    XRAM[34375] = 8'b0;
    XRAM[34376] = 8'b0;
    XRAM[34377] = 8'b0;
    XRAM[34378] = 8'b0;
    XRAM[34379] = 8'b0;
    XRAM[34380] = 8'b0;
    XRAM[34381] = 8'b0;
    XRAM[34382] = 8'b0;
    XRAM[34383] = 8'b0;
    XRAM[34384] = 8'b0;
    XRAM[34385] = 8'b0;
    XRAM[34386] = 8'b0;
    XRAM[34387] = 8'b0;
    XRAM[34388] = 8'b0;
    XRAM[34389] = 8'b0;
    XRAM[34390] = 8'b0;
    XRAM[34391] = 8'b0;
    XRAM[34392] = 8'b0;
    XRAM[34393] = 8'b0;
    XRAM[34394] = 8'b0;
    XRAM[34395] = 8'b0;
    XRAM[34396] = 8'b0;
    XRAM[34397] = 8'b0;
    XRAM[34398] = 8'b0;
    XRAM[34399] = 8'b0;
    XRAM[34400] = 8'b0;
    XRAM[34401] = 8'b0;
    XRAM[34402] = 8'b0;
    XRAM[34403] = 8'b0;
    XRAM[34404] = 8'b0;
    XRAM[34405] = 8'b0;
    XRAM[34406] = 8'b0;
    XRAM[34407] = 8'b0;
    XRAM[34408] = 8'b0;
    XRAM[34409] = 8'b0;
    XRAM[34410] = 8'b0;
    XRAM[34411] = 8'b0;
    XRAM[34412] = 8'b0;
    XRAM[34413] = 8'b0;
    XRAM[34414] = 8'b0;
    XRAM[34415] = 8'b0;
    XRAM[34416] = 8'b0;
    XRAM[34417] = 8'b0;
    XRAM[34418] = 8'b0;
    XRAM[34419] = 8'b0;
    XRAM[34420] = 8'b0;
    XRAM[34421] = 8'b0;
    XRAM[34422] = 8'b0;
    XRAM[34423] = 8'b0;
    XRAM[34424] = 8'b0;
    XRAM[34425] = 8'b0;
    XRAM[34426] = 8'b0;
    XRAM[34427] = 8'b0;
    XRAM[34428] = 8'b0;
    XRAM[34429] = 8'b0;
    XRAM[34430] = 8'b0;
    XRAM[34431] = 8'b0;
    XRAM[34432] = 8'b0;
    XRAM[34433] = 8'b0;
    XRAM[34434] = 8'b0;
    XRAM[34435] = 8'b0;
    XRAM[34436] = 8'b0;
    XRAM[34437] = 8'b0;
    XRAM[34438] = 8'b0;
    XRAM[34439] = 8'b0;
    XRAM[34440] = 8'b0;
    XRAM[34441] = 8'b0;
    XRAM[34442] = 8'b0;
    XRAM[34443] = 8'b0;
    XRAM[34444] = 8'b0;
    XRAM[34445] = 8'b0;
    XRAM[34446] = 8'b0;
    XRAM[34447] = 8'b0;
    XRAM[34448] = 8'b0;
    XRAM[34449] = 8'b0;
    XRAM[34450] = 8'b0;
    XRAM[34451] = 8'b0;
    XRAM[34452] = 8'b0;
    XRAM[34453] = 8'b0;
    XRAM[34454] = 8'b0;
    XRAM[34455] = 8'b0;
    XRAM[34456] = 8'b0;
    XRAM[34457] = 8'b0;
    XRAM[34458] = 8'b0;
    XRAM[34459] = 8'b0;
    XRAM[34460] = 8'b0;
    XRAM[34461] = 8'b0;
    XRAM[34462] = 8'b0;
    XRAM[34463] = 8'b0;
    XRAM[34464] = 8'b0;
    XRAM[34465] = 8'b0;
    XRAM[34466] = 8'b0;
    XRAM[34467] = 8'b0;
    XRAM[34468] = 8'b0;
    XRAM[34469] = 8'b0;
    XRAM[34470] = 8'b0;
    XRAM[34471] = 8'b0;
    XRAM[34472] = 8'b0;
    XRAM[34473] = 8'b0;
    XRAM[34474] = 8'b0;
    XRAM[34475] = 8'b0;
    XRAM[34476] = 8'b0;
    XRAM[34477] = 8'b0;
    XRAM[34478] = 8'b0;
    XRAM[34479] = 8'b0;
    XRAM[34480] = 8'b0;
    XRAM[34481] = 8'b0;
    XRAM[34482] = 8'b0;
    XRAM[34483] = 8'b0;
    XRAM[34484] = 8'b0;
    XRAM[34485] = 8'b0;
    XRAM[34486] = 8'b0;
    XRAM[34487] = 8'b0;
    XRAM[34488] = 8'b0;
    XRAM[34489] = 8'b0;
    XRAM[34490] = 8'b0;
    XRAM[34491] = 8'b0;
    XRAM[34492] = 8'b0;
    XRAM[34493] = 8'b0;
    XRAM[34494] = 8'b0;
    XRAM[34495] = 8'b0;
    XRAM[34496] = 8'b0;
    XRAM[34497] = 8'b0;
    XRAM[34498] = 8'b0;
    XRAM[34499] = 8'b0;
    XRAM[34500] = 8'b0;
    XRAM[34501] = 8'b0;
    XRAM[34502] = 8'b0;
    XRAM[34503] = 8'b0;
    XRAM[34504] = 8'b0;
    XRAM[34505] = 8'b0;
    XRAM[34506] = 8'b0;
    XRAM[34507] = 8'b0;
    XRAM[34508] = 8'b0;
    XRAM[34509] = 8'b0;
    XRAM[34510] = 8'b0;
    XRAM[34511] = 8'b0;
    XRAM[34512] = 8'b0;
    XRAM[34513] = 8'b0;
    XRAM[34514] = 8'b0;
    XRAM[34515] = 8'b0;
    XRAM[34516] = 8'b0;
    XRAM[34517] = 8'b0;
    XRAM[34518] = 8'b0;
    XRAM[34519] = 8'b0;
    XRAM[34520] = 8'b0;
    XRAM[34521] = 8'b0;
    XRAM[34522] = 8'b0;
    XRAM[34523] = 8'b0;
    XRAM[34524] = 8'b0;
    XRAM[34525] = 8'b0;
    XRAM[34526] = 8'b0;
    XRAM[34527] = 8'b0;
    XRAM[34528] = 8'b0;
    XRAM[34529] = 8'b0;
    XRAM[34530] = 8'b0;
    XRAM[34531] = 8'b0;
    XRAM[34532] = 8'b0;
    XRAM[34533] = 8'b0;
    XRAM[34534] = 8'b0;
    XRAM[34535] = 8'b0;
    XRAM[34536] = 8'b0;
    XRAM[34537] = 8'b0;
    XRAM[34538] = 8'b0;
    XRAM[34539] = 8'b0;
    XRAM[34540] = 8'b0;
    XRAM[34541] = 8'b0;
    XRAM[34542] = 8'b0;
    XRAM[34543] = 8'b0;
    XRAM[34544] = 8'b0;
    XRAM[34545] = 8'b0;
    XRAM[34546] = 8'b0;
    XRAM[34547] = 8'b0;
    XRAM[34548] = 8'b0;
    XRAM[34549] = 8'b0;
    XRAM[34550] = 8'b0;
    XRAM[34551] = 8'b0;
    XRAM[34552] = 8'b0;
    XRAM[34553] = 8'b0;
    XRAM[34554] = 8'b0;
    XRAM[34555] = 8'b0;
    XRAM[34556] = 8'b0;
    XRAM[34557] = 8'b0;
    XRAM[34558] = 8'b0;
    XRAM[34559] = 8'b0;
    XRAM[34560] = 8'b0;
    XRAM[34561] = 8'b0;
    XRAM[34562] = 8'b0;
    XRAM[34563] = 8'b0;
    XRAM[34564] = 8'b0;
    XRAM[34565] = 8'b0;
    XRAM[34566] = 8'b0;
    XRAM[34567] = 8'b0;
    XRAM[34568] = 8'b0;
    XRAM[34569] = 8'b0;
    XRAM[34570] = 8'b0;
    XRAM[34571] = 8'b0;
    XRAM[34572] = 8'b0;
    XRAM[34573] = 8'b0;
    XRAM[34574] = 8'b0;
    XRAM[34575] = 8'b0;
    XRAM[34576] = 8'b0;
    XRAM[34577] = 8'b0;
    XRAM[34578] = 8'b0;
    XRAM[34579] = 8'b0;
    XRAM[34580] = 8'b0;
    XRAM[34581] = 8'b0;
    XRAM[34582] = 8'b0;
    XRAM[34583] = 8'b0;
    XRAM[34584] = 8'b0;
    XRAM[34585] = 8'b0;
    XRAM[34586] = 8'b0;
    XRAM[34587] = 8'b0;
    XRAM[34588] = 8'b0;
    XRAM[34589] = 8'b0;
    XRAM[34590] = 8'b0;
    XRAM[34591] = 8'b0;
    XRAM[34592] = 8'b0;
    XRAM[34593] = 8'b0;
    XRAM[34594] = 8'b0;
    XRAM[34595] = 8'b0;
    XRAM[34596] = 8'b0;
    XRAM[34597] = 8'b0;
    XRAM[34598] = 8'b0;
    XRAM[34599] = 8'b0;
    XRAM[34600] = 8'b0;
    XRAM[34601] = 8'b0;
    XRAM[34602] = 8'b0;
    XRAM[34603] = 8'b0;
    XRAM[34604] = 8'b0;
    XRAM[34605] = 8'b0;
    XRAM[34606] = 8'b0;
    XRAM[34607] = 8'b0;
    XRAM[34608] = 8'b0;
    XRAM[34609] = 8'b0;
    XRAM[34610] = 8'b0;
    XRAM[34611] = 8'b0;
    XRAM[34612] = 8'b0;
    XRAM[34613] = 8'b0;
    XRAM[34614] = 8'b0;
    XRAM[34615] = 8'b0;
    XRAM[34616] = 8'b0;
    XRAM[34617] = 8'b0;
    XRAM[34618] = 8'b0;
    XRAM[34619] = 8'b0;
    XRAM[34620] = 8'b0;
    XRAM[34621] = 8'b0;
    XRAM[34622] = 8'b0;
    XRAM[34623] = 8'b0;
    XRAM[34624] = 8'b0;
    XRAM[34625] = 8'b0;
    XRAM[34626] = 8'b0;
    XRAM[34627] = 8'b0;
    XRAM[34628] = 8'b0;
    XRAM[34629] = 8'b0;
    XRAM[34630] = 8'b0;
    XRAM[34631] = 8'b0;
    XRAM[34632] = 8'b0;
    XRAM[34633] = 8'b0;
    XRAM[34634] = 8'b0;
    XRAM[34635] = 8'b0;
    XRAM[34636] = 8'b0;
    XRAM[34637] = 8'b0;
    XRAM[34638] = 8'b0;
    XRAM[34639] = 8'b0;
    XRAM[34640] = 8'b0;
    XRAM[34641] = 8'b0;
    XRAM[34642] = 8'b0;
    XRAM[34643] = 8'b0;
    XRAM[34644] = 8'b0;
    XRAM[34645] = 8'b0;
    XRAM[34646] = 8'b0;
    XRAM[34647] = 8'b0;
    XRAM[34648] = 8'b0;
    XRAM[34649] = 8'b0;
    XRAM[34650] = 8'b0;
    XRAM[34651] = 8'b0;
    XRAM[34652] = 8'b0;
    XRAM[34653] = 8'b0;
    XRAM[34654] = 8'b0;
    XRAM[34655] = 8'b0;
    XRAM[34656] = 8'b0;
    XRAM[34657] = 8'b0;
    XRAM[34658] = 8'b0;
    XRAM[34659] = 8'b0;
    XRAM[34660] = 8'b0;
    XRAM[34661] = 8'b0;
    XRAM[34662] = 8'b0;
    XRAM[34663] = 8'b0;
    XRAM[34664] = 8'b0;
    XRAM[34665] = 8'b0;
    XRAM[34666] = 8'b0;
    XRAM[34667] = 8'b0;
    XRAM[34668] = 8'b0;
    XRAM[34669] = 8'b0;
    XRAM[34670] = 8'b0;
    XRAM[34671] = 8'b0;
    XRAM[34672] = 8'b0;
    XRAM[34673] = 8'b0;
    XRAM[34674] = 8'b0;
    XRAM[34675] = 8'b0;
    XRAM[34676] = 8'b0;
    XRAM[34677] = 8'b0;
    XRAM[34678] = 8'b0;
    XRAM[34679] = 8'b0;
    XRAM[34680] = 8'b0;
    XRAM[34681] = 8'b0;
    XRAM[34682] = 8'b0;
    XRAM[34683] = 8'b0;
    XRAM[34684] = 8'b0;
    XRAM[34685] = 8'b0;
    XRAM[34686] = 8'b0;
    XRAM[34687] = 8'b0;
    XRAM[34688] = 8'b0;
    XRAM[34689] = 8'b0;
    XRAM[34690] = 8'b0;
    XRAM[34691] = 8'b0;
    XRAM[34692] = 8'b0;
    XRAM[34693] = 8'b0;
    XRAM[34694] = 8'b0;
    XRAM[34695] = 8'b0;
    XRAM[34696] = 8'b0;
    XRAM[34697] = 8'b0;
    XRAM[34698] = 8'b0;
    XRAM[34699] = 8'b0;
    XRAM[34700] = 8'b0;
    XRAM[34701] = 8'b0;
    XRAM[34702] = 8'b0;
    XRAM[34703] = 8'b0;
    XRAM[34704] = 8'b0;
    XRAM[34705] = 8'b0;
    XRAM[34706] = 8'b0;
    XRAM[34707] = 8'b0;
    XRAM[34708] = 8'b0;
    XRAM[34709] = 8'b0;
    XRAM[34710] = 8'b0;
    XRAM[34711] = 8'b0;
    XRAM[34712] = 8'b0;
    XRAM[34713] = 8'b0;
    XRAM[34714] = 8'b0;
    XRAM[34715] = 8'b0;
    XRAM[34716] = 8'b0;
    XRAM[34717] = 8'b0;
    XRAM[34718] = 8'b0;
    XRAM[34719] = 8'b0;
    XRAM[34720] = 8'b0;
    XRAM[34721] = 8'b0;
    XRAM[34722] = 8'b0;
    XRAM[34723] = 8'b0;
    XRAM[34724] = 8'b0;
    XRAM[34725] = 8'b0;
    XRAM[34726] = 8'b0;
    XRAM[34727] = 8'b0;
    XRAM[34728] = 8'b0;
    XRAM[34729] = 8'b0;
    XRAM[34730] = 8'b0;
    XRAM[34731] = 8'b0;
    XRAM[34732] = 8'b0;
    XRAM[34733] = 8'b0;
    XRAM[34734] = 8'b0;
    XRAM[34735] = 8'b0;
    XRAM[34736] = 8'b0;
    XRAM[34737] = 8'b0;
    XRAM[34738] = 8'b0;
    XRAM[34739] = 8'b0;
    XRAM[34740] = 8'b0;
    XRAM[34741] = 8'b0;
    XRAM[34742] = 8'b0;
    XRAM[34743] = 8'b0;
    XRAM[34744] = 8'b0;
    XRAM[34745] = 8'b0;
    XRAM[34746] = 8'b0;
    XRAM[34747] = 8'b0;
    XRAM[34748] = 8'b0;
    XRAM[34749] = 8'b0;
    XRAM[34750] = 8'b0;
    XRAM[34751] = 8'b0;
    XRAM[34752] = 8'b0;
    XRAM[34753] = 8'b0;
    XRAM[34754] = 8'b0;
    XRAM[34755] = 8'b0;
    XRAM[34756] = 8'b0;
    XRAM[34757] = 8'b0;
    XRAM[34758] = 8'b0;
    XRAM[34759] = 8'b0;
    XRAM[34760] = 8'b0;
    XRAM[34761] = 8'b0;
    XRAM[34762] = 8'b0;
    XRAM[34763] = 8'b0;
    XRAM[34764] = 8'b0;
    XRAM[34765] = 8'b0;
    XRAM[34766] = 8'b0;
    XRAM[34767] = 8'b0;
    XRAM[34768] = 8'b0;
    XRAM[34769] = 8'b0;
    XRAM[34770] = 8'b0;
    XRAM[34771] = 8'b0;
    XRAM[34772] = 8'b0;
    XRAM[34773] = 8'b0;
    XRAM[34774] = 8'b0;
    XRAM[34775] = 8'b0;
    XRAM[34776] = 8'b0;
    XRAM[34777] = 8'b0;
    XRAM[34778] = 8'b0;
    XRAM[34779] = 8'b0;
    XRAM[34780] = 8'b0;
    XRAM[34781] = 8'b0;
    XRAM[34782] = 8'b0;
    XRAM[34783] = 8'b0;
    XRAM[34784] = 8'b0;
    XRAM[34785] = 8'b0;
    XRAM[34786] = 8'b0;
    XRAM[34787] = 8'b0;
    XRAM[34788] = 8'b0;
    XRAM[34789] = 8'b0;
    XRAM[34790] = 8'b0;
    XRAM[34791] = 8'b0;
    XRAM[34792] = 8'b0;
    XRAM[34793] = 8'b0;
    XRAM[34794] = 8'b0;
    XRAM[34795] = 8'b0;
    XRAM[34796] = 8'b0;
    XRAM[34797] = 8'b0;
    XRAM[34798] = 8'b0;
    XRAM[34799] = 8'b0;
    XRAM[34800] = 8'b0;
    XRAM[34801] = 8'b0;
    XRAM[34802] = 8'b0;
    XRAM[34803] = 8'b0;
    XRAM[34804] = 8'b0;
    XRAM[34805] = 8'b0;
    XRAM[34806] = 8'b0;
    XRAM[34807] = 8'b0;
    XRAM[34808] = 8'b0;
    XRAM[34809] = 8'b0;
    XRAM[34810] = 8'b0;
    XRAM[34811] = 8'b0;
    XRAM[34812] = 8'b0;
    XRAM[34813] = 8'b0;
    XRAM[34814] = 8'b0;
    XRAM[34815] = 8'b0;
    XRAM[34816] = 8'b0;
    XRAM[34817] = 8'b0;
    XRAM[34818] = 8'b0;
    XRAM[34819] = 8'b0;
    XRAM[34820] = 8'b0;
    XRAM[34821] = 8'b0;
    XRAM[34822] = 8'b0;
    XRAM[34823] = 8'b0;
    XRAM[34824] = 8'b0;
    XRAM[34825] = 8'b0;
    XRAM[34826] = 8'b0;
    XRAM[34827] = 8'b0;
    XRAM[34828] = 8'b0;
    XRAM[34829] = 8'b0;
    XRAM[34830] = 8'b0;
    XRAM[34831] = 8'b0;
    XRAM[34832] = 8'b0;
    XRAM[34833] = 8'b0;
    XRAM[34834] = 8'b0;
    XRAM[34835] = 8'b0;
    XRAM[34836] = 8'b0;
    XRAM[34837] = 8'b0;
    XRAM[34838] = 8'b0;
    XRAM[34839] = 8'b0;
    XRAM[34840] = 8'b0;
    XRAM[34841] = 8'b0;
    XRAM[34842] = 8'b0;
    XRAM[34843] = 8'b0;
    XRAM[34844] = 8'b0;
    XRAM[34845] = 8'b0;
    XRAM[34846] = 8'b0;
    XRAM[34847] = 8'b0;
    XRAM[34848] = 8'b0;
    XRAM[34849] = 8'b0;
    XRAM[34850] = 8'b0;
    XRAM[34851] = 8'b0;
    XRAM[34852] = 8'b0;
    XRAM[34853] = 8'b0;
    XRAM[34854] = 8'b0;
    XRAM[34855] = 8'b0;
    XRAM[34856] = 8'b0;
    XRAM[34857] = 8'b0;
    XRAM[34858] = 8'b0;
    XRAM[34859] = 8'b0;
    XRAM[34860] = 8'b0;
    XRAM[34861] = 8'b0;
    XRAM[34862] = 8'b0;
    XRAM[34863] = 8'b0;
    XRAM[34864] = 8'b0;
    XRAM[34865] = 8'b0;
    XRAM[34866] = 8'b0;
    XRAM[34867] = 8'b0;
    XRAM[34868] = 8'b0;
    XRAM[34869] = 8'b0;
    XRAM[34870] = 8'b0;
    XRAM[34871] = 8'b0;
    XRAM[34872] = 8'b0;
    XRAM[34873] = 8'b0;
    XRAM[34874] = 8'b0;
    XRAM[34875] = 8'b0;
    XRAM[34876] = 8'b0;
    XRAM[34877] = 8'b0;
    XRAM[34878] = 8'b0;
    XRAM[34879] = 8'b0;
    XRAM[34880] = 8'b0;
    XRAM[34881] = 8'b0;
    XRAM[34882] = 8'b0;
    XRAM[34883] = 8'b0;
    XRAM[34884] = 8'b0;
    XRAM[34885] = 8'b0;
    XRAM[34886] = 8'b0;
    XRAM[34887] = 8'b0;
    XRAM[34888] = 8'b0;
    XRAM[34889] = 8'b0;
    XRAM[34890] = 8'b0;
    XRAM[34891] = 8'b0;
    XRAM[34892] = 8'b0;
    XRAM[34893] = 8'b0;
    XRAM[34894] = 8'b0;
    XRAM[34895] = 8'b0;
    XRAM[34896] = 8'b0;
    XRAM[34897] = 8'b0;
    XRAM[34898] = 8'b0;
    XRAM[34899] = 8'b0;
    XRAM[34900] = 8'b0;
    XRAM[34901] = 8'b0;
    XRAM[34902] = 8'b0;
    XRAM[34903] = 8'b0;
    XRAM[34904] = 8'b0;
    XRAM[34905] = 8'b0;
    XRAM[34906] = 8'b0;
    XRAM[34907] = 8'b0;
    XRAM[34908] = 8'b0;
    XRAM[34909] = 8'b0;
    XRAM[34910] = 8'b0;
    XRAM[34911] = 8'b0;
    XRAM[34912] = 8'b0;
    XRAM[34913] = 8'b0;
    XRAM[34914] = 8'b0;
    XRAM[34915] = 8'b0;
    XRAM[34916] = 8'b0;
    XRAM[34917] = 8'b0;
    XRAM[34918] = 8'b0;
    XRAM[34919] = 8'b0;
    XRAM[34920] = 8'b0;
    XRAM[34921] = 8'b0;
    XRAM[34922] = 8'b0;
    XRAM[34923] = 8'b0;
    XRAM[34924] = 8'b0;
    XRAM[34925] = 8'b0;
    XRAM[34926] = 8'b0;
    XRAM[34927] = 8'b0;
    XRAM[34928] = 8'b0;
    XRAM[34929] = 8'b0;
    XRAM[34930] = 8'b0;
    XRAM[34931] = 8'b0;
    XRAM[34932] = 8'b0;
    XRAM[34933] = 8'b0;
    XRAM[34934] = 8'b0;
    XRAM[34935] = 8'b0;
    XRAM[34936] = 8'b0;
    XRAM[34937] = 8'b0;
    XRAM[34938] = 8'b0;
    XRAM[34939] = 8'b0;
    XRAM[34940] = 8'b0;
    XRAM[34941] = 8'b0;
    XRAM[34942] = 8'b0;
    XRAM[34943] = 8'b0;
    XRAM[34944] = 8'b0;
    XRAM[34945] = 8'b0;
    XRAM[34946] = 8'b0;
    XRAM[34947] = 8'b0;
    XRAM[34948] = 8'b0;
    XRAM[34949] = 8'b0;
    XRAM[34950] = 8'b0;
    XRAM[34951] = 8'b0;
    XRAM[34952] = 8'b0;
    XRAM[34953] = 8'b0;
    XRAM[34954] = 8'b0;
    XRAM[34955] = 8'b0;
    XRAM[34956] = 8'b0;
    XRAM[34957] = 8'b0;
    XRAM[34958] = 8'b0;
    XRAM[34959] = 8'b0;
    XRAM[34960] = 8'b0;
    XRAM[34961] = 8'b0;
    XRAM[34962] = 8'b0;
    XRAM[34963] = 8'b0;
    XRAM[34964] = 8'b0;
    XRAM[34965] = 8'b0;
    XRAM[34966] = 8'b0;
    XRAM[34967] = 8'b0;
    XRAM[34968] = 8'b0;
    XRAM[34969] = 8'b0;
    XRAM[34970] = 8'b0;
    XRAM[34971] = 8'b0;
    XRAM[34972] = 8'b0;
    XRAM[34973] = 8'b0;
    XRAM[34974] = 8'b0;
    XRAM[34975] = 8'b0;
    XRAM[34976] = 8'b0;
    XRAM[34977] = 8'b0;
    XRAM[34978] = 8'b0;
    XRAM[34979] = 8'b0;
    XRAM[34980] = 8'b0;
    XRAM[34981] = 8'b0;
    XRAM[34982] = 8'b0;
    XRAM[34983] = 8'b0;
    XRAM[34984] = 8'b0;
    XRAM[34985] = 8'b0;
    XRAM[34986] = 8'b0;
    XRAM[34987] = 8'b0;
    XRAM[34988] = 8'b0;
    XRAM[34989] = 8'b0;
    XRAM[34990] = 8'b0;
    XRAM[34991] = 8'b0;
    XRAM[34992] = 8'b0;
    XRAM[34993] = 8'b0;
    XRAM[34994] = 8'b0;
    XRAM[34995] = 8'b0;
    XRAM[34996] = 8'b0;
    XRAM[34997] = 8'b0;
    XRAM[34998] = 8'b0;
    XRAM[34999] = 8'b0;
    XRAM[35000] = 8'b0;
    XRAM[35001] = 8'b0;
    XRAM[35002] = 8'b0;
    XRAM[35003] = 8'b0;
    XRAM[35004] = 8'b0;
    XRAM[35005] = 8'b0;
    XRAM[35006] = 8'b0;
    XRAM[35007] = 8'b0;
    XRAM[35008] = 8'b0;
    XRAM[35009] = 8'b0;
    XRAM[35010] = 8'b0;
    XRAM[35011] = 8'b0;
    XRAM[35012] = 8'b0;
    XRAM[35013] = 8'b0;
    XRAM[35014] = 8'b0;
    XRAM[35015] = 8'b0;
    XRAM[35016] = 8'b0;
    XRAM[35017] = 8'b0;
    XRAM[35018] = 8'b0;
    XRAM[35019] = 8'b0;
    XRAM[35020] = 8'b0;
    XRAM[35021] = 8'b0;
    XRAM[35022] = 8'b0;
    XRAM[35023] = 8'b0;
    XRAM[35024] = 8'b0;
    XRAM[35025] = 8'b0;
    XRAM[35026] = 8'b0;
    XRAM[35027] = 8'b0;
    XRAM[35028] = 8'b0;
    XRAM[35029] = 8'b0;
    XRAM[35030] = 8'b0;
    XRAM[35031] = 8'b0;
    XRAM[35032] = 8'b0;
    XRAM[35033] = 8'b0;
    XRAM[35034] = 8'b0;
    XRAM[35035] = 8'b0;
    XRAM[35036] = 8'b0;
    XRAM[35037] = 8'b0;
    XRAM[35038] = 8'b0;
    XRAM[35039] = 8'b0;
    XRAM[35040] = 8'b0;
    XRAM[35041] = 8'b0;
    XRAM[35042] = 8'b0;
    XRAM[35043] = 8'b0;
    XRAM[35044] = 8'b0;
    XRAM[35045] = 8'b0;
    XRAM[35046] = 8'b0;
    XRAM[35047] = 8'b0;
    XRAM[35048] = 8'b0;
    XRAM[35049] = 8'b0;
    XRAM[35050] = 8'b0;
    XRAM[35051] = 8'b0;
    XRAM[35052] = 8'b0;
    XRAM[35053] = 8'b0;
    XRAM[35054] = 8'b0;
    XRAM[35055] = 8'b0;
    XRAM[35056] = 8'b0;
    XRAM[35057] = 8'b0;
    XRAM[35058] = 8'b0;
    XRAM[35059] = 8'b0;
    XRAM[35060] = 8'b0;
    XRAM[35061] = 8'b0;
    XRAM[35062] = 8'b0;
    XRAM[35063] = 8'b0;
    XRAM[35064] = 8'b0;
    XRAM[35065] = 8'b0;
    XRAM[35066] = 8'b0;
    XRAM[35067] = 8'b0;
    XRAM[35068] = 8'b0;
    XRAM[35069] = 8'b0;
    XRAM[35070] = 8'b0;
    XRAM[35071] = 8'b0;
    XRAM[35072] = 8'b0;
    XRAM[35073] = 8'b0;
    XRAM[35074] = 8'b0;
    XRAM[35075] = 8'b0;
    XRAM[35076] = 8'b0;
    XRAM[35077] = 8'b0;
    XRAM[35078] = 8'b0;
    XRAM[35079] = 8'b0;
    XRAM[35080] = 8'b0;
    XRAM[35081] = 8'b0;
    XRAM[35082] = 8'b0;
    XRAM[35083] = 8'b0;
    XRAM[35084] = 8'b0;
    XRAM[35085] = 8'b0;
    XRAM[35086] = 8'b0;
    XRAM[35087] = 8'b0;
    XRAM[35088] = 8'b0;
    XRAM[35089] = 8'b0;
    XRAM[35090] = 8'b0;
    XRAM[35091] = 8'b0;
    XRAM[35092] = 8'b0;
    XRAM[35093] = 8'b0;
    XRAM[35094] = 8'b0;
    XRAM[35095] = 8'b0;
    XRAM[35096] = 8'b0;
    XRAM[35097] = 8'b0;
    XRAM[35098] = 8'b0;
    XRAM[35099] = 8'b0;
    XRAM[35100] = 8'b0;
    XRAM[35101] = 8'b0;
    XRAM[35102] = 8'b0;
    XRAM[35103] = 8'b0;
    XRAM[35104] = 8'b0;
    XRAM[35105] = 8'b0;
    XRAM[35106] = 8'b0;
    XRAM[35107] = 8'b0;
    XRAM[35108] = 8'b0;
    XRAM[35109] = 8'b0;
    XRAM[35110] = 8'b0;
    XRAM[35111] = 8'b0;
    XRAM[35112] = 8'b0;
    XRAM[35113] = 8'b0;
    XRAM[35114] = 8'b0;
    XRAM[35115] = 8'b0;
    XRAM[35116] = 8'b0;
    XRAM[35117] = 8'b0;
    XRAM[35118] = 8'b0;
    XRAM[35119] = 8'b0;
    XRAM[35120] = 8'b0;
    XRAM[35121] = 8'b0;
    XRAM[35122] = 8'b0;
    XRAM[35123] = 8'b0;
    XRAM[35124] = 8'b0;
    XRAM[35125] = 8'b0;
    XRAM[35126] = 8'b0;
    XRAM[35127] = 8'b0;
    XRAM[35128] = 8'b0;
    XRAM[35129] = 8'b0;
    XRAM[35130] = 8'b0;
    XRAM[35131] = 8'b0;
    XRAM[35132] = 8'b0;
    XRAM[35133] = 8'b0;
    XRAM[35134] = 8'b0;
    XRAM[35135] = 8'b0;
    XRAM[35136] = 8'b0;
    XRAM[35137] = 8'b0;
    XRAM[35138] = 8'b0;
    XRAM[35139] = 8'b0;
    XRAM[35140] = 8'b0;
    XRAM[35141] = 8'b0;
    XRAM[35142] = 8'b0;
    XRAM[35143] = 8'b0;
    XRAM[35144] = 8'b0;
    XRAM[35145] = 8'b0;
    XRAM[35146] = 8'b0;
    XRAM[35147] = 8'b0;
    XRAM[35148] = 8'b0;
    XRAM[35149] = 8'b0;
    XRAM[35150] = 8'b0;
    XRAM[35151] = 8'b0;
    XRAM[35152] = 8'b0;
    XRAM[35153] = 8'b0;
    XRAM[35154] = 8'b0;
    XRAM[35155] = 8'b0;
    XRAM[35156] = 8'b0;
    XRAM[35157] = 8'b0;
    XRAM[35158] = 8'b0;
    XRAM[35159] = 8'b0;
    XRAM[35160] = 8'b0;
    XRAM[35161] = 8'b0;
    XRAM[35162] = 8'b0;
    XRAM[35163] = 8'b0;
    XRAM[35164] = 8'b0;
    XRAM[35165] = 8'b0;
    XRAM[35166] = 8'b0;
    XRAM[35167] = 8'b0;
    XRAM[35168] = 8'b0;
    XRAM[35169] = 8'b0;
    XRAM[35170] = 8'b0;
    XRAM[35171] = 8'b0;
    XRAM[35172] = 8'b0;
    XRAM[35173] = 8'b0;
    XRAM[35174] = 8'b0;
    XRAM[35175] = 8'b0;
    XRAM[35176] = 8'b0;
    XRAM[35177] = 8'b0;
    XRAM[35178] = 8'b0;
    XRAM[35179] = 8'b0;
    XRAM[35180] = 8'b0;
    XRAM[35181] = 8'b0;
    XRAM[35182] = 8'b0;
    XRAM[35183] = 8'b0;
    XRAM[35184] = 8'b0;
    XRAM[35185] = 8'b0;
    XRAM[35186] = 8'b0;
    XRAM[35187] = 8'b0;
    XRAM[35188] = 8'b0;
    XRAM[35189] = 8'b0;
    XRAM[35190] = 8'b0;
    XRAM[35191] = 8'b0;
    XRAM[35192] = 8'b0;
    XRAM[35193] = 8'b0;
    XRAM[35194] = 8'b0;
    XRAM[35195] = 8'b0;
    XRAM[35196] = 8'b0;
    XRAM[35197] = 8'b0;
    XRAM[35198] = 8'b0;
    XRAM[35199] = 8'b0;
    XRAM[35200] = 8'b0;
    XRAM[35201] = 8'b0;
    XRAM[35202] = 8'b0;
    XRAM[35203] = 8'b0;
    XRAM[35204] = 8'b0;
    XRAM[35205] = 8'b0;
    XRAM[35206] = 8'b0;
    XRAM[35207] = 8'b0;
    XRAM[35208] = 8'b0;
    XRAM[35209] = 8'b0;
    XRAM[35210] = 8'b0;
    XRAM[35211] = 8'b0;
    XRAM[35212] = 8'b0;
    XRAM[35213] = 8'b0;
    XRAM[35214] = 8'b0;
    XRAM[35215] = 8'b0;
    XRAM[35216] = 8'b0;
    XRAM[35217] = 8'b0;
    XRAM[35218] = 8'b0;
    XRAM[35219] = 8'b0;
    XRAM[35220] = 8'b0;
    XRAM[35221] = 8'b0;
    XRAM[35222] = 8'b0;
    XRAM[35223] = 8'b0;
    XRAM[35224] = 8'b0;
    XRAM[35225] = 8'b0;
    XRAM[35226] = 8'b0;
    XRAM[35227] = 8'b0;
    XRAM[35228] = 8'b0;
    XRAM[35229] = 8'b0;
    XRAM[35230] = 8'b0;
    XRAM[35231] = 8'b0;
    XRAM[35232] = 8'b0;
    XRAM[35233] = 8'b0;
    XRAM[35234] = 8'b0;
    XRAM[35235] = 8'b0;
    XRAM[35236] = 8'b0;
    XRAM[35237] = 8'b0;
    XRAM[35238] = 8'b0;
    XRAM[35239] = 8'b0;
    XRAM[35240] = 8'b0;
    XRAM[35241] = 8'b0;
    XRAM[35242] = 8'b0;
    XRAM[35243] = 8'b0;
    XRAM[35244] = 8'b0;
    XRAM[35245] = 8'b0;
    XRAM[35246] = 8'b0;
    XRAM[35247] = 8'b0;
    XRAM[35248] = 8'b0;
    XRAM[35249] = 8'b0;
    XRAM[35250] = 8'b0;
    XRAM[35251] = 8'b0;
    XRAM[35252] = 8'b0;
    XRAM[35253] = 8'b0;
    XRAM[35254] = 8'b0;
    XRAM[35255] = 8'b0;
    XRAM[35256] = 8'b0;
    XRAM[35257] = 8'b0;
    XRAM[35258] = 8'b0;
    XRAM[35259] = 8'b0;
    XRAM[35260] = 8'b0;
    XRAM[35261] = 8'b0;
    XRAM[35262] = 8'b0;
    XRAM[35263] = 8'b0;
    XRAM[35264] = 8'b0;
    XRAM[35265] = 8'b0;
    XRAM[35266] = 8'b0;
    XRAM[35267] = 8'b0;
    XRAM[35268] = 8'b0;
    XRAM[35269] = 8'b0;
    XRAM[35270] = 8'b0;
    XRAM[35271] = 8'b0;
    XRAM[35272] = 8'b0;
    XRAM[35273] = 8'b0;
    XRAM[35274] = 8'b0;
    XRAM[35275] = 8'b0;
    XRAM[35276] = 8'b0;
    XRAM[35277] = 8'b0;
    XRAM[35278] = 8'b0;
    XRAM[35279] = 8'b0;
    XRAM[35280] = 8'b0;
    XRAM[35281] = 8'b0;
    XRAM[35282] = 8'b0;
    XRAM[35283] = 8'b0;
    XRAM[35284] = 8'b0;
    XRAM[35285] = 8'b0;
    XRAM[35286] = 8'b0;
    XRAM[35287] = 8'b0;
    XRAM[35288] = 8'b0;
    XRAM[35289] = 8'b0;
    XRAM[35290] = 8'b0;
    XRAM[35291] = 8'b0;
    XRAM[35292] = 8'b0;
    XRAM[35293] = 8'b0;
    XRAM[35294] = 8'b0;
    XRAM[35295] = 8'b0;
    XRAM[35296] = 8'b0;
    XRAM[35297] = 8'b0;
    XRAM[35298] = 8'b0;
    XRAM[35299] = 8'b0;
    XRAM[35300] = 8'b0;
    XRAM[35301] = 8'b0;
    XRAM[35302] = 8'b0;
    XRAM[35303] = 8'b0;
    XRAM[35304] = 8'b0;
    XRAM[35305] = 8'b0;
    XRAM[35306] = 8'b0;
    XRAM[35307] = 8'b0;
    XRAM[35308] = 8'b0;
    XRAM[35309] = 8'b0;
    XRAM[35310] = 8'b0;
    XRAM[35311] = 8'b0;
    XRAM[35312] = 8'b0;
    XRAM[35313] = 8'b0;
    XRAM[35314] = 8'b0;
    XRAM[35315] = 8'b0;
    XRAM[35316] = 8'b0;
    XRAM[35317] = 8'b0;
    XRAM[35318] = 8'b0;
    XRAM[35319] = 8'b0;
    XRAM[35320] = 8'b0;
    XRAM[35321] = 8'b0;
    XRAM[35322] = 8'b0;
    XRAM[35323] = 8'b0;
    XRAM[35324] = 8'b0;
    XRAM[35325] = 8'b0;
    XRAM[35326] = 8'b0;
    XRAM[35327] = 8'b0;
    XRAM[35328] = 8'b0;
    XRAM[35329] = 8'b0;
    XRAM[35330] = 8'b0;
    XRAM[35331] = 8'b0;
    XRAM[35332] = 8'b0;
    XRAM[35333] = 8'b0;
    XRAM[35334] = 8'b0;
    XRAM[35335] = 8'b0;
    XRAM[35336] = 8'b0;
    XRAM[35337] = 8'b0;
    XRAM[35338] = 8'b0;
    XRAM[35339] = 8'b0;
    XRAM[35340] = 8'b0;
    XRAM[35341] = 8'b0;
    XRAM[35342] = 8'b0;
    XRAM[35343] = 8'b0;
    XRAM[35344] = 8'b0;
    XRAM[35345] = 8'b0;
    XRAM[35346] = 8'b0;
    XRAM[35347] = 8'b0;
    XRAM[35348] = 8'b0;
    XRAM[35349] = 8'b0;
    XRAM[35350] = 8'b0;
    XRAM[35351] = 8'b0;
    XRAM[35352] = 8'b0;
    XRAM[35353] = 8'b0;
    XRAM[35354] = 8'b0;
    XRAM[35355] = 8'b0;
    XRAM[35356] = 8'b0;
    XRAM[35357] = 8'b0;
    XRAM[35358] = 8'b0;
    XRAM[35359] = 8'b0;
    XRAM[35360] = 8'b0;
    XRAM[35361] = 8'b0;
    XRAM[35362] = 8'b0;
    XRAM[35363] = 8'b0;
    XRAM[35364] = 8'b0;
    XRAM[35365] = 8'b0;
    XRAM[35366] = 8'b0;
    XRAM[35367] = 8'b0;
    XRAM[35368] = 8'b0;
    XRAM[35369] = 8'b0;
    XRAM[35370] = 8'b0;
    XRAM[35371] = 8'b0;
    XRAM[35372] = 8'b0;
    XRAM[35373] = 8'b0;
    XRAM[35374] = 8'b0;
    XRAM[35375] = 8'b0;
    XRAM[35376] = 8'b0;
    XRAM[35377] = 8'b0;
    XRAM[35378] = 8'b0;
    XRAM[35379] = 8'b0;
    XRAM[35380] = 8'b0;
    XRAM[35381] = 8'b0;
    XRAM[35382] = 8'b0;
    XRAM[35383] = 8'b0;
    XRAM[35384] = 8'b0;
    XRAM[35385] = 8'b0;
    XRAM[35386] = 8'b0;
    XRAM[35387] = 8'b0;
    XRAM[35388] = 8'b0;
    XRAM[35389] = 8'b0;
    XRAM[35390] = 8'b0;
    XRAM[35391] = 8'b0;
    XRAM[35392] = 8'b0;
    XRAM[35393] = 8'b0;
    XRAM[35394] = 8'b0;
    XRAM[35395] = 8'b0;
    XRAM[35396] = 8'b0;
    XRAM[35397] = 8'b0;
    XRAM[35398] = 8'b0;
    XRAM[35399] = 8'b0;
    XRAM[35400] = 8'b0;
    XRAM[35401] = 8'b0;
    XRAM[35402] = 8'b0;
    XRAM[35403] = 8'b0;
    XRAM[35404] = 8'b0;
    XRAM[35405] = 8'b0;
    XRAM[35406] = 8'b0;
    XRAM[35407] = 8'b0;
    XRAM[35408] = 8'b0;
    XRAM[35409] = 8'b0;
    XRAM[35410] = 8'b0;
    XRAM[35411] = 8'b0;
    XRAM[35412] = 8'b0;
    XRAM[35413] = 8'b0;
    XRAM[35414] = 8'b0;
    XRAM[35415] = 8'b0;
    XRAM[35416] = 8'b0;
    XRAM[35417] = 8'b0;
    XRAM[35418] = 8'b0;
    XRAM[35419] = 8'b0;
    XRAM[35420] = 8'b0;
    XRAM[35421] = 8'b0;
    XRAM[35422] = 8'b0;
    XRAM[35423] = 8'b0;
    XRAM[35424] = 8'b0;
    XRAM[35425] = 8'b0;
    XRAM[35426] = 8'b0;
    XRAM[35427] = 8'b0;
    XRAM[35428] = 8'b0;
    XRAM[35429] = 8'b0;
    XRAM[35430] = 8'b0;
    XRAM[35431] = 8'b0;
    XRAM[35432] = 8'b0;
    XRAM[35433] = 8'b0;
    XRAM[35434] = 8'b0;
    XRAM[35435] = 8'b0;
    XRAM[35436] = 8'b0;
    XRAM[35437] = 8'b0;
    XRAM[35438] = 8'b0;
    XRAM[35439] = 8'b0;
    XRAM[35440] = 8'b0;
    XRAM[35441] = 8'b0;
    XRAM[35442] = 8'b0;
    XRAM[35443] = 8'b0;
    XRAM[35444] = 8'b0;
    XRAM[35445] = 8'b0;
    XRAM[35446] = 8'b0;
    XRAM[35447] = 8'b0;
    XRAM[35448] = 8'b0;
    XRAM[35449] = 8'b0;
    XRAM[35450] = 8'b0;
    XRAM[35451] = 8'b0;
    XRAM[35452] = 8'b0;
    XRAM[35453] = 8'b0;
    XRAM[35454] = 8'b0;
    XRAM[35455] = 8'b0;
    XRAM[35456] = 8'b0;
    XRAM[35457] = 8'b0;
    XRAM[35458] = 8'b0;
    XRAM[35459] = 8'b0;
    XRAM[35460] = 8'b0;
    XRAM[35461] = 8'b0;
    XRAM[35462] = 8'b0;
    XRAM[35463] = 8'b0;
    XRAM[35464] = 8'b0;
    XRAM[35465] = 8'b0;
    XRAM[35466] = 8'b0;
    XRAM[35467] = 8'b0;
    XRAM[35468] = 8'b0;
    XRAM[35469] = 8'b0;
    XRAM[35470] = 8'b0;
    XRAM[35471] = 8'b0;
    XRAM[35472] = 8'b0;
    XRAM[35473] = 8'b0;
    XRAM[35474] = 8'b0;
    XRAM[35475] = 8'b0;
    XRAM[35476] = 8'b0;
    XRAM[35477] = 8'b0;
    XRAM[35478] = 8'b0;
    XRAM[35479] = 8'b0;
    XRAM[35480] = 8'b0;
    XRAM[35481] = 8'b0;
    XRAM[35482] = 8'b0;
    XRAM[35483] = 8'b0;
    XRAM[35484] = 8'b0;
    XRAM[35485] = 8'b0;
    XRAM[35486] = 8'b0;
    XRAM[35487] = 8'b0;
    XRAM[35488] = 8'b0;
    XRAM[35489] = 8'b0;
    XRAM[35490] = 8'b0;
    XRAM[35491] = 8'b0;
    XRAM[35492] = 8'b0;
    XRAM[35493] = 8'b0;
    XRAM[35494] = 8'b0;
    XRAM[35495] = 8'b0;
    XRAM[35496] = 8'b0;
    XRAM[35497] = 8'b0;
    XRAM[35498] = 8'b0;
    XRAM[35499] = 8'b0;
    XRAM[35500] = 8'b0;
    XRAM[35501] = 8'b0;
    XRAM[35502] = 8'b0;
    XRAM[35503] = 8'b0;
    XRAM[35504] = 8'b0;
    XRAM[35505] = 8'b0;
    XRAM[35506] = 8'b0;
    XRAM[35507] = 8'b0;
    XRAM[35508] = 8'b0;
    XRAM[35509] = 8'b0;
    XRAM[35510] = 8'b0;
    XRAM[35511] = 8'b0;
    XRAM[35512] = 8'b0;
    XRAM[35513] = 8'b0;
    XRAM[35514] = 8'b0;
    XRAM[35515] = 8'b0;
    XRAM[35516] = 8'b0;
    XRAM[35517] = 8'b0;
    XRAM[35518] = 8'b0;
    XRAM[35519] = 8'b0;
    XRAM[35520] = 8'b0;
    XRAM[35521] = 8'b0;
    XRAM[35522] = 8'b0;
    XRAM[35523] = 8'b0;
    XRAM[35524] = 8'b0;
    XRAM[35525] = 8'b0;
    XRAM[35526] = 8'b0;
    XRAM[35527] = 8'b0;
    XRAM[35528] = 8'b0;
    XRAM[35529] = 8'b0;
    XRAM[35530] = 8'b0;
    XRAM[35531] = 8'b0;
    XRAM[35532] = 8'b0;
    XRAM[35533] = 8'b0;
    XRAM[35534] = 8'b0;
    XRAM[35535] = 8'b0;
    XRAM[35536] = 8'b0;
    XRAM[35537] = 8'b0;
    XRAM[35538] = 8'b0;
    XRAM[35539] = 8'b0;
    XRAM[35540] = 8'b0;
    XRAM[35541] = 8'b0;
    XRAM[35542] = 8'b0;
    XRAM[35543] = 8'b0;
    XRAM[35544] = 8'b0;
    XRAM[35545] = 8'b0;
    XRAM[35546] = 8'b0;
    XRAM[35547] = 8'b0;
    XRAM[35548] = 8'b0;
    XRAM[35549] = 8'b0;
    XRAM[35550] = 8'b0;
    XRAM[35551] = 8'b0;
    XRAM[35552] = 8'b0;
    XRAM[35553] = 8'b0;
    XRAM[35554] = 8'b0;
    XRAM[35555] = 8'b0;
    XRAM[35556] = 8'b0;
    XRAM[35557] = 8'b0;
    XRAM[35558] = 8'b0;
    XRAM[35559] = 8'b0;
    XRAM[35560] = 8'b0;
    XRAM[35561] = 8'b0;
    XRAM[35562] = 8'b0;
    XRAM[35563] = 8'b0;
    XRAM[35564] = 8'b0;
    XRAM[35565] = 8'b0;
    XRAM[35566] = 8'b0;
    XRAM[35567] = 8'b0;
    XRAM[35568] = 8'b0;
    XRAM[35569] = 8'b0;
    XRAM[35570] = 8'b0;
    XRAM[35571] = 8'b0;
    XRAM[35572] = 8'b0;
    XRAM[35573] = 8'b0;
    XRAM[35574] = 8'b0;
    XRAM[35575] = 8'b0;
    XRAM[35576] = 8'b0;
    XRAM[35577] = 8'b0;
    XRAM[35578] = 8'b0;
    XRAM[35579] = 8'b0;
    XRAM[35580] = 8'b0;
    XRAM[35581] = 8'b0;
    XRAM[35582] = 8'b0;
    XRAM[35583] = 8'b0;
    XRAM[35584] = 8'b0;
    XRAM[35585] = 8'b0;
    XRAM[35586] = 8'b0;
    XRAM[35587] = 8'b0;
    XRAM[35588] = 8'b0;
    XRAM[35589] = 8'b0;
    XRAM[35590] = 8'b0;
    XRAM[35591] = 8'b0;
    XRAM[35592] = 8'b0;
    XRAM[35593] = 8'b0;
    XRAM[35594] = 8'b0;
    XRAM[35595] = 8'b0;
    XRAM[35596] = 8'b0;
    XRAM[35597] = 8'b0;
    XRAM[35598] = 8'b0;
    XRAM[35599] = 8'b0;
    XRAM[35600] = 8'b0;
    XRAM[35601] = 8'b0;
    XRAM[35602] = 8'b0;
    XRAM[35603] = 8'b0;
    XRAM[35604] = 8'b0;
    XRAM[35605] = 8'b0;
    XRAM[35606] = 8'b0;
    XRAM[35607] = 8'b0;
    XRAM[35608] = 8'b0;
    XRAM[35609] = 8'b0;
    XRAM[35610] = 8'b0;
    XRAM[35611] = 8'b0;
    XRAM[35612] = 8'b0;
    XRAM[35613] = 8'b0;
    XRAM[35614] = 8'b0;
    XRAM[35615] = 8'b0;
    XRAM[35616] = 8'b0;
    XRAM[35617] = 8'b0;
    XRAM[35618] = 8'b0;
    XRAM[35619] = 8'b0;
    XRAM[35620] = 8'b0;
    XRAM[35621] = 8'b0;
    XRAM[35622] = 8'b0;
    XRAM[35623] = 8'b0;
    XRAM[35624] = 8'b0;
    XRAM[35625] = 8'b0;
    XRAM[35626] = 8'b0;
    XRAM[35627] = 8'b0;
    XRAM[35628] = 8'b0;
    XRAM[35629] = 8'b0;
    XRAM[35630] = 8'b0;
    XRAM[35631] = 8'b0;
    XRAM[35632] = 8'b0;
    XRAM[35633] = 8'b0;
    XRAM[35634] = 8'b0;
    XRAM[35635] = 8'b0;
    XRAM[35636] = 8'b0;
    XRAM[35637] = 8'b0;
    XRAM[35638] = 8'b0;
    XRAM[35639] = 8'b0;
    XRAM[35640] = 8'b0;
    XRAM[35641] = 8'b0;
    XRAM[35642] = 8'b0;
    XRAM[35643] = 8'b0;
    XRAM[35644] = 8'b0;
    XRAM[35645] = 8'b0;
    XRAM[35646] = 8'b0;
    XRAM[35647] = 8'b0;
    XRAM[35648] = 8'b0;
    XRAM[35649] = 8'b0;
    XRAM[35650] = 8'b0;
    XRAM[35651] = 8'b0;
    XRAM[35652] = 8'b0;
    XRAM[35653] = 8'b0;
    XRAM[35654] = 8'b0;
    XRAM[35655] = 8'b0;
    XRAM[35656] = 8'b0;
    XRAM[35657] = 8'b0;
    XRAM[35658] = 8'b0;
    XRAM[35659] = 8'b0;
    XRAM[35660] = 8'b0;
    XRAM[35661] = 8'b0;
    XRAM[35662] = 8'b0;
    XRAM[35663] = 8'b0;
    XRAM[35664] = 8'b0;
    XRAM[35665] = 8'b0;
    XRAM[35666] = 8'b0;
    XRAM[35667] = 8'b0;
    XRAM[35668] = 8'b0;
    XRAM[35669] = 8'b0;
    XRAM[35670] = 8'b0;
    XRAM[35671] = 8'b0;
    XRAM[35672] = 8'b0;
    XRAM[35673] = 8'b0;
    XRAM[35674] = 8'b0;
    XRAM[35675] = 8'b0;
    XRAM[35676] = 8'b0;
    XRAM[35677] = 8'b0;
    XRAM[35678] = 8'b0;
    XRAM[35679] = 8'b0;
    XRAM[35680] = 8'b0;
    XRAM[35681] = 8'b0;
    XRAM[35682] = 8'b0;
    XRAM[35683] = 8'b0;
    XRAM[35684] = 8'b0;
    XRAM[35685] = 8'b0;
    XRAM[35686] = 8'b0;
    XRAM[35687] = 8'b0;
    XRAM[35688] = 8'b0;
    XRAM[35689] = 8'b0;
    XRAM[35690] = 8'b0;
    XRAM[35691] = 8'b0;
    XRAM[35692] = 8'b0;
    XRAM[35693] = 8'b0;
    XRAM[35694] = 8'b0;
    XRAM[35695] = 8'b0;
    XRAM[35696] = 8'b0;
    XRAM[35697] = 8'b0;
    XRAM[35698] = 8'b0;
    XRAM[35699] = 8'b0;
    XRAM[35700] = 8'b0;
    XRAM[35701] = 8'b0;
    XRAM[35702] = 8'b0;
    XRAM[35703] = 8'b0;
    XRAM[35704] = 8'b0;
    XRAM[35705] = 8'b0;
    XRAM[35706] = 8'b0;
    XRAM[35707] = 8'b0;
    XRAM[35708] = 8'b0;
    XRAM[35709] = 8'b0;
    XRAM[35710] = 8'b0;
    XRAM[35711] = 8'b0;
    XRAM[35712] = 8'b0;
    XRAM[35713] = 8'b0;
    XRAM[35714] = 8'b0;
    XRAM[35715] = 8'b0;
    XRAM[35716] = 8'b0;
    XRAM[35717] = 8'b0;
    XRAM[35718] = 8'b0;
    XRAM[35719] = 8'b0;
    XRAM[35720] = 8'b0;
    XRAM[35721] = 8'b0;
    XRAM[35722] = 8'b0;
    XRAM[35723] = 8'b0;
    XRAM[35724] = 8'b0;
    XRAM[35725] = 8'b0;
    XRAM[35726] = 8'b0;
    XRAM[35727] = 8'b0;
    XRAM[35728] = 8'b0;
    XRAM[35729] = 8'b0;
    XRAM[35730] = 8'b0;
    XRAM[35731] = 8'b0;
    XRAM[35732] = 8'b0;
    XRAM[35733] = 8'b0;
    XRAM[35734] = 8'b0;
    XRAM[35735] = 8'b0;
    XRAM[35736] = 8'b0;
    XRAM[35737] = 8'b0;
    XRAM[35738] = 8'b0;
    XRAM[35739] = 8'b0;
    XRAM[35740] = 8'b0;
    XRAM[35741] = 8'b0;
    XRAM[35742] = 8'b0;
    XRAM[35743] = 8'b0;
    XRAM[35744] = 8'b0;
    XRAM[35745] = 8'b0;
    XRAM[35746] = 8'b0;
    XRAM[35747] = 8'b0;
    XRAM[35748] = 8'b0;
    XRAM[35749] = 8'b0;
    XRAM[35750] = 8'b0;
    XRAM[35751] = 8'b0;
    XRAM[35752] = 8'b0;
    XRAM[35753] = 8'b0;
    XRAM[35754] = 8'b0;
    XRAM[35755] = 8'b0;
    XRAM[35756] = 8'b0;
    XRAM[35757] = 8'b0;
    XRAM[35758] = 8'b0;
    XRAM[35759] = 8'b0;
    XRAM[35760] = 8'b0;
    XRAM[35761] = 8'b0;
    XRAM[35762] = 8'b0;
    XRAM[35763] = 8'b0;
    XRAM[35764] = 8'b0;
    XRAM[35765] = 8'b0;
    XRAM[35766] = 8'b0;
    XRAM[35767] = 8'b0;
    XRAM[35768] = 8'b0;
    XRAM[35769] = 8'b0;
    XRAM[35770] = 8'b0;
    XRAM[35771] = 8'b0;
    XRAM[35772] = 8'b0;
    XRAM[35773] = 8'b0;
    XRAM[35774] = 8'b0;
    XRAM[35775] = 8'b0;
    XRAM[35776] = 8'b0;
    XRAM[35777] = 8'b0;
    XRAM[35778] = 8'b0;
    XRAM[35779] = 8'b0;
    XRAM[35780] = 8'b0;
    XRAM[35781] = 8'b0;
    XRAM[35782] = 8'b0;
    XRAM[35783] = 8'b0;
    XRAM[35784] = 8'b0;
    XRAM[35785] = 8'b0;
    XRAM[35786] = 8'b0;
    XRAM[35787] = 8'b0;
    XRAM[35788] = 8'b0;
    XRAM[35789] = 8'b0;
    XRAM[35790] = 8'b0;
    XRAM[35791] = 8'b0;
    XRAM[35792] = 8'b0;
    XRAM[35793] = 8'b0;
    XRAM[35794] = 8'b0;
    XRAM[35795] = 8'b0;
    XRAM[35796] = 8'b0;
    XRAM[35797] = 8'b0;
    XRAM[35798] = 8'b0;
    XRAM[35799] = 8'b0;
    XRAM[35800] = 8'b0;
    XRAM[35801] = 8'b0;
    XRAM[35802] = 8'b0;
    XRAM[35803] = 8'b0;
    XRAM[35804] = 8'b0;
    XRAM[35805] = 8'b0;
    XRAM[35806] = 8'b0;
    XRAM[35807] = 8'b0;
    XRAM[35808] = 8'b0;
    XRAM[35809] = 8'b0;
    XRAM[35810] = 8'b0;
    XRAM[35811] = 8'b0;
    XRAM[35812] = 8'b0;
    XRAM[35813] = 8'b0;
    XRAM[35814] = 8'b0;
    XRAM[35815] = 8'b0;
    XRAM[35816] = 8'b0;
    XRAM[35817] = 8'b0;
    XRAM[35818] = 8'b0;
    XRAM[35819] = 8'b0;
    XRAM[35820] = 8'b0;
    XRAM[35821] = 8'b0;
    XRAM[35822] = 8'b0;
    XRAM[35823] = 8'b0;
    XRAM[35824] = 8'b0;
    XRAM[35825] = 8'b0;
    XRAM[35826] = 8'b0;
    XRAM[35827] = 8'b0;
    XRAM[35828] = 8'b0;
    XRAM[35829] = 8'b0;
    XRAM[35830] = 8'b0;
    XRAM[35831] = 8'b0;
    XRAM[35832] = 8'b0;
    XRAM[35833] = 8'b0;
    XRAM[35834] = 8'b0;
    XRAM[35835] = 8'b0;
    XRAM[35836] = 8'b0;
    XRAM[35837] = 8'b0;
    XRAM[35838] = 8'b0;
    XRAM[35839] = 8'b0;
    XRAM[35840] = 8'b0;
    XRAM[35841] = 8'b0;
    XRAM[35842] = 8'b0;
    XRAM[35843] = 8'b0;
    XRAM[35844] = 8'b0;
    XRAM[35845] = 8'b0;
    XRAM[35846] = 8'b0;
    XRAM[35847] = 8'b0;
    XRAM[35848] = 8'b0;
    XRAM[35849] = 8'b0;
    XRAM[35850] = 8'b0;
    XRAM[35851] = 8'b0;
    XRAM[35852] = 8'b0;
    XRAM[35853] = 8'b0;
    XRAM[35854] = 8'b0;
    XRAM[35855] = 8'b0;
    XRAM[35856] = 8'b0;
    XRAM[35857] = 8'b0;
    XRAM[35858] = 8'b0;
    XRAM[35859] = 8'b0;
    XRAM[35860] = 8'b0;
    XRAM[35861] = 8'b0;
    XRAM[35862] = 8'b0;
    XRAM[35863] = 8'b0;
    XRAM[35864] = 8'b0;
    XRAM[35865] = 8'b0;
    XRAM[35866] = 8'b0;
    XRAM[35867] = 8'b0;
    XRAM[35868] = 8'b0;
    XRAM[35869] = 8'b0;
    XRAM[35870] = 8'b0;
    XRAM[35871] = 8'b0;
    XRAM[35872] = 8'b0;
    XRAM[35873] = 8'b0;
    XRAM[35874] = 8'b0;
    XRAM[35875] = 8'b0;
    XRAM[35876] = 8'b0;
    XRAM[35877] = 8'b0;
    XRAM[35878] = 8'b0;
    XRAM[35879] = 8'b0;
    XRAM[35880] = 8'b0;
    XRAM[35881] = 8'b0;
    XRAM[35882] = 8'b0;
    XRAM[35883] = 8'b0;
    XRAM[35884] = 8'b0;
    XRAM[35885] = 8'b0;
    XRAM[35886] = 8'b0;
    XRAM[35887] = 8'b0;
    XRAM[35888] = 8'b0;
    XRAM[35889] = 8'b0;
    XRAM[35890] = 8'b0;
    XRAM[35891] = 8'b0;
    XRAM[35892] = 8'b0;
    XRAM[35893] = 8'b0;
    XRAM[35894] = 8'b0;
    XRAM[35895] = 8'b0;
    XRAM[35896] = 8'b0;
    XRAM[35897] = 8'b0;
    XRAM[35898] = 8'b0;
    XRAM[35899] = 8'b0;
    XRAM[35900] = 8'b0;
    XRAM[35901] = 8'b0;
    XRAM[35902] = 8'b0;
    XRAM[35903] = 8'b0;
    XRAM[35904] = 8'b0;
    XRAM[35905] = 8'b0;
    XRAM[35906] = 8'b0;
    XRAM[35907] = 8'b0;
    XRAM[35908] = 8'b0;
    XRAM[35909] = 8'b0;
    XRAM[35910] = 8'b0;
    XRAM[35911] = 8'b0;
    XRAM[35912] = 8'b0;
    XRAM[35913] = 8'b0;
    XRAM[35914] = 8'b0;
    XRAM[35915] = 8'b0;
    XRAM[35916] = 8'b0;
    XRAM[35917] = 8'b0;
    XRAM[35918] = 8'b0;
    XRAM[35919] = 8'b0;
    XRAM[35920] = 8'b0;
    XRAM[35921] = 8'b0;
    XRAM[35922] = 8'b0;
    XRAM[35923] = 8'b0;
    XRAM[35924] = 8'b0;
    XRAM[35925] = 8'b0;
    XRAM[35926] = 8'b0;
    XRAM[35927] = 8'b0;
    XRAM[35928] = 8'b0;
    XRAM[35929] = 8'b0;
    XRAM[35930] = 8'b0;
    XRAM[35931] = 8'b0;
    XRAM[35932] = 8'b0;
    XRAM[35933] = 8'b0;
    XRAM[35934] = 8'b0;
    XRAM[35935] = 8'b0;
    XRAM[35936] = 8'b0;
    XRAM[35937] = 8'b0;
    XRAM[35938] = 8'b0;
    XRAM[35939] = 8'b0;
    XRAM[35940] = 8'b0;
    XRAM[35941] = 8'b0;
    XRAM[35942] = 8'b0;
    XRAM[35943] = 8'b0;
    XRAM[35944] = 8'b0;
    XRAM[35945] = 8'b0;
    XRAM[35946] = 8'b0;
    XRAM[35947] = 8'b0;
    XRAM[35948] = 8'b0;
    XRAM[35949] = 8'b0;
    XRAM[35950] = 8'b0;
    XRAM[35951] = 8'b0;
    XRAM[35952] = 8'b0;
    XRAM[35953] = 8'b0;
    XRAM[35954] = 8'b0;
    XRAM[35955] = 8'b0;
    XRAM[35956] = 8'b0;
    XRAM[35957] = 8'b0;
    XRAM[35958] = 8'b0;
    XRAM[35959] = 8'b0;
    XRAM[35960] = 8'b0;
    XRAM[35961] = 8'b0;
    XRAM[35962] = 8'b0;
    XRAM[35963] = 8'b0;
    XRAM[35964] = 8'b0;
    XRAM[35965] = 8'b0;
    XRAM[35966] = 8'b0;
    XRAM[35967] = 8'b0;
    XRAM[35968] = 8'b0;
    XRAM[35969] = 8'b0;
    XRAM[35970] = 8'b0;
    XRAM[35971] = 8'b0;
    XRAM[35972] = 8'b0;
    XRAM[35973] = 8'b0;
    XRAM[35974] = 8'b0;
    XRAM[35975] = 8'b0;
    XRAM[35976] = 8'b0;
    XRAM[35977] = 8'b0;
    XRAM[35978] = 8'b0;
    XRAM[35979] = 8'b0;
    XRAM[35980] = 8'b0;
    XRAM[35981] = 8'b0;
    XRAM[35982] = 8'b0;
    XRAM[35983] = 8'b0;
    XRAM[35984] = 8'b0;
    XRAM[35985] = 8'b0;
    XRAM[35986] = 8'b0;
    XRAM[35987] = 8'b0;
    XRAM[35988] = 8'b0;
    XRAM[35989] = 8'b0;
    XRAM[35990] = 8'b0;
    XRAM[35991] = 8'b0;
    XRAM[35992] = 8'b0;
    XRAM[35993] = 8'b0;
    XRAM[35994] = 8'b0;
    XRAM[35995] = 8'b0;
    XRAM[35996] = 8'b0;
    XRAM[35997] = 8'b0;
    XRAM[35998] = 8'b0;
    XRAM[35999] = 8'b0;
    XRAM[36000] = 8'b0;
    XRAM[36001] = 8'b0;
    XRAM[36002] = 8'b0;
    XRAM[36003] = 8'b0;
    XRAM[36004] = 8'b0;
    XRAM[36005] = 8'b0;
    XRAM[36006] = 8'b0;
    XRAM[36007] = 8'b0;
    XRAM[36008] = 8'b0;
    XRAM[36009] = 8'b0;
    XRAM[36010] = 8'b0;
    XRAM[36011] = 8'b0;
    XRAM[36012] = 8'b0;
    XRAM[36013] = 8'b0;
    XRAM[36014] = 8'b0;
    XRAM[36015] = 8'b0;
    XRAM[36016] = 8'b0;
    XRAM[36017] = 8'b0;
    XRAM[36018] = 8'b0;
    XRAM[36019] = 8'b0;
    XRAM[36020] = 8'b0;
    XRAM[36021] = 8'b0;
    XRAM[36022] = 8'b0;
    XRAM[36023] = 8'b0;
    XRAM[36024] = 8'b0;
    XRAM[36025] = 8'b0;
    XRAM[36026] = 8'b0;
    XRAM[36027] = 8'b0;
    XRAM[36028] = 8'b0;
    XRAM[36029] = 8'b0;
    XRAM[36030] = 8'b0;
    XRAM[36031] = 8'b0;
    XRAM[36032] = 8'b0;
    XRAM[36033] = 8'b0;
    XRAM[36034] = 8'b0;
    XRAM[36035] = 8'b0;
    XRAM[36036] = 8'b0;
    XRAM[36037] = 8'b0;
    XRAM[36038] = 8'b0;
    XRAM[36039] = 8'b0;
    XRAM[36040] = 8'b0;
    XRAM[36041] = 8'b0;
    XRAM[36042] = 8'b0;
    XRAM[36043] = 8'b0;
    XRAM[36044] = 8'b0;
    XRAM[36045] = 8'b0;
    XRAM[36046] = 8'b0;
    XRAM[36047] = 8'b0;
    XRAM[36048] = 8'b0;
    XRAM[36049] = 8'b0;
    XRAM[36050] = 8'b0;
    XRAM[36051] = 8'b0;
    XRAM[36052] = 8'b0;
    XRAM[36053] = 8'b0;
    XRAM[36054] = 8'b0;
    XRAM[36055] = 8'b0;
    XRAM[36056] = 8'b0;
    XRAM[36057] = 8'b0;
    XRAM[36058] = 8'b0;
    XRAM[36059] = 8'b0;
    XRAM[36060] = 8'b0;
    XRAM[36061] = 8'b0;
    XRAM[36062] = 8'b0;
    XRAM[36063] = 8'b0;
    XRAM[36064] = 8'b0;
    XRAM[36065] = 8'b0;
    XRAM[36066] = 8'b0;
    XRAM[36067] = 8'b0;
    XRAM[36068] = 8'b0;
    XRAM[36069] = 8'b0;
    XRAM[36070] = 8'b0;
    XRAM[36071] = 8'b0;
    XRAM[36072] = 8'b0;
    XRAM[36073] = 8'b0;
    XRAM[36074] = 8'b0;
    XRAM[36075] = 8'b0;
    XRAM[36076] = 8'b0;
    XRAM[36077] = 8'b0;
    XRAM[36078] = 8'b0;
    XRAM[36079] = 8'b0;
    XRAM[36080] = 8'b0;
    XRAM[36081] = 8'b0;
    XRAM[36082] = 8'b0;
    XRAM[36083] = 8'b0;
    XRAM[36084] = 8'b0;
    XRAM[36085] = 8'b0;
    XRAM[36086] = 8'b0;
    XRAM[36087] = 8'b0;
    XRAM[36088] = 8'b0;
    XRAM[36089] = 8'b0;
    XRAM[36090] = 8'b0;
    XRAM[36091] = 8'b0;
    XRAM[36092] = 8'b0;
    XRAM[36093] = 8'b0;
    XRAM[36094] = 8'b0;
    XRAM[36095] = 8'b0;
    XRAM[36096] = 8'b0;
    XRAM[36097] = 8'b0;
    XRAM[36098] = 8'b0;
    XRAM[36099] = 8'b0;
    XRAM[36100] = 8'b0;
    XRAM[36101] = 8'b0;
    XRAM[36102] = 8'b0;
    XRAM[36103] = 8'b0;
    XRAM[36104] = 8'b0;
    XRAM[36105] = 8'b0;
    XRAM[36106] = 8'b0;
    XRAM[36107] = 8'b0;
    XRAM[36108] = 8'b0;
    XRAM[36109] = 8'b0;
    XRAM[36110] = 8'b0;
    XRAM[36111] = 8'b0;
    XRAM[36112] = 8'b0;
    XRAM[36113] = 8'b0;
    XRAM[36114] = 8'b0;
    XRAM[36115] = 8'b0;
    XRAM[36116] = 8'b0;
    XRAM[36117] = 8'b0;
    XRAM[36118] = 8'b0;
    XRAM[36119] = 8'b0;
    XRAM[36120] = 8'b0;
    XRAM[36121] = 8'b0;
    XRAM[36122] = 8'b0;
    XRAM[36123] = 8'b0;
    XRAM[36124] = 8'b0;
    XRAM[36125] = 8'b0;
    XRAM[36126] = 8'b0;
    XRAM[36127] = 8'b0;
    XRAM[36128] = 8'b0;
    XRAM[36129] = 8'b0;
    XRAM[36130] = 8'b0;
    XRAM[36131] = 8'b0;
    XRAM[36132] = 8'b0;
    XRAM[36133] = 8'b0;
    XRAM[36134] = 8'b0;
    XRAM[36135] = 8'b0;
    XRAM[36136] = 8'b0;
    XRAM[36137] = 8'b0;
    XRAM[36138] = 8'b0;
    XRAM[36139] = 8'b0;
    XRAM[36140] = 8'b0;
    XRAM[36141] = 8'b0;
    XRAM[36142] = 8'b0;
    XRAM[36143] = 8'b0;
    XRAM[36144] = 8'b0;
    XRAM[36145] = 8'b0;
    XRAM[36146] = 8'b0;
    XRAM[36147] = 8'b0;
    XRAM[36148] = 8'b0;
    XRAM[36149] = 8'b0;
    XRAM[36150] = 8'b0;
    XRAM[36151] = 8'b0;
    XRAM[36152] = 8'b0;
    XRAM[36153] = 8'b0;
    XRAM[36154] = 8'b0;
    XRAM[36155] = 8'b0;
    XRAM[36156] = 8'b0;
    XRAM[36157] = 8'b0;
    XRAM[36158] = 8'b0;
    XRAM[36159] = 8'b0;
    XRAM[36160] = 8'b0;
    XRAM[36161] = 8'b0;
    XRAM[36162] = 8'b0;
    XRAM[36163] = 8'b0;
    XRAM[36164] = 8'b0;
    XRAM[36165] = 8'b0;
    XRAM[36166] = 8'b0;
    XRAM[36167] = 8'b0;
    XRAM[36168] = 8'b0;
    XRAM[36169] = 8'b0;
    XRAM[36170] = 8'b0;
    XRAM[36171] = 8'b0;
    XRAM[36172] = 8'b0;
    XRAM[36173] = 8'b0;
    XRAM[36174] = 8'b0;
    XRAM[36175] = 8'b0;
    XRAM[36176] = 8'b0;
    XRAM[36177] = 8'b0;
    XRAM[36178] = 8'b0;
    XRAM[36179] = 8'b0;
    XRAM[36180] = 8'b0;
    XRAM[36181] = 8'b0;
    XRAM[36182] = 8'b0;
    XRAM[36183] = 8'b0;
    XRAM[36184] = 8'b0;
    XRAM[36185] = 8'b0;
    XRAM[36186] = 8'b0;
    XRAM[36187] = 8'b0;
    XRAM[36188] = 8'b0;
    XRAM[36189] = 8'b0;
    XRAM[36190] = 8'b0;
    XRAM[36191] = 8'b0;
    XRAM[36192] = 8'b0;
    XRAM[36193] = 8'b0;
    XRAM[36194] = 8'b0;
    XRAM[36195] = 8'b0;
    XRAM[36196] = 8'b0;
    XRAM[36197] = 8'b0;
    XRAM[36198] = 8'b0;
    XRAM[36199] = 8'b0;
    XRAM[36200] = 8'b0;
    XRAM[36201] = 8'b0;
    XRAM[36202] = 8'b0;
    XRAM[36203] = 8'b0;
    XRAM[36204] = 8'b0;
    XRAM[36205] = 8'b0;
    XRAM[36206] = 8'b0;
    XRAM[36207] = 8'b0;
    XRAM[36208] = 8'b0;
    XRAM[36209] = 8'b0;
    XRAM[36210] = 8'b0;
    XRAM[36211] = 8'b0;
    XRAM[36212] = 8'b0;
    XRAM[36213] = 8'b0;
    XRAM[36214] = 8'b0;
    XRAM[36215] = 8'b0;
    XRAM[36216] = 8'b0;
    XRAM[36217] = 8'b0;
    XRAM[36218] = 8'b0;
    XRAM[36219] = 8'b0;
    XRAM[36220] = 8'b0;
    XRAM[36221] = 8'b0;
    XRAM[36222] = 8'b0;
    XRAM[36223] = 8'b0;
    XRAM[36224] = 8'b0;
    XRAM[36225] = 8'b0;
    XRAM[36226] = 8'b0;
    XRAM[36227] = 8'b0;
    XRAM[36228] = 8'b0;
    XRAM[36229] = 8'b0;
    XRAM[36230] = 8'b0;
    XRAM[36231] = 8'b0;
    XRAM[36232] = 8'b0;
    XRAM[36233] = 8'b0;
    XRAM[36234] = 8'b0;
    XRAM[36235] = 8'b0;
    XRAM[36236] = 8'b0;
    XRAM[36237] = 8'b0;
    XRAM[36238] = 8'b0;
    XRAM[36239] = 8'b0;
    XRAM[36240] = 8'b0;
    XRAM[36241] = 8'b0;
    XRAM[36242] = 8'b0;
    XRAM[36243] = 8'b0;
    XRAM[36244] = 8'b0;
    XRAM[36245] = 8'b0;
    XRAM[36246] = 8'b0;
    XRAM[36247] = 8'b0;
    XRAM[36248] = 8'b0;
    XRAM[36249] = 8'b0;
    XRAM[36250] = 8'b0;
    XRAM[36251] = 8'b0;
    XRAM[36252] = 8'b0;
    XRAM[36253] = 8'b0;
    XRAM[36254] = 8'b0;
    XRAM[36255] = 8'b0;
    XRAM[36256] = 8'b0;
    XRAM[36257] = 8'b0;
    XRAM[36258] = 8'b0;
    XRAM[36259] = 8'b0;
    XRAM[36260] = 8'b0;
    XRAM[36261] = 8'b0;
    XRAM[36262] = 8'b0;
    XRAM[36263] = 8'b0;
    XRAM[36264] = 8'b0;
    XRAM[36265] = 8'b0;
    XRAM[36266] = 8'b0;
    XRAM[36267] = 8'b0;
    XRAM[36268] = 8'b0;
    XRAM[36269] = 8'b0;
    XRAM[36270] = 8'b0;
    XRAM[36271] = 8'b0;
    XRAM[36272] = 8'b0;
    XRAM[36273] = 8'b0;
    XRAM[36274] = 8'b0;
    XRAM[36275] = 8'b0;
    XRAM[36276] = 8'b0;
    XRAM[36277] = 8'b0;
    XRAM[36278] = 8'b0;
    XRAM[36279] = 8'b0;
    XRAM[36280] = 8'b0;
    XRAM[36281] = 8'b0;
    XRAM[36282] = 8'b0;
    XRAM[36283] = 8'b0;
    XRAM[36284] = 8'b0;
    XRAM[36285] = 8'b0;
    XRAM[36286] = 8'b0;
    XRAM[36287] = 8'b0;
    XRAM[36288] = 8'b0;
    XRAM[36289] = 8'b0;
    XRAM[36290] = 8'b0;
    XRAM[36291] = 8'b0;
    XRAM[36292] = 8'b0;
    XRAM[36293] = 8'b0;
    XRAM[36294] = 8'b0;
    XRAM[36295] = 8'b0;
    XRAM[36296] = 8'b0;
    XRAM[36297] = 8'b0;
    XRAM[36298] = 8'b0;
    XRAM[36299] = 8'b0;
    XRAM[36300] = 8'b0;
    XRAM[36301] = 8'b0;
    XRAM[36302] = 8'b0;
    XRAM[36303] = 8'b0;
    XRAM[36304] = 8'b0;
    XRAM[36305] = 8'b0;
    XRAM[36306] = 8'b0;
    XRAM[36307] = 8'b0;
    XRAM[36308] = 8'b0;
    XRAM[36309] = 8'b0;
    XRAM[36310] = 8'b0;
    XRAM[36311] = 8'b0;
    XRAM[36312] = 8'b0;
    XRAM[36313] = 8'b0;
    XRAM[36314] = 8'b0;
    XRAM[36315] = 8'b0;
    XRAM[36316] = 8'b0;
    XRAM[36317] = 8'b0;
    XRAM[36318] = 8'b0;
    XRAM[36319] = 8'b0;
    XRAM[36320] = 8'b0;
    XRAM[36321] = 8'b0;
    XRAM[36322] = 8'b0;
    XRAM[36323] = 8'b0;
    XRAM[36324] = 8'b0;
    XRAM[36325] = 8'b0;
    XRAM[36326] = 8'b0;
    XRAM[36327] = 8'b0;
    XRAM[36328] = 8'b0;
    XRAM[36329] = 8'b0;
    XRAM[36330] = 8'b0;
    XRAM[36331] = 8'b0;
    XRAM[36332] = 8'b0;
    XRAM[36333] = 8'b0;
    XRAM[36334] = 8'b0;
    XRAM[36335] = 8'b0;
    XRAM[36336] = 8'b0;
    XRAM[36337] = 8'b0;
    XRAM[36338] = 8'b0;
    XRAM[36339] = 8'b0;
    XRAM[36340] = 8'b0;
    XRAM[36341] = 8'b0;
    XRAM[36342] = 8'b0;
    XRAM[36343] = 8'b0;
    XRAM[36344] = 8'b0;
    XRAM[36345] = 8'b0;
    XRAM[36346] = 8'b0;
    XRAM[36347] = 8'b0;
    XRAM[36348] = 8'b0;
    XRAM[36349] = 8'b0;
    XRAM[36350] = 8'b0;
    XRAM[36351] = 8'b0;
    XRAM[36352] = 8'b0;
    XRAM[36353] = 8'b0;
    XRAM[36354] = 8'b0;
    XRAM[36355] = 8'b0;
    XRAM[36356] = 8'b0;
    XRAM[36357] = 8'b0;
    XRAM[36358] = 8'b0;
    XRAM[36359] = 8'b0;
    XRAM[36360] = 8'b0;
    XRAM[36361] = 8'b0;
    XRAM[36362] = 8'b0;
    XRAM[36363] = 8'b0;
    XRAM[36364] = 8'b0;
    XRAM[36365] = 8'b0;
    XRAM[36366] = 8'b0;
    XRAM[36367] = 8'b0;
    XRAM[36368] = 8'b0;
    XRAM[36369] = 8'b0;
    XRAM[36370] = 8'b0;
    XRAM[36371] = 8'b0;
    XRAM[36372] = 8'b0;
    XRAM[36373] = 8'b0;
    XRAM[36374] = 8'b0;
    XRAM[36375] = 8'b0;
    XRAM[36376] = 8'b0;
    XRAM[36377] = 8'b0;
    XRAM[36378] = 8'b0;
    XRAM[36379] = 8'b0;
    XRAM[36380] = 8'b0;
    XRAM[36381] = 8'b0;
    XRAM[36382] = 8'b0;
    XRAM[36383] = 8'b0;
    XRAM[36384] = 8'b0;
    XRAM[36385] = 8'b0;
    XRAM[36386] = 8'b0;
    XRAM[36387] = 8'b0;
    XRAM[36388] = 8'b0;
    XRAM[36389] = 8'b0;
    XRAM[36390] = 8'b0;
    XRAM[36391] = 8'b0;
    XRAM[36392] = 8'b0;
    XRAM[36393] = 8'b0;
    XRAM[36394] = 8'b0;
    XRAM[36395] = 8'b0;
    XRAM[36396] = 8'b0;
    XRAM[36397] = 8'b0;
    XRAM[36398] = 8'b0;
    XRAM[36399] = 8'b0;
    XRAM[36400] = 8'b0;
    XRAM[36401] = 8'b0;
    XRAM[36402] = 8'b0;
    XRAM[36403] = 8'b0;
    XRAM[36404] = 8'b0;
    XRAM[36405] = 8'b0;
    XRAM[36406] = 8'b0;
    XRAM[36407] = 8'b0;
    XRAM[36408] = 8'b0;
    XRAM[36409] = 8'b0;
    XRAM[36410] = 8'b0;
    XRAM[36411] = 8'b0;
    XRAM[36412] = 8'b0;
    XRAM[36413] = 8'b0;
    XRAM[36414] = 8'b0;
    XRAM[36415] = 8'b0;
    XRAM[36416] = 8'b0;
    XRAM[36417] = 8'b0;
    XRAM[36418] = 8'b0;
    XRAM[36419] = 8'b0;
    XRAM[36420] = 8'b0;
    XRAM[36421] = 8'b0;
    XRAM[36422] = 8'b0;
    XRAM[36423] = 8'b0;
    XRAM[36424] = 8'b0;
    XRAM[36425] = 8'b0;
    XRAM[36426] = 8'b0;
    XRAM[36427] = 8'b0;
    XRAM[36428] = 8'b0;
    XRAM[36429] = 8'b0;
    XRAM[36430] = 8'b0;
    XRAM[36431] = 8'b0;
    XRAM[36432] = 8'b0;
    XRAM[36433] = 8'b0;
    XRAM[36434] = 8'b0;
    XRAM[36435] = 8'b0;
    XRAM[36436] = 8'b0;
    XRAM[36437] = 8'b0;
    XRAM[36438] = 8'b0;
    XRAM[36439] = 8'b0;
    XRAM[36440] = 8'b0;
    XRAM[36441] = 8'b0;
    XRAM[36442] = 8'b0;
    XRAM[36443] = 8'b0;
    XRAM[36444] = 8'b0;
    XRAM[36445] = 8'b0;
    XRAM[36446] = 8'b0;
    XRAM[36447] = 8'b0;
    XRAM[36448] = 8'b0;
    XRAM[36449] = 8'b0;
    XRAM[36450] = 8'b0;
    XRAM[36451] = 8'b0;
    XRAM[36452] = 8'b0;
    XRAM[36453] = 8'b0;
    XRAM[36454] = 8'b0;
    XRAM[36455] = 8'b0;
    XRAM[36456] = 8'b0;
    XRAM[36457] = 8'b0;
    XRAM[36458] = 8'b0;
    XRAM[36459] = 8'b0;
    XRAM[36460] = 8'b0;
    XRAM[36461] = 8'b0;
    XRAM[36462] = 8'b0;
    XRAM[36463] = 8'b0;
    XRAM[36464] = 8'b0;
    XRAM[36465] = 8'b0;
    XRAM[36466] = 8'b0;
    XRAM[36467] = 8'b0;
    XRAM[36468] = 8'b0;
    XRAM[36469] = 8'b0;
    XRAM[36470] = 8'b0;
    XRAM[36471] = 8'b0;
    XRAM[36472] = 8'b0;
    XRAM[36473] = 8'b0;
    XRAM[36474] = 8'b0;
    XRAM[36475] = 8'b0;
    XRAM[36476] = 8'b0;
    XRAM[36477] = 8'b0;
    XRAM[36478] = 8'b0;
    XRAM[36479] = 8'b0;
    XRAM[36480] = 8'b0;
    XRAM[36481] = 8'b0;
    XRAM[36482] = 8'b0;
    XRAM[36483] = 8'b0;
    XRAM[36484] = 8'b0;
    XRAM[36485] = 8'b0;
    XRAM[36486] = 8'b0;
    XRAM[36487] = 8'b0;
    XRAM[36488] = 8'b0;
    XRAM[36489] = 8'b0;
    XRAM[36490] = 8'b0;
    XRAM[36491] = 8'b0;
    XRAM[36492] = 8'b0;
    XRAM[36493] = 8'b0;
    XRAM[36494] = 8'b0;
    XRAM[36495] = 8'b0;
    XRAM[36496] = 8'b0;
    XRAM[36497] = 8'b0;
    XRAM[36498] = 8'b0;
    XRAM[36499] = 8'b0;
    XRAM[36500] = 8'b0;
    XRAM[36501] = 8'b0;
    XRAM[36502] = 8'b0;
    XRAM[36503] = 8'b0;
    XRAM[36504] = 8'b0;
    XRAM[36505] = 8'b0;
    XRAM[36506] = 8'b0;
    XRAM[36507] = 8'b0;
    XRAM[36508] = 8'b0;
    XRAM[36509] = 8'b0;
    XRAM[36510] = 8'b0;
    XRAM[36511] = 8'b0;
    XRAM[36512] = 8'b0;
    XRAM[36513] = 8'b0;
    XRAM[36514] = 8'b0;
    XRAM[36515] = 8'b0;
    XRAM[36516] = 8'b0;
    XRAM[36517] = 8'b0;
    XRAM[36518] = 8'b0;
    XRAM[36519] = 8'b0;
    XRAM[36520] = 8'b0;
    XRAM[36521] = 8'b0;
    XRAM[36522] = 8'b0;
    XRAM[36523] = 8'b0;
    XRAM[36524] = 8'b0;
    XRAM[36525] = 8'b0;
    XRAM[36526] = 8'b0;
    XRAM[36527] = 8'b0;
    XRAM[36528] = 8'b0;
    XRAM[36529] = 8'b0;
    XRAM[36530] = 8'b0;
    XRAM[36531] = 8'b0;
    XRAM[36532] = 8'b0;
    XRAM[36533] = 8'b0;
    XRAM[36534] = 8'b0;
    XRAM[36535] = 8'b0;
    XRAM[36536] = 8'b0;
    XRAM[36537] = 8'b0;
    XRAM[36538] = 8'b0;
    XRAM[36539] = 8'b0;
    XRAM[36540] = 8'b0;
    XRAM[36541] = 8'b0;
    XRAM[36542] = 8'b0;
    XRAM[36543] = 8'b0;
    XRAM[36544] = 8'b0;
    XRAM[36545] = 8'b0;
    XRAM[36546] = 8'b0;
    XRAM[36547] = 8'b0;
    XRAM[36548] = 8'b0;
    XRAM[36549] = 8'b0;
    XRAM[36550] = 8'b0;
    XRAM[36551] = 8'b0;
    XRAM[36552] = 8'b0;
    XRAM[36553] = 8'b0;
    XRAM[36554] = 8'b0;
    XRAM[36555] = 8'b0;
    XRAM[36556] = 8'b0;
    XRAM[36557] = 8'b0;
    XRAM[36558] = 8'b0;
    XRAM[36559] = 8'b0;
    XRAM[36560] = 8'b0;
    XRAM[36561] = 8'b0;
    XRAM[36562] = 8'b0;
    XRAM[36563] = 8'b0;
    XRAM[36564] = 8'b0;
    XRAM[36565] = 8'b0;
    XRAM[36566] = 8'b0;
    XRAM[36567] = 8'b0;
    XRAM[36568] = 8'b0;
    XRAM[36569] = 8'b0;
    XRAM[36570] = 8'b0;
    XRAM[36571] = 8'b0;
    XRAM[36572] = 8'b0;
    XRAM[36573] = 8'b0;
    XRAM[36574] = 8'b0;
    XRAM[36575] = 8'b0;
    XRAM[36576] = 8'b0;
    XRAM[36577] = 8'b0;
    XRAM[36578] = 8'b0;
    XRAM[36579] = 8'b0;
    XRAM[36580] = 8'b0;
    XRAM[36581] = 8'b0;
    XRAM[36582] = 8'b0;
    XRAM[36583] = 8'b0;
    XRAM[36584] = 8'b0;
    XRAM[36585] = 8'b0;
    XRAM[36586] = 8'b0;
    XRAM[36587] = 8'b0;
    XRAM[36588] = 8'b0;
    XRAM[36589] = 8'b0;
    XRAM[36590] = 8'b0;
    XRAM[36591] = 8'b0;
    XRAM[36592] = 8'b0;
    XRAM[36593] = 8'b0;
    XRAM[36594] = 8'b0;
    XRAM[36595] = 8'b0;
    XRAM[36596] = 8'b0;
    XRAM[36597] = 8'b0;
    XRAM[36598] = 8'b0;
    XRAM[36599] = 8'b0;
    XRAM[36600] = 8'b0;
    XRAM[36601] = 8'b0;
    XRAM[36602] = 8'b0;
    XRAM[36603] = 8'b0;
    XRAM[36604] = 8'b0;
    XRAM[36605] = 8'b0;
    XRAM[36606] = 8'b0;
    XRAM[36607] = 8'b0;
    XRAM[36608] = 8'b0;
    XRAM[36609] = 8'b0;
    XRAM[36610] = 8'b0;
    XRAM[36611] = 8'b0;
    XRAM[36612] = 8'b0;
    XRAM[36613] = 8'b0;
    XRAM[36614] = 8'b0;
    XRAM[36615] = 8'b0;
    XRAM[36616] = 8'b0;
    XRAM[36617] = 8'b0;
    XRAM[36618] = 8'b0;
    XRAM[36619] = 8'b0;
    XRAM[36620] = 8'b0;
    XRAM[36621] = 8'b0;
    XRAM[36622] = 8'b0;
    XRAM[36623] = 8'b0;
    XRAM[36624] = 8'b0;
    XRAM[36625] = 8'b0;
    XRAM[36626] = 8'b0;
    XRAM[36627] = 8'b0;
    XRAM[36628] = 8'b0;
    XRAM[36629] = 8'b0;
    XRAM[36630] = 8'b0;
    XRAM[36631] = 8'b0;
    XRAM[36632] = 8'b0;
    XRAM[36633] = 8'b0;
    XRAM[36634] = 8'b0;
    XRAM[36635] = 8'b0;
    XRAM[36636] = 8'b0;
    XRAM[36637] = 8'b0;
    XRAM[36638] = 8'b0;
    XRAM[36639] = 8'b0;
    XRAM[36640] = 8'b0;
    XRAM[36641] = 8'b0;
    XRAM[36642] = 8'b0;
    XRAM[36643] = 8'b0;
    XRAM[36644] = 8'b0;
    XRAM[36645] = 8'b0;
    XRAM[36646] = 8'b0;
    XRAM[36647] = 8'b0;
    XRAM[36648] = 8'b0;
    XRAM[36649] = 8'b0;
    XRAM[36650] = 8'b0;
    XRAM[36651] = 8'b0;
    XRAM[36652] = 8'b0;
    XRAM[36653] = 8'b0;
    XRAM[36654] = 8'b0;
    XRAM[36655] = 8'b0;
    XRAM[36656] = 8'b0;
    XRAM[36657] = 8'b0;
    XRAM[36658] = 8'b0;
    XRAM[36659] = 8'b0;
    XRAM[36660] = 8'b0;
    XRAM[36661] = 8'b0;
    XRAM[36662] = 8'b0;
    XRAM[36663] = 8'b0;
    XRAM[36664] = 8'b0;
    XRAM[36665] = 8'b0;
    XRAM[36666] = 8'b0;
    XRAM[36667] = 8'b0;
    XRAM[36668] = 8'b0;
    XRAM[36669] = 8'b0;
    XRAM[36670] = 8'b0;
    XRAM[36671] = 8'b0;
    XRAM[36672] = 8'b0;
    XRAM[36673] = 8'b0;
    XRAM[36674] = 8'b0;
    XRAM[36675] = 8'b0;
    XRAM[36676] = 8'b0;
    XRAM[36677] = 8'b0;
    XRAM[36678] = 8'b0;
    XRAM[36679] = 8'b0;
    XRAM[36680] = 8'b0;
    XRAM[36681] = 8'b0;
    XRAM[36682] = 8'b0;
    XRAM[36683] = 8'b0;
    XRAM[36684] = 8'b0;
    XRAM[36685] = 8'b0;
    XRAM[36686] = 8'b0;
    XRAM[36687] = 8'b0;
    XRAM[36688] = 8'b0;
    XRAM[36689] = 8'b0;
    XRAM[36690] = 8'b0;
    XRAM[36691] = 8'b0;
    XRAM[36692] = 8'b0;
    XRAM[36693] = 8'b0;
    XRAM[36694] = 8'b0;
    XRAM[36695] = 8'b0;
    XRAM[36696] = 8'b0;
    XRAM[36697] = 8'b0;
    XRAM[36698] = 8'b0;
    XRAM[36699] = 8'b0;
    XRAM[36700] = 8'b0;
    XRAM[36701] = 8'b0;
    XRAM[36702] = 8'b0;
    XRAM[36703] = 8'b0;
    XRAM[36704] = 8'b0;
    XRAM[36705] = 8'b0;
    XRAM[36706] = 8'b0;
    XRAM[36707] = 8'b0;
    XRAM[36708] = 8'b0;
    XRAM[36709] = 8'b0;
    XRAM[36710] = 8'b0;
    XRAM[36711] = 8'b0;
    XRAM[36712] = 8'b0;
    XRAM[36713] = 8'b0;
    XRAM[36714] = 8'b0;
    XRAM[36715] = 8'b0;
    XRAM[36716] = 8'b0;
    XRAM[36717] = 8'b0;
    XRAM[36718] = 8'b0;
    XRAM[36719] = 8'b0;
    XRAM[36720] = 8'b0;
    XRAM[36721] = 8'b0;
    XRAM[36722] = 8'b0;
    XRAM[36723] = 8'b0;
    XRAM[36724] = 8'b0;
    XRAM[36725] = 8'b0;
    XRAM[36726] = 8'b0;
    XRAM[36727] = 8'b0;
    XRAM[36728] = 8'b0;
    XRAM[36729] = 8'b0;
    XRAM[36730] = 8'b0;
    XRAM[36731] = 8'b0;
    XRAM[36732] = 8'b0;
    XRAM[36733] = 8'b0;
    XRAM[36734] = 8'b0;
    XRAM[36735] = 8'b0;
    XRAM[36736] = 8'b0;
    XRAM[36737] = 8'b0;
    XRAM[36738] = 8'b0;
    XRAM[36739] = 8'b0;
    XRAM[36740] = 8'b0;
    XRAM[36741] = 8'b0;
    XRAM[36742] = 8'b0;
    XRAM[36743] = 8'b0;
    XRAM[36744] = 8'b0;
    XRAM[36745] = 8'b0;
    XRAM[36746] = 8'b0;
    XRAM[36747] = 8'b0;
    XRAM[36748] = 8'b0;
    XRAM[36749] = 8'b0;
    XRAM[36750] = 8'b0;
    XRAM[36751] = 8'b0;
    XRAM[36752] = 8'b0;
    XRAM[36753] = 8'b0;
    XRAM[36754] = 8'b0;
    XRAM[36755] = 8'b0;
    XRAM[36756] = 8'b0;
    XRAM[36757] = 8'b0;
    XRAM[36758] = 8'b0;
    XRAM[36759] = 8'b0;
    XRAM[36760] = 8'b0;
    XRAM[36761] = 8'b0;
    XRAM[36762] = 8'b0;
    XRAM[36763] = 8'b0;
    XRAM[36764] = 8'b0;
    XRAM[36765] = 8'b0;
    XRAM[36766] = 8'b0;
    XRAM[36767] = 8'b0;
    XRAM[36768] = 8'b0;
    XRAM[36769] = 8'b0;
    XRAM[36770] = 8'b0;
    XRAM[36771] = 8'b0;
    XRAM[36772] = 8'b0;
    XRAM[36773] = 8'b0;
    XRAM[36774] = 8'b0;
    XRAM[36775] = 8'b0;
    XRAM[36776] = 8'b0;
    XRAM[36777] = 8'b0;
    XRAM[36778] = 8'b0;
    XRAM[36779] = 8'b0;
    XRAM[36780] = 8'b0;
    XRAM[36781] = 8'b0;
    XRAM[36782] = 8'b0;
    XRAM[36783] = 8'b0;
    XRAM[36784] = 8'b0;
    XRAM[36785] = 8'b0;
    XRAM[36786] = 8'b0;
    XRAM[36787] = 8'b0;
    XRAM[36788] = 8'b0;
    XRAM[36789] = 8'b0;
    XRAM[36790] = 8'b0;
    XRAM[36791] = 8'b0;
    XRAM[36792] = 8'b0;
    XRAM[36793] = 8'b0;
    XRAM[36794] = 8'b0;
    XRAM[36795] = 8'b0;
    XRAM[36796] = 8'b0;
    XRAM[36797] = 8'b0;
    XRAM[36798] = 8'b0;
    XRAM[36799] = 8'b0;
    XRAM[36800] = 8'b0;
    XRAM[36801] = 8'b0;
    XRAM[36802] = 8'b0;
    XRAM[36803] = 8'b0;
    XRAM[36804] = 8'b0;
    XRAM[36805] = 8'b0;
    XRAM[36806] = 8'b0;
    XRAM[36807] = 8'b0;
    XRAM[36808] = 8'b0;
    XRAM[36809] = 8'b0;
    XRAM[36810] = 8'b0;
    XRAM[36811] = 8'b0;
    XRAM[36812] = 8'b0;
    XRAM[36813] = 8'b0;
    XRAM[36814] = 8'b0;
    XRAM[36815] = 8'b0;
    XRAM[36816] = 8'b0;
    XRAM[36817] = 8'b0;
    XRAM[36818] = 8'b0;
    XRAM[36819] = 8'b0;
    XRAM[36820] = 8'b0;
    XRAM[36821] = 8'b0;
    XRAM[36822] = 8'b0;
    XRAM[36823] = 8'b0;
    XRAM[36824] = 8'b0;
    XRAM[36825] = 8'b0;
    XRAM[36826] = 8'b0;
    XRAM[36827] = 8'b0;
    XRAM[36828] = 8'b0;
    XRAM[36829] = 8'b0;
    XRAM[36830] = 8'b0;
    XRAM[36831] = 8'b0;
    XRAM[36832] = 8'b0;
    XRAM[36833] = 8'b0;
    XRAM[36834] = 8'b0;
    XRAM[36835] = 8'b0;
    XRAM[36836] = 8'b0;
    XRAM[36837] = 8'b0;
    XRAM[36838] = 8'b0;
    XRAM[36839] = 8'b0;
    XRAM[36840] = 8'b0;
    XRAM[36841] = 8'b0;
    XRAM[36842] = 8'b0;
    XRAM[36843] = 8'b0;
    XRAM[36844] = 8'b0;
    XRAM[36845] = 8'b0;
    XRAM[36846] = 8'b0;
    XRAM[36847] = 8'b0;
    XRAM[36848] = 8'b0;
    XRAM[36849] = 8'b0;
    XRAM[36850] = 8'b0;
    XRAM[36851] = 8'b0;
    XRAM[36852] = 8'b0;
    XRAM[36853] = 8'b0;
    XRAM[36854] = 8'b0;
    XRAM[36855] = 8'b0;
    XRAM[36856] = 8'b0;
    XRAM[36857] = 8'b0;
    XRAM[36858] = 8'b0;
    XRAM[36859] = 8'b0;
    XRAM[36860] = 8'b0;
    XRAM[36861] = 8'b0;
    XRAM[36862] = 8'b0;
    XRAM[36863] = 8'b0;
    XRAM[36864] = 8'b0;
    XRAM[36865] = 8'b0;
    XRAM[36866] = 8'b0;
    XRAM[36867] = 8'b0;
    XRAM[36868] = 8'b0;
    XRAM[36869] = 8'b0;
    XRAM[36870] = 8'b0;
    XRAM[36871] = 8'b0;
    XRAM[36872] = 8'b0;
    XRAM[36873] = 8'b0;
    XRAM[36874] = 8'b0;
    XRAM[36875] = 8'b0;
    XRAM[36876] = 8'b0;
    XRAM[36877] = 8'b0;
    XRAM[36878] = 8'b0;
    XRAM[36879] = 8'b0;
    XRAM[36880] = 8'b0;
    XRAM[36881] = 8'b0;
    XRAM[36882] = 8'b0;
    XRAM[36883] = 8'b0;
    XRAM[36884] = 8'b0;
    XRAM[36885] = 8'b0;
    XRAM[36886] = 8'b0;
    XRAM[36887] = 8'b0;
    XRAM[36888] = 8'b0;
    XRAM[36889] = 8'b0;
    XRAM[36890] = 8'b0;
    XRAM[36891] = 8'b0;
    XRAM[36892] = 8'b0;
    XRAM[36893] = 8'b0;
    XRAM[36894] = 8'b0;
    XRAM[36895] = 8'b0;
    XRAM[36896] = 8'b0;
    XRAM[36897] = 8'b0;
    XRAM[36898] = 8'b0;
    XRAM[36899] = 8'b0;
    XRAM[36900] = 8'b0;
    XRAM[36901] = 8'b0;
    XRAM[36902] = 8'b0;
    XRAM[36903] = 8'b0;
    XRAM[36904] = 8'b0;
    XRAM[36905] = 8'b0;
    XRAM[36906] = 8'b0;
    XRAM[36907] = 8'b0;
    XRAM[36908] = 8'b0;
    XRAM[36909] = 8'b0;
    XRAM[36910] = 8'b0;
    XRAM[36911] = 8'b0;
    XRAM[36912] = 8'b0;
    XRAM[36913] = 8'b0;
    XRAM[36914] = 8'b0;
    XRAM[36915] = 8'b0;
    XRAM[36916] = 8'b0;
    XRAM[36917] = 8'b0;
    XRAM[36918] = 8'b0;
    XRAM[36919] = 8'b0;
    XRAM[36920] = 8'b0;
    XRAM[36921] = 8'b0;
    XRAM[36922] = 8'b0;
    XRAM[36923] = 8'b0;
    XRAM[36924] = 8'b0;
    XRAM[36925] = 8'b0;
    XRAM[36926] = 8'b0;
    XRAM[36927] = 8'b0;
    XRAM[36928] = 8'b0;
    XRAM[36929] = 8'b0;
    XRAM[36930] = 8'b0;
    XRAM[36931] = 8'b0;
    XRAM[36932] = 8'b0;
    XRAM[36933] = 8'b0;
    XRAM[36934] = 8'b0;
    XRAM[36935] = 8'b0;
    XRAM[36936] = 8'b0;
    XRAM[36937] = 8'b0;
    XRAM[36938] = 8'b0;
    XRAM[36939] = 8'b0;
    XRAM[36940] = 8'b0;
    XRAM[36941] = 8'b0;
    XRAM[36942] = 8'b0;
    XRAM[36943] = 8'b0;
    XRAM[36944] = 8'b0;
    XRAM[36945] = 8'b0;
    XRAM[36946] = 8'b0;
    XRAM[36947] = 8'b0;
    XRAM[36948] = 8'b0;
    XRAM[36949] = 8'b0;
    XRAM[36950] = 8'b0;
    XRAM[36951] = 8'b0;
    XRAM[36952] = 8'b0;
    XRAM[36953] = 8'b0;
    XRAM[36954] = 8'b0;
    XRAM[36955] = 8'b0;
    XRAM[36956] = 8'b0;
    XRAM[36957] = 8'b0;
    XRAM[36958] = 8'b0;
    XRAM[36959] = 8'b0;
    XRAM[36960] = 8'b0;
    XRAM[36961] = 8'b0;
    XRAM[36962] = 8'b0;
    XRAM[36963] = 8'b0;
    XRAM[36964] = 8'b0;
    XRAM[36965] = 8'b0;
    XRAM[36966] = 8'b0;
    XRAM[36967] = 8'b0;
    XRAM[36968] = 8'b0;
    XRAM[36969] = 8'b0;
    XRAM[36970] = 8'b0;
    XRAM[36971] = 8'b0;
    XRAM[36972] = 8'b0;
    XRAM[36973] = 8'b0;
    XRAM[36974] = 8'b0;
    XRAM[36975] = 8'b0;
    XRAM[36976] = 8'b0;
    XRAM[36977] = 8'b0;
    XRAM[36978] = 8'b0;
    XRAM[36979] = 8'b0;
    XRAM[36980] = 8'b0;
    XRAM[36981] = 8'b0;
    XRAM[36982] = 8'b0;
    XRAM[36983] = 8'b0;
    XRAM[36984] = 8'b0;
    XRAM[36985] = 8'b0;
    XRAM[36986] = 8'b0;
    XRAM[36987] = 8'b0;
    XRAM[36988] = 8'b0;
    XRAM[36989] = 8'b0;
    XRAM[36990] = 8'b0;
    XRAM[36991] = 8'b0;
    XRAM[36992] = 8'b0;
    XRAM[36993] = 8'b0;
    XRAM[36994] = 8'b0;
    XRAM[36995] = 8'b0;
    XRAM[36996] = 8'b0;
    XRAM[36997] = 8'b0;
    XRAM[36998] = 8'b0;
    XRAM[36999] = 8'b0;
    XRAM[37000] = 8'b0;
    XRAM[37001] = 8'b0;
    XRAM[37002] = 8'b0;
    XRAM[37003] = 8'b0;
    XRAM[37004] = 8'b0;
    XRAM[37005] = 8'b0;
    XRAM[37006] = 8'b0;
    XRAM[37007] = 8'b0;
    XRAM[37008] = 8'b0;
    XRAM[37009] = 8'b0;
    XRAM[37010] = 8'b0;
    XRAM[37011] = 8'b0;
    XRAM[37012] = 8'b0;
    XRAM[37013] = 8'b0;
    XRAM[37014] = 8'b0;
    XRAM[37015] = 8'b0;
    XRAM[37016] = 8'b0;
    XRAM[37017] = 8'b0;
    XRAM[37018] = 8'b0;
    XRAM[37019] = 8'b0;
    XRAM[37020] = 8'b0;
    XRAM[37021] = 8'b0;
    XRAM[37022] = 8'b0;
    XRAM[37023] = 8'b0;
    XRAM[37024] = 8'b0;
    XRAM[37025] = 8'b0;
    XRAM[37026] = 8'b0;
    XRAM[37027] = 8'b0;
    XRAM[37028] = 8'b0;
    XRAM[37029] = 8'b0;
    XRAM[37030] = 8'b0;
    XRAM[37031] = 8'b0;
    XRAM[37032] = 8'b0;
    XRAM[37033] = 8'b0;
    XRAM[37034] = 8'b0;
    XRAM[37035] = 8'b0;
    XRAM[37036] = 8'b0;
    XRAM[37037] = 8'b0;
    XRAM[37038] = 8'b0;
    XRAM[37039] = 8'b0;
    XRAM[37040] = 8'b0;
    XRAM[37041] = 8'b0;
    XRAM[37042] = 8'b0;
    XRAM[37043] = 8'b0;
    XRAM[37044] = 8'b0;
    XRAM[37045] = 8'b0;
    XRAM[37046] = 8'b0;
    XRAM[37047] = 8'b0;
    XRAM[37048] = 8'b0;
    XRAM[37049] = 8'b0;
    XRAM[37050] = 8'b0;
    XRAM[37051] = 8'b0;
    XRAM[37052] = 8'b0;
    XRAM[37053] = 8'b0;
    XRAM[37054] = 8'b0;
    XRAM[37055] = 8'b0;
    XRAM[37056] = 8'b0;
    XRAM[37057] = 8'b0;
    XRAM[37058] = 8'b0;
    XRAM[37059] = 8'b0;
    XRAM[37060] = 8'b0;
    XRAM[37061] = 8'b0;
    XRAM[37062] = 8'b0;
    XRAM[37063] = 8'b0;
    XRAM[37064] = 8'b0;
    XRAM[37065] = 8'b0;
    XRAM[37066] = 8'b0;
    XRAM[37067] = 8'b0;
    XRAM[37068] = 8'b0;
    XRAM[37069] = 8'b0;
    XRAM[37070] = 8'b0;
    XRAM[37071] = 8'b0;
    XRAM[37072] = 8'b0;
    XRAM[37073] = 8'b0;
    XRAM[37074] = 8'b0;
    XRAM[37075] = 8'b0;
    XRAM[37076] = 8'b0;
    XRAM[37077] = 8'b0;
    XRAM[37078] = 8'b0;
    XRAM[37079] = 8'b0;
    XRAM[37080] = 8'b0;
    XRAM[37081] = 8'b0;
    XRAM[37082] = 8'b0;
    XRAM[37083] = 8'b0;
    XRAM[37084] = 8'b0;
    XRAM[37085] = 8'b0;
    XRAM[37086] = 8'b0;
    XRAM[37087] = 8'b0;
    XRAM[37088] = 8'b0;
    XRAM[37089] = 8'b0;
    XRAM[37090] = 8'b0;
    XRAM[37091] = 8'b0;
    XRAM[37092] = 8'b0;
    XRAM[37093] = 8'b0;
    XRAM[37094] = 8'b0;
    XRAM[37095] = 8'b0;
    XRAM[37096] = 8'b0;
    XRAM[37097] = 8'b0;
    XRAM[37098] = 8'b0;
    XRAM[37099] = 8'b0;
    XRAM[37100] = 8'b0;
    XRAM[37101] = 8'b0;
    XRAM[37102] = 8'b0;
    XRAM[37103] = 8'b0;
    XRAM[37104] = 8'b0;
    XRAM[37105] = 8'b0;
    XRAM[37106] = 8'b0;
    XRAM[37107] = 8'b0;
    XRAM[37108] = 8'b0;
    XRAM[37109] = 8'b0;
    XRAM[37110] = 8'b0;
    XRAM[37111] = 8'b0;
    XRAM[37112] = 8'b0;
    XRAM[37113] = 8'b0;
    XRAM[37114] = 8'b0;
    XRAM[37115] = 8'b0;
    XRAM[37116] = 8'b0;
    XRAM[37117] = 8'b0;
    XRAM[37118] = 8'b0;
    XRAM[37119] = 8'b0;
    XRAM[37120] = 8'b0;
    XRAM[37121] = 8'b0;
    XRAM[37122] = 8'b0;
    XRAM[37123] = 8'b0;
    XRAM[37124] = 8'b0;
    XRAM[37125] = 8'b0;
    XRAM[37126] = 8'b0;
    XRAM[37127] = 8'b0;
    XRAM[37128] = 8'b0;
    XRAM[37129] = 8'b0;
    XRAM[37130] = 8'b0;
    XRAM[37131] = 8'b0;
    XRAM[37132] = 8'b0;
    XRAM[37133] = 8'b0;
    XRAM[37134] = 8'b0;
    XRAM[37135] = 8'b0;
    XRAM[37136] = 8'b0;
    XRAM[37137] = 8'b0;
    XRAM[37138] = 8'b0;
    XRAM[37139] = 8'b0;
    XRAM[37140] = 8'b0;
    XRAM[37141] = 8'b0;
    XRAM[37142] = 8'b0;
    XRAM[37143] = 8'b0;
    XRAM[37144] = 8'b0;
    XRAM[37145] = 8'b0;
    XRAM[37146] = 8'b0;
    XRAM[37147] = 8'b0;
    XRAM[37148] = 8'b0;
    XRAM[37149] = 8'b0;
    XRAM[37150] = 8'b0;
    XRAM[37151] = 8'b0;
    XRAM[37152] = 8'b0;
    XRAM[37153] = 8'b0;
    XRAM[37154] = 8'b0;
    XRAM[37155] = 8'b0;
    XRAM[37156] = 8'b0;
    XRAM[37157] = 8'b0;
    XRAM[37158] = 8'b0;
    XRAM[37159] = 8'b0;
    XRAM[37160] = 8'b0;
    XRAM[37161] = 8'b0;
    XRAM[37162] = 8'b0;
    XRAM[37163] = 8'b0;
    XRAM[37164] = 8'b0;
    XRAM[37165] = 8'b0;
    XRAM[37166] = 8'b0;
    XRAM[37167] = 8'b0;
    XRAM[37168] = 8'b0;
    XRAM[37169] = 8'b0;
    XRAM[37170] = 8'b0;
    XRAM[37171] = 8'b0;
    XRAM[37172] = 8'b0;
    XRAM[37173] = 8'b0;
    XRAM[37174] = 8'b0;
    XRAM[37175] = 8'b0;
    XRAM[37176] = 8'b0;
    XRAM[37177] = 8'b0;
    XRAM[37178] = 8'b0;
    XRAM[37179] = 8'b0;
    XRAM[37180] = 8'b0;
    XRAM[37181] = 8'b0;
    XRAM[37182] = 8'b0;
    XRAM[37183] = 8'b0;
    XRAM[37184] = 8'b0;
    XRAM[37185] = 8'b0;
    XRAM[37186] = 8'b0;
    XRAM[37187] = 8'b0;
    XRAM[37188] = 8'b0;
    XRAM[37189] = 8'b0;
    XRAM[37190] = 8'b0;
    XRAM[37191] = 8'b0;
    XRAM[37192] = 8'b0;
    XRAM[37193] = 8'b0;
    XRAM[37194] = 8'b0;
    XRAM[37195] = 8'b0;
    XRAM[37196] = 8'b0;
    XRAM[37197] = 8'b0;
    XRAM[37198] = 8'b0;
    XRAM[37199] = 8'b0;
    XRAM[37200] = 8'b0;
    XRAM[37201] = 8'b0;
    XRAM[37202] = 8'b0;
    XRAM[37203] = 8'b0;
    XRAM[37204] = 8'b0;
    XRAM[37205] = 8'b0;
    XRAM[37206] = 8'b0;
    XRAM[37207] = 8'b0;
    XRAM[37208] = 8'b0;
    XRAM[37209] = 8'b0;
    XRAM[37210] = 8'b0;
    XRAM[37211] = 8'b0;
    XRAM[37212] = 8'b0;
    XRAM[37213] = 8'b0;
    XRAM[37214] = 8'b0;
    XRAM[37215] = 8'b0;
    XRAM[37216] = 8'b0;
    XRAM[37217] = 8'b0;
    XRAM[37218] = 8'b0;
    XRAM[37219] = 8'b0;
    XRAM[37220] = 8'b0;
    XRAM[37221] = 8'b0;
    XRAM[37222] = 8'b0;
    XRAM[37223] = 8'b0;
    XRAM[37224] = 8'b0;
    XRAM[37225] = 8'b0;
    XRAM[37226] = 8'b0;
    XRAM[37227] = 8'b0;
    XRAM[37228] = 8'b0;
    XRAM[37229] = 8'b0;
    XRAM[37230] = 8'b0;
    XRAM[37231] = 8'b0;
    XRAM[37232] = 8'b0;
    XRAM[37233] = 8'b0;
    XRAM[37234] = 8'b0;
    XRAM[37235] = 8'b0;
    XRAM[37236] = 8'b0;
    XRAM[37237] = 8'b0;
    XRAM[37238] = 8'b0;
    XRAM[37239] = 8'b0;
    XRAM[37240] = 8'b0;
    XRAM[37241] = 8'b0;
    XRAM[37242] = 8'b0;
    XRAM[37243] = 8'b0;
    XRAM[37244] = 8'b0;
    XRAM[37245] = 8'b0;
    XRAM[37246] = 8'b0;
    XRAM[37247] = 8'b0;
    XRAM[37248] = 8'b0;
    XRAM[37249] = 8'b0;
    XRAM[37250] = 8'b0;
    XRAM[37251] = 8'b0;
    XRAM[37252] = 8'b0;
    XRAM[37253] = 8'b0;
    XRAM[37254] = 8'b0;
    XRAM[37255] = 8'b0;
    XRAM[37256] = 8'b0;
    XRAM[37257] = 8'b0;
    XRAM[37258] = 8'b0;
    XRAM[37259] = 8'b0;
    XRAM[37260] = 8'b0;
    XRAM[37261] = 8'b0;
    XRAM[37262] = 8'b0;
    XRAM[37263] = 8'b0;
    XRAM[37264] = 8'b0;
    XRAM[37265] = 8'b0;
    XRAM[37266] = 8'b0;
    XRAM[37267] = 8'b0;
    XRAM[37268] = 8'b0;
    XRAM[37269] = 8'b0;
    XRAM[37270] = 8'b0;
    XRAM[37271] = 8'b0;
    XRAM[37272] = 8'b0;
    XRAM[37273] = 8'b0;
    XRAM[37274] = 8'b0;
    XRAM[37275] = 8'b0;
    XRAM[37276] = 8'b0;
    XRAM[37277] = 8'b0;
    XRAM[37278] = 8'b0;
    XRAM[37279] = 8'b0;
    XRAM[37280] = 8'b0;
    XRAM[37281] = 8'b0;
    XRAM[37282] = 8'b0;
    XRAM[37283] = 8'b0;
    XRAM[37284] = 8'b0;
    XRAM[37285] = 8'b0;
    XRAM[37286] = 8'b0;
    XRAM[37287] = 8'b0;
    XRAM[37288] = 8'b0;
    XRAM[37289] = 8'b0;
    XRAM[37290] = 8'b0;
    XRAM[37291] = 8'b0;
    XRAM[37292] = 8'b0;
    XRAM[37293] = 8'b0;
    XRAM[37294] = 8'b0;
    XRAM[37295] = 8'b0;
    XRAM[37296] = 8'b0;
    XRAM[37297] = 8'b0;
    XRAM[37298] = 8'b0;
    XRAM[37299] = 8'b0;
    XRAM[37300] = 8'b0;
    XRAM[37301] = 8'b0;
    XRAM[37302] = 8'b0;
    XRAM[37303] = 8'b0;
    XRAM[37304] = 8'b0;
    XRAM[37305] = 8'b0;
    XRAM[37306] = 8'b0;
    XRAM[37307] = 8'b0;
    XRAM[37308] = 8'b0;
    XRAM[37309] = 8'b0;
    XRAM[37310] = 8'b0;
    XRAM[37311] = 8'b0;
    XRAM[37312] = 8'b0;
    XRAM[37313] = 8'b0;
    XRAM[37314] = 8'b0;
    XRAM[37315] = 8'b0;
    XRAM[37316] = 8'b0;
    XRAM[37317] = 8'b0;
    XRAM[37318] = 8'b0;
    XRAM[37319] = 8'b0;
    XRAM[37320] = 8'b0;
    XRAM[37321] = 8'b0;
    XRAM[37322] = 8'b0;
    XRAM[37323] = 8'b0;
    XRAM[37324] = 8'b0;
    XRAM[37325] = 8'b0;
    XRAM[37326] = 8'b0;
    XRAM[37327] = 8'b0;
    XRAM[37328] = 8'b0;
    XRAM[37329] = 8'b0;
    XRAM[37330] = 8'b0;
    XRAM[37331] = 8'b0;
    XRAM[37332] = 8'b0;
    XRAM[37333] = 8'b0;
    XRAM[37334] = 8'b0;
    XRAM[37335] = 8'b0;
    XRAM[37336] = 8'b0;
    XRAM[37337] = 8'b0;
    XRAM[37338] = 8'b0;
    XRAM[37339] = 8'b0;
    XRAM[37340] = 8'b0;
    XRAM[37341] = 8'b0;
    XRAM[37342] = 8'b0;
    XRAM[37343] = 8'b0;
    XRAM[37344] = 8'b0;
    XRAM[37345] = 8'b0;
    XRAM[37346] = 8'b0;
    XRAM[37347] = 8'b0;
    XRAM[37348] = 8'b0;
    XRAM[37349] = 8'b0;
    XRAM[37350] = 8'b0;
    XRAM[37351] = 8'b0;
    XRAM[37352] = 8'b0;
    XRAM[37353] = 8'b0;
    XRAM[37354] = 8'b0;
    XRAM[37355] = 8'b0;
    XRAM[37356] = 8'b0;
    XRAM[37357] = 8'b0;
    XRAM[37358] = 8'b0;
    XRAM[37359] = 8'b0;
    XRAM[37360] = 8'b0;
    XRAM[37361] = 8'b0;
    XRAM[37362] = 8'b0;
    XRAM[37363] = 8'b0;
    XRAM[37364] = 8'b0;
    XRAM[37365] = 8'b0;
    XRAM[37366] = 8'b0;
    XRAM[37367] = 8'b0;
    XRAM[37368] = 8'b0;
    XRAM[37369] = 8'b0;
    XRAM[37370] = 8'b0;
    XRAM[37371] = 8'b0;
    XRAM[37372] = 8'b0;
    XRAM[37373] = 8'b0;
    XRAM[37374] = 8'b0;
    XRAM[37375] = 8'b0;
    XRAM[37376] = 8'b0;
    XRAM[37377] = 8'b0;
    XRAM[37378] = 8'b0;
    XRAM[37379] = 8'b0;
    XRAM[37380] = 8'b0;
    XRAM[37381] = 8'b0;
    XRAM[37382] = 8'b0;
    XRAM[37383] = 8'b0;
    XRAM[37384] = 8'b0;
    XRAM[37385] = 8'b0;
    XRAM[37386] = 8'b0;
    XRAM[37387] = 8'b0;
    XRAM[37388] = 8'b0;
    XRAM[37389] = 8'b0;
    XRAM[37390] = 8'b0;
    XRAM[37391] = 8'b0;
    XRAM[37392] = 8'b0;
    XRAM[37393] = 8'b0;
    XRAM[37394] = 8'b0;
    XRAM[37395] = 8'b0;
    XRAM[37396] = 8'b0;
    XRAM[37397] = 8'b0;
    XRAM[37398] = 8'b0;
    XRAM[37399] = 8'b0;
    XRAM[37400] = 8'b0;
    XRAM[37401] = 8'b0;
    XRAM[37402] = 8'b0;
    XRAM[37403] = 8'b0;
    XRAM[37404] = 8'b0;
    XRAM[37405] = 8'b0;
    XRAM[37406] = 8'b0;
    XRAM[37407] = 8'b0;
    XRAM[37408] = 8'b0;
    XRAM[37409] = 8'b0;
    XRAM[37410] = 8'b0;
    XRAM[37411] = 8'b0;
    XRAM[37412] = 8'b0;
    XRAM[37413] = 8'b0;
    XRAM[37414] = 8'b0;
    XRAM[37415] = 8'b0;
    XRAM[37416] = 8'b0;
    XRAM[37417] = 8'b0;
    XRAM[37418] = 8'b0;
    XRAM[37419] = 8'b0;
    XRAM[37420] = 8'b0;
    XRAM[37421] = 8'b0;
    XRAM[37422] = 8'b0;
    XRAM[37423] = 8'b0;
    XRAM[37424] = 8'b0;
    XRAM[37425] = 8'b0;
    XRAM[37426] = 8'b0;
    XRAM[37427] = 8'b0;
    XRAM[37428] = 8'b0;
    XRAM[37429] = 8'b0;
    XRAM[37430] = 8'b0;
    XRAM[37431] = 8'b0;
    XRAM[37432] = 8'b0;
    XRAM[37433] = 8'b0;
    XRAM[37434] = 8'b0;
    XRAM[37435] = 8'b0;
    XRAM[37436] = 8'b0;
    XRAM[37437] = 8'b0;
    XRAM[37438] = 8'b0;
    XRAM[37439] = 8'b0;
    XRAM[37440] = 8'b0;
    XRAM[37441] = 8'b0;
    XRAM[37442] = 8'b0;
    XRAM[37443] = 8'b0;
    XRAM[37444] = 8'b0;
    XRAM[37445] = 8'b0;
    XRAM[37446] = 8'b0;
    XRAM[37447] = 8'b0;
    XRAM[37448] = 8'b0;
    XRAM[37449] = 8'b0;
    XRAM[37450] = 8'b0;
    XRAM[37451] = 8'b0;
    XRAM[37452] = 8'b0;
    XRAM[37453] = 8'b0;
    XRAM[37454] = 8'b0;
    XRAM[37455] = 8'b0;
    XRAM[37456] = 8'b0;
    XRAM[37457] = 8'b0;
    XRAM[37458] = 8'b0;
    XRAM[37459] = 8'b0;
    XRAM[37460] = 8'b0;
    XRAM[37461] = 8'b0;
    XRAM[37462] = 8'b0;
    XRAM[37463] = 8'b0;
    XRAM[37464] = 8'b0;
    XRAM[37465] = 8'b0;
    XRAM[37466] = 8'b0;
    XRAM[37467] = 8'b0;
    XRAM[37468] = 8'b0;
    XRAM[37469] = 8'b0;
    XRAM[37470] = 8'b0;
    XRAM[37471] = 8'b0;
    XRAM[37472] = 8'b0;
    XRAM[37473] = 8'b0;
    XRAM[37474] = 8'b0;
    XRAM[37475] = 8'b0;
    XRAM[37476] = 8'b0;
    XRAM[37477] = 8'b0;
    XRAM[37478] = 8'b0;
    XRAM[37479] = 8'b0;
    XRAM[37480] = 8'b0;
    XRAM[37481] = 8'b0;
    XRAM[37482] = 8'b0;
    XRAM[37483] = 8'b0;
    XRAM[37484] = 8'b0;
    XRAM[37485] = 8'b0;
    XRAM[37486] = 8'b0;
    XRAM[37487] = 8'b0;
    XRAM[37488] = 8'b0;
    XRAM[37489] = 8'b0;
    XRAM[37490] = 8'b0;
    XRAM[37491] = 8'b0;
    XRAM[37492] = 8'b0;
    XRAM[37493] = 8'b0;
    XRAM[37494] = 8'b0;
    XRAM[37495] = 8'b0;
    XRAM[37496] = 8'b0;
    XRAM[37497] = 8'b0;
    XRAM[37498] = 8'b0;
    XRAM[37499] = 8'b0;
    XRAM[37500] = 8'b0;
    XRAM[37501] = 8'b0;
    XRAM[37502] = 8'b0;
    XRAM[37503] = 8'b0;
    XRAM[37504] = 8'b0;
    XRAM[37505] = 8'b0;
    XRAM[37506] = 8'b0;
    XRAM[37507] = 8'b0;
    XRAM[37508] = 8'b0;
    XRAM[37509] = 8'b0;
    XRAM[37510] = 8'b0;
    XRAM[37511] = 8'b0;
    XRAM[37512] = 8'b0;
    XRAM[37513] = 8'b0;
    XRAM[37514] = 8'b0;
    XRAM[37515] = 8'b0;
    XRAM[37516] = 8'b0;
    XRAM[37517] = 8'b0;
    XRAM[37518] = 8'b0;
    XRAM[37519] = 8'b0;
    XRAM[37520] = 8'b0;
    XRAM[37521] = 8'b0;
    XRAM[37522] = 8'b0;
    XRAM[37523] = 8'b0;
    XRAM[37524] = 8'b0;
    XRAM[37525] = 8'b0;
    XRAM[37526] = 8'b0;
    XRAM[37527] = 8'b0;
    XRAM[37528] = 8'b0;
    XRAM[37529] = 8'b0;
    XRAM[37530] = 8'b0;
    XRAM[37531] = 8'b0;
    XRAM[37532] = 8'b0;
    XRAM[37533] = 8'b0;
    XRAM[37534] = 8'b0;
    XRAM[37535] = 8'b0;
    XRAM[37536] = 8'b0;
    XRAM[37537] = 8'b0;
    XRAM[37538] = 8'b0;
    XRAM[37539] = 8'b0;
    XRAM[37540] = 8'b0;
    XRAM[37541] = 8'b0;
    XRAM[37542] = 8'b0;
    XRAM[37543] = 8'b0;
    XRAM[37544] = 8'b0;
    XRAM[37545] = 8'b0;
    XRAM[37546] = 8'b0;
    XRAM[37547] = 8'b0;
    XRAM[37548] = 8'b0;
    XRAM[37549] = 8'b0;
    XRAM[37550] = 8'b0;
    XRAM[37551] = 8'b0;
    XRAM[37552] = 8'b0;
    XRAM[37553] = 8'b0;
    XRAM[37554] = 8'b0;
    XRAM[37555] = 8'b0;
    XRAM[37556] = 8'b0;
    XRAM[37557] = 8'b0;
    XRAM[37558] = 8'b0;
    XRAM[37559] = 8'b0;
    XRAM[37560] = 8'b0;
    XRAM[37561] = 8'b0;
    XRAM[37562] = 8'b0;
    XRAM[37563] = 8'b0;
    XRAM[37564] = 8'b0;
    XRAM[37565] = 8'b0;
    XRAM[37566] = 8'b0;
    XRAM[37567] = 8'b0;
    XRAM[37568] = 8'b0;
    XRAM[37569] = 8'b0;
    XRAM[37570] = 8'b0;
    XRAM[37571] = 8'b0;
    XRAM[37572] = 8'b0;
    XRAM[37573] = 8'b0;
    XRAM[37574] = 8'b0;
    XRAM[37575] = 8'b0;
    XRAM[37576] = 8'b0;
    XRAM[37577] = 8'b0;
    XRAM[37578] = 8'b0;
    XRAM[37579] = 8'b0;
    XRAM[37580] = 8'b0;
    XRAM[37581] = 8'b0;
    XRAM[37582] = 8'b0;
    XRAM[37583] = 8'b0;
    XRAM[37584] = 8'b0;
    XRAM[37585] = 8'b0;
    XRAM[37586] = 8'b0;
    XRAM[37587] = 8'b0;
    XRAM[37588] = 8'b0;
    XRAM[37589] = 8'b0;
    XRAM[37590] = 8'b0;
    XRAM[37591] = 8'b0;
    XRAM[37592] = 8'b0;
    XRAM[37593] = 8'b0;
    XRAM[37594] = 8'b0;
    XRAM[37595] = 8'b0;
    XRAM[37596] = 8'b0;
    XRAM[37597] = 8'b0;
    XRAM[37598] = 8'b0;
    XRAM[37599] = 8'b0;
    XRAM[37600] = 8'b0;
    XRAM[37601] = 8'b0;
    XRAM[37602] = 8'b0;
    XRAM[37603] = 8'b0;
    XRAM[37604] = 8'b0;
    XRAM[37605] = 8'b0;
    XRAM[37606] = 8'b0;
    XRAM[37607] = 8'b0;
    XRAM[37608] = 8'b0;
    XRAM[37609] = 8'b0;
    XRAM[37610] = 8'b0;
    XRAM[37611] = 8'b0;
    XRAM[37612] = 8'b0;
    XRAM[37613] = 8'b0;
    XRAM[37614] = 8'b0;
    XRAM[37615] = 8'b0;
    XRAM[37616] = 8'b0;
    XRAM[37617] = 8'b0;
    XRAM[37618] = 8'b0;
    XRAM[37619] = 8'b0;
    XRAM[37620] = 8'b0;
    XRAM[37621] = 8'b0;
    XRAM[37622] = 8'b0;
    XRAM[37623] = 8'b0;
    XRAM[37624] = 8'b0;
    XRAM[37625] = 8'b0;
    XRAM[37626] = 8'b0;
    XRAM[37627] = 8'b0;
    XRAM[37628] = 8'b0;
    XRAM[37629] = 8'b0;
    XRAM[37630] = 8'b0;
    XRAM[37631] = 8'b0;
    XRAM[37632] = 8'b0;
    XRAM[37633] = 8'b0;
    XRAM[37634] = 8'b0;
    XRAM[37635] = 8'b0;
    XRAM[37636] = 8'b0;
    XRAM[37637] = 8'b0;
    XRAM[37638] = 8'b0;
    XRAM[37639] = 8'b0;
    XRAM[37640] = 8'b0;
    XRAM[37641] = 8'b0;
    XRAM[37642] = 8'b0;
    XRAM[37643] = 8'b0;
    XRAM[37644] = 8'b0;
    XRAM[37645] = 8'b0;
    XRAM[37646] = 8'b0;
    XRAM[37647] = 8'b0;
    XRAM[37648] = 8'b0;
    XRAM[37649] = 8'b0;
    XRAM[37650] = 8'b0;
    XRAM[37651] = 8'b0;
    XRAM[37652] = 8'b0;
    XRAM[37653] = 8'b0;
    XRAM[37654] = 8'b0;
    XRAM[37655] = 8'b0;
    XRAM[37656] = 8'b0;
    XRAM[37657] = 8'b0;
    XRAM[37658] = 8'b0;
    XRAM[37659] = 8'b0;
    XRAM[37660] = 8'b0;
    XRAM[37661] = 8'b0;
    XRAM[37662] = 8'b0;
    XRAM[37663] = 8'b0;
    XRAM[37664] = 8'b0;
    XRAM[37665] = 8'b0;
    XRAM[37666] = 8'b0;
    XRAM[37667] = 8'b0;
    XRAM[37668] = 8'b0;
    XRAM[37669] = 8'b0;
    XRAM[37670] = 8'b0;
    XRAM[37671] = 8'b0;
    XRAM[37672] = 8'b0;
    XRAM[37673] = 8'b0;
    XRAM[37674] = 8'b0;
    XRAM[37675] = 8'b0;
    XRAM[37676] = 8'b0;
    XRAM[37677] = 8'b0;
    XRAM[37678] = 8'b0;
    XRAM[37679] = 8'b0;
    XRAM[37680] = 8'b0;
    XRAM[37681] = 8'b0;
    XRAM[37682] = 8'b0;
    XRAM[37683] = 8'b0;
    XRAM[37684] = 8'b0;
    XRAM[37685] = 8'b0;
    XRAM[37686] = 8'b0;
    XRAM[37687] = 8'b0;
    XRAM[37688] = 8'b0;
    XRAM[37689] = 8'b0;
    XRAM[37690] = 8'b0;
    XRAM[37691] = 8'b0;
    XRAM[37692] = 8'b0;
    XRAM[37693] = 8'b0;
    XRAM[37694] = 8'b0;
    XRAM[37695] = 8'b0;
    XRAM[37696] = 8'b0;
    XRAM[37697] = 8'b0;
    XRAM[37698] = 8'b0;
    XRAM[37699] = 8'b0;
    XRAM[37700] = 8'b0;
    XRAM[37701] = 8'b0;
    XRAM[37702] = 8'b0;
    XRAM[37703] = 8'b0;
    XRAM[37704] = 8'b0;
    XRAM[37705] = 8'b0;
    XRAM[37706] = 8'b0;
    XRAM[37707] = 8'b0;
    XRAM[37708] = 8'b0;
    XRAM[37709] = 8'b0;
    XRAM[37710] = 8'b0;
    XRAM[37711] = 8'b0;
    XRAM[37712] = 8'b0;
    XRAM[37713] = 8'b0;
    XRAM[37714] = 8'b0;
    XRAM[37715] = 8'b0;
    XRAM[37716] = 8'b0;
    XRAM[37717] = 8'b0;
    XRAM[37718] = 8'b0;
    XRAM[37719] = 8'b0;
    XRAM[37720] = 8'b0;
    XRAM[37721] = 8'b0;
    XRAM[37722] = 8'b0;
    XRAM[37723] = 8'b0;
    XRAM[37724] = 8'b0;
    XRAM[37725] = 8'b0;
    XRAM[37726] = 8'b0;
    XRAM[37727] = 8'b0;
    XRAM[37728] = 8'b0;
    XRAM[37729] = 8'b0;
    XRAM[37730] = 8'b0;
    XRAM[37731] = 8'b0;
    XRAM[37732] = 8'b0;
    XRAM[37733] = 8'b0;
    XRAM[37734] = 8'b0;
    XRAM[37735] = 8'b0;
    XRAM[37736] = 8'b0;
    XRAM[37737] = 8'b0;
    XRAM[37738] = 8'b0;
    XRAM[37739] = 8'b0;
    XRAM[37740] = 8'b0;
    XRAM[37741] = 8'b0;
    XRAM[37742] = 8'b0;
    XRAM[37743] = 8'b0;
    XRAM[37744] = 8'b0;
    XRAM[37745] = 8'b0;
    XRAM[37746] = 8'b0;
    XRAM[37747] = 8'b0;
    XRAM[37748] = 8'b0;
    XRAM[37749] = 8'b0;
    XRAM[37750] = 8'b0;
    XRAM[37751] = 8'b0;
    XRAM[37752] = 8'b0;
    XRAM[37753] = 8'b0;
    XRAM[37754] = 8'b0;
    XRAM[37755] = 8'b0;
    XRAM[37756] = 8'b0;
    XRAM[37757] = 8'b0;
    XRAM[37758] = 8'b0;
    XRAM[37759] = 8'b0;
    XRAM[37760] = 8'b0;
    XRAM[37761] = 8'b0;
    XRAM[37762] = 8'b0;
    XRAM[37763] = 8'b0;
    XRAM[37764] = 8'b0;
    XRAM[37765] = 8'b0;
    XRAM[37766] = 8'b0;
    XRAM[37767] = 8'b0;
    XRAM[37768] = 8'b0;
    XRAM[37769] = 8'b0;
    XRAM[37770] = 8'b0;
    XRAM[37771] = 8'b0;
    XRAM[37772] = 8'b0;
    XRAM[37773] = 8'b0;
    XRAM[37774] = 8'b0;
    XRAM[37775] = 8'b0;
    XRAM[37776] = 8'b0;
    XRAM[37777] = 8'b0;
    XRAM[37778] = 8'b0;
    XRAM[37779] = 8'b0;
    XRAM[37780] = 8'b0;
    XRAM[37781] = 8'b0;
    XRAM[37782] = 8'b0;
    XRAM[37783] = 8'b0;
    XRAM[37784] = 8'b0;
    XRAM[37785] = 8'b0;
    XRAM[37786] = 8'b0;
    XRAM[37787] = 8'b0;
    XRAM[37788] = 8'b0;
    XRAM[37789] = 8'b0;
    XRAM[37790] = 8'b0;
    XRAM[37791] = 8'b0;
    XRAM[37792] = 8'b0;
    XRAM[37793] = 8'b0;
    XRAM[37794] = 8'b0;
    XRAM[37795] = 8'b0;
    XRAM[37796] = 8'b0;
    XRAM[37797] = 8'b0;
    XRAM[37798] = 8'b0;
    XRAM[37799] = 8'b0;
    XRAM[37800] = 8'b0;
    XRAM[37801] = 8'b0;
    XRAM[37802] = 8'b0;
    XRAM[37803] = 8'b0;
    XRAM[37804] = 8'b0;
    XRAM[37805] = 8'b0;
    XRAM[37806] = 8'b0;
    XRAM[37807] = 8'b0;
    XRAM[37808] = 8'b0;
    XRAM[37809] = 8'b0;
    XRAM[37810] = 8'b0;
    XRAM[37811] = 8'b0;
    XRAM[37812] = 8'b0;
    XRAM[37813] = 8'b0;
    XRAM[37814] = 8'b0;
    XRAM[37815] = 8'b0;
    XRAM[37816] = 8'b0;
    XRAM[37817] = 8'b0;
    XRAM[37818] = 8'b0;
    XRAM[37819] = 8'b0;
    XRAM[37820] = 8'b0;
    XRAM[37821] = 8'b0;
    XRAM[37822] = 8'b0;
    XRAM[37823] = 8'b0;
    XRAM[37824] = 8'b0;
    XRAM[37825] = 8'b0;
    XRAM[37826] = 8'b0;
    XRAM[37827] = 8'b0;
    XRAM[37828] = 8'b0;
    XRAM[37829] = 8'b0;
    XRAM[37830] = 8'b0;
    XRAM[37831] = 8'b0;
    XRAM[37832] = 8'b0;
    XRAM[37833] = 8'b0;
    XRAM[37834] = 8'b0;
    XRAM[37835] = 8'b0;
    XRAM[37836] = 8'b0;
    XRAM[37837] = 8'b0;
    XRAM[37838] = 8'b0;
    XRAM[37839] = 8'b0;
    XRAM[37840] = 8'b0;
    XRAM[37841] = 8'b0;
    XRAM[37842] = 8'b0;
    XRAM[37843] = 8'b0;
    XRAM[37844] = 8'b0;
    XRAM[37845] = 8'b0;
    XRAM[37846] = 8'b0;
    XRAM[37847] = 8'b0;
    XRAM[37848] = 8'b0;
    XRAM[37849] = 8'b0;
    XRAM[37850] = 8'b0;
    XRAM[37851] = 8'b0;
    XRAM[37852] = 8'b0;
    XRAM[37853] = 8'b0;
    XRAM[37854] = 8'b0;
    XRAM[37855] = 8'b0;
    XRAM[37856] = 8'b0;
    XRAM[37857] = 8'b0;
    XRAM[37858] = 8'b0;
    XRAM[37859] = 8'b0;
    XRAM[37860] = 8'b0;
    XRAM[37861] = 8'b0;
    XRAM[37862] = 8'b0;
    XRAM[37863] = 8'b0;
    XRAM[37864] = 8'b0;
    XRAM[37865] = 8'b0;
    XRAM[37866] = 8'b0;
    XRAM[37867] = 8'b0;
    XRAM[37868] = 8'b0;
    XRAM[37869] = 8'b0;
    XRAM[37870] = 8'b0;
    XRAM[37871] = 8'b0;
    XRAM[37872] = 8'b0;
    XRAM[37873] = 8'b0;
    XRAM[37874] = 8'b0;
    XRAM[37875] = 8'b0;
    XRAM[37876] = 8'b0;
    XRAM[37877] = 8'b0;
    XRAM[37878] = 8'b0;
    XRAM[37879] = 8'b0;
    XRAM[37880] = 8'b0;
    XRAM[37881] = 8'b0;
    XRAM[37882] = 8'b0;
    XRAM[37883] = 8'b0;
    XRAM[37884] = 8'b0;
    XRAM[37885] = 8'b0;
    XRAM[37886] = 8'b0;
    XRAM[37887] = 8'b0;
    XRAM[37888] = 8'b0;
    XRAM[37889] = 8'b0;
    XRAM[37890] = 8'b0;
    XRAM[37891] = 8'b0;
    XRAM[37892] = 8'b0;
    XRAM[37893] = 8'b0;
    XRAM[37894] = 8'b0;
    XRAM[37895] = 8'b0;
    XRAM[37896] = 8'b0;
    XRAM[37897] = 8'b0;
    XRAM[37898] = 8'b0;
    XRAM[37899] = 8'b0;
    XRAM[37900] = 8'b0;
    XRAM[37901] = 8'b0;
    XRAM[37902] = 8'b0;
    XRAM[37903] = 8'b0;
    XRAM[37904] = 8'b0;
    XRAM[37905] = 8'b0;
    XRAM[37906] = 8'b0;
    XRAM[37907] = 8'b0;
    XRAM[37908] = 8'b0;
    XRAM[37909] = 8'b0;
    XRAM[37910] = 8'b0;
    XRAM[37911] = 8'b0;
    XRAM[37912] = 8'b0;
    XRAM[37913] = 8'b0;
    XRAM[37914] = 8'b0;
    XRAM[37915] = 8'b0;
    XRAM[37916] = 8'b0;
    XRAM[37917] = 8'b0;
    XRAM[37918] = 8'b0;
    XRAM[37919] = 8'b0;
    XRAM[37920] = 8'b0;
    XRAM[37921] = 8'b0;
    XRAM[37922] = 8'b0;
    XRAM[37923] = 8'b0;
    XRAM[37924] = 8'b0;
    XRAM[37925] = 8'b0;
    XRAM[37926] = 8'b0;
    XRAM[37927] = 8'b0;
    XRAM[37928] = 8'b0;
    XRAM[37929] = 8'b0;
    XRAM[37930] = 8'b0;
    XRAM[37931] = 8'b0;
    XRAM[37932] = 8'b0;
    XRAM[37933] = 8'b0;
    XRAM[37934] = 8'b0;
    XRAM[37935] = 8'b0;
    XRAM[37936] = 8'b0;
    XRAM[37937] = 8'b0;
    XRAM[37938] = 8'b0;
    XRAM[37939] = 8'b0;
    XRAM[37940] = 8'b0;
    XRAM[37941] = 8'b0;
    XRAM[37942] = 8'b0;
    XRAM[37943] = 8'b0;
    XRAM[37944] = 8'b0;
    XRAM[37945] = 8'b0;
    XRAM[37946] = 8'b0;
    XRAM[37947] = 8'b0;
    XRAM[37948] = 8'b0;
    XRAM[37949] = 8'b0;
    XRAM[37950] = 8'b0;
    XRAM[37951] = 8'b0;
    XRAM[37952] = 8'b0;
    XRAM[37953] = 8'b0;
    XRAM[37954] = 8'b0;
    XRAM[37955] = 8'b0;
    XRAM[37956] = 8'b0;
    XRAM[37957] = 8'b0;
    XRAM[37958] = 8'b0;
    XRAM[37959] = 8'b0;
    XRAM[37960] = 8'b0;
    XRAM[37961] = 8'b0;
    XRAM[37962] = 8'b0;
    XRAM[37963] = 8'b0;
    XRAM[37964] = 8'b0;
    XRAM[37965] = 8'b0;
    XRAM[37966] = 8'b0;
    XRAM[37967] = 8'b0;
    XRAM[37968] = 8'b0;
    XRAM[37969] = 8'b0;
    XRAM[37970] = 8'b0;
    XRAM[37971] = 8'b0;
    XRAM[37972] = 8'b0;
    XRAM[37973] = 8'b0;
    XRAM[37974] = 8'b0;
    XRAM[37975] = 8'b0;
    XRAM[37976] = 8'b0;
    XRAM[37977] = 8'b0;
    XRAM[37978] = 8'b0;
    XRAM[37979] = 8'b0;
    XRAM[37980] = 8'b0;
    XRAM[37981] = 8'b0;
    XRAM[37982] = 8'b0;
    XRAM[37983] = 8'b0;
    XRAM[37984] = 8'b0;
    XRAM[37985] = 8'b0;
    XRAM[37986] = 8'b0;
    XRAM[37987] = 8'b0;
    XRAM[37988] = 8'b0;
    XRAM[37989] = 8'b0;
    XRAM[37990] = 8'b0;
    XRAM[37991] = 8'b0;
    XRAM[37992] = 8'b0;
    XRAM[37993] = 8'b0;
    XRAM[37994] = 8'b0;
    XRAM[37995] = 8'b0;
    XRAM[37996] = 8'b0;
    XRAM[37997] = 8'b0;
    XRAM[37998] = 8'b0;
    XRAM[37999] = 8'b0;
    XRAM[38000] = 8'b0;
    XRAM[38001] = 8'b0;
    XRAM[38002] = 8'b0;
    XRAM[38003] = 8'b0;
    XRAM[38004] = 8'b0;
    XRAM[38005] = 8'b0;
    XRAM[38006] = 8'b0;
    XRAM[38007] = 8'b0;
    XRAM[38008] = 8'b0;
    XRAM[38009] = 8'b0;
    XRAM[38010] = 8'b0;
    XRAM[38011] = 8'b0;
    XRAM[38012] = 8'b0;
    XRAM[38013] = 8'b0;
    XRAM[38014] = 8'b0;
    XRAM[38015] = 8'b0;
    XRAM[38016] = 8'b0;
    XRAM[38017] = 8'b0;
    XRAM[38018] = 8'b0;
    XRAM[38019] = 8'b0;
    XRAM[38020] = 8'b0;
    XRAM[38021] = 8'b0;
    XRAM[38022] = 8'b0;
    XRAM[38023] = 8'b0;
    XRAM[38024] = 8'b0;
    XRAM[38025] = 8'b0;
    XRAM[38026] = 8'b0;
    XRAM[38027] = 8'b0;
    XRAM[38028] = 8'b0;
    XRAM[38029] = 8'b0;
    XRAM[38030] = 8'b0;
    XRAM[38031] = 8'b0;
    XRAM[38032] = 8'b0;
    XRAM[38033] = 8'b0;
    XRAM[38034] = 8'b0;
    XRAM[38035] = 8'b0;
    XRAM[38036] = 8'b0;
    XRAM[38037] = 8'b0;
    XRAM[38038] = 8'b0;
    XRAM[38039] = 8'b0;
    XRAM[38040] = 8'b0;
    XRAM[38041] = 8'b0;
    XRAM[38042] = 8'b0;
    XRAM[38043] = 8'b0;
    XRAM[38044] = 8'b0;
    XRAM[38045] = 8'b0;
    XRAM[38046] = 8'b0;
    XRAM[38047] = 8'b0;
    XRAM[38048] = 8'b0;
    XRAM[38049] = 8'b0;
    XRAM[38050] = 8'b0;
    XRAM[38051] = 8'b0;
    XRAM[38052] = 8'b0;
    XRAM[38053] = 8'b0;
    XRAM[38054] = 8'b0;
    XRAM[38055] = 8'b0;
    XRAM[38056] = 8'b0;
    XRAM[38057] = 8'b0;
    XRAM[38058] = 8'b0;
    XRAM[38059] = 8'b0;
    XRAM[38060] = 8'b0;
    XRAM[38061] = 8'b0;
    XRAM[38062] = 8'b0;
    XRAM[38063] = 8'b0;
    XRAM[38064] = 8'b0;
    XRAM[38065] = 8'b0;
    XRAM[38066] = 8'b0;
    XRAM[38067] = 8'b0;
    XRAM[38068] = 8'b0;
    XRAM[38069] = 8'b0;
    XRAM[38070] = 8'b0;
    XRAM[38071] = 8'b0;
    XRAM[38072] = 8'b0;
    XRAM[38073] = 8'b0;
    XRAM[38074] = 8'b0;
    XRAM[38075] = 8'b0;
    XRAM[38076] = 8'b0;
    XRAM[38077] = 8'b0;
    XRAM[38078] = 8'b0;
    XRAM[38079] = 8'b0;
    XRAM[38080] = 8'b0;
    XRAM[38081] = 8'b0;
    XRAM[38082] = 8'b0;
    XRAM[38083] = 8'b0;
    XRAM[38084] = 8'b0;
    XRAM[38085] = 8'b0;
    XRAM[38086] = 8'b0;
    XRAM[38087] = 8'b0;
    XRAM[38088] = 8'b0;
    XRAM[38089] = 8'b0;
    XRAM[38090] = 8'b0;
    XRAM[38091] = 8'b0;
    XRAM[38092] = 8'b0;
    XRAM[38093] = 8'b0;
    XRAM[38094] = 8'b0;
    XRAM[38095] = 8'b0;
    XRAM[38096] = 8'b0;
    XRAM[38097] = 8'b0;
    XRAM[38098] = 8'b0;
    XRAM[38099] = 8'b0;
    XRAM[38100] = 8'b0;
    XRAM[38101] = 8'b0;
    XRAM[38102] = 8'b0;
    XRAM[38103] = 8'b0;
    XRAM[38104] = 8'b0;
    XRAM[38105] = 8'b0;
    XRAM[38106] = 8'b0;
    XRAM[38107] = 8'b0;
    XRAM[38108] = 8'b0;
    XRAM[38109] = 8'b0;
    XRAM[38110] = 8'b0;
    XRAM[38111] = 8'b0;
    XRAM[38112] = 8'b0;
    XRAM[38113] = 8'b0;
    XRAM[38114] = 8'b0;
    XRAM[38115] = 8'b0;
    XRAM[38116] = 8'b0;
    XRAM[38117] = 8'b0;
    XRAM[38118] = 8'b0;
    XRAM[38119] = 8'b0;
    XRAM[38120] = 8'b0;
    XRAM[38121] = 8'b0;
    XRAM[38122] = 8'b0;
    XRAM[38123] = 8'b0;
    XRAM[38124] = 8'b0;
    XRAM[38125] = 8'b0;
    XRAM[38126] = 8'b0;
    XRAM[38127] = 8'b0;
    XRAM[38128] = 8'b0;
    XRAM[38129] = 8'b0;
    XRAM[38130] = 8'b0;
    XRAM[38131] = 8'b0;
    XRAM[38132] = 8'b0;
    XRAM[38133] = 8'b0;
    XRAM[38134] = 8'b0;
    XRAM[38135] = 8'b0;
    XRAM[38136] = 8'b0;
    XRAM[38137] = 8'b0;
    XRAM[38138] = 8'b0;
    XRAM[38139] = 8'b0;
    XRAM[38140] = 8'b0;
    XRAM[38141] = 8'b0;
    XRAM[38142] = 8'b0;
    XRAM[38143] = 8'b0;
    XRAM[38144] = 8'b0;
    XRAM[38145] = 8'b0;
    XRAM[38146] = 8'b0;
    XRAM[38147] = 8'b0;
    XRAM[38148] = 8'b0;
    XRAM[38149] = 8'b0;
    XRAM[38150] = 8'b0;
    XRAM[38151] = 8'b0;
    XRAM[38152] = 8'b0;
    XRAM[38153] = 8'b0;
    XRAM[38154] = 8'b0;
    XRAM[38155] = 8'b0;
    XRAM[38156] = 8'b0;
    XRAM[38157] = 8'b0;
    XRAM[38158] = 8'b0;
    XRAM[38159] = 8'b0;
    XRAM[38160] = 8'b0;
    XRAM[38161] = 8'b0;
    XRAM[38162] = 8'b0;
    XRAM[38163] = 8'b0;
    XRAM[38164] = 8'b0;
    XRAM[38165] = 8'b0;
    XRAM[38166] = 8'b0;
    XRAM[38167] = 8'b0;
    XRAM[38168] = 8'b0;
    XRAM[38169] = 8'b0;
    XRAM[38170] = 8'b0;
    XRAM[38171] = 8'b0;
    XRAM[38172] = 8'b0;
    XRAM[38173] = 8'b0;
    XRAM[38174] = 8'b0;
    XRAM[38175] = 8'b0;
    XRAM[38176] = 8'b0;
    XRAM[38177] = 8'b0;
    XRAM[38178] = 8'b0;
    XRAM[38179] = 8'b0;
    XRAM[38180] = 8'b0;
    XRAM[38181] = 8'b0;
    XRAM[38182] = 8'b0;
    XRAM[38183] = 8'b0;
    XRAM[38184] = 8'b0;
    XRAM[38185] = 8'b0;
    XRAM[38186] = 8'b0;
    XRAM[38187] = 8'b0;
    XRAM[38188] = 8'b0;
    XRAM[38189] = 8'b0;
    XRAM[38190] = 8'b0;
    XRAM[38191] = 8'b0;
    XRAM[38192] = 8'b0;
    XRAM[38193] = 8'b0;
    XRAM[38194] = 8'b0;
    XRAM[38195] = 8'b0;
    XRAM[38196] = 8'b0;
    XRAM[38197] = 8'b0;
    XRAM[38198] = 8'b0;
    XRAM[38199] = 8'b0;
    XRAM[38200] = 8'b0;
    XRAM[38201] = 8'b0;
    XRAM[38202] = 8'b0;
    XRAM[38203] = 8'b0;
    XRAM[38204] = 8'b0;
    XRAM[38205] = 8'b0;
    XRAM[38206] = 8'b0;
    XRAM[38207] = 8'b0;
    XRAM[38208] = 8'b0;
    XRAM[38209] = 8'b0;
    XRAM[38210] = 8'b0;
    XRAM[38211] = 8'b0;
    XRAM[38212] = 8'b0;
    XRAM[38213] = 8'b0;
    XRAM[38214] = 8'b0;
    XRAM[38215] = 8'b0;
    XRAM[38216] = 8'b0;
    XRAM[38217] = 8'b0;
    XRAM[38218] = 8'b0;
    XRAM[38219] = 8'b0;
    XRAM[38220] = 8'b0;
    XRAM[38221] = 8'b0;
    XRAM[38222] = 8'b0;
    XRAM[38223] = 8'b0;
    XRAM[38224] = 8'b0;
    XRAM[38225] = 8'b0;
    XRAM[38226] = 8'b0;
    XRAM[38227] = 8'b0;
    XRAM[38228] = 8'b0;
    XRAM[38229] = 8'b0;
    XRAM[38230] = 8'b0;
    XRAM[38231] = 8'b0;
    XRAM[38232] = 8'b0;
    XRAM[38233] = 8'b0;
    XRAM[38234] = 8'b0;
    XRAM[38235] = 8'b0;
    XRAM[38236] = 8'b0;
    XRAM[38237] = 8'b0;
    XRAM[38238] = 8'b0;
    XRAM[38239] = 8'b0;
    XRAM[38240] = 8'b0;
    XRAM[38241] = 8'b0;
    XRAM[38242] = 8'b0;
    XRAM[38243] = 8'b0;
    XRAM[38244] = 8'b0;
    XRAM[38245] = 8'b0;
    XRAM[38246] = 8'b0;
    XRAM[38247] = 8'b0;
    XRAM[38248] = 8'b0;
    XRAM[38249] = 8'b0;
    XRAM[38250] = 8'b0;
    XRAM[38251] = 8'b0;
    XRAM[38252] = 8'b0;
    XRAM[38253] = 8'b0;
    XRAM[38254] = 8'b0;
    XRAM[38255] = 8'b0;
    XRAM[38256] = 8'b0;
    XRAM[38257] = 8'b0;
    XRAM[38258] = 8'b0;
    XRAM[38259] = 8'b0;
    XRAM[38260] = 8'b0;
    XRAM[38261] = 8'b0;
    XRAM[38262] = 8'b0;
    XRAM[38263] = 8'b0;
    XRAM[38264] = 8'b0;
    XRAM[38265] = 8'b0;
    XRAM[38266] = 8'b0;
    XRAM[38267] = 8'b0;
    XRAM[38268] = 8'b0;
    XRAM[38269] = 8'b0;
    XRAM[38270] = 8'b0;
    XRAM[38271] = 8'b0;
    XRAM[38272] = 8'b0;
    XRAM[38273] = 8'b0;
    XRAM[38274] = 8'b0;
    XRAM[38275] = 8'b0;
    XRAM[38276] = 8'b0;
    XRAM[38277] = 8'b0;
    XRAM[38278] = 8'b0;
    XRAM[38279] = 8'b0;
    XRAM[38280] = 8'b0;
    XRAM[38281] = 8'b0;
    XRAM[38282] = 8'b0;
    XRAM[38283] = 8'b0;
    XRAM[38284] = 8'b0;
    XRAM[38285] = 8'b0;
    XRAM[38286] = 8'b0;
    XRAM[38287] = 8'b0;
    XRAM[38288] = 8'b0;
    XRAM[38289] = 8'b0;
    XRAM[38290] = 8'b0;
    XRAM[38291] = 8'b0;
    XRAM[38292] = 8'b0;
    XRAM[38293] = 8'b0;
    XRAM[38294] = 8'b0;
    XRAM[38295] = 8'b0;
    XRAM[38296] = 8'b0;
    XRAM[38297] = 8'b0;
    XRAM[38298] = 8'b0;
    XRAM[38299] = 8'b0;
    XRAM[38300] = 8'b0;
    XRAM[38301] = 8'b0;
    XRAM[38302] = 8'b0;
    XRAM[38303] = 8'b0;
    XRAM[38304] = 8'b0;
    XRAM[38305] = 8'b0;
    XRAM[38306] = 8'b0;
    XRAM[38307] = 8'b0;
    XRAM[38308] = 8'b0;
    XRAM[38309] = 8'b0;
    XRAM[38310] = 8'b0;
    XRAM[38311] = 8'b0;
    XRAM[38312] = 8'b0;
    XRAM[38313] = 8'b0;
    XRAM[38314] = 8'b0;
    XRAM[38315] = 8'b0;
    XRAM[38316] = 8'b0;
    XRAM[38317] = 8'b0;
    XRAM[38318] = 8'b0;
    XRAM[38319] = 8'b0;
    XRAM[38320] = 8'b0;
    XRAM[38321] = 8'b0;
    XRAM[38322] = 8'b0;
    XRAM[38323] = 8'b0;
    XRAM[38324] = 8'b0;
    XRAM[38325] = 8'b0;
    XRAM[38326] = 8'b0;
    XRAM[38327] = 8'b0;
    XRAM[38328] = 8'b0;
    XRAM[38329] = 8'b0;
    XRAM[38330] = 8'b0;
    XRAM[38331] = 8'b0;
    XRAM[38332] = 8'b0;
    XRAM[38333] = 8'b0;
    XRAM[38334] = 8'b0;
    XRAM[38335] = 8'b0;
    XRAM[38336] = 8'b0;
    XRAM[38337] = 8'b0;
    XRAM[38338] = 8'b0;
    XRAM[38339] = 8'b0;
    XRAM[38340] = 8'b0;
    XRAM[38341] = 8'b0;
    XRAM[38342] = 8'b0;
    XRAM[38343] = 8'b0;
    XRAM[38344] = 8'b0;
    XRAM[38345] = 8'b0;
    XRAM[38346] = 8'b0;
    XRAM[38347] = 8'b0;
    XRAM[38348] = 8'b0;
    XRAM[38349] = 8'b0;
    XRAM[38350] = 8'b0;
    XRAM[38351] = 8'b0;
    XRAM[38352] = 8'b0;
    XRAM[38353] = 8'b0;
    XRAM[38354] = 8'b0;
    XRAM[38355] = 8'b0;
    XRAM[38356] = 8'b0;
    XRAM[38357] = 8'b0;
    XRAM[38358] = 8'b0;
    XRAM[38359] = 8'b0;
    XRAM[38360] = 8'b0;
    XRAM[38361] = 8'b0;
    XRAM[38362] = 8'b0;
    XRAM[38363] = 8'b0;
    XRAM[38364] = 8'b0;
    XRAM[38365] = 8'b0;
    XRAM[38366] = 8'b0;
    XRAM[38367] = 8'b0;
    XRAM[38368] = 8'b0;
    XRAM[38369] = 8'b0;
    XRAM[38370] = 8'b0;
    XRAM[38371] = 8'b0;
    XRAM[38372] = 8'b0;
    XRAM[38373] = 8'b0;
    XRAM[38374] = 8'b0;
    XRAM[38375] = 8'b0;
    XRAM[38376] = 8'b0;
    XRAM[38377] = 8'b0;
    XRAM[38378] = 8'b0;
    XRAM[38379] = 8'b0;
    XRAM[38380] = 8'b0;
    XRAM[38381] = 8'b0;
    XRAM[38382] = 8'b0;
    XRAM[38383] = 8'b0;
    XRAM[38384] = 8'b0;
    XRAM[38385] = 8'b0;
    XRAM[38386] = 8'b0;
    XRAM[38387] = 8'b0;
    XRAM[38388] = 8'b0;
    XRAM[38389] = 8'b0;
    XRAM[38390] = 8'b0;
    XRAM[38391] = 8'b0;
    XRAM[38392] = 8'b0;
    XRAM[38393] = 8'b0;
    XRAM[38394] = 8'b0;
    XRAM[38395] = 8'b0;
    XRAM[38396] = 8'b0;
    XRAM[38397] = 8'b0;
    XRAM[38398] = 8'b0;
    XRAM[38399] = 8'b0;
    XRAM[38400] = 8'b0;
    XRAM[38401] = 8'b0;
    XRAM[38402] = 8'b0;
    XRAM[38403] = 8'b0;
    XRAM[38404] = 8'b0;
    XRAM[38405] = 8'b0;
    XRAM[38406] = 8'b0;
    XRAM[38407] = 8'b0;
    XRAM[38408] = 8'b0;
    XRAM[38409] = 8'b0;
    XRAM[38410] = 8'b0;
    XRAM[38411] = 8'b0;
    XRAM[38412] = 8'b0;
    XRAM[38413] = 8'b0;
    XRAM[38414] = 8'b0;
    XRAM[38415] = 8'b0;
    XRAM[38416] = 8'b0;
    XRAM[38417] = 8'b0;
    XRAM[38418] = 8'b0;
    XRAM[38419] = 8'b0;
    XRAM[38420] = 8'b0;
    XRAM[38421] = 8'b0;
    XRAM[38422] = 8'b0;
    XRAM[38423] = 8'b0;
    XRAM[38424] = 8'b0;
    XRAM[38425] = 8'b0;
    XRAM[38426] = 8'b0;
    XRAM[38427] = 8'b0;
    XRAM[38428] = 8'b0;
    XRAM[38429] = 8'b0;
    XRAM[38430] = 8'b0;
    XRAM[38431] = 8'b0;
    XRAM[38432] = 8'b0;
    XRAM[38433] = 8'b0;
    XRAM[38434] = 8'b0;
    XRAM[38435] = 8'b0;
    XRAM[38436] = 8'b0;
    XRAM[38437] = 8'b0;
    XRAM[38438] = 8'b0;
    XRAM[38439] = 8'b0;
    XRAM[38440] = 8'b0;
    XRAM[38441] = 8'b0;
    XRAM[38442] = 8'b0;
    XRAM[38443] = 8'b0;
    XRAM[38444] = 8'b0;
    XRAM[38445] = 8'b0;
    XRAM[38446] = 8'b0;
    XRAM[38447] = 8'b0;
    XRAM[38448] = 8'b0;
    XRAM[38449] = 8'b0;
    XRAM[38450] = 8'b0;
    XRAM[38451] = 8'b0;
    XRAM[38452] = 8'b0;
    XRAM[38453] = 8'b0;
    XRAM[38454] = 8'b0;
    XRAM[38455] = 8'b0;
    XRAM[38456] = 8'b0;
    XRAM[38457] = 8'b0;
    XRAM[38458] = 8'b0;
    XRAM[38459] = 8'b0;
    XRAM[38460] = 8'b0;
    XRAM[38461] = 8'b0;
    XRAM[38462] = 8'b0;
    XRAM[38463] = 8'b0;
    XRAM[38464] = 8'b0;
    XRAM[38465] = 8'b0;
    XRAM[38466] = 8'b0;
    XRAM[38467] = 8'b0;
    XRAM[38468] = 8'b0;
    XRAM[38469] = 8'b0;
    XRAM[38470] = 8'b0;
    XRAM[38471] = 8'b0;
    XRAM[38472] = 8'b0;
    XRAM[38473] = 8'b0;
    XRAM[38474] = 8'b0;
    XRAM[38475] = 8'b0;
    XRAM[38476] = 8'b0;
    XRAM[38477] = 8'b0;
    XRAM[38478] = 8'b0;
    XRAM[38479] = 8'b0;
    XRAM[38480] = 8'b0;
    XRAM[38481] = 8'b0;
    XRAM[38482] = 8'b0;
    XRAM[38483] = 8'b0;
    XRAM[38484] = 8'b0;
    XRAM[38485] = 8'b0;
    XRAM[38486] = 8'b0;
    XRAM[38487] = 8'b0;
    XRAM[38488] = 8'b0;
    XRAM[38489] = 8'b0;
    XRAM[38490] = 8'b0;
    XRAM[38491] = 8'b0;
    XRAM[38492] = 8'b0;
    XRAM[38493] = 8'b0;
    XRAM[38494] = 8'b0;
    XRAM[38495] = 8'b0;
    XRAM[38496] = 8'b0;
    XRAM[38497] = 8'b0;
    XRAM[38498] = 8'b0;
    XRAM[38499] = 8'b0;
    XRAM[38500] = 8'b0;
    XRAM[38501] = 8'b0;
    XRAM[38502] = 8'b0;
    XRAM[38503] = 8'b0;
    XRAM[38504] = 8'b0;
    XRAM[38505] = 8'b0;
    XRAM[38506] = 8'b0;
    XRAM[38507] = 8'b0;
    XRAM[38508] = 8'b0;
    XRAM[38509] = 8'b0;
    XRAM[38510] = 8'b0;
    XRAM[38511] = 8'b0;
    XRAM[38512] = 8'b0;
    XRAM[38513] = 8'b0;
    XRAM[38514] = 8'b0;
    XRAM[38515] = 8'b0;
    XRAM[38516] = 8'b0;
    XRAM[38517] = 8'b0;
    XRAM[38518] = 8'b0;
    XRAM[38519] = 8'b0;
    XRAM[38520] = 8'b0;
    XRAM[38521] = 8'b0;
    XRAM[38522] = 8'b0;
    XRAM[38523] = 8'b0;
    XRAM[38524] = 8'b0;
    XRAM[38525] = 8'b0;
    XRAM[38526] = 8'b0;
    XRAM[38527] = 8'b0;
    XRAM[38528] = 8'b0;
    XRAM[38529] = 8'b0;
    XRAM[38530] = 8'b0;
    XRAM[38531] = 8'b0;
    XRAM[38532] = 8'b0;
    XRAM[38533] = 8'b0;
    XRAM[38534] = 8'b0;
    XRAM[38535] = 8'b0;
    XRAM[38536] = 8'b0;
    XRAM[38537] = 8'b0;
    XRAM[38538] = 8'b0;
    XRAM[38539] = 8'b0;
    XRAM[38540] = 8'b0;
    XRAM[38541] = 8'b0;
    XRAM[38542] = 8'b0;
    XRAM[38543] = 8'b0;
    XRAM[38544] = 8'b0;
    XRAM[38545] = 8'b0;
    XRAM[38546] = 8'b0;
    XRAM[38547] = 8'b0;
    XRAM[38548] = 8'b0;
    XRAM[38549] = 8'b0;
    XRAM[38550] = 8'b0;
    XRAM[38551] = 8'b0;
    XRAM[38552] = 8'b0;
    XRAM[38553] = 8'b0;
    XRAM[38554] = 8'b0;
    XRAM[38555] = 8'b0;
    XRAM[38556] = 8'b0;
    XRAM[38557] = 8'b0;
    XRAM[38558] = 8'b0;
    XRAM[38559] = 8'b0;
    XRAM[38560] = 8'b0;
    XRAM[38561] = 8'b0;
    XRAM[38562] = 8'b0;
    XRAM[38563] = 8'b0;
    XRAM[38564] = 8'b0;
    XRAM[38565] = 8'b0;
    XRAM[38566] = 8'b0;
    XRAM[38567] = 8'b0;
    XRAM[38568] = 8'b0;
    XRAM[38569] = 8'b0;
    XRAM[38570] = 8'b0;
    XRAM[38571] = 8'b0;
    XRAM[38572] = 8'b0;
    XRAM[38573] = 8'b0;
    XRAM[38574] = 8'b0;
    XRAM[38575] = 8'b0;
    XRAM[38576] = 8'b0;
    XRAM[38577] = 8'b0;
    XRAM[38578] = 8'b0;
    XRAM[38579] = 8'b0;
    XRAM[38580] = 8'b0;
    XRAM[38581] = 8'b0;
    XRAM[38582] = 8'b0;
    XRAM[38583] = 8'b0;
    XRAM[38584] = 8'b0;
    XRAM[38585] = 8'b0;
    XRAM[38586] = 8'b0;
    XRAM[38587] = 8'b0;
    XRAM[38588] = 8'b0;
    XRAM[38589] = 8'b0;
    XRAM[38590] = 8'b0;
    XRAM[38591] = 8'b0;
    XRAM[38592] = 8'b0;
    XRAM[38593] = 8'b0;
    XRAM[38594] = 8'b0;
    XRAM[38595] = 8'b0;
    XRAM[38596] = 8'b0;
    XRAM[38597] = 8'b0;
    XRAM[38598] = 8'b0;
    XRAM[38599] = 8'b0;
    XRAM[38600] = 8'b0;
    XRAM[38601] = 8'b0;
    XRAM[38602] = 8'b0;
    XRAM[38603] = 8'b0;
    XRAM[38604] = 8'b0;
    XRAM[38605] = 8'b0;
    XRAM[38606] = 8'b0;
    XRAM[38607] = 8'b0;
    XRAM[38608] = 8'b0;
    XRAM[38609] = 8'b0;
    XRAM[38610] = 8'b0;
    XRAM[38611] = 8'b0;
    XRAM[38612] = 8'b0;
    XRAM[38613] = 8'b0;
    XRAM[38614] = 8'b0;
    XRAM[38615] = 8'b0;
    XRAM[38616] = 8'b0;
    XRAM[38617] = 8'b0;
    XRAM[38618] = 8'b0;
    XRAM[38619] = 8'b0;
    XRAM[38620] = 8'b0;
    XRAM[38621] = 8'b0;
    XRAM[38622] = 8'b0;
    XRAM[38623] = 8'b0;
    XRAM[38624] = 8'b0;
    XRAM[38625] = 8'b0;
    XRAM[38626] = 8'b0;
    XRAM[38627] = 8'b0;
    XRAM[38628] = 8'b0;
    XRAM[38629] = 8'b0;
    XRAM[38630] = 8'b0;
    XRAM[38631] = 8'b0;
    XRAM[38632] = 8'b0;
    XRAM[38633] = 8'b0;
    XRAM[38634] = 8'b0;
    XRAM[38635] = 8'b0;
    XRAM[38636] = 8'b0;
    XRAM[38637] = 8'b0;
    XRAM[38638] = 8'b0;
    XRAM[38639] = 8'b0;
    XRAM[38640] = 8'b0;
    XRAM[38641] = 8'b0;
    XRAM[38642] = 8'b0;
    XRAM[38643] = 8'b0;
    XRAM[38644] = 8'b0;
    XRAM[38645] = 8'b0;
    XRAM[38646] = 8'b0;
    XRAM[38647] = 8'b0;
    XRAM[38648] = 8'b0;
    XRAM[38649] = 8'b0;
    XRAM[38650] = 8'b0;
    XRAM[38651] = 8'b0;
    XRAM[38652] = 8'b0;
    XRAM[38653] = 8'b0;
    XRAM[38654] = 8'b0;
    XRAM[38655] = 8'b0;
    XRAM[38656] = 8'b0;
    XRAM[38657] = 8'b0;
    XRAM[38658] = 8'b0;
    XRAM[38659] = 8'b0;
    XRAM[38660] = 8'b0;
    XRAM[38661] = 8'b0;
    XRAM[38662] = 8'b0;
    XRAM[38663] = 8'b0;
    XRAM[38664] = 8'b0;
    XRAM[38665] = 8'b0;
    XRAM[38666] = 8'b0;
    XRAM[38667] = 8'b0;
    XRAM[38668] = 8'b0;
    XRAM[38669] = 8'b0;
    XRAM[38670] = 8'b0;
    XRAM[38671] = 8'b0;
    XRAM[38672] = 8'b0;
    XRAM[38673] = 8'b0;
    XRAM[38674] = 8'b0;
    XRAM[38675] = 8'b0;
    XRAM[38676] = 8'b0;
    XRAM[38677] = 8'b0;
    XRAM[38678] = 8'b0;
    XRAM[38679] = 8'b0;
    XRAM[38680] = 8'b0;
    XRAM[38681] = 8'b0;
    XRAM[38682] = 8'b0;
    XRAM[38683] = 8'b0;
    XRAM[38684] = 8'b0;
    XRAM[38685] = 8'b0;
    XRAM[38686] = 8'b0;
    XRAM[38687] = 8'b0;
    XRAM[38688] = 8'b0;
    XRAM[38689] = 8'b0;
    XRAM[38690] = 8'b0;
    XRAM[38691] = 8'b0;
    XRAM[38692] = 8'b0;
    XRAM[38693] = 8'b0;
    XRAM[38694] = 8'b0;
    XRAM[38695] = 8'b0;
    XRAM[38696] = 8'b0;
    XRAM[38697] = 8'b0;
    XRAM[38698] = 8'b0;
    XRAM[38699] = 8'b0;
    XRAM[38700] = 8'b0;
    XRAM[38701] = 8'b0;
    XRAM[38702] = 8'b0;
    XRAM[38703] = 8'b0;
    XRAM[38704] = 8'b0;
    XRAM[38705] = 8'b0;
    XRAM[38706] = 8'b0;
    XRAM[38707] = 8'b0;
    XRAM[38708] = 8'b0;
    XRAM[38709] = 8'b0;
    XRAM[38710] = 8'b0;
    XRAM[38711] = 8'b0;
    XRAM[38712] = 8'b0;
    XRAM[38713] = 8'b0;
    XRAM[38714] = 8'b0;
    XRAM[38715] = 8'b0;
    XRAM[38716] = 8'b0;
    XRAM[38717] = 8'b0;
    XRAM[38718] = 8'b0;
    XRAM[38719] = 8'b0;
    XRAM[38720] = 8'b0;
    XRAM[38721] = 8'b0;
    XRAM[38722] = 8'b0;
    XRAM[38723] = 8'b0;
    XRAM[38724] = 8'b0;
    XRAM[38725] = 8'b0;
    XRAM[38726] = 8'b0;
    XRAM[38727] = 8'b0;
    XRAM[38728] = 8'b0;
    XRAM[38729] = 8'b0;
    XRAM[38730] = 8'b0;
    XRAM[38731] = 8'b0;
    XRAM[38732] = 8'b0;
    XRAM[38733] = 8'b0;
    XRAM[38734] = 8'b0;
    XRAM[38735] = 8'b0;
    XRAM[38736] = 8'b0;
    XRAM[38737] = 8'b0;
    XRAM[38738] = 8'b0;
    XRAM[38739] = 8'b0;
    XRAM[38740] = 8'b0;
    XRAM[38741] = 8'b0;
    XRAM[38742] = 8'b0;
    XRAM[38743] = 8'b0;
    XRAM[38744] = 8'b0;
    XRAM[38745] = 8'b0;
    XRAM[38746] = 8'b0;
    XRAM[38747] = 8'b0;
    XRAM[38748] = 8'b0;
    XRAM[38749] = 8'b0;
    XRAM[38750] = 8'b0;
    XRAM[38751] = 8'b0;
    XRAM[38752] = 8'b0;
    XRAM[38753] = 8'b0;
    XRAM[38754] = 8'b0;
    XRAM[38755] = 8'b0;
    XRAM[38756] = 8'b0;
    XRAM[38757] = 8'b0;
    XRAM[38758] = 8'b0;
    XRAM[38759] = 8'b0;
    XRAM[38760] = 8'b0;
    XRAM[38761] = 8'b0;
    XRAM[38762] = 8'b0;
    XRAM[38763] = 8'b0;
    XRAM[38764] = 8'b0;
    XRAM[38765] = 8'b0;
    XRAM[38766] = 8'b0;
    XRAM[38767] = 8'b0;
    XRAM[38768] = 8'b0;
    XRAM[38769] = 8'b0;
    XRAM[38770] = 8'b0;
    XRAM[38771] = 8'b0;
    XRAM[38772] = 8'b0;
    XRAM[38773] = 8'b0;
    XRAM[38774] = 8'b0;
    XRAM[38775] = 8'b0;
    XRAM[38776] = 8'b0;
    XRAM[38777] = 8'b0;
    XRAM[38778] = 8'b0;
    XRAM[38779] = 8'b0;
    XRAM[38780] = 8'b0;
    XRAM[38781] = 8'b0;
    XRAM[38782] = 8'b0;
    XRAM[38783] = 8'b0;
    XRAM[38784] = 8'b0;
    XRAM[38785] = 8'b0;
    XRAM[38786] = 8'b0;
    XRAM[38787] = 8'b0;
    XRAM[38788] = 8'b0;
    XRAM[38789] = 8'b0;
    XRAM[38790] = 8'b0;
    XRAM[38791] = 8'b0;
    XRAM[38792] = 8'b0;
    XRAM[38793] = 8'b0;
    XRAM[38794] = 8'b0;
    XRAM[38795] = 8'b0;
    XRAM[38796] = 8'b0;
    XRAM[38797] = 8'b0;
    XRAM[38798] = 8'b0;
    XRAM[38799] = 8'b0;
    XRAM[38800] = 8'b0;
    XRAM[38801] = 8'b0;
    XRAM[38802] = 8'b0;
    XRAM[38803] = 8'b0;
    XRAM[38804] = 8'b0;
    XRAM[38805] = 8'b0;
    XRAM[38806] = 8'b0;
    XRAM[38807] = 8'b0;
    XRAM[38808] = 8'b0;
    XRAM[38809] = 8'b0;
    XRAM[38810] = 8'b0;
    XRAM[38811] = 8'b0;
    XRAM[38812] = 8'b0;
    XRAM[38813] = 8'b0;
    XRAM[38814] = 8'b0;
    XRAM[38815] = 8'b0;
    XRAM[38816] = 8'b0;
    XRAM[38817] = 8'b0;
    XRAM[38818] = 8'b0;
    XRAM[38819] = 8'b0;
    XRAM[38820] = 8'b0;
    XRAM[38821] = 8'b0;
    XRAM[38822] = 8'b0;
    XRAM[38823] = 8'b0;
    XRAM[38824] = 8'b0;
    XRAM[38825] = 8'b0;
    XRAM[38826] = 8'b0;
    XRAM[38827] = 8'b0;
    XRAM[38828] = 8'b0;
    XRAM[38829] = 8'b0;
    XRAM[38830] = 8'b0;
    XRAM[38831] = 8'b0;
    XRAM[38832] = 8'b0;
    XRAM[38833] = 8'b0;
    XRAM[38834] = 8'b0;
    XRAM[38835] = 8'b0;
    XRAM[38836] = 8'b0;
    XRAM[38837] = 8'b0;
    XRAM[38838] = 8'b0;
    XRAM[38839] = 8'b0;
    XRAM[38840] = 8'b0;
    XRAM[38841] = 8'b0;
    XRAM[38842] = 8'b0;
    XRAM[38843] = 8'b0;
    XRAM[38844] = 8'b0;
    XRAM[38845] = 8'b0;
    XRAM[38846] = 8'b0;
    XRAM[38847] = 8'b0;
    XRAM[38848] = 8'b0;
    XRAM[38849] = 8'b0;
    XRAM[38850] = 8'b0;
    XRAM[38851] = 8'b0;
    XRAM[38852] = 8'b0;
    XRAM[38853] = 8'b0;
    XRAM[38854] = 8'b0;
    XRAM[38855] = 8'b0;
    XRAM[38856] = 8'b0;
    XRAM[38857] = 8'b0;
    XRAM[38858] = 8'b0;
    XRAM[38859] = 8'b0;
    XRAM[38860] = 8'b0;
    XRAM[38861] = 8'b0;
    XRAM[38862] = 8'b0;
    XRAM[38863] = 8'b0;
    XRAM[38864] = 8'b0;
    XRAM[38865] = 8'b0;
    XRAM[38866] = 8'b0;
    XRAM[38867] = 8'b0;
    XRAM[38868] = 8'b0;
    XRAM[38869] = 8'b0;
    XRAM[38870] = 8'b0;
    XRAM[38871] = 8'b0;
    XRAM[38872] = 8'b0;
    XRAM[38873] = 8'b0;
    XRAM[38874] = 8'b0;
    XRAM[38875] = 8'b0;
    XRAM[38876] = 8'b0;
    XRAM[38877] = 8'b0;
    XRAM[38878] = 8'b0;
    XRAM[38879] = 8'b0;
    XRAM[38880] = 8'b0;
    XRAM[38881] = 8'b0;
    XRAM[38882] = 8'b0;
    XRAM[38883] = 8'b0;
    XRAM[38884] = 8'b0;
    XRAM[38885] = 8'b0;
    XRAM[38886] = 8'b0;
    XRAM[38887] = 8'b0;
    XRAM[38888] = 8'b0;
    XRAM[38889] = 8'b0;
    XRAM[38890] = 8'b0;
    XRAM[38891] = 8'b0;
    XRAM[38892] = 8'b0;
    XRAM[38893] = 8'b0;
    XRAM[38894] = 8'b0;
    XRAM[38895] = 8'b0;
    XRAM[38896] = 8'b0;
    XRAM[38897] = 8'b0;
    XRAM[38898] = 8'b0;
    XRAM[38899] = 8'b0;
    XRAM[38900] = 8'b0;
    XRAM[38901] = 8'b0;
    XRAM[38902] = 8'b0;
    XRAM[38903] = 8'b0;
    XRAM[38904] = 8'b0;
    XRAM[38905] = 8'b0;
    XRAM[38906] = 8'b0;
    XRAM[38907] = 8'b0;
    XRAM[38908] = 8'b0;
    XRAM[38909] = 8'b0;
    XRAM[38910] = 8'b0;
    XRAM[38911] = 8'b0;
    XRAM[38912] = 8'b0;
    XRAM[38913] = 8'b0;
    XRAM[38914] = 8'b0;
    XRAM[38915] = 8'b0;
    XRAM[38916] = 8'b0;
    XRAM[38917] = 8'b0;
    XRAM[38918] = 8'b0;
    XRAM[38919] = 8'b0;
    XRAM[38920] = 8'b0;
    XRAM[38921] = 8'b0;
    XRAM[38922] = 8'b0;
    XRAM[38923] = 8'b0;
    XRAM[38924] = 8'b0;
    XRAM[38925] = 8'b0;
    XRAM[38926] = 8'b0;
    XRAM[38927] = 8'b0;
    XRAM[38928] = 8'b0;
    XRAM[38929] = 8'b0;
    XRAM[38930] = 8'b0;
    XRAM[38931] = 8'b0;
    XRAM[38932] = 8'b0;
    XRAM[38933] = 8'b0;
    XRAM[38934] = 8'b0;
    XRAM[38935] = 8'b0;
    XRAM[38936] = 8'b0;
    XRAM[38937] = 8'b0;
    XRAM[38938] = 8'b0;
    XRAM[38939] = 8'b0;
    XRAM[38940] = 8'b0;
    XRAM[38941] = 8'b0;
    XRAM[38942] = 8'b0;
    XRAM[38943] = 8'b0;
    XRAM[38944] = 8'b0;
    XRAM[38945] = 8'b0;
    XRAM[38946] = 8'b0;
    XRAM[38947] = 8'b0;
    XRAM[38948] = 8'b0;
    XRAM[38949] = 8'b0;
    XRAM[38950] = 8'b0;
    XRAM[38951] = 8'b0;
    XRAM[38952] = 8'b0;
    XRAM[38953] = 8'b0;
    XRAM[38954] = 8'b0;
    XRAM[38955] = 8'b0;
    XRAM[38956] = 8'b0;
    XRAM[38957] = 8'b0;
    XRAM[38958] = 8'b0;
    XRAM[38959] = 8'b0;
    XRAM[38960] = 8'b0;
    XRAM[38961] = 8'b0;
    XRAM[38962] = 8'b0;
    XRAM[38963] = 8'b0;
    XRAM[38964] = 8'b0;
    XRAM[38965] = 8'b0;
    XRAM[38966] = 8'b0;
    XRAM[38967] = 8'b0;
    XRAM[38968] = 8'b0;
    XRAM[38969] = 8'b0;
    XRAM[38970] = 8'b0;
    XRAM[38971] = 8'b0;
    XRAM[38972] = 8'b0;
    XRAM[38973] = 8'b0;
    XRAM[38974] = 8'b0;
    XRAM[38975] = 8'b0;
    XRAM[38976] = 8'b0;
    XRAM[38977] = 8'b0;
    XRAM[38978] = 8'b0;
    XRAM[38979] = 8'b0;
    XRAM[38980] = 8'b0;
    XRAM[38981] = 8'b0;
    XRAM[38982] = 8'b0;
    XRAM[38983] = 8'b0;
    XRAM[38984] = 8'b0;
    XRAM[38985] = 8'b0;
    XRAM[38986] = 8'b0;
    XRAM[38987] = 8'b0;
    XRAM[38988] = 8'b0;
    XRAM[38989] = 8'b0;
    XRAM[38990] = 8'b0;
    XRAM[38991] = 8'b0;
    XRAM[38992] = 8'b0;
    XRAM[38993] = 8'b0;
    XRAM[38994] = 8'b0;
    XRAM[38995] = 8'b0;
    XRAM[38996] = 8'b0;
    XRAM[38997] = 8'b0;
    XRAM[38998] = 8'b0;
    XRAM[38999] = 8'b0;
    XRAM[39000] = 8'b0;
    XRAM[39001] = 8'b0;
    XRAM[39002] = 8'b0;
    XRAM[39003] = 8'b0;
    XRAM[39004] = 8'b0;
    XRAM[39005] = 8'b0;
    XRAM[39006] = 8'b0;
    XRAM[39007] = 8'b0;
    XRAM[39008] = 8'b0;
    XRAM[39009] = 8'b0;
    XRAM[39010] = 8'b0;
    XRAM[39011] = 8'b0;
    XRAM[39012] = 8'b0;
    XRAM[39013] = 8'b0;
    XRAM[39014] = 8'b0;
    XRAM[39015] = 8'b0;
    XRAM[39016] = 8'b0;
    XRAM[39017] = 8'b0;
    XRAM[39018] = 8'b0;
    XRAM[39019] = 8'b0;
    XRAM[39020] = 8'b0;
    XRAM[39021] = 8'b0;
    XRAM[39022] = 8'b0;
    XRAM[39023] = 8'b0;
    XRAM[39024] = 8'b0;
    XRAM[39025] = 8'b0;
    XRAM[39026] = 8'b0;
    XRAM[39027] = 8'b0;
    XRAM[39028] = 8'b0;
    XRAM[39029] = 8'b0;
    XRAM[39030] = 8'b0;
    XRAM[39031] = 8'b0;
    XRAM[39032] = 8'b0;
    XRAM[39033] = 8'b0;
    XRAM[39034] = 8'b0;
    XRAM[39035] = 8'b0;
    XRAM[39036] = 8'b0;
    XRAM[39037] = 8'b0;
    XRAM[39038] = 8'b0;
    XRAM[39039] = 8'b0;
    XRAM[39040] = 8'b0;
    XRAM[39041] = 8'b0;
    XRAM[39042] = 8'b0;
    XRAM[39043] = 8'b0;
    XRAM[39044] = 8'b0;
    XRAM[39045] = 8'b0;
    XRAM[39046] = 8'b0;
    XRAM[39047] = 8'b0;
    XRAM[39048] = 8'b0;
    XRAM[39049] = 8'b0;
    XRAM[39050] = 8'b0;
    XRAM[39051] = 8'b0;
    XRAM[39052] = 8'b0;
    XRAM[39053] = 8'b0;
    XRAM[39054] = 8'b0;
    XRAM[39055] = 8'b0;
    XRAM[39056] = 8'b0;
    XRAM[39057] = 8'b0;
    XRAM[39058] = 8'b0;
    XRAM[39059] = 8'b0;
    XRAM[39060] = 8'b0;
    XRAM[39061] = 8'b0;
    XRAM[39062] = 8'b0;
    XRAM[39063] = 8'b0;
    XRAM[39064] = 8'b0;
    XRAM[39065] = 8'b0;
    XRAM[39066] = 8'b0;
    XRAM[39067] = 8'b0;
    XRAM[39068] = 8'b0;
    XRAM[39069] = 8'b0;
    XRAM[39070] = 8'b0;
    XRAM[39071] = 8'b0;
    XRAM[39072] = 8'b0;
    XRAM[39073] = 8'b0;
    XRAM[39074] = 8'b0;
    XRAM[39075] = 8'b0;
    XRAM[39076] = 8'b0;
    XRAM[39077] = 8'b0;
    XRAM[39078] = 8'b0;
    XRAM[39079] = 8'b0;
    XRAM[39080] = 8'b0;
    XRAM[39081] = 8'b0;
    XRAM[39082] = 8'b0;
    XRAM[39083] = 8'b0;
    XRAM[39084] = 8'b0;
    XRAM[39085] = 8'b0;
    XRAM[39086] = 8'b0;
    XRAM[39087] = 8'b0;
    XRAM[39088] = 8'b0;
    XRAM[39089] = 8'b0;
    XRAM[39090] = 8'b0;
    XRAM[39091] = 8'b0;
    XRAM[39092] = 8'b0;
    XRAM[39093] = 8'b0;
    XRAM[39094] = 8'b0;
    XRAM[39095] = 8'b0;
    XRAM[39096] = 8'b0;
    XRAM[39097] = 8'b0;
    XRAM[39098] = 8'b0;
    XRAM[39099] = 8'b0;
    XRAM[39100] = 8'b0;
    XRAM[39101] = 8'b0;
    XRAM[39102] = 8'b0;
    XRAM[39103] = 8'b0;
    XRAM[39104] = 8'b0;
    XRAM[39105] = 8'b0;
    XRAM[39106] = 8'b0;
    XRAM[39107] = 8'b0;
    XRAM[39108] = 8'b0;
    XRAM[39109] = 8'b0;
    XRAM[39110] = 8'b0;
    XRAM[39111] = 8'b0;
    XRAM[39112] = 8'b0;
    XRAM[39113] = 8'b0;
    XRAM[39114] = 8'b0;
    XRAM[39115] = 8'b0;
    XRAM[39116] = 8'b0;
    XRAM[39117] = 8'b0;
    XRAM[39118] = 8'b0;
    XRAM[39119] = 8'b0;
    XRAM[39120] = 8'b0;
    XRAM[39121] = 8'b0;
    XRAM[39122] = 8'b0;
    XRAM[39123] = 8'b0;
    XRAM[39124] = 8'b0;
    XRAM[39125] = 8'b0;
    XRAM[39126] = 8'b0;
    XRAM[39127] = 8'b0;
    XRAM[39128] = 8'b0;
    XRAM[39129] = 8'b0;
    XRAM[39130] = 8'b0;
    XRAM[39131] = 8'b0;
    XRAM[39132] = 8'b0;
    XRAM[39133] = 8'b0;
    XRAM[39134] = 8'b0;
    XRAM[39135] = 8'b0;
    XRAM[39136] = 8'b0;
    XRAM[39137] = 8'b0;
    XRAM[39138] = 8'b0;
    XRAM[39139] = 8'b0;
    XRAM[39140] = 8'b0;
    XRAM[39141] = 8'b0;
    XRAM[39142] = 8'b0;
    XRAM[39143] = 8'b0;
    XRAM[39144] = 8'b0;
    XRAM[39145] = 8'b0;
    XRAM[39146] = 8'b0;
    XRAM[39147] = 8'b0;
    XRAM[39148] = 8'b0;
    XRAM[39149] = 8'b0;
    XRAM[39150] = 8'b0;
    XRAM[39151] = 8'b0;
    XRAM[39152] = 8'b0;
    XRAM[39153] = 8'b0;
    XRAM[39154] = 8'b0;
    XRAM[39155] = 8'b0;
    XRAM[39156] = 8'b0;
    XRAM[39157] = 8'b0;
    XRAM[39158] = 8'b0;
    XRAM[39159] = 8'b0;
    XRAM[39160] = 8'b0;
    XRAM[39161] = 8'b0;
    XRAM[39162] = 8'b0;
    XRAM[39163] = 8'b0;
    XRAM[39164] = 8'b0;
    XRAM[39165] = 8'b0;
    XRAM[39166] = 8'b0;
    XRAM[39167] = 8'b0;
    XRAM[39168] = 8'b0;
    XRAM[39169] = 8'b0;
    XRAM[39170] = 8'b0;
    XRAM[39171] = 8'b0;
    XRAM[39172] = 8'b0;
    XRAM[39173] = 8'b0;
    XRAM[39174] = 8'b0;
    XRAM[39175] = 8'b0;
    XRAM[39176] = 8'b0;
    XRAM[39177] = 8'b0;
    XRAM[39178] = 8'b0;
    XRAM[39179] = 8'b0;
    XRAM[39180] = 8'b0;
    XRAM[39181] = 8'b0;
    XRAM[39182] = 8'b0;
    XRAM[39183] = 8'b0;
    XRAM[39184] = 8'b0;
    XRAM[39185] = 8'b0;
    XRAM[39186] = 8'b0;
    XRAM[39187] = 8'b0;
    XRAM[39188] = 8'b0;
    XRAM[39189] = 8'b0;
    XRAM[39190] = 8'b0;
    XRAM[39191] = 8'b0;
    XRAM[39192] = 8'b0;
    XRAM[39193] = 8'b0;
    XRAM[39194] = 8'b0;
    XRAM[39195] = 8'b0;
    XRAM[39196] = 8'b0;
    XRAM[39197] = 8'b0;
    XRAM[39198] = 8'b0;
    XRAM[39199] = 8'b0;
    XRAM[39200] = 8'b0;
    XRAM[39201] = 8'b0;
    XRAM[39202] = 8'b0;
    XRAM[39203] = 8'b0;
    XRAM[39204] = 8'b0;
    XRAM[39205] = 8'b0;
    XRAM[39206] = 8'b0;
    XRAM[39207] = 8'b0;
    XRAM[39208] = 8'b0;
    XRAM[39209] = 8'b0;
    XRAM[39210] = 8'b0;
    XRAM[39211] = 8'b0;
    XRAM[39212] = 8'b0;
    XRAM[39213] = 8'b0;
    XRAM[39214] = 8'b0;
    XRAM[39215] = 8'b0;
    XRAM[39216] = 8'b0;
    XRAM[39217] = 8'b0;
    XRAM[39218] = 8'b0;
    XRAM[39219] = 8'b0;
    XRAM[39220] = 8'b0;
    XRAM[39221] = 8'b0;
    XRAM[39222] = 8'b0;
    XRAM[39223] = 8'b0;
    XRAM[39224] = 8'b0;
    XRAM[39225] = 8'b0;
    XRAM[39226] = 8'b0;
    XRAM[39227] = 8'b0;
    XRAM[39228] = 8'b0;
    XRAM[39229] = 8'b0;
    XRAM[39230] = 8'b0;
    XRAM[39231] = 8'b0;
    XRAM[39232] = 8'b0;
    XRAM[39233] = 8'b0;
    XRAM[39234] = 8'b0;
    XRAM[39235] = 8'b0;
    XRAM[39236] = 8'b0;
    XRAM[39237] = 8'b0;
    XRAM[39238] = 8'b0;
    XRAM[39239] = 8'b0;
    XRAM[39240] = 8'b0;
    XRAM[39241] = 8'b0;
    XRAM[39242] = 8'b0;
    XRAM[39243] = 8'b0;
    XRAM[39244] = 8'b0;
    XRAM[39245] = 8'b0;
    XRAM[39246] = 8'b0;
    XRAM[39247] = 8'b0;
    XRAM[39248] = 8'b0;
    XRAM[39249] = 8'b0;
    XRAM[39250] = 8'b0;
    XRAM[39251] = 8'b0;
    XRAM[39252] = 8'b0;
    XRAM[39253] = 8'b0;
    XRAM[39254] = 8'b0;
    XRAM[39255] = 8'b0;
    XRAM[39256] = 8'b0;
    XRAM[39257] = 8'b0;
    XRAM[39258] = 8'b0;
    XRAM[39259] = 8'b0;
    XRAM[39260] = 8'b0;
    XRAM[39261] = 8'b0;
    XRAM[39262] = 8'b0;
    XRAM[39263] = 8'b0;
    XRAM[39264] = 8'b0;
    XRAM[39265] = 8'b0;
    XRAM[39266] = 8'b0;
    XRAM[39267] = 8'b0;
    XRAM[39268] = 8'b0;
    XRAM[39269] = 8'b0;
    XRAM[39270] = 8'b0;
    XRAM[39271] = 8'b0;
    XRAM[39272] = 8'b0;
    XRAM[39273] = 8'b0;
    XRAM[39274] = 8'b0;
    XRAM[39275] = 8'b0;
    XRAM[39276] = 8'b0;
    XRAM[39277] = 8'b0;
    XRAM[39278] = 8'b0;
    XRAM[39279] = 8'b0;
    XRAM[39280] = 8'b0;
    XRAM[39281] = 8'b0;
    XRAM[39282] = 8'b0;
    XRAM[39283] = 8'b0;
    XRAM[39284] = 8'b0;
    XRAM[39285] = 8'b0;
    XRAM[39286] = 8'b0;
    XRAM[39287] = 8'b0;
    XRAM[39288] = 8'b0;
    XRAM[39289] = 8'b0;
    XRAM[39290] = 8'b0;
    XRAM[39291] = 8'b0;
    XRAM[39292] = 8'b0;
    XRAM[39293] = 8'b0;
    XRAM[39294] = 8'b0;
    XRAM[39295] = 8'b0;
    XRAM[39296] = 8'b0;
    XRAM[39297] = 8'b0;
    XRAM[39298] = 8'b0;
    XRAM[39299] = 8'b0;
    XRAM[39300] = 8'b0;
    XRAM[39301] = 8'b0;
    XRAM[39302] = 8'b0;
    XRAM[39303] = 8'b0;
    XRAM[39304] = 8'b0;
    XRAM[39305] = 8'b0;
    XRAM[39306] = 8'b0;
    XRAM[39307] = 8'b0;
    XRAM[39308] = 8'b0;
    XRAM[39309] = 8'b0;
    XRAM[39310] = 8'b0;
    XRAM[39311] = 8'b0;
    XRAM[39312] = 8'b0;
    XRAM[39313] = 8'b0;
    XRAM[39314] = 8'b0;
    XRAM[39315] = 8'b0;
    XRAM[39316] = 8'b0;
    XRAM[39317] = 8'b0;
    XRAM[39318] = 8'b0;
    XRAM[39319] = 8'b0;
    XRAM[39320] = 8'b0;
    XRAM[39321] = 8'b0;
    XRAM[39322] = 8'b0;
    XRAM[39323] = 8'b0;
    XRAM[39324] = 8'b0;
    XRAM[39325] = 8'b0;
    XRAM[39326] = 8'b0;
    XRAM[39327] = 8'b0;
    XRAM[39328] = 8'b0;
    XRAM[39329] = 8'b0;
    XRAM[39330] = 8'b0;
    XRAM[39331] = 8'b0;
    XRAM[39332] = 8'b0;
    XRAM[39333] = 8'b0;
    XRAM[39334] = 8'b0;
    XRAM[39335] = 8'b0;
    XRAM[39336] = 8'b0;
    XRAM[39337] = 8'b0;
    XRAM[39338] = 8'b0;
    XRAM[39339] = 8'b0;
    XRAM[39340] = 8'b0;
    XRAM[39341] = 8'b0;
    XRAM[39342] = 8'b0;
    XRAM[39343] = 8'b0;
    XRAM[39344] = 8'b0;
    XRAM[39345] = 8'b0;
    XRAM[39346] = 8'b0;
    XRAM[39347] = 8'b0;
    XRAM[39348] = 8'b0;
    XRAM[39349] = 8'b0;
    XRAM[39350] = 8'b0;
    XRAM[39351] = 8'b0;
    XRAM[39352] = 8'b0;
    XRAM[39353] = 8'b0;
    XRAM[39354] = 8'b0;
    XRAM[39355] = 8'b0;
    XRAM[39356] = 8'b0;
    XRAM[39357] = 8'b0;
    XRAM[39358] = 8'b0;
    XRAM[39359] = 8'b0;
    XRAM[39360] = 8'b0;
    XRAM[39361] = 8'b0;
    XRAM[39362] = 8'b0;
    XRAM[39363] = 8'b0;
    XRAM[39364] = 8'b0;
    XRAM[39365] = 8'b0;
    XRAM[39366] = 8'b0;
    XRAM[39367] = 8'b0;
    XRAM[39368] = 8'b0;
    XRAM[39369] = 8'b0;
    XRAM[39370] = 8'b0;
    XRAM[39371] = 8'b0;
    XRAM[39372] = 8'b0;
    XRAM[39373] = 8'b0;
    XRAM[39374] = 8'b0;
    XRAM[39375] = 8'b0;
    XRAM[39376] = 8'b0;
    XRAM[39377] = 8'b0;
    XRAM[39378] = 8'b0;
    XRAM[39379] = 8'b0;
    XRAM[39380] = 8'b0;
    XRAM[39381] = 8'b0;
    XRAM[39382] = 8'b0;
    XRAM[39383] = 8'b0;
    XRAM[39384] = 8'b0;
    XRAM[39385] = 8'b0;
    XRAM[39386] = 8'b0;
    XRAM[39387] = 8'b0;
    XRAM[39388] = 8'b0;
    XRAM[39389] = 8'b0;
    XRAM[39390] = 8'b0;
    XRAM[39391] = 8'b0;
    XRAM[39392] = 8'b0;
    XRAM[39393] = 8'b0;
    XRAM[39394] = 8'b0;
    XRAM[39395] = 8'b0;
    XRAM[39396] = 8'b0;
    XRAM[39397] = 8'b0;
    XRAM[39398] = 8'b0;
    XRAM[39399] = 8'b0;
    XRAM[39400] = 8'b0;
    XRAM[39401] = 8'b0;
    XRAM[39402] = 8'b0;
    XRAM[39403] = 8'b0;
    XRAM[39404] = 8'b0;
    XRAM[39405] = 8'b0;
    XRAM[39406] = 8'b0;
    XRAM[39407] = 8'b0;
    XRAM[39408] = 8'b0;
    XRAM[39409] = 8'b0;
    XRAM[39410] = 8'b0;
    XRAM[39411] = 8'b0;
    XRAM[39412] = 8'b0;
    XRAM[39413] = 8'b0;
    XRAM[39414] = 8'b0;
    XRAM[39415] = 8'b0;
    XRAM[39416] = 8'b0;
    XRAM[39417] = 8'b0;
    XRAM[39418] = 8'b0;
    XRAM[39419] = 8'b0;
    XRAM[39420] = 8'b0;
    XRAM[39421] = 8'b0;
    XRAM[39422] = 8'b0;
    XRAM[39423] = 8'b0;
    XRAM[39424] = 8'b0;
    XRAM[39425] = 8'b0;
    XRAM[39426] = 8'b0;
    XRAM[39427] = 8'b0;
    XRAM[39428] = 8'b0;
    XRAM[39429] = 8'b0;
    XRAM[39430] = 8'b0;
    XRAM[39431] = 8'b0;
    XRAM[39432] = 8'b0;
    XRAM[39433] = 8'b0;
    XRAM[39434] = 8'b0;
    XRAM[39435] = 8'b0;
    XRAM[39436] = 8'b0;
    XRAM[39437] = 8'b0;
    XRAM[39438] = 8'b0;
    XRAM[39439] = 8'b0;
    XRAM[39440] = 8'b0;
    XRAM[39441] = 8'b0;
    XRAM[39442] = 8'b0;
    XRAM[39443] = 8'b0;
    XRAM[39444] = 8'b0;
    XRAM[39445] = 8'b0;
    XRAM[39446] = 8'b0;
    XRAM[39447] = 8'b0;
    XRAM[39448] = 8'b0;
    XRAM[39449] = 8'b0;
    XRAM[39450] = 8'b0;
    XRAM[39451] = 8'b0;
    XRAM[39452] = 8'b0;
    XRAM[39453] = 8'b0;
    XRAM[39454] = 8'b0;
    XRAM[39455] = 8'b0;
    XRAM[39456] = 8'b0;
    XRAM[39457] = 8'b0;
    XRAM[39458] = 8'b0;
    XRAM[39459] = 8'b0;
    XRAM[39460] = 8'b0;
    XRAM[39461] = 8'b0;
    XRAM[39462] = 8'b0;
    XRAM[39463] = 8'b0;
    XRAM[39464] = 8'b0;
    XRAM[39465] = 8'b0;
    XRAM[39466] = 8'b0;
    XRAM[39467] = 8'b0;
    XRAM[39468] = 8'b0;
    XRAM[39469] = 8'b0;
    XRAM[39470] = 8'b0;
    XRAM[39471] = 8'b0;
    XRAM[39472] = 8'b0;
    XRAM[39473] = 8'b0;
    XRAM[39474] = 8'b0;
    XRAM[39475] = 8'b0;
    XRAM[39476] = 8'b0;
    XRAM[39477] = 8'b0;
    XRAM[39478] = 8'b0;
    XRAM[39479] = 8'b0;
    XRAM[39480] = 8'b0;
    XRAM[39481] = 8'b0;
    XRAM[39482] = 8'b0;
    XRAM[39483] = 8'b0;
    XRAM[39484] = 8'b0;
    XRAM[39485] = 8'b0;
    XRAM[39486] = 8'b0;
    XRAM[39487] = 8'b0;
    XRAM[39488] = 8'b0;
    XRAM[39489] = 8'b0;
    XRAM[39490] = 8'b0;
    XRAM[39491] = 8'b0;
    XRAM[39492] = 8'b0;
    XRAM[39493] = 8'b0;
    XRAM[39494] = 8'b0;
    XRAM[39495] = 8'b0;
    XRAM[39496] = 8'b0;
    XRAM[39497] = 8'b0;
    XRAM[39498] = 8'b0;
    XRAM[39499] = 8'b0;
    XRAM[39500] = 8'b0;
    XRAM[39501] = 8'b0;
    XRAM[39502] = 8'b0;
    XRAM[39503] = 8'b0;
    XRAM[39504] = 8'b0;
    XRAM[39505] = 8'b0;
    XRAM[39506] = 8'b0;
    XRAM[39507] = 8'b0;
    XRAM[39508] = 8'b0;
    XRAM[39509] = 8'b0;
    XRAM[39510] = 8'b0;
    XRAM[39511] = 8'b0;
    XRAM[39512] = 8'b0;
    XRAM[39513] = 8'b0;
    XRAM[39514] = 8'b0;
    XRAM[39515] = 8'b0;
    XRAM[39516] = 8'b0;
    XRAM[39517] = 8'b0;
    XRAM[39518] = 8'b0;
    XRAM[39519] = 8'b0;
    XRAM[39520] = 8'b0;
    XRAM[39521] = 8'b0;
    XRAM[39522] = 8'b0;
    XRAM[39523] = 8'b0;
    XRAM[39524] = 8'b0;
    XRAM[39525] = 8'b0;
    XRAM[39526] = 8'b0;
    XRAM[39527] = 8'b0;
    XRAM[39528] = 8'b0;
    XRAM[39529] = 8'b0;
    XRAM[39530] = 8'b0;
    XRAM[39531] = 8'b0;
    XRAM[39532] = 8'b0;
    XRAM[39533] = 8'b0;
    XRAM[39534] = 8'b0;
    XRAM[39535] = 8'b0;
    XRAM[39536] = 8'b0;
    XRAM[39537] = 8'b0;
    XRAM[39538] = 8'b0;
    XRAM[39539] = 8'b0;
    XRAM[39540] = 8'b0;
    XRAM[39541] = 8'b0;
    XRAM[39542] = 8'b0;
    XRAM[39543] = 8'b0;
    XRAM[39544] = 8'b0;
    XRAM[39545] = 8'b0;
    XRAM[39546] = 8'b0;
    XRAM[39547] = 8'b0;
    XRAM[39548] = 8'b0;
    XRAM[39549] = 8'b0;
    XRAM[39550] = 8'b0;
    XRAM[39551] = 8'b0;
    XRAM[39552] = 8'b0;
    XRAM[39553] = 8'b0;
    XRAM[39554] = 8'b0;
    XRAM[39555] = 8'b0;
    XRAM[39556] = 8'b0;
    XRAM[39557] = 8'b0;
    XRAM[39558] = 8'b0;
    XRAM[39559] = 8'b0;
    XRAM[39560] = 8'b0;
    XRAM[39561] = 8'b0;
    XRAM[39562] = 8'b0;
    XRAM[39563] = 8'b0;
    XRAM[39564] = 8'b0;
    XRAM[39565] = 8'b0;
    XRAM[39566] = 8'b0;
    XRAM[39567] = 8'b0;
    XRAM[39568] = 8'b0;
    XRAM[39569] = 8'b0;
    XRAM[39570] = 8'b0;
    XRAM[39571] = 8'b0;
    XRAM[39572] = 8'b0;
    XRAM[39573] = 8'b0;
    XRAM[39574] = 8'b0;
    XRAM[39575] = 8'b0;
    XRAM[39576] = 8'b0;
    XRAM[39577] = 8'b0;
    XRAM[39578] = 8'b0;
    XRAM[39579] = 8'b0;
    XRAM[39580] = 8'b0;
    XRAM[39581] = 8'b0;
    XRAM[39582] = 8'b0;
    XRAM[39583] = 8'b0;
    XRAM[39584] = 8'b0;
    XRAM[39585] = 8'b0;
    XRAM[39586] = 8'b0;
    XRAM[39587] = 8'b0;
    XRAM[39588] = 8'b0;
    XRAM[39589] = 8'b0;
    XRAM[39590] = 8'b0;
    XRAM[39591] = 8'b0;
    XRAM[39592] = 8'b0;
    XRAM[39593] = 8'b0;
    XRAM[39594] = 8'b0;
    XRAM[39595] = 8'b0;
    XRAM[39596] = 8'b0;
    XRAM[39597] = 8'b0;
    XRAM[39598] = 8'b0;
    XRAM[39599] = 8'b0;
    XRAM[39600] = 8'b0;
    XRAM[39601] = 8'b0;
    XRAM[39602] = 8'b0;
    XRAM[39603] = 8'b0;
    XRAM[39604] = 8'b0;
    XRAM[39605] = 8'b0;
    XRAM[39606] = 8'b0;
    XRAM[39607] = 8'b0;
    XRAM[39608] = 8'b0;
    XRAM[39609] = 8'b0;
    XRAM[39610] = 8'b0;
    XRAM[39611] = 8'b0;
    XRAM[39612] = 8'b0;
    XRAM[39613] = 8'b0;
    XRAM[39614] = 8'b0;
    XRAM[39615] = 8'b0;
    XRAM[39616] = 8'b0;
    XRAM[39617] = 8'b0;
    XRAM[39618] = 8'b0;
    XRAM[39619] = 8'b0;
    XRAM[39620] = 8'b0;
    XRAM[39621] = 8'b0;
    XRAM[39622] = 8'b0;
    XRAM[39623] = 8'b0;
    XRAM[39624] = 8'b0;
    XRAM[39625] = 8'b0;
    XRAM[39626] = 8'b0;
    XRAM[39627] = 8'b0;
    XRAM[39628] = 8'b0;
    XRAM[39629] = 8'b0;
    XRAM[39630] = 8'b0;
    XRAM[39631] = 8'b0;
    XRAM[39632] = 8'b0;
    XRAM[39633] = 8'b0;
    XRAM[39634] = 8'b0;
    XRAM[39635] = 8'b0;
    XRAM[39636] = 8'b0;
    XRAM[39637] = 8'b0;
    XRAM[39638] = 8'b0;
    XRAM[39639] = 8'b0;
    XRAM[39640] = 8'b0;
    XRAM[39641] = 8'b0;
    XRAM[39642] = 8'b0;
    XRAM[39643] = 8'b0;
    XRAM[39644] = 8'b0;
    XRAM[39645] = 8'b0;
    XRAM[39646] = 8'b0;
    XRAM[39647] = 8'b0;
    XRAM[39648] = 8'b0;
    XRAM[39649] = 8'b0;
    XRAM[39650] = 8'b0;
    XRAM[39651] = 8'b0;
    XRAM[39652] = 8'b0;
    XRAM[39653] = 8'b0;
    XRAM[39654] = 8'b0;
    XRAM[39655] = 8'b0;
    XRAM[39656] = 8'b0;
    XRAM[39657] = 8'b0;
    XRAM[39658] = 8'b0;
    XRAM[39659] = 8'b0;
    XRAM[39660] = 8'b0;
    XRAM[39661] = 8'b0;
    XRAM[39662] = 8'b0;
    XRAM[39663] = 8'b0;
    XRAM[39664] = 8'b0;
    XRAM[39665] = 8'b0;
    XRAM[39666] = 8'b0;
    XRAM[39667] = 8'b0;
    XRAM[39668] = 8'b0;
    XRAM[39669] = 8'b0;
    XRAM[39670] = 8'b0;
    XRAM[39671] = 8'b0;
    XRAM[39672] = 8'b0;
    XRAM[39673] = 8'b0;
    XRAM[39674] = 8'b0;
    XRAM[39675] = 8'b0;
    XRAM[39676] = 8'b0;
    XRAM[39677] = 8'b0;
    XRAM[39678] = 8'b0;
    XRAM[39679] = 8'b0;
    XRAM[39680] = 8'b0;
    XRAM[39681] = 8'b0;
    XRAM[39682] = 8'b0;
    XRAM[39683] = 8'b0;
    XRAM[39684] = 8'b0;
    XRAM[39685] = 8'b0;
    XRAM[39686] = 8'b0;
    XRAM[39687] = 8'b0;
    XRAM[39688] = 8'b0;
    XRAM[39689] = 8'b0;
    XRAM[39690] = 8'b0;
    XRAM[39691] = 8'b0;
    XRAM[39692] = 8'b0;
    XRAM[39693] = 8'b0;
    XRAM[39694] = 8'b0;
    XRAM[39695] = 8'b0;
    XRAM[39696] = 8'b0;
    XRAM[39697] = 8'b0;
    XRAM[39698] = 8'b0;
    XRAM[39699] = 8'b0;
    XRAM[39700] = 8'b0;
    XRAM[39701] = 8'b0;
    XRAM[39702] = 8'b0;
    XRAM[39703] = 8'b0;
    XRAM[39704] = 8'b0;
    XRAM[39705] = 8'b0;
    XRAM[39706] = 8'b0;
    XRAM[39707] = 8'b0;
    XRAM[39708] = 8'b0;
    XRAM[39709] = 8'b0;
    XRAM[39710] = 8'b0;
    XRAM[39711] = 8'b0;
    XRAM[39712] = 8'b0;
    XRAM[39713] = 8'b0;
    XRAM[39714] = 8'b0;
    XRAM[39715] = 8'b0;
    XRAM[39716] = 8'b0;
    XRAM[39717] = 8'b0;
    XRAM[39718] = 8'b0;
    XRAM[39719] = 8'b0;
    XRAM[39720] = 8'b0;
    XRAM[39721] = 8'b0;
    XRAM[39722] = 8'b0;
    XRAM[39723] = 8'b0;
    XRAM[39724] = 8'b0;
    XRAM[39725] = 8'b0;
    XRAM[39726] = 8'b0;
    XRAM[39727] = 8'b0;
    XRAM[39728] = 8'b0;
    XRAM[39729] = 8'b0;
    XRAM[39730] = 8'b0;
    XRAM[39731] = 8'b0;
    XRAM[39732] = 8'b0;
    XRAM[39733] = 8'b0;
    XRAM[39734] = 8'b0;
    XRAM[39735] = 8'b0;
    XRAM[39736] = 8'b0;
    XRAM[39737] = 8'b0;
    XRAM[39738] = 8'b0;
    XRAM[39739] = 8'b0;
    XRAM[39740] = 8'b0;
    XRAM[39741] = 8'b0;
    XRAM[39742] = 8'b0;
    XRAM[39743] = 8'b0;
    XRAM[39744] = 8'b0;
    XRAM[39745] = 8'b0;
    XRAM[39746] = 8'b0;
    XRAM[39747] = 8'b0;
    XRAM[39748] = 8'b0;
    XRAM[39749] = 8'b0;
    XRAM[39750] = 8'b0;
    XRAM[39751] = 8'b0;
    XRAM[39752] = 8'b0;
    XRAM[39753] = 8'b0;
    XRAM[39754] = 8'b0;
    XRAM[39755] = 8'b0;
    XRAM[39756] = 8'b0;
    XRAM[39757] = 8'b0;
    XRAM[39758] = 8'b0;
    XRAM[39759] = 8'b0;
    XRAM[39760] = 8'b0;
    XRAM[39761] = 8'b0;
    XRAM[39762] = 8'b0;
    XRAM[39763] = 8'b0;
    XRAM[39764] = 8'b0;
    XRAM[39765] = 8'b0;
    XRAM[39766] = 8'b0;
    XRAM[39767] = 8'b0;
    XRAM[39768] = 8'b0;
    XRAM[39769] = 8'b0;
    XRAM[39770] = 8'b0;
    XRAM[39771] = 8'b0;
    XRAM[39772] = 8'b0;
    XRAM[39773] = 8'b0;
    XRAM[39774] = 8'b0;
    XRAM[39775] = 8'b0;
    XRAM[39776] = 8'b0;
    XRAM[39777] = 8'b0;
    XRAM[39778] = 8'b0;
    XRAM[39779] = 8'b0;
    XRAM[39780] = 8'b0;
    XRAM[39781] = 8'b0;
    XRAM[39782] = 8'b0;
    XRAM[39783] = 8'b0;
    XRAM[39784] = 8'b0;
    XRAM[39785] = 8'b0;
    XRAM[39786] = 8'b0;
    XRAM[39787] = 8'b0;
    XRAM[39788] = 8'b0;
    XRAM[39789] = 8'b0;
    XRAM[39790] = 8'b0;
    XRAM[39791] = 8'b0;
    XRAM[39792] = 8'b0;
    XRAM[39793] = 8'b0;
    XRAM[39794] = 8'b0;
    XRAM[39795] = 8'b0;
    XRAM[39796] = 8'b0;
    XRAM[39797] = 8'b0;
    XRAM[39798] = 8'b0;
    XRAM[39799] = 8'b0;
    XRAM[39800] = 8'b0;
    XRAM[39801] = 8'b0;
    XRAM[39802] = 8'b0;
    XRAM[39803] = 8'b0;
    XRAM[39804] = 8'b0;
    XRAM[39805] = 8'b0;
    XRAM[39806] = 8'b0;
    XRAM[39807] = 8'b0;
    XRAM[39808] = 8'b0;
    XRAM[39809] = 8'b0;
    XRAM[39810] = 8'b0;
    XRAM[39811] = 8'b0;
    XRAM[39812] = 8'b0;
    XRAM[39813] = 8'b0;
    XRAM[39814] = 8'b0;
    XRAM[39815] = 8'b0;
    XRAM[39816] = 8'b0;
    XRAM[39817] = 8'b0;
    XRAM[39818] = 8'b0;
    XRAM[39819] = 8'b0;
    XRAM[39820] = 8'b0;
    XRAM[39821] = 8'b0;
    XRAM[39822] = 8'b0;
    XRAM[39823] = 8'b0;
    XRAM[39824] = 8'b0;
    XRAM[39825] = 8'b0;
    XRAM[39826] = 8'b0;
    XRAM[39827] = 8'b0;
    XRAM[39828] = 8'b0;
    XRAM[39829] = 8'b0;
    XRAM[39830] = 8'b0;
    XRAM[39831] = 8'b0;
    XRAM[39832] = 8'b0;
    XRAM[39833] = 8'b0;
    XRAM[39834] = 8'b0;
    XRAM[39835] = 8'b0;
    XRAM[39836] = 8'b0;
    XRAM[39837] = 8'b0;
    XRAM[39838] = 8'b0;
    XRAM[39839] = 8'b0;
    XRAM[39840] = 8'b0;
    XRAM[39841] = 8'b0;
    XRAM[39842] = 8'b0;
    XRAM[39843] = 8'b0;
    XRAM[39844] = 8'b0;
    XRAM[39845] = 8'b0;
    XRAM[39846] = 8'b0;
    XRAM[39847] = 8'b0;
    XRAM[39848] = 8'b0;
    XRAM[39849] = 8'b0;
    XRAM[39850] = 8'b0;
    XRAM[39851] = 8'b0;
    XRAM[39852] = 8'b0;
    XRAM[39853] = 8'b0;
    XRAM[39854] = 8'b0;
    XRAM[39855] = 8'b0;
    XRAM[39856] = 8'b0;
    XRAM[39857] = 8'b0;
    XRAM[39858] = 8'b0;
    XRAM[39859] = 8'b0;
    XRAM[39860] = 8'b0;
    XRAM[39861] = 8'b0;
    XRAM[39862] = 8'b0;
    XRAM[39863] = 8'b0;
    XRAM[39864] = 8'b0;
    XRAM[39865] = 8'b0;
    XRAM[39866] = 8'b0;
    XRAM[39867] = 8'b0;
    XRAM[39868] = 8'b0;
    XRAM[39869] = 8'b0;
    XRAM[39870] = 8'b0;
    XRAM[39871] = 8'b0;
    XRAM[39872] = 8'b0;
    XRAM[39873] = 8'b0;
    XRAM[39874] = 8'b0;
    XRAM[39875] = 8'b0;
    XRAM[39876] = 8'b0;
    XRAM[39877] = 8'b0;
    XRAM[39878] = 8'b0;
    XRAM[39879] = 8'b0;
    XRAM[39880] = 8'b0;
    XRAM[39881] = 8'b0;
    XRAM[39882] = 8'b0;
    XRAM[39883] = 8'b0;
    XRAM[39884] = 8'b0;
    XRAM[39885] = 8'b0;
    XRAM[39886] = 8'b0;
    XRAM[39887] = 8'b0;
    XRAM[39888] = 8'b0;
    XRAM[39889] = 8'b0;
    XRAM[39890] = 8'b0;
    XRAM[39891] = 8'b0;
    XRAM[39892] = 8'b0;
    XRAM[39893] = 8'b0;
    XRAM[39894] = 8'b0;
    XRAM[39895] = 8'b0;
    XRAM[39896] = 8'b0;
    XRAM[39897] = 8'b0;
    XRAM[39898] = 8'b0;
    XRAM[39899] = 8'b0;
    XRAM[39900] = 8'b0;
    XRAM[39901] = 8'b0;
    XRAM[39902] = 8'b0;
    XRAM[39903] = 8'b0;
    XRAM[39904] = 8'b0;
    XRAM[39905] = 8'b0;
    XRAM[39906] = 8'b0;
    XRAM[39907] = 8'b0;
    XRAM[39908] = 8'b0;
    XRAM[39909] = 8'b0;
    XRAM[39910] = 8'b0;
    XRAM[39911] = 8'b0;
    XRAM[39912] = 8'b0;
    XRAM[39913] = 8'b0;
    XRAM[39914] = 8'b0;
    XRAM[39915] = 8'b0;
    XRAM[39916] = 8'b0;
    XRAM[39917] = 8'b0;
    XRAM[39918] = 8'b0;
    XRAM[39919] = 8'b0;
    XRAM[39920] = 8'b0;
    XRAM[39921] = 8'b0;
    XRAM[39922] = 8'b0;
    XRAM[39923] = 8'b0;
    XRAM[39924] = 8'b0;
    XRAM[39925] = 8'b0;
    XRAM[39926] = 8'b0;
    XRAM[39927] = 8'b0;
    XRAM[39928] = 8'b0;
    XRAM[39929] = 8'b0;
    XRAM[39930] = 8'b0;
    XRAM[39931] = 8'b0;
    XRAM[39932] = 8'b0;
    XRAM[39933] = 8'b0;
    XRAM[39934] = 8'b0;
    XRAM[39935] = 8'b0;
    XRAM[39936] = 8'b0;
    XRAM[39937] = 8'b0;
    XRAM[39938] = 8'b0;
    XRAM[39939] = 8'b0;
    XRAM[39940] = 8'b0;
    XRAM[39941] = 8'b0;
    XRAM[39942] = 8'b0;
    XRAM[39943] = 8'b0;
    XRAM[39944] = 8'b0;
    XRAM[39945] = 8'b0;
    XRAM[39946] = 8'b0;
    XRAM[39947] = 8'b0;
    XRAM[39948] = 8'b0;
    XRAM[39949] = 8'b0;
    XRAM[39950] = 8'b0;
    XRAM[39951] = 8'b0;
    XRAM[39952] = 8'b0;
    XRAM[39953] = 8'b0;
    XRAM[39954] = 8'b0;
    XRAM[39955] = 8'b0;
    XRAM[39956] = 8'b0;
    XRAM[39957] = 8'b0;
    XRAM[39958] = 8'b0;
    XRAM[39959] = 8'b0;
    XRAM[39960] = 8'b0;
    XRAM[39961] = 8'b0;
    XRAM[39962] = 8'b0;
    XRAM[39963] = 8'b0;
    XRAM[39964] = 8'b0;
    XRAM[39965] = 8'b0;
    XRAM[39966] = 8'b0;
    XRAM[39967] = 8'b0;
    XRAM[39968] = 8'b0;
    XRAM[39969] = 8'b0;
    XRAM[39970] = 8'b0;
    XRAM[39971] = 8'b0;
    XRAM[39972] = 8'b0;
    XRAM[39973] = 8'b0;
    XRAM[39974] = 8'b0;
    XRAM[39975] = 8'b0;
    XRAM[39976] = 8'b0;
    XRAM[39977] = 8'b0;
    XRAM[39978] = 8'b0;
    XRAM[39979] = 8'b0;
    XRAM[39980] = 8'b0;
    XRAM[39981] = 8'b0;
    XRAM[39982] = 8'b0;
    XRAM[39983] = 8'b0;
    XRAM[39984] = 8'b0;
    XRAM[39985] = 8'b0;
    XRAM[39986] = 8'b0;
    XRAM[39987] = 8'b0;
    XRAM[39988] = 8'b0;
    XRAM[39989] = 8'b0;
    XRAM[39990] = 8'b0;
    XRAM[39991] = 8'b0;
    XRAM[39992] = 8'b0;
    XRAM[39993] = 8'b0;
    XRAM[39994] = 8'b0;
    XRAM[39995] = 8'b0;
    XRAM[39996] = 8'b0;
    XRAM[39997] = 8'b0;
    XRAM[39998] = 8'b0;
    XRAM[39999] = 8'b0;
    XRAM[40000] = 8'b0;
    XRAM[40001] = 8'b0;
    XRAM[40002] = 8'b0;
    XRAM[40003] = 8'b0;
    XRAM[40004] = 8'b0;
    XRAM[40005] = 8'b0;
    XRAM[40006] = 8'b0;
    XRAM[40007] = 8'b0;
    XRAM[40008] = 8'b0;
    XRAM[40009] = 8'b0;
    XRAM[40010] = 8'b0;
    XRAM[40011] = 8'b0;
    XRAM[40012] = 8'b0;
    XRAM[40013] = 8'b0;
    XRAM[40014] = 8'b0;
    XRAM[40015] = 8'b0;
    XRAM[40016] = 8'b0;
    XRAM[40017] = 8'b0;
    XRAM[40018] = 8'b0;
    XRAM[40019] = 8'b0;
    XRAM[40020] = 8'b0;
    XRAM[40021] = 8'b0;
    XRAM[40022] = 8'b0;
    XRAM[40023] = 8'b0;
    XRAM[40024] = 8'b0;
    XRAM[40025] = 8'b0;
    XRAM[40026] = 8'b0;
    XRAM[40027] = 8'b0;
    XRAM[40028] = 8'b0;
    XRAM[40029] = 8'b0;
    XRAM[40030] = 8'b0;
    XRAM[40031] = 8'b0;
    XRAM[40032] = 8'b0;
    XRAM[40033] = 8'b0;
    XRAM[40034] = 8'b0;
    XRAM[40035] = 8'b0;
    XRAM[40036] = 8'b0;
    XRAM[40037] = 8'b0;
    XRAM[40038] = 8'b0;
    XRAM[40039] = 8'b0;
    XRAM[40040] = 8'b0;
    XRAM[40041] = 8'b0;
    XRAM[40042] = 8'b0;
    XRAM[40043] = 8'b0;
    XRAM[40044] = 8'b0;
    XRAM[40045] = 8'b0;
    XRAM[40046] = 8'b0;
    XRAM[40047] = 8'b0;
    XRAM[40048] = 8'b0;
    XRAM[40049] = 8'b0;
    XRAM[40050] = 8'b0;
    XRAM[40051] = 8'b0;
    XRAM[40052] = 8'b0;
    XRAM[40053] = 8'b0;
    XRAM[40054] = 8'b0;
    XRAM[40055] = 8'b0;
    XRAM[40056] = 8'b0;
    XRAM[40057] = 8'b0;
    XRAM[40058] = 8'b0;
    XRAM[40059] = 8'b0;
    XRAM[40060] = 8'b0;
    XRAM[40061] = 8'b0;
    XRAM[40062] = 8'b0;
    XRAM[40063] = 8'b0;
    XRAM[40064] = 8'b0;
    XRAM[40065] = 8'b0;
    XRAM[40066] = 8'b0;
    XRAM[40067] = 8'b0;
    XRAM[40068] = 8'b0;
    XRAM[40069] = 8'b0;
    XRAM[40070] = 8'b0;
    XRAM[40071] = 8'b0;
    XRAM[40072] = 8'b0;
    XRAM[40073] = 8'b0;
    XRAM[40074] = 8'b0;
    XRAM[40075] = 8'b0;
    XRAM[40076] = 8'b0;
    XRAM[40077] = 8'b0;
    XRAM[40078] = 8'b0;
    XRAM[40079] = 8'b0;
    XRAM[40080] = 8'b0;
    XRAM[40081] = 8'b0;
    XRAM[40082] = 8'b0;
    XRAM[40083] = 8'b0;
    XRAM[40084] = 8'b0;
    XRAM[40085] = 8'b0;
    XRAM[40086] = 8'b0;
    XRAM[40087] = 8'b0;
    XRAM[40088] = 8'b0;
    XRAM[40089] = 8'b0;
    XRAM[40090] = 8'b0;
    XRAM[40091] = 8'b0;
    XRAM[40092] = 8'b0;
    XRAM[40093] = 8'b0;
    XRAM[40094] = 8'b0;
    XRAM[40095] = 8'b0;
    XRAM[40096] = 8'b0;
    XRAM[40097] = 8'b0;
    XRAM[40098] = 8'b0;
    XRAM[40099] = 8'b0;
    XRAM[40100] = 8'b0;
    XRAM[40101] = 8'b0;
    XRAM[40102] = 8'b0;
    XRAM[40103] = 8'b0;
    XRAM[40104] = 8'b0;
    XRAM[40105] = 8'b0;
    XRAM[40106] = 8'b0;
    XRAM[40107] = 8'b0;
    XRAM[40108] = 8'b0;
    XRAM[40109] = 8'b0;
    XRAM[40110] = 8'b0;
    XRAM[40111] = 8'b0;
    XRAM[40112] = 8'b0;
    XRAM[40113] = 8'b0;
    XRAM[40114] = 8'b0;
    XRAM[40115] = 8'b0;
    XRAM[40116] = 8'b0;
    XRAM[40117] = 8'b0;
    XRAM[40118] = 8'b0;
    XRAM[40119] = 8'b0;
    XRAM[40120] = 8'b0;
    XRAM[40121] = 8'b0;
    XRAM[40122] = 8'b0;
    XRAM[40123] = 8'b0;
    XRAM[40124] = 8'b0;
    XRAM[40125] = 8'b0;
    XRAM[40126] = 8'b0;
    XRAM[40127] = 8'b0;
    XRAM[40128] = 8'b0;
    XRAM[40129] = 8'b0;
    XRAM[40130] = 8'b0;
    XRAM[40131] = 8'b0;
    XRAM[40132] = 8'b0;
    XRAM[40133] = 8'b0;
    XRAM[40134] = 8'b0;
    XRAM[40135] = 8'b0;
    XRAM[40136] = 8'b0;
    XRAM[40137] = 8'b0;
    XRAM[40138] = 8'b0;
    XRAM[40139] = 8'b0;
    XRAM[40140] = 8'b0;
    XRAM[40141] = 8'b0;
    XRAM[40142] = 8'b0;
    XRAM[40143] = 8'b0;
    XRAM[40144] = 8'b0;
    XRAM[40145] = 8'b0;
    XRAM[40146] = 8'b0;
    XRAM[40147] = 8'b0;
    XRAM[40148] = 8'b0;
    XRAM[40149] = 8'b0;
    XRAM[40150] = 8'b0;
    XRAM[40151] = 8'b0;
    XRAM[40152] = 8'b0;
    XRAM[40153] = 8'b0;
    XRAM[40154] = 8'b0;
    XRAM[40155] = 8'b0;
    XRAM[40156] = 8'b0;
    XRAM[40157] = 8'b0;
    XRAM[40158] = 8'b0;
    XRAM[40159] = 8'b0;
    XRAM[40160] = 8'b0;
    XRAM[40161] = 8'b0;
    XRAM[40162] = 8'b0;
    XRAM[40163] = 8'b0;
    XRAM[40164] = 8'b0;
    XRAM[40165] = 8'b0;
    XRAM[40166] = 8'b0;
    XRAM[40167] = 8'b0;
    XRAM[40168] = 8'b0;
    XRAM[40169] = 8'b0;
    XRAM[40170] = 8'b0;
    XRAM[40171] = 8'b0;
    XRAM[40172] = 8'b0;
    XRAM[40173] = 8'b0;
    XRAM[40174] = 8'b0;
    XRAM[40175] = 8'b0;
    XRAM[40176] = 8'b0;
    XRAM[40177] = 8'b0;
    XRAM[40178] = 8'b0;
    XRAM[40179] = 8'b0;
    XRAM[40180] = 8'b0;
    XRAM[40181] = 8'b0;
    XRAM[40182] = 8'b0;
    XRAM[40183] = 8'b0;
    XRAM[40184] = 8'b0;
    XRAM[40185] = 8'b0;
    XRAM[40186] = 8'b0;
    XRAM[40187] = 8'b0;
    XRAM[40188] = 8'b0;
    XRAM[40189] = 8'b0;
    XRAM[40190] = 8'b0;
    XRAM[40191] = 8'b0;
    XRAM[40192] = 8'b0;
    XRAM[40193] = 8'b0;
    XRAM[40194] = 8'b0;
    XRAM[40195] = 8'b0;
    XRAM[40196] = 8'b0;
    XRAM[40197] = 8'b0;
    XRAM[40198] = 8'b0;
    XRAM[40199] = 8'b0;
    XRAM[40200] = 8'b0;
    XRAM[40201] = 8'b0;
    XRAM[40202] = 8'b0;
    XRAM[40203] = 8'b0;
    XRAM[40204] = 8'b0;
    XRAM[40205] = 8'b0;
    XRAM[40206] = 8'b0;
    XRAM[40207] = 8'b0;
    XRAM[40208] = 8'b0;
    XRAM[40209] = 8'b0;
    XRAM[40210] = 8'b0;
    XRAM[40211] = 8'b0;
    XRAM[40212] = 8'b0;
    XRAM[40213] = 8'b0;
    XRAM[40214] = 8'b0;
    XRAM[40215] = 8'b0;
    XRAM[40216] = 8'b0;
    XRAM[40217] = 8'b0;
    XRAM[40218] = 8'b0;
    XRAM[40219] = 8'b0;
    XRAM[40220] = 8'b0;
    XRAM[40221] = 8'b0;
    XRAM[40222] = 8'b0;
    XRAM[40223] = 8'b0;
    XRAM[40224] = 8'b0;
    XRAM[40225] = 8'b0;
    XRAM[40226] = 8'b0;
    XRAM[40227] = 8'b0;
    XRAM[40228] = 8'b0;
    XRAM[40229] = 8'b0;
    XRAM[40230] = 8'b0;
    XRAM[40231] = 8'b0;
    XRAM[40232] = 8'b0;
    XRAM[40233] = 8'b0;
    XRAM[40234] = 8'b0;
    XRAM[40235] = 8'b0;
    XRAM[40236] = 8'b0;
    XRAM[40237] = 8'b0;
    XRAM[40238] = 8'b0;
    XRAM[40239] = 8'b0;
    XRAM[40240] = 8'b0;
    XRAM[40241] = 8'b0;
    XRAM[40242] = 8'b0;
    XRAM[40243] = 8'b0;
    XRAM[40244] = 8'b0;
    XRAM[40245] = 8'b0;
    XRAM[40246] = 8'b0;
    XRAM[40247] = 8'b0;
    XRAM[40248] = 8'b0;
    XRAM[40249] = 8'b0;
    XRAM[40250] = 8'b0;
    XRAM[40251] = 8'b0;
    XRAM[40252] = 8'b0;
    XRAM[40253] = 8'b0;
    XRAM[40254] = 8'b0;
    XRAM[40255] = 8'b0;
    XRAM[40256] = 8'b0;
    XRAM[40257] = 8'b0;
    XRAM[40258] = 8'b0;
    XRAM[40259] = 8'b0;
    XRAM[40260] = 8'b0;
    XRAM[40261] = 8'b0;
    XRAM[40262] = 8'b0;
    XRAM[40263] = 8'b0;
    XRAM[40264] = 8'b0;
    XRAM[40265] = 8'b0;
    XRAM[40266] = 8'b0;
    XRAM[40267] = 8'b0;
    XRAM[40268] = 8'b0;
    XRAM[40269] = 8'b0;
    XRAM[40270] = 8'b0;
    XRAM[40271] = 8'b0;
    XRAM[40272] = 8'b0;
    XRAM[40273] = 8'b0;
    XRAM[40274] = 8'b0;
    XRAM[40275] = 8'b0;
    XRAM[40276] = 8'b0;
    XRAM[40277] = 8'b0;
    XRAM[40278] = 8'b0;
    XRAM[40279] = 8'b0;
    XRAM[40280] = 8'b0;
    XRAM[40281] = 8'b0;
    XRAM[40282] = 8'b0;
    XRAM[40283] = 8'b0;
    XRAM[40284] = 8'b0;
    XRAM[40285] = 8'b0;
    XRAM[40286] = 8'b0;
    XRAM[40287] = 8'b0;
    XRAM[40288] = 8'b0;
    XRAM[40289] = 8'b0;
    XRAM[40290] = 8'b0;
    XRAM[40291] = 8'b0;
    XRAM[40292] = 8'b0;
    XRAM[40293] = 8'b0;
    XRAM[40294] = 8'b0;
    XRAM[40295] = 8'b0;
    XRAM[40296] = 8'b0;
    XRAM[40297] = 8'b0;
    XRAM[40298] = 8'b0;
    XRAM[40299] = 8'b0;
    XRAM[40300] = 8'b0;
    XRAM[40301] = 8'b0;
    XRAM[40302] = 8'b0;
    XRAM[40303] = 8'b0;
    XRAM[40304] = 8'b0;
    XRAM[40305] = 8'b0;
    XRAM[40306] = 8'b0;
    XRAM[40307] = 8'b0;
    XRAM[40308] = 8'b0;
    XRAM[40309] = 8'b0;
    XRAM[40310] = 8'b0;
    XRAM[40311] = 8'b0;
    XRAM[40312] = 8'b0;
    XRAM[40313] = 8'b0;
    XRAM[40314] = 8'b0;
    XRAM[40315] = 8'b0;
    XRAM[40316] = 8'b0;
    XRAM[40317] = 8'b0;
    XRAM[40318] = 8'b0;
    XRAM[40319] = 8'b0;
    XRAM[40320] = 8'b0;
    XRAM[40321] = 8'b0;
    XRAM[40322] = 8'b0;
    XRAM[40323] = 8'b0;
    XRAM[40324] = 8'b0;
    XRAM[40325] = 8'b0;
    XRAM[40326] = 8'b0;
    XRAM[40327] = 8'b0;
    XRAM[40328] = 8'b0;
    XRAM[40329] = 8'b0;
    XRAM[40330] = 8'b0;
    XRAM[40331] = 8'b0;
    XRAM[40332] = 8'b0;
    XRAM[40333] = 8'b0;
    XRAM[40334] = 8'b0;
    XRAM[40335] = 8'b0;
    XRAM[40336] = 8'b0;
    XRAM[40337] = 8'b0;
    XRAM[40338] = 8'b0;
    XRAM[40339] = 8'b0;
    XRAM[40340] = 8'b0;
    XRAM[40341] = 8'b0;
    XRAM[40342] = 8'b0;
    XRAM[40343] = 8'b0;
    XRAM[40344] = 8'b0;
    XRAM[40345] = 8'b0;
    XRAM[40346] = 8'b0;
    XRAM[40347] = 8'b0;
    XRAM[40348] = 8'b0;
    XRAM[40349] = 8'b0;
    XRAM[40350] = 8'b0;
    XRAM[40351] = 8'b0;
    XRAM[40352] = 8'b0;
    XRAM[40353] = 8'b0;
    XRAM[40354] = 8'b0;
    XRAM[40355] = 8'b0;
    XRAM[40356] = 8'b0;
    XRAM[40357] = 8'b0;
    XRAM[40358] = 8'b0;
    XRAM[40359] = 8'b0;
    XRAM[40360] = 8'b0;
    XRAM[40361] = 8'b0;
    XRAM[40362] = 8'b0;
    XRAM[40363] = 8'b0;
    XRAM[40364] = 8'b0;
    XRAM[40365] = 8'b0;
    XRAM[40366] = 8'b0;
    XRAM[40367] = 8'b0;
    XRAM[40368] = 8'b0;
    XRAM[40369] = 8'b0;
    XRAM[40370] = 8'b0;
    XRAM[40371] = 8'b0;
    XRAM[40372] = 8'b0;
    XRAM[40373] = 8'b0;
    XRAM[40374] = 8'b0;
    XRAM[40375] = 8'b0;
    XRAM[40376] = 8'b0;
    XRAM[40377] = 8'b0;
    XRAM[40378] = 8'b0;
    XRAM[40379] = 8'b0;
    XRAM[40380] = 8'b0;
    XRAM[40381] = 8'b0;
    XRAM[40382] = 8'b0;
    XRAM[40383] = 8'b0;
    XRAM[40384] = 8'b0;
    XRAM[40385] = 8'b0;
    XRAM[40386] = 8'b0;
    XRAM[40387] = 8'b0;
    XRAM[40388] = 8'b0;
    XRAM[40389] = 8'b0;
    XRAM[40390] = 8'b0;
    XRAM[40391] = 8'b0;
    XRAM[40392] = 8'b0;
    XRAM[40393] = 8'b0;
    XRAM[40394] = 8'b0;
    XRAM[40395] = 8'b0;
    XRAM[40396] = 8'b0;
    XRAM[40397] = 8'b0;
    XRAM[40398] = 8'b0;
    XRAM[40399] = 8'b0;
    XRAM[40400] = 8'b0;
    XRAM[40401] = 8'b0;
    XRAM[40402] = 8'b0;
    XRAM[40403] = 8'b0;
    XRAM[40404] = 8'b0;
    XRAM[40405] = 8'b0;
    XRAM[40406] = 8'b0;
    XRAM[40407] = 8'b0;
    XRAM[40408] = 8'b0;
    XRAM[40409] = 8'b0;
    XRAM[40410] = 8'b0;
    XRAM[40411] = 8'b0;
    XRAM[40412] = 8'b0;
    XRAM[40413] = 8'b0;
    XRAM[40414] = 8'b0;
    XRAM[40415] = 8'b0;
    XRAM[40416] = 8'b0;
    XRAM[40417] = 8'b0;
    XRAM[40418] = 8'b0;
    XRAM[40419] = 8'b0;
    XRAM[40420] = 8'b0;
    XRAM[40421] = 8'b0;
    XRAM[40422] = 8'b0;
    XRAM[40423] = 8'b0;
    XRAM[40424] = 8'b0;
    XRAM[40425] = 8'b0;
    XRAM[40426] = 8'b0;
    XRAM[40427] = 8'b0;
    XRAM[40428] = 8'b0;
    XRAM[40429] = 8'b0;
    XRAM[40430] = 8'b0;
    XRAM[40431] = 8'b0;
    XRAM[40432] = 8'b0;
    XRAM[40433] = 8'b0;
    XRAM[40434] = 8'b0;
    XRAM[40435] = 8'b0;
    XRAM[40436] = 8'b0;
    XRAM[40437] = 8'b0;
    XRAM[40438] = 8'b0;
    XRAM[40439] = 8'b0;
    XRAM[40440] = 8'b0;
    XRAM[40441] = 8'b0;
    XRAM[40442] = 8'b0;
    XRAM[40443] = 8'b0;
    XRAM[40444] = 8'b0;
    XRAM[40445] = 8'b0;
    XRAM[40446] = 8'b0;
    XRAM[40447] = 8'b0;
    XRAM[40448] = 8'b0;
    XRAM[40449] = 8'b0;
    XRAM[40450] = 8'b0;
    XRAM[40451] = 8'b0;
    XRAM[40452] = 8'b0;
    XRAM[40453] = 8'b0;
    XRAM[40454] = 8'b0;
    XRAM[40455] = 8'b0;
    XRAM[40456] = 8'b0;
    XRAM[40457] = 8'b0;
    XRAM[40458] = 8'b0;
    XRAM[40459] = 8'b0;
    XRAM[40460] = 8'b0;
    XRAM[40461] = 8'b0;
    XRAM[40462] = 8'b0;
    XRAM[40463] = 8'b0;
    XRAM[40464] = 8'b0;
    XRAM[40465] = 8'b0;
    XRAM[40466] = 8'b0;
    XRAM[40467] = 8'b0;
    XRAM[40468] = 8'b0;
    XRAM[40469] = 8'b0;
    XRAM[40470] = 8'b0;
    XRAM[40471] = 8'b0;
    XRAM[40472] = 8'b0;
    XRAM[40473] = 8'b0;
    XRAM[40474] = 8'b0;
    XRAM[40475] = 8'b0;
    XRAM[40476] = 8'b0;
    XRAM[40477] = 8'b0;
    XRAM[40478] = 8'b0;
    XRAM[40479] = 8'b0;
    XRAM[40480] = 8'b0;
    XRAM[40481] = 8'b0;
    XRAM[40482] = 8'b0;
    XRAM[40483] = 8'b0;
    XRAM[40484] = 8'b0;
    XRAM[40485] = 8'b0;
    XRAM[40486] = 8'b0;
    XRAM[40487] = 8'b0;
    XRAM[40488] = 8'b0;
    XRAM[40489] = 8'b0;
    XRAM[40490] = 8'b0;
    XRAM[40491] = 8'b0;
    XRAM[40492] = 8'b0;
    XRAM[40493] = 8'b0;
    XRAM[40494] = 8'b0;
    XRAM[40495] = 8'b0;
    XRAM[40496] = 8'b0;
    XRAM[40497] = 8'b0;
    XRAM[40498] = 8'b0;
    XRAM[40499] = 8'b0;
    XRAM[40500] = 8'b0;
    XRAM[40501] = 8'b0;
    XRAM[40502] = 8'b0;
    XRAM[40503] = 8'b0;
    XRAM[40504] = 8'b0;
    XRAM[40505] = 8'b0;
    XRAM[40506] = 8'b0;
    XRAM[40507] = 8'b0;
    XRAM[40508] = 8'b0;
    XRAM[40509] = 8'b0;
    XRAM[40510] = 8'b0;
    XRAM[40511] = 8'b0;
    XRAM[40512] = 8'b0;
    XRAM[40513] = 8'b0;
    XRAM[40514] = 8'b0;
    XRAM[40515] = 8'b0;
    XRAM[40516] = 8'b0;
    XRAM[40517] = 8'b0;
    XRAM[40518] = 8'b0;
    XRAM[40519] = 8'b0;
    XRAM[40520] = 8'b0;
    XRAM[40521] = 8'b0;
    XRAM[40522] = 8'b0;
    XRAM[40523] = 8'b0;
    XRAM[40524] = 8'b0;
    XRAM[40525] = 8'b0;
    XRAM[40526] = 8'b0;
    XRAM[40527] = 8'b0;
    XRAM[40528] = 8'b0;
    XRAM[40529] = 8'b0;
    XRAM[40530] = 8'b0;
    XRAM[40531] = 8'b0;
    XRAM[40532] = 8'b0;
    XRAM[40533] = 8'b0;
    XRAM[40534] = 8'b0;
    XRAM[40535] = 8'b0;
    XRAM[40536] = 8'b0;
    XRAM[40537] = 8'b0;
    XRAM[40538] = 8'b0;
    XRAM[40539] = 8'b0;
    XRAM[40540] = 8'b0;
    XRAM[40541] = 8'b0;
    XRAM[40542] = 8'b0;
    XRAM[40543] = 8'b0;
    XRAM[40544] = 8'b0;
    XRAM[40545] = 8'b0;
    XRAM[40546] = 8'b0;
    XRAM[40547] = 8'b0;
    XRAM[40548] = 8'b0;
    XRAM[40549] = 8'b0;
    XRAM[40550] = 8'b0;
    XRAM[40551] = 8'b0;
    XRAM[40552] = 8'b0;
    XRAM[40553] = 8'b0;
    XRAM[40554] = 8'b0;
    XRAM[40555] = 8'b0;
    XRAM[40556] = 8'b0;
    XRAM[40557] = 8'b0;
    XRAM[40558] = 8'b0;
    XRAM[40559] = 8'b0;
    XRAM[40560] = 8'b0;
    XRAM[40561] = 8'b0;
    XRAM[40562] = 8'b0;
    XRAM[40563] = 8'b0;
    XRAM[40564] = 8'b0;
    XRAM[40565] = 8'b0;
    XRAM[40566] = 8'b0;
    XRAM[40567] = 8'b0;
    XRAM[40568] = 8'b0;
    XRAM[40569] = 8'b0;
    XRAM[40570] = 8'b0;
    XRAM[40571] = 8'b0;
    XRAM[40572] = 8'b0;
    XRAM[40573] = 8'b0;
    XRAM[40574] = 8'b0;
    XRAM[40575] = 8'b0;
    XRAM[40576] = 8'b0;
    XRAM[40577] = 8'b0;
    XRAM[40578] = 8'b0;
    XRAM[40579] = 8'b0;
    XRAM[40580] = 8'b0;
    XRAM[40581] = 8'b0;
    XRAM[40582] = 8'b0;
    XRAM[40583] = 8'b0;
    XRAM[40584] = 8'b0;
    XRAM[40585] = 8'b0;
    XRAM[40586] = 8'b0;
    XRAM[40587] = 8'b0;
    XRAM[40588] = 8'b0;
    XRAM[40589] = 8'b0;
    XRAM[40590] = 8'b0;
    XRAM[40591] = 8'b0;
    XRAM[40592] = 8'b0;
    XRAM[40593] = 8'b0;
    XRAM[40594] = 8'b0;
    XRAM[40595] = 8'b0;
    XRAM[40596] = 8'b0;
    XRAM[40597] = 8'b0;
    XRAM[40598] = 8'b0;
    XRAM[40599] = 8'b0;
    XRAM[40600] = 8'b0;
    XRAM[40601] = 8'b0;
    XRAM[40602] = 8'b0;
    XRAM[40603] = 8'b0;
    XRAM[40604] = 8'b0;
    XRAM[40605] = 8'b0;
    XRAM[40606] = 8'b0;
    XRAM[40607] = 8'b0;
    XRAM[40608] = 8'b0;
    XRAM[40609] = 8'b0;
    XRAM[40610] = 8'b0;
    XRAM[40611] = 8'b0;
    XRAM[40612] = 8'b0;
    XRAM[40613] = 8'b0;
    XRAM[40614] = 8'b0;
    XRAM[40615] = 8'b0;
    XRAM[40616] = 8'b0;
    XRAM[40617] = 8'b0;
    XRAM[40618] = 8'b0;
    XRAM[40619] = 8'b0;
    XRAM[40620] = 8'b0;
    XRAM[40621] = 8'b0;
    XRAM[40622] = 8'b0;
    XRAM[40623] = 8'b0;
    XRAM[40624] = 8'b0;
    XRAM[40625] = 8'b0;
    XRAM[40626] = 8'b0;
    XRAM[40627] = 8'b0;
    XRAM[40628] = 8'b0;
    XRAM[40629] = 8'b0;
    XRAM[40630] = 8'b0;
    XRAM[40631] = 8'b0;
    XRAM[40632] = 8'b0;
    XRAM[40633] = 8'b0;
    XRAM[40634] = 8'b0;
    XRAM[40635] = 8'b0;
    XRAM[40636] = 8'b0;
    XRAM[40637] = 8'b0;
    XRAM[40638] = 8'b0;
    XRAM[40639] = 8'b0;
    XRAM[40640] = 8'b0;
    XRAM[40641] = 8'b0;
    XRAM[40642] = 8'b0;
    XRAM[40643] = 8'b0;
    XRAM[40644] = 8'b0;
    XRAM[40645] = 8'b0;
    XRAM[40646] = 8'b0;
    XRAM[40647] = 8'b0;
    XRAM[40648] = 8'b0;
    XRAM[40649] = 8'b0;
    XRAM[40650] = 8'b0;
    XRAM[40651] = 8'b0;
    XRAM[40652] = 8'b0;
    XRAM[40653] = 8'b0;
    XRAM[40654] = 8'b0;
    XRAM[40655] = 8'b0;
    XRAM[40656] = 8'b0;
    XRAM[40657] = 8'b0;
    XRAM[40658] = 8'b0;
    XRAM[40659] = 8'b0;
    XRAM[40660] = 8'b0;
    XRAM[40661] = 8'b0;
    XRAM[40662] = 8'b0;
    XRAM[40663] = 8'b0;
    XRAM[40664] = 8'b0;
    XRAM[40665] = 8'b0;
    XRAM[40666] = 8'b0;
    XRAM[40667] = 8'b0;
    XRAM[40668] = 8'b0;
    XRAM[40669] = 8'b0;
    XRAM[40670] = 8'b0;
    XRAM[40671] = 8'b0;
    XRAM[40672] = 8'b0;
    XRAM[40673] = 8'b0;
    XRAM[40674] = 8'b0;
    XRAM[40675] = 8'b0;
    XRAM[40676] = 8'b0;
    XRAM[40677] = 8'b0;
    XRAM[40678] = 8'b0;
    XRAM[40679] = 8'b0;
    XRAM[40680] = 8'b0;
    XRAM[40681] = 8'b0;
    XRAM[40682] = 8'b0;
    XRAM[40683] = 8'b0;
    XRAM[40684] = 8'b0;
    XRAM[40685] = 8'b0;
    XRAM[40686] = 8'b0;
    XRAM[40687] = 8'b0;
    XRAM[40688] = 8'b0;
    XRAM[40689] = 8'b0;
    XRAM[40690] = 8'b0;
    XRAM[40691] = 8'b0;
    XRAM[40692] = 8'b0;
    XRAM[40693] = 8'b0;
    XRAM[40694] = 8'b0;
    XRAM[40695] = 8'b0;
    XRAM[40696] = 8'b0;
    XRAM[40697] = 8'b0;
    XRAM[40698] = 8'b0;
    XRAM[40699] = 8'b0;
    XRAM[40700] = 8'b0;
    XRAM[40701] = 8'b0;
    XRAM[40702] = 8'b0;
    XRAM[40703] = 8'b0;
    XRAM[40704] = 8'b0;
    XRAM[40705] = 8'b0;
    XRAM[40706] = 8'b0;
    XRAM[40707] = 8'b0;
    XRAM[40708] = 8'b0;
    XRAM[40709] = 8'b0;
    XRAM[40710] = 8'b0;
    XRAM[40711] = 8'b0;
    XRAM[40712] = 8'b0;
    XRAM[40713] = 8'b0;
    XRAM[40714] = 8'b0;
    XRAM[40715] = 8'b0;
    XRAM[40716] = 8'b0;
    XRAM[40717] = 8'b0;
    XRAM[40718] = 8'b0;
    XRAM[40719] = 8'b0;
    XRAM[40720] = 8'b0;
    XRAM[40721] = 8'b0;
    XRAM[40722] = 8'b0;
    XRAM[40723] = 8'b0;
    XRAM[40724] = 8'b0;
    XRAM[40725] = 8'b0;
    XRAM[40726] = 8'b0;
    XRAM[40727] = 8'b0;
    XRAM[40728] = 8'b0;
    XRAM[40729] = 8'b0;
    XRAM[40730] = 8'b0;
    XRAM[40731] = 8'b0;
    XRAM[40732] = 8'b0;
    XRAM[40733] = 8'b0;
    XRAM[40734] = 8'b0;
    XRAM[40735] = 8'b0;
    XRAM[40736] = 8'b0;
    XRAM[40737] = 8'b0;
    XRAM[40738] = 8'b0;
    XRAM[40739] = 8'b0;
    XRAM[40740] = 8'b0;
    XRAM[40741] = 8'b0;
    XRAM[40742] = 8'b0;
    XRAM[40743] = 8'b0;
    XRAM[40744] = 8'b0;
    XRAM[40745] = 8'b0;
    XRAM[40746] = 8'b0;
    XRAM[40747] = 8'b0;
    XRAM[40748] = 8'b0;
    XRAM[40749] = 8'b0;
    XRAM[40750] = 8'b0;
    XRAM[40751] = 8'b0;
    XRAM[40752] = 8'b0;
    XRAM[40753] = 8'b0;
    XRAM[40754] = 8'b0;
    XRAM[40755] = 8'b0;
    XRAM[40756] = 8'b0;
    XRAM[40757] = 8'b0;
    XRAM[40758] = 8'b0;
    XRAM[40759] = 8'b0;
    XRAM[40760] = 8'b0;
    XRAM[40761] = 8'b0;
    XRAM[40762] = 8'b0;
    XRAM[40763] = 8'b0;
    XRAM[40764] = 8'b0;
    XRAM[40765] = 8'b0;
    XRAM[40766] = 8'b0;
    XRAM[40767] = 8'b0;
    XRAM[40768] = 8'b0;
    XRAM[40769] = 8'b0;
    XRAM[40770] = 8'b0;
    XRAM[40771] = 8'b0;
    XRAM[40772] = 8'b0;
    XRAM[40773] = 8'b0;
    XRAM[40774] = 8'b0;
    XRAM[40775] = 8'b0;
    XRAM[40776] = 8'b0;
    XRAM[40777] = 8'b0;
    XRAM[40778] = 8'b0;
    XRAM[40779] = 8'b0;
    XRAM[40780] = 8'b0;
    XRAM[40781] = 8'b0;
    XRAM[40782] = 8'b0;
    XRAM[40783] = 8'b0;
    XRAM[40784] = 8'b0;
    XRAM[40785] = 8'b0;
    XRAM[40786] = 8'b0;
    XRAM[40787] = 8'b0;
    XRAM[40788] = 8'b0;
    XRAM[40789] = 8'b0;
    XRAM[40790] = 8'b0;
    XRAM[40791] = 8'b0;
    XRAM[40792] = 8'b0;
    XRAM[40793] = 8'b0;
    XRAM[40794] = 8'b0;
    XRAM[40795] = 8'b0;
    XRAM[40796] = 8'b0;
    XRAM[40797] = 8'b0;
    XRAM[40798] = 8'b0;
    XRAM[40799] = 8'b0;
    XRAM[40800] = 8'b0;
    XRAM[40801] = 8'b0;
    XRAM[40802] = 8'b0;
    XRAM[40803] = 8'b0;
    XRAM[40804] = 8'b0;
    XRAM[40805] = 8'b0;
    XRAM[40806] = 8'b0;
    XRAM[40807] = 8'b0;
    XRAM[40808] = 8'b0;
    XRAM[40809] = 8'b0;
    XRAM[40810] = 8'b0;
    XRAM[40811] = 8'b0;
    XRAM[40812] = 8'b0;
    XRAM[40813] = 8'b0;
    XRAM[40814] = 8'b0;
    XRAM[40815] = 8'b0;
    XRAM[40816] = 8'b0;
    XRAM[40817] = 8'b0;
    XRAM[40818] = 8'b0;
    XRAM[40819] = 8'b0;
    XRAM[40820] = 8'b0;
    XRAM[40821] = 8'b0;
    XRAM[40822] = 8'b0;
    XRAM[40823] = 8'b0;
    XRAM[40824] = 8'b0;
    XRAM[40825] = 8'b0;
    XRAM[40826] = 8'b0;
    XRAM[40827] = 8'b0;
    XRAM[40828] = 8'b0;
    XRAM[40829] = 8'b0;
    XRAM[40830] = 8'b0;
    XRAM[40831] = 8'b0;
    XRAM[40832] = 8'b0;
    XRAM[40833] = 8'b0;
    XRAM[40834] = 8'b0;
    XRAM[40835] = 8'b0;
    XRAM[40836] = 8'b0;
    XRAM[40837] = 8'b0;
    XRAM[40838] = 8'b0;
    XRAM[40839] = 8'b0;
    XRAM[40840] = 8'b0;
    XRAM[40841] = 8'b0;
    XRAM[40842] = 8'b0;
    XRAM[40843] = 8'b0;
    XRAM[40844] = 8'b0;
    XRAM[40845] = 8'b0;
    XRAM[40846] = 8'b0;
    XRAM[40847] = 8'b0;
    XRAM[40848] = 8'b0;
    XRAM[40849] = 8'b0;
    XRAM[40850] = 8'b0;
    XRAM[40851] = 8'b0;
    XRAM[40852] = 8'b0;
    XRAM[40853] = 8'b0;
    XRAM[40854] = 8'b0;
    XRAM[40855] = 8'b0;
    XRAM[40856] = 8'b0;
    XRAM[40857] = 8'b0;
    XRAM[40858] = 8'b0;
    XRAM[40859] = 8'b0;
    XRAM[40860] = 8'b0;
    XRAM[40861] = 8'b0;
    XRAM[40862] = 8'b0;
    XRAM[40863] = 8'b0;
    XRAM[40864] = 8'b0;
    XRAM[40865] = 8'b0;
    XRAM[40866] = 8'b0;
    XRAM[40867] = 8'b0;
    XRAM[40868] = 8'b0;
    XRAM[40869] = 8'b0;
    XRAM[40870] = 8'b0;
    XRAM[40871] = 8'b0;
    XRAM[40872] = 8'b0;
    XRAM[40873] = 8'b0;
    XRAM[40874] = 8'b0;
    XRAM[40875] = 8'b0;
    XRAM[40876] = 8'b0;
    XRAM[40877] = 8'b0;
    XRAM[40878] = 8'b0;
    XRAM[40879] = 8'b0;
    XRAM[40880] = 8'b0;
    XRAM[40881] = 8'b0;
    XRAM[40882] = 8'b0;
    XRAM[40883] = 8'b0;
    XRAM[40884] = 8'b0;
    XRAM[40885] = 8'b0;
    XRAM[40886] = 8'b0;
    XRAM[40887] = 8'b0;
    XRAM[40888] = 8'b0;
    XRAM[40889] = 8'b0;
    XRAM[40890] = 8'b0;
    XRAM[40891] = 8'b0;
    XRAM[40892] = 8'b0;
    XRAM[40893] = 8'b0;
    XRAM[40894] = 8'b0;
    XRAM[40895] = 8'b0;
    XRAM[40896] = 8'b0;
    XRAM[40897] = 8'b0;
    XRAM[40898] = 8'b0;
    XRAM[40899] = 8'b0;
    XRAM[40900] = 8'b0;
    XRAM[40901] = 8'b0;
    XRAM[40902] = 8'b0;
    XRAM[40903] = 8'b0;
    XRAM[40904] = 8'b0;
    XRAM[40905] = 8'b0;
    XRAM[40906] = 8'b0;
    XRAM[40907] = 8'b0;
    XRAM[40908] = 8'b0;
    XRAM[40909] = 8'b0;
    XRAM[40910] = 8'b0;
    XRAM[40911] = 8'b0;
    XRAM[40912] = 8'b0;
    XRAM[40913] = 8'b0;
    XRAM[40914] = 8'b0;
    XRAM[40915] = 8'b0;
    XRAM[40916] = 8'b0;
    XRAM[40917] = 8'b0;
    XRAM[40918] = 8'b0;
    XRAM[40919] = 8'b0;
    XRAM[40920] = 8'b0;
    XRAM[40921] = 8'b0;
    XRAM[40922] = 8'b0;
    XRAM[40923] = 8'b0;
    XRAM[40924] = 8'b0;
    XRAM[40925] = 8'b0;
    XRAM[40926] = 8'b0;
    XRAM[40927] = 8'b0;
    XRAM[40928] = 8'b0;
    XRAM[40929] = 8'b0;
    XRAM[40930] = 8'b0;
    XRAM[40931] = 8'b0;
    XRAM[40932] = 8'b0;
    XRAM[40933] = 8'b0;
    XRAM[40934] = 8'b0;
    XRAM[40935] = 8'b0;
    XRAM[40936] = 8'b0;
    XRAM[40937] = 8'b0;
    XRAM[40938] = 8'b0;
    XRAM[40939] = 8'b0;
    XRAM[40940] = 8'b0;
    XRAM[40941] = 8'b0;
    XRAM[40942] = 8'b0;
    XRAM[40943] = 8'b0;
    XRAM[40944] = 8'b0;
    XRAM[40945] = 8'b0;
    XRAM[40946] = 8'b0;
    XRAM[40947] = 8'b0;
    XRAM[40948] = 8'b0;
    XRAM[40949] = 8'b0;
    XRAM[40950] = 8'b0;
    XRAM[40951] = 8'b0;
    XRAM[40952] = 8'b0;
    XRAM[40953] = 8'b0;
    XRAM[40954] = 8'b0;
    XRAM[40955] = 8'b0;
    XRAM[40956] = 8'b0;
    XRAM[40957] = 8'b0;
    XRAM[40958] = 8'b0;
    XRAM[40959] = 8'b0;
    XRAM[40960] = 8'b0;
    XRAM[40961] = 8'b0;
    XRAM[40962] = 8'b0;
    XRAM[40963] = 8'b0;
    XRAM[40964] = 8'b0;
    XRAM[40965] = 8'b0;
    XRAM[40966] = 8'b0;
    XRAM[40967] = 8'b0;
    XRAM[40968] = 8'b0;
    XRAM[40969] = 8'b0;
    XRAM[40970] = 8'b0;
    XRAM[40971] = 8'b0;
    XRAM[40972] = 8'b0;
    XRAM[40973] = 8'b0;
    XRAM[40974] = 8'b0;
    XRAM[40975] = 8'b0;
    XRAM[40976] = 8'b0;
    XRAM[40977] = 8'b0;
    XRAM[40978] = 8'b0;
    XRAM[40979] = 8'b0;
    XRAM[40980] = 8'b0;
    XRAM[40981] = 8'b0;
    XRAM[40982] = 8'b0;
    XRAM[40983] = 8'b0;
    XRAM[40984] = 8'b0;
    XRAM[40985] = 8'b0;
    XRAM[40986] = 8'b0;
    XRAM[40987] = 8'b0;
    XRAM[40988] = 8'b0;
    XRAM[40989] = 8'b0;
    XRAM[40990] = 8'b0;
    XRAM[40991] = 8'b0;
    XRAM[40992] = 8'b0;
    XRAM[40993] = 8'b0;
    XRAM[40994] = 8'b0;
    XRAM[40995] = 8'b0;
    XRAM[40996] = 8'b0;
    XRAM[40997] = 8'b0;
    XRAM[40998] = 8'b0;
    XRAM[40999] = 8'b0;
    XRAM[41000] = 8'b0;
    XRAM[41001] = 8'b0;
    XRAM[41002] = 8'b0;
    XRAM[41003] = 8'b0;
    XRAM[41004] = 8'b0;
    XRAM[41005] = 8'b0;
    XRAM[41006] = 8'b0;
    XRAM[41007] = 8'b0;
    XRAM[41008] = 8'b0;
    XRAM[41009] = 8'b0;
    XRAM[41010] = 8'b0;
    XRAM[41011] = 8'b0;
    XRAM[41012] = 8'b0;
    XRAM[41013] = 8'b0;
    XRAM[41014] = 8'b0;
    XRAM[41015] = 8'b0;
    XRAM[41016] = 8'b0;
    XRAM[41017] = 8'b0;
    XRAM[41018] = 8'b0;
    XRAM[41019] = 8'b0;
    XRAM[41020] = 8'b0;
    XRAM[41021] = 8'b0;
    XRAM[41022] = 8'b0;
    XRAM[41023] = 8'b0;
    XRAM[41024] = 8'b0;
    XRAM[41025] = 8'b0;
    XRAM[41026] = 8'b0;
    XRAM[41027] = 8'b0;
    XRAM[41028] = 8'b0;
    XRAM[41029] = 8'b0;
    XRAM[41030] = 8'b0;
    XRAM[41031] = 8'b0;
    XRAM[41032] = 8'b0;
    XRAM[41033] = 8'b0;
    XRAM[41034] = 8'b0;
    XRAM[41035] = 8'b0;
    XRAM[41036] = 8'b0;
    XRAM[41037] = 8'b0;
    XRAM[41038] = 8'b0;
    XRAM[41039] = 8'b0;
    XRAM[41040] = 8'b0;
    XRAM[41041] = 8'b0;
    XRAM[41042] = 8'b0;
    XRAM[41043] = 8'b0;
    XRAM[41044] = 8'b0;
    XRAM[41045] = 8'b0;
    XRAM[41046] = 8'b0;
    XRAM[41047] = 8'b0;
    XRAM[41048] = 8'b0;
    XRAM[41049] = 8'b0;
    XRAM[41050] = 8'b0;
    XRAM[41051] = 8'b0;
    XRAM[41052] = 8'b0;
    XRAM[41053] = 8'b0;
    XRAM[41054] = 8'b0;
    XRAM[41055] = 8'b0;
    XRAM[41056] = 8'b0;
    XRAM[41057] = 8'b0;
    XRAM[41058] = 8'b0;
    XRAM[41059] = 8'b0;
    XRAM[41060] = 8'b0;
    XRAM[41061] = 8'b0;
    XRAM[41062] = 8'b0;
    XRAM[41063] = 8'b0;
    XRAM[41064] = 8'b0;
    XRAM[41065] = 8'b0;
    XRAM[41066] = 8'b0;
    XRAM[41067] = 8'b0;
    XRAM[41068] = 8'b0;
    XRAM[41069] = 8'b0;
    XRAM[41070] = 8'b0;
    XRAM[41071] = 8'b0;
    XRAM[41072] = 8'b0;
    XRAM[41073] = 8'b0;
    XRAM[41074] = 8'b0;
    XRAM[41075] = 8'b0;
    XRAM[41076] = 8'b0;
    XRAM[41077] = 8'b0;
    XRAM[41078] = 8'b0;
    XRAM[41079] = 8'b0;
    XRAM[41080] = 8'b0;
    XRAM[41081] = 8'b0;
    XRAM[41082] = 8'b0;
    XRAM[41083] = 8'b0;
    XRAM[41084] = 8'b0;
    XRAM[41085] = 8'b0;
    XRAM[41086] = 8'b0;
    XRAM[41087] = 8'b0;
    XRAM[41088] = 8'b0;
    XRAM[41089] = 8'b0;
    XRAM[41090] = 8'b0;
    XRAM[41091] = 8'b0;
    XRAM[41092] = 8'b0;
    XRAM[41093] = 8'b0;
    XRAM[41094] = 8'b0;
    XRAM[41095] = 8'b0;
    XRAM[41096] = 8'b0;
    XRAM[41097] = 8'b0;
    XRAM[41098] = 8'b0;
    XRAM[41099] = 8'b0;
    XRAM[41100] = 8'b0;
    XRAM[41101] = 8'b0;
    XRAM[41102] = 8'b0;
    XRAM[41103] = 8'b0;
    XRAM[41104] = 8'b0;
    XRAM[41105] = 8'b0;
    XRAM[41106] = 8'b0;
    XRAM[41107] = 8'b0;
    XRAM[41108] = 8'b0;
    XRAM[41109] = 8'b0;
    XRAM[41110] = 8'b0;
    XRAM[41111] = 8'b0;
    XRAM[41112] = 8'b0;
    XRAM[41113] = 8'b0;
    XRAM[41114] = 8'b0;
    XRAM[41115] = 8'b0;
    XRAM[41116] = 8'b0;
    XRAM[41117] = 8'b0;
    XRAM[41118] = 8'b0;
    XRAM[41119] = 8'b0;
    XRAM[41120] = 8'b0;
    XRAM[41121] = 8'b0;
    XRAM[41122] = 8'b0;
    XRAM[41123] = 8'b0;
    XRAM[41124] = 8'b0;
    XRAM[41125] = 8'b0;
    XRAM[41126] = 8'b0;
    XRAM[41127] = 8'b0;
    XRAM[41128] = 8'b0;
    XRAM[41129] = 8'b0;
    XRAM[41130] = 8'b0;
    XRAM[41131] = 8'b0;
    XRAM[41132] = 8'b0;
    XRAM[41133] = 8'b0;
    XRAM[41134] = 8'b0;
    XRAM[41135] = 8'b0;
    XRAM[41136] = 8'b0;
    XRAM[41137] = 8'b0;
    XRAM[41138] = 8'b0;
    XRAM[41139] = 8'b0;
    XRAM[41140] = 8'b0;
    XRAM[41141] = 8'b0;
    XRAM[41142] = 8'b0;
    XRAM[41143] = 8'b0;
    XRAM[41144] = 8'b0;
    XRAM[41145] = 8'b0;
    XRAM[41146] = 8'b0;
    XRAM[41147] = 8'b0;
    XRAM[41148] = 8'b0;
    XRAM[41149] = 8'b0;
    XRAM[41150] = 8'b0;
    XRAM[41151] = 8'b0;
    XRAM[41152] = 8'b0;
    XRAM[41153] = 8'b0;
    XRAM[41154] = 8'b0;
    XRAM[41155] = 8'b0;
    XRAM[41156] = 8'b0;
    XRAM[41157] = 8'b0;
    XRAM[41158] = 8'b0;
    XRAM[41159] = 8'b0;
    XRAM[41160] = 8'b0;
    XRAM[41161] = 8'b0;
    XRAM[41162] = 8'b0;
    XRAM[41163] = 8'b0;
    XRAM[41164] = 8'b0;
    XRAM[41165] = 8'b0;
    XRAM[41166] = 8'b0;
    XRAM[41167] = 8'b0;
    XRAM[41168] = 8'b0;
    XRAM[41169] = 8'b0;
    XRAM[41170] = 8'b0;
    XRAM[41171] = 8'b0;
    XRAM[41172] = 8'b0;
    XRAM[41173] = 8'b0;
    XRAM[41174] = 8'b0;
    XRAM[41175] = 8'b0;
    XRAM[41176] = 8'b0;
    XRAM[41177] = 8'b0;
    XRAM[41178] = 8'b0;
    XRAM[41179] = 8'b0;
    XRAM[41180] = 8'b0;
    XRAM[41181] = 8'b0;
    XRAM[41182] = 8'b0;
    XRAM[41183] = 8'b0;
    XRAM[41184] = 8'b0;
    XRAM[41185] = 8'b0;
    XRAM[41186] = 8'b0;
    XRAM[41187] = 8'b0;
    XRAM[41188] = 8'b0;
    XRAM[41189] = 8'b0;
    XRAM[41190] = 8'b0;
    XRAM[41191] = 8'b0;
    XRAM[41192] = 8'b0;
    XRAM[41193] = 8'b0;
    XRAM[41194] = 8'b0;
    XRAM[41195] = 8'b0;
    XRAM[41196] = 8'b0;
    XRAM[41197] = 8'b0;
    XRAM[41198] = 8'b0;
    XRAM[41199] = 8'b0;
    XRAM[41200] = 8'b0;
    XRAM[41201] = 8'b0;
    XRAM[41202] = 8'b0;
    XRAM[41203] = 8'b0;
    XRAM[41204] = 8'b0;
    XRAM[41205] = 8'b0;
    XRAM[41206] = 8'b0;
    XRAM[41207] = 8'b0;
    XRAM[41208] = 8'b0;
    XRAM[41209] = 8'b0;
    XRAM[41210] = 8'b0;
    XRAM[41211] = 8'b0;
    XRAM[41212] = 8'b0;
    XRAM[41213] = 8'b0;
    XRAM[41214] = 8'b0;
    XRAM[41215] = 8'b0;
    XRAM[41216] = 8'b0;
    XRAM[41217] = 8'b0;
    XRAM[41218] = 8'b0;
    XRAM[41219] = 8'b0;
    XRAM[41220] = 8'b0;
    XRAM[41221] = 8'b0;
    XRAM[41222] = 8'b0;
    XRAM[41223] = 8'b0;
    XRAM[41224] = 8'b0;
    XRAM[41225] = 8'b0;
    XRAM[41226] = 8'b0;
    XRAM[41227] = 8'b0;
    XRAM[41228] = 8'b0;
    XRAM[41229] = 8'b0;
    XRAM[41230] = 8'b0;
    XRAM[41231] = 8'b0;
    XRAM[41232] = 8'b0;
    XRAM[41233] = 8'b0;
    XRAM[41234] = 8'b0;
    XRAM[41235] = 8'b0;
    XRAM[41236] = 8'b0;
    XRAM[41237] = 8'b0;
    XRAM[41238] = 8'b0;
    XRAM[41239] = 8'b0;
    XRAM[41240] = 8'b0;
    XRAM[41241] = 8'b0;
    XRAM[41242] = 8'b0;
    XRAM[41243] = 8'b0;
    XRAM[41244] = 8'b0;
    XRAM[41245] = 8'b0;
    XRAM[41246] = 8'b0;
    XRAM[41247] = 8'b0;
    XRAM[41248] = 8'b0;
    XRAM[41249] = 8'b0;
    XRAM[41250] = 8'b0;
    XRAM[41251] = 8'b0;
    XRAM[41252] = 8'b0;
    XRAM[41253] = 8'b0;
    XRAM[41254] = 8'b0;
    XRAM[41255] = 8'b0;
    XRAM[41256] = 8'b0;
    XRAM[41257] = 8'b0;
    XRAM[41258] = 8'b0;
    XRAM[41259] = 8'b0;
    XRAM[41260] = 8'b0;
    XRAM[41261] = 8'b0;
    XRAM[41262] = 8'b0;
    XRAM[41263] = 8'b0;
    XRAM[41264] = 8'b0;
    XRAM[41265] = 8'b0;
    XRAM[41266] = 8'b0;
    XRAM[41267] = 8'b0;
    XRAM[41268] = 8'b0;
    XRAM[41269] = 8'b0;
    XRAM[41270] = 8'b0;
    XRAM[41271] = 8'b0;
    XRAM[41272] = 8'b0;
    XRAM[41273] = 8'b0;
    XRAM[41274] = 8'b0;
    XRAM[41275] = 8'b0;
    XRAM[41276] = 8'b0;
    XRAM[41277] = 8'b0;
    XRAM[41278] = 8'b0;
    XRAM[41279] = 8'b0;
    XRAM[41280] = 8'b0;
    XRAM[41281] = 8'b0;
    XRAM[41282] = 8'b0;
    XRAM[41283] = 8'b0;
    XRAM[41284] = 8'b0;
    XRAM[41285] = 8'b0;
    XRAM[41286] = 8'b0;
    XRAM[41287] = 8'b0;
    XRAM[41288] = 8'b0;
    XRAM[41289] = 8'b0;
    XRAM[41290] = 8'b0;
    XRAM[41291] = 8'b0;
    XRAM[41292] = 8'b0;
    XRAM[41293] = 8'b0;
    XRAM[41294] = 8'b0;
    XRAM[41295] = 8'b0;
    XRAM[41296] = 8'b0;
    XRAM[41297] = 8'b0;
    XRAM[41298] = 8'b0;
    XRAM[41299] = 8'b0;
    XRAM[41300] = 8'b0;
    XRAM[41301] = 8'b0;
    XRAM[41302] = 8'b0;
    XRAM[41303] = 8'b0;
    XRAM[41304] = 8'b0;
    XRAM[41305] = 8'b0;
    XRAM[41306] = 8'b0;
    XRAM[41307] = 8'b0;
    XRAM[41308] = 8'b0;
    XRAM[41309] = 8'b0;
    XRAM[41310] = 8'b0;
    XRAM[41311] = 8'b0;
    XRAM[41312] = 8'b0;
    XRAM[41313] = 8'b0;
    XRAM[41314] = 8'b0;
    XRAM[41315] = 8'b0;
    XRAM[41316] = 8'b0;
    XRAM[41317] = 8'b0;
    XRAM[41318] = 8'b0;
    XRAM[41319] = 8'b0;
    XRAM[41320] = 8'b0;
    XRAM[41321] = 8'b0;
    XRAM[41322] = 8'b0;
    XRAM[41323] = 8'b0;
    XRAM[41324] = 8'b0;
    XRAM[41325] = 8'b0;
    XRAM[41326] = 8'b0;
    XRAM[41327] = 8'b0;
    XRAM[41328] = 8'b0;
    XRAM[41329] = 8'b0;
    XRAM[41330] = 8'b0;
    XRAM[41331] = 8'b0;
    XRAM[41332] = 8'b0;
    XRAM[41333] = 8'b0;
    XRAM[41334] = 8'b0;
    XRAM[41335] = 8'b0;
    XRAM[41336] = 8'b0;
    XRAM[41337] = 8'b0;
    XRAM[41338] = 8'b0;
    XRAM[41339] = 8'b0;
    XRAM[41340] = 8'b0;
    XRAM[41341] = 8'b0;
    XRAM[41342] = 8'b0;
    XRAM[41343] = 8'b0;
    XRAM[41344] = 8'b0;
    XRAM[41345] = 8'b0;
    XRAM[41346] = 8'b0;
    XRAM[41347] = 8'b0;
    XRAM[41348] = 8'b0;
    XRAM[41349] = 8'b0;
    XRAM[41350] = 8'b0;
    XRAM[41351] = 8'b0;
    XRAM[41352] = 8'b0;
    XRAM[41353] = 8'b0;
    XRAM[41354] = 8'b0;
    XRAM[41355] = 8'b0;
    XRAM[41356] = 8'b0;
    XRAM[41357] = 8'b0;
    XRAM[41358] = 8'b0;
    XRAM[41359] = 8'b0;
    XRAM[41360] = 8'b0;
    XRAM[41361] = 8'b0;
    XRAM[41362] = 8'b0;
    XRAM[41363] = 8'b0;
    XRAM[41364] = 8'b0;
    XRAM[41365] = 8'b0;
    XRAM[41366] = 8'b0;
    XRAM[41367] = 8'b0;
    XRAM[41368] = 8'b0;
    XRAM[41369] = 8'b0;
    XRAM[41370] = 8'b0;
    XRAM[41371] = 8'b0;
    XRAM[41372] = 8'b0;
    XRAM[41373] = 8'b0;
    XRAM[41374] = 8'b0;
    XRAM[41375] = 8'b0;
    XRAM[41376] = 8'b0;
    XRAM[41377] = 8'b0;
    XRAM[41378] = 8'b0;
    XRAM[41379] = 8'b0;
    XRAM[41380] = 8'b0;
    XRAM[41381] = 8'b0;
    XRAM[41382] = 8'b0;
    XRAM[41383] = 8'b0;
    XRAM[41384] = 8'b0;
    XRAM[41385] = 8'b0;
    XRAM[41386] = 8'b0;
    XRAM[41387] = 8'b0;
    XRAM[41388] = 8'b0;
    XRAM[41389] = 8'b0;
    XRAM[41390] = 8'b0;
    XRAM[41391] = 8'b0;
    XRAM[41392] = 8'b0;
    XRAM[41393] = 8'b0;
    XRAM[41394] = 8'b0;
    XRAM[41395] = 8'b0;
    XRAM[41396] = 8'b0;
    XRAM[41397] = 8'b0;
    XRAM[41398] = 8'b0;
    XRAM[41399] = 8'b0;
    XRAM[41400] = 8'b0;
    XRAM[41401] = 8'b0;
    XRAM[41402] = 8'b0;
    XRAM[41403] = 8'b0;
    XRAM[41404] = 8'b0;
    XRAM[41405] = 8'b0;
    XRAM[41406] = 8'b0;
    XRAM[41407] = 8'b0;
    XRAM[41408] = 8'b0;
    XRAM[41409] = 8'b0;
    XRAM[41410] = 8'b0;
    XRAM[41411] = 8'b0;
    XRAM[41412] = 8'b0;
    XRAM[41413] = 8'b0;
    XRAM[41414] = 8'b0;
    XRAM[41415] = 8'b0;
    XRAM[41416] = 8'b0;
    XRAM[41417] = 8'b0;
    XRAM[41418] = 8'b0;
    XRAM[41419] = 8'b0;
    XRAM[41420] = 8'b0;
    XRAM[41421] = 8'b0;
    XRAM[41422] = 8'b0;
    XRAM[41423] = 8'b0;
    XRAM[41424] = 8'b0;
    XRAM[41425] = 8'b0;
    XRAM[41426] = 8'b0;
    XRAM[41427] = 8'b0;
    XRAM[41428] = 8'b0;
    XRAM[41429] = 8'b0;
    XRAM[41430] = 8'b0;
    XRAM[41431] = 8'b0;
    XRAM[41432] = 8'b0;
    XRAM[41433] = 8'b0;
    XRAM[41434] = 8'b0;
    XRAM[41435] = 8'b0;
    XRAM[41436] = 8'b0;
    XRAM[41437] = 8'b0;
    XRAM[41438] = 8'b0;
    XRAM[41439] = 8'b0;
    XRAM[41440] = 8'b0;
    XRAM[41441] = 8'b0;
    XRAM[41442] = 8'b0;
    XRAM[41443] = 8'b0;
    XRAM[41444] = 8'b0;
    XRAM[41445] = 8'b0;
    XRAM[41446] = 8'b0;
    XRAM[41447] = 8'b0;
    XRAM[41448] = 8'b0;
    XRAM[41449] = 8'b0;
    XRAM[41450] = 8'b0;
    XRAM[41451] = 8'b0;
    XRAM[41452] = 8'b0;
    XRAM[41453] = 8'b0;
    XRAM[41454] = 8'b0;
    XRAM[41455] = 8'b0;
    XRAM[41456] = 8'b0;
    XRAM[41457] = 8'b0;
    XRAM[41458] = 8'b0;
    XRAM[41459] = 8'b0;
    XRAM[41460] = 8'b0;
    XRAM[41461] = 8'b0;
    XRAM[41462] = 8'b0;
    XRAM[41463] = 8'b0;
    XRAM[41464] = 8'b0;
    XRAM[41465] = 8'b0;
    XRAM[41466] = 8'b0;
    XRAM[41467] = 8'b0;
    XRAM[41468] = 8'b0;
    XRAM[41469] = 8'b0;
    XRAM[41470] = 8'b0;
    XRAM[41471] = 8'b0;
    XRAM[41472] = 8'b0;
    XRAM[41473] = 8'b0;
    XRAM[41474] = 8'b0;
    XRAM[41475] = 8'b0;
    XRAM[41476] = 8'b0;
    XRAM[41477] = 8'b0;
    XRAM[41478] = 8'b0;
    XRAM[41479] = 8'b0;
    XRAM[41480] = 8'b0;
    XRAM[41481] = 8'b0;
    XRAM[41482] = 8'b0;
    XRAM[41483] = 8'b0;
    XRAM[41484] = 8'b0;
    XRAM[41485] = 8'b0;
    XRAM[41486] = 8'b0;
    XRAM[41487] = 8'b0;
    XRAM[41488] = 8'b0;
    XRAM[41489] = 8'b0;
    XRAM[41490] = 8'b0;
    XRAM[41491] = 8'b0;
    XRAM[41492] = 8'b0;
    XRAM[41493] = 8'b0;
    XRAM[41494] = 8'b0;
    XRAM[41495] = 8'b0;
    XRAM[41496] = 8'b0;
    XRAM[41497] = 8'b0;
    XRAM[41498] = 8'b0;
    XRAM[41499] = 8'b0;
    XRAM[41500] = 8'b0;
    XRAM[41501] = 8'b0;
    XRAM[41502] = 8'b0;
    XRAM[41503] = 8'b0;
    XRAM[41504] = 8'b0;
    XRAM[41505] = 8'b0;
    XRAM[41506] = 8'b0;
    XRAM[41507] = 8'b0;
    XRAM[41508] = 8'b0;
    XRAM[41509] = 8'b0;
    XRAM[41510] = 8'b0;
    XRAM[41511] = 8'b0;
    XRAM[41512] = 8'b0;
    XRAM[41513] = 8'b0;
    XRAM[41514] = 8'b0;
    XRAM[41515] = 8'b0;
    XRAM[41516] = 8'b0;
    XRAM[41517] = 8'b0;
    XRAM[41518] = 8'b0;
    XRAM[41519] = 8'b0;
    XRAM[41520] = 8'b0;
    XRAM[41521] = 8'b0;
    XRAM[41522] = 8'b0;
    XRAM[41523] = 8'b0;
    XRAM[41524] = 8'b0;
    XRAM[41525] = 8'b0;
    XRAM[41526] = 8'b0;
    XRAM[41527] = 8'b0;
    XRAM[41528] = 8'b0;
    XRAM[41529] = 8'b0;
    XRAM[41530] = 8'b0;
    XRAM[41531] = 8'b0;
    XRAM[41532] = 8'b0;
    XRAM[41533] = 8'b0;
    XRAM[41534] = 8'b0;
    XRAM[41535] = 8'b0;
    XRAM[41536] = 8'b0;
    XRAM[41537] = 8'b0;
    XRAM[41538] = 8'b0;
    XRAM[41539] = 8'b0;
    XRAM[41540] = 8'b0;
    XRAM[41541] = 8'b0;
    XRAM[41542] = 8'b0;
    XRAM[41543] = 8'b0;
    XRAM[41544] = 8'b0;
    XRAM[41545] = 8'b0;
    XRAM[41546] = 8'b0;
    XRAM[41547] = 8'b0;
    XRAM[41548] = 8'b0;
    XRAM[41549] = 8'b0;
    XRAM[41550] = 8'b0;
    XRAM[41551] = 8'b0;
    XRAM[41552] = 8'b0;
    XRAM[41553] = 8'b0;
    XRAM[41554] = 8'b0;
    XRAM[41555] = 8'b0;
    XRAM[41556] = 8'b0;
    XRAM[41557] = 8'b0;
    XRAM[41558] = 8'b0;
    XRAM[41559] = 8'b0;
    XRAM[41560] = 8'b0;
    XRAM[41561] = 8'b0;
    XRAM[41562] = 8'b0;
    XRAM[41563] = 8'b0;
    XRAM[41564] = 8'b0;
    XRAM[41565] = 8'b0;
    XRAM[41566] = 8'b0;
    XRAM[41567] = 8'b0;
    XRAM[41568] = 8'b0;
    XRAM[41569] = 8'b0;
    XRAM[41570] = 8'b0;
    XRAM[41571] = 8'b0;
    XRAM[41572] = 8'b0;
    XRAM[41573] = 8'b0;
    XRAM[41574] = 8'b0;
    XRAM[41575] = 8'b0;
    XRAM[41576] = 8'b0;
    XRAM[41577] = 8'b0;
    XRAM[41578] = 8'b0;
    XRAM[41579] = 8'b0;
    XRAM[41580] = 8'b0;
    XRAM[41581] = 8'b0;
    XRAM[41582] = 8'b0;
    XRAM[41583] = 8'b0;
    XRAM[41584] = 8'b0;
    XRAM[41585] = 8'b0;
    XRAM[41586] = 8'b0;
    XRAM[41587] = 8'b0;
    XRAM[41588] = 8'b0;
    XRAM[41589] = 8'b0;
    XRAM[41590] = 8'b0;
    XRAM[41591] = 8'b0;
    XRAM[41592] = 8'b0;
    XRAM[41593] = 8'b0;
    XRAM[41594] = 8'b0;
    XRAM[41595] = 8'b0;
    XRAM[41596] = 8'b0;
    XRAM[41597] = 8'b0;
    XRAM[41598] = 8'b0;
    XRAM[41599] = 8'b0;
    XRAM[41600] = 8'b0;
    XRAM[41601] = 8'b0;
    XRAM[41602] = 8'b0;
    XRAM[41603] = 8'b0;
    XRAM[41604] = 8'b0;
    XRAM[41605] = 8'b0;
    XRAM[41606] = 8'b0;
    XRAM[41607] = 8'b0;
    XRAM[41608] = 8'b0;
    XRAM[41609] = 8'b0;
    XRAM[41610] = 8'b0;
    XRAM[41611] = 8'b0;
    XRAM[41612] = 8'b0;
    XRAM[41613] = 8'b0;
    XRAM[41614] = 8'b0;
    XRAM[41615] = 8'b0;
    XRAM[41616] = 8'b0;
    XRAM[41617] = 8'b0;
    XRAM[41618] = 8'b0;
    XRAM[41619] = 8'b0;
    XRAM[41620] = 8'b0;
    XRAM[41621] = 8'b0;
    XRAM[41622] = 8'b0;
    XRAM[41623] = 8'b0;
    XRAM[41624] = 8'b0;
    XRAM[41625] = 8'b0;
    XRAM[41626] = 8'b0;
    XRAM[41627] = 8'b0;
    XRAM[41628] = 8'b0;
    XRAM[41629] = 8'b0;
    XRAM[41630] = 8'b0;
    XRAM[41631] = 8'b0;
    XRAM[41632] = 8'b0;
    XRAM[41633] = 8'b0;
    XRAM[41634] = 8'b0;
    XRAM[41635] = 8'b0;
    XRAM[41636] = 8'b0;
    XRAM[41637] = 8'b0;
    XRAM[41638] = 8'b0;
    XRAM[41639] = 8'b0;
    XRAM[41640] = 8'b0;
    XRAM[41641] = 8'b0;
    XRAM[41642] = 8'b0;
    XRAM[41643] = 8'b0;
    XRAM[41644] = 8'b0;
    XRAM[41645] = 8'b0;
    XRAM[41646] = 8'b0;
    XRAM[41647] = 8'b0;
    XRAM[41648] = 8'b0;
    XRAM[41649] = 8'b0;
    XRAM[41650] = 8'b0;
    XRAM[41651] = 8'b0;
    XRAM[41652] = 8'b0;
    XRAM[41653] = 8'b0;
    XRAM[41654] = 8'b0;
    XRAM[41655] = 8'b0;
    XRAM[41656] = 8'b0;
    XRAM[41657] = 8'b0;
    XRAM[41658] = 8'b0;
    XRAM[41659] = 8'b0;
    XRAM[41660] = 8'b0;
    XRAM[41661] = 8'b0;
    XRAM[41662] = 8'b0;
    XRAM[41663] = 8'b0;
    XRAM[41664] = 8'b0;
    XRAM[41665] = 8'b0;
    XRAM[41666] = 8'b0;
    XRAM[41667] = 8'b0;
    XRAM[41668] = 8'b0;
    XRAM[41669] = 8'b0;
    XRAM[41670] = 8'b0;
    XRAM[41671] = 8'b0;
    XRAM[41672] = 8'b0;
    XRAM[41673] = 8'b0;
    XRAM[41674] = 8'b0;
    XRAM[41675] = 8'b0;
    XRAM[41676] = 8'b0;
    XRAM[41677] = 8'b0;
    XRAM[41678] = 8'b0;
    XRAM[41679] = 8'b0;
    XRAM[41680] = 8'b0;
    XRAM[41681] = 8'b0;
    XRAM[41682] = 8'b0;
    XRAM[41683] = 8'b0;
    XRAM[41684] = 8'b0;
    XRAM[41685] = 8'b0;
    XRAM[41686] = 8'b0;
    XRAM[41687] = 8'b0;
    XRAM[41688] = 8'b0;
    XRAM[41689] = 8'b0;
    XRAM[41690] = 8'b0;
    XRAM[41691] = 8'b0;
    XRAM[41692] = 8'b0;
    XRAM[41693] = 8'b0;
    XRAM[41694] = 8'b0;
    XRAM[41695] = 8'b0;
    XRAM[41696] = 8'b0;
    XRAM[41697] = 8'b0;
    XRAM[41698] = 8'b0;
    XRAM[41699] = 8'b0;
    XRAM[41700] = 8'b0;
    XRAM[41701] = 8'b0;
    XRAM[41702] = 8'b0;
    XRAM[41703] = 8'b0;
    XRAM[41704] = 8'b0;
    XRAM[41705] = 8'b0;
    XRAM[41706] = 8'b0;
    XRAM[41707] = 8'b0;
    XRAM[41708] = 8'b0;
    XRAM[41709] = 8'b0;
    XRAM[41710] = 8'b0;
    XRAM[41711] = 8'b0;
    XRAM[41712] = 8'b0;
    XRAM[41713] = 8'b0;
    XRAM[41714] = 8'b0;
    XRAM[41715] = 8'b0;
    XRAM[41716] = 8'b0;
    XRAM[41717] = 8'b0;
    XRAM[41718] = 8'b0;
    XRAM[41719] = 8'b0;
    XRAM[41720] = 8'b0;
    XRAM[41721] = 8'b0;
    XRAM[41722] = 8'b0;
    XRAM[41723] = 8'b0;
    XRAM[41724] = 8'b0;
    XRAM[41725] = 8'b0;
    XRAM[41726] = 8'b0;
    XRAM[41727] = 8'b0;
    XRAM[41728] = 8'b0;
    XRAM[41729] = 8'b0;
    XRAM[41730] = 8'b0;
    XRAM[41731] = 8'b0;
    XRAM[41732] = 8'b0;
    XRAM[41733] = 8'b0;
    XRAM[41734] = 8'b0;
    XRAM[41735] = 8'b0;
    XRAM[41736] = 8'b0;
    XRAM[41737] = 8'b0;
    XRAM[41738] = 8'b0;
    XRAM[41739] = 8'b0;
    XRAM[41740] = 8'b0;
    XRAM[41741] = 8'b0;
    XRAM[41742] = 8'b0;
    XRAM[41743] = 8'b0;
    XRAM[41744] = 8'b0;
    XRAM[41745] = 8'b0;
    XRAM[41746] = 8'b0;
    XRAM[41747] = 8'b0;
    XRAM[41748] = 8'b0;
    XRAM[41749] = 8'b0;
    XRAM[41750] = 8'b0;
    XRAM[41751] = 8'b0;
    XRAM[41752] = 8'b0;
    XRAM[41753] = 8'b0;
    XRAM[41754] = 8'b0;
    XRAM[41755] = 8'b0;
    XRAM[41756] = 8'b0;
    XRAM[41757] = 8'b0;
    XRAM[41758] = 8'b0;
    XRAM[41759] = 8'b0;
    XRAM[41760] = 8'b0;
    XRAM[41761] = 8'b0;
    XRAM[41762] = 8'b0;
    XRAM[41763] = 8'b0;
    XRAM[41764] = 8'b0;
    XRAM[41765] = 8'b0;
    XRAM[41766] = 8'b0;
    XRAM[41767] = 8'b0;
    XRAM[41768] = 8'b0;
    XRAM[41769] = 8'b0;
    XRAM[41770] = 8'b0;
    XRAM[41771] = 8'b0;
    XRAM[41772] = 8'b0;
    XRAM[41773] = 8'b0;
    XRAM[41774] = 8'b0;
    XRAM[41775] = 8'b0;
    XRAM[41776] = 8'b0;
    XRAM[41777] = 8'b0;
    XRAM[41778] = 8'b0;
    XRAM[41779] = 8'b0;
    XRAM[41780] = 8'b0;
    XRAM[41781] = 8'b0;
    XRAM[41782] = 8'b0;
    XRAM[41783] = 8'b0;
    XRAM[41784] = 8'b0;
    XRAM[41785] = 8'b0;
    XRAM[41786] = 8'b0;
    XRAM[41787] = 8'b0;
    XRAM[41788] = 8'b0;
    XRAM[41789] = 8'b0;
    XRAM[41790] = 8'b0;
    XRAM[41791] = 8'b0;
    XRAM[41792] = 8'b0;
    XRAM[41793] = 8'b0;
    XRAM[41794] = 8'b0;
    XRAM[41795] = 8'b0;
    XRAM[41796] = 8'b0;
    XRAM[41797] = 8'b0;
    XRAM[41798] = 8'b0;
    XRAM[41799] = 8'b0;
    XRAM[41800] = 8'b0;
    XRAM[41801] = 8'b0;
    XRAM[41802] = 8'b0;
    XRAM[41803] = 8'b0;
    XRAM[41804] = 8'b0;
    XRAM[41805] = 8'b0;
    XRAM[41806] = 8'b0;
    XRAM[41807] = 8'b0;
    XRAM[41808] = 8'b0;
    XRAM[41809] = 8'b0;
    XRAM[41810] = 8'b0;
    XRAM[41811] = 8'b0;
    XRAM[41812] = 8'b0;
    XRAM[41813] = 8'b0;
    XRAM[41814] = 8'b0;
    XRAM[41815] = 8'b0;
    XRAM[41816] = 8'b0;
    XRAM[41817] = 8'b0;
    XRAM[41818] = 8'b0;
    XRAM[41819] = 8'b0;
    XRAM[41820] = 8'b0;
    XRAM[41821] = 8'b0;
    XRAM[41822] = 8'b0;
    XRAM[41823] = 8'b0;
    XRAM[41824] = 8'b0;
    XRAM[41825] = 8'b0;
    XRAM[41826] = 8'b0;
    XRAM[41827] = 8'b0;
    XRAM[41828] = 8'b0;
    XRAM[41829] = 8'b0;
    XRAM[41830] = 8'b0;
    XRAM[41831] = 8'b0;
    XRAM[41832] = 8'b0;
    XRAM[41833] = 8'b0;
    XRAM[41834] = 8'b0;
    XRAM[41835] = 8'b0;
    XRAM[41836] = 8'b0;
    XRAM[41837] = 8'b0;
    XRAM[41838] = 8'b0;
    XRAM[41839] = 8'b0;
    XRAM[41840] = 8'b0;
    XRAM[41841] = 8'b0;
    XRAM[41842] = 8'b0;
    XRAM[41843] = 8'b0;
    XRAM[41844] = 8'b0;
    XRAM[41845] = 8'b0;
    XRAM[41846] = 8'b0;
    XRAM[41847] = 8'b0;
    XRAM[41848] = 8'b0;
    XRAM[41849] = 8'b0;
    XRAM[41850] = 8'b0;
    XRAM[41851] = 8'b0;
    XRAM[41852] = 8'b0;
    XRAM[41853] = 8'b0;
    XRAM[41854] = 8'b0;
    XRAM[41855] = 8'b0;
    XRAM[41856] = 8'b0;
    XRAM[41857] = 8'b0;
    XRAM[41858] = 8'b0;
    XRAM[41859] = 8'b0;
    XRAM[41860] = 8'b0;
    XRAM[41861] = 8'b0;
    XRAM[41862] = 8'b0;
    XRAM[41863] = 8'b0;
    XRAM[41864] = 8'b0;
    XRAM[41865] = 8'b0;
    XRAM[41866] = 8'b0;
    XRAM[41867] = 8'b0;
    XRAM[41868] = 8'b0;
    XRAM[41869] = 8'b0;
    XRAM[41870] = 8'b0;
    XRAM[41871] = 8'b0;
    XRAM[41872] = 8'b0;
    XRAM[41873] = 8'b0;
    XRAM[41874] = 8'b0;
    XRAM[41875] = 8'b0;
    XRAM[41876] = 8'b0;
    XRAM[41877] = 8'b0;
    XRAM[41878] = 8'b0;
    XRAM[41879] = 8'b0;
    XRAM[41880] = 8'b0;
    XRAM[41881] = 8'b0;
    XRAM[41882] = 8'b0;
    XRAM[41883] = 8'b0;
    XRAM[41884] = 8'b0;
    XRAM[41885] = 8'b0;
    XRAM[41886] = 8'b0;
    XRAM[41887] = 8'b0;
    XRAM[41888] = 8'b0;
    XRAM[41889] = 8'b0;
    XRAM[41890] = 8'b0;
    XRAM[41891] = 8'b0;
    XRAM[41892] = 8'b0;
    XRAM[41893] = 8'b0;
    XRAM[41894] = 8'b0;
    XRAM[41895] = 8'b0;
    XRAM[41896] = 8'b0;
    XRAM[41897] = 8'b0;
    XRAM[41898] = 8'b0;
    XRAM[41899] = 8'b0;
    XRAM[41900] = 8'b0;
    XRAM[41901] = 8'b0;
    XRAM[41902] = 8'b0;
    XRAM[41903] = 8'b0;
    XRAM[41904] = 8'b0;
    XRAM[41905] = 8'b0;
    XRAM[41906] = 8'b0;
    XRAM[41907] = 8'b0;
    XRAM[41908] = 8'b0;
    XRAM[41909] = 8'b0;
    XRAM[41910] = 8'b0;
    XRAM[41911] = 8'b0;
    XRAM[41912] = 8'b0;
    XRAM[41913] = 8'b0;
    XRAM[41914] = 8'b0;
    XRAM[41915] = 8'b0;
    XRAM[41916] = 8'b0;
    XRAM[41917] = 8'b0;
    XRAM[41918] = 8'b0;
    XRAM[41919] = 8'b0;
    XRAM[41920] = 8'b0;
    XRAM[41921] = 8'b0;
    XRAM[41922] = 8'b0;
    XRAM[41923] = 8'b0;
    XRAM[41924] = 8'b0;
    XRAM[41925] = 8'b0;
    XRAM[41926] = 8'b0;
    XRAM[41927] = 8'b0;
    XRAM[41928] = 8'b0;
    XRAM[41929] = 8'b0;
    XRAM[41930] = 8'b0;
    XRAM[41931] = 8'b0;
    XRAM[41932] = 8'b0;
    XRAM[41933] = 8'b0;
    XRAM[41934] = 8'b0;
    XRAM[41935] = 8'b0;
    XRAM[41936] = 8'b0;
    XRAM[41937] = 8'b0;
    XRAM[41938] = 8'b0;
    XRAM[41939] = 8'b0;
    XRAM[41940] = 8'b0;
    XRAM[41941] = 8'b0;
    XRAM[41942] = 8'b0;
    XRAM[41943] = 8'b0;
    XRAM[41944] = 8'b0;
    XRAM[41945] = 8'b0;
    XRAM[41946] = 8'b0;
    XRAM[41947] = 8'b0;
    XRAM[41948] = 8'b0;
    XRAM[41949] = 8'b0;
    XRAM[41950] = 8'b0;
    XRAM[41951] = 8'b0;
    XRAM[41952] = 8'b0;
    XRAM[41953] = 8'b0;
    XRAM[41954] = 8'b0;
    XRAM[41955] = 8'b0;
    XRAM[41956] = 8'b0;
    XRAM[41957] = 8'b0;
    XRAM[41958] = 8'b0;
    XRAM[41959] = 8'b0;
    XRAM[41960] = 8'b0;
    XRAM[41961] = 8'b0;
    XRAM[41962] = 8'b0;
    XRAM[41963] = 8'b0;
    XRAM[41964] = 8'b0;
    XRAM[41965] = 8'b0;
    XRAM[41966] = 8'b0;
    XRAM[41967] = 8'b0;
    XRAM[41968] = 8'b0;
    XRAM[41969] = 8'b0;
    XRAM[41970] = 8'b0;
    XRAM[41971] = 8'b0;
    XRAM[41972] = 8'b0;
    XRAM[41973] = 8'b0;
    XRAM[41974] = 8'b0;
    XRAM[41975] = 8'b0;
    XRAM[41976] = 8'b0;
    XRAM[41977] = 8'b0;
    XRAM[41978] = 8'b0;
    XRAM[41979] = 8'b0;
    XRAM[41980] = 8'b0;
    XRAM[41981] = 8'b0;
    XRAM[41982] = 8'b0;
    XRAM[41983] = 8'b0;
    XRAM[41984] = 8'b0;
    XRAM[41985] = 8'b0;
    XRAM[41986] = 8'b0;
    XRAM[41987] = 8'b0;
    XRAM[41988] = 8'b0;
    XRAM[41989] = 8'b0;
    XRAM[41990] = 8'b0;
    XRAM[41991] = 8'b0;
    XRAM[41992] = 8'b0;
    XRAM[41993] = 8'b0;
    XRAM[41994] = 8'b0;
    XRAM[41995] = 8'b0;
    XRAM[41996] = 8'b0;
    XRAM[41997] = 8'b0;
    XRAM[41998] = 8'b0;
    XRAM[41999] = 8'b0;
    XRAM[42000] = 8'b0;
    XRAM[42001] = 8'b0;
    XRAM[42002] = 8'b0;
    XRAM[42003] = 8'b0;
    XRAM[42004] = 8'b0;
    XRAM[42005] = 8'b0;
    XRAM[42006] = 8'b0;
    XRAM[42007] = 8'b0;
    XRAM[42008] = 8'b0;
    XRAM[42009] = 8'b0;
    XRAM[42010] = 8'b0;
    XRAM[42011] = 8'b0;
    XRAM[42012] = 8'b0;
    XRAM[42013] = 8'b0;
    XRAM[42014] = 8'b0;
    XRAM[42015] = 8'b0;
    XRAM[42016] = 8'b0;
    XRAM[42017] = 8'b0;
    XRAM[42018] = 8'b0;
    XRAM[42019] = 8'b0;
    XRAM[42020] = 8'b0;
    XRAM[42021] = 8'b0;
    XRAM[42022] = 8'b0;
    XRAM[42023] = 8'b0;
    XRAM[42024] = 8'b0;
    XRAM[42025] = 8'b0;
    XRAM[42026] = 8'b0;
    XRAM[42027] = 8'b0;
    XRAM[42028] = 8'b0;
    XRAM[42029] = 8'b0;
    XRAM[42030] = 8'b0;
    XRAM[42031] = 8'b0;
    XRAM[42032] = 8'b0;
    XRAM[42033] = 8'b0;
    XRAM[42034] = 8'b0;
    XRAM[42035] = 8'b0;
    XRAM[42036] = 8'b0;
    XRAM[42037] = 8'b0;
    XRAM[42038] = 8'b0;
    XRAM[42039] = 8'b0;
    XRAM[42040] = 8'b0;
    XRAM[42041] = 8'b0;
    XRAM[42042] = 8'b0;
    XRAM[42043] = 8'b0;
    XRAM[42044] = 8'b0;
    XRAM[42045] = 8'b0;
    XRAM[42046] = 8'b0;
    XRAM[42047] = 8'b0;
    XRAM[42048] = 8'b0;
    XRAM[42049] = 8'b0;
    XRAM[42050] = 8'b0;
    XRAM[42051] = 8'b0;
    XRAM[42052] = 8'b0;
    XRAM[42053] = 8'b0;
    XRAM[42054] = 8'b0;
    XRAM[42055] = 8'b0;
    XRAM[42056] = 8'b0;
    XRAM[42057] = 8'b0;
    XRAM[42058] = 8'b0;
    XRAM[42059] = 8'b0;
    XRAM[42060] = 8'b0;
    XRAM[42061] = 8'b0;
    XRAM[42062] = 8'b0;
    XRAM[42063] = 8'b0;
    XRAM[42064] = 8'b0;
    XRAM[42065] = 8'b0;
    XRAM[42066] = 8'b0;
    XRAM[42067] = 8'b0;
    XRAM[42068] = 8'b0;
    XRAM[42069] = 8'b0;
    XRAM[42070] = 8'b0;
    XRAM[42071] = 8'b0;
    XRAM[42072] = 8'b0;
    XRAM[42073] = 8'b0;
    XRAM[42074] = 8'b0;
    XRAM[42075] = 8'b0;
    XRAM[42076] = 8'b0;
    XRAM[42077] = 8'b0;
    XRAM[42078] = 8'b0;
    XRAM[42079] = 8'b0;
    XRAM[42080] = 8'b0;
    XRAM[42081] = 8'b0;
    XRAM[42082] = 8'b0;
    XRAM[42083] = 8'b0;
    XRAM[42084] = 8'b0;
    XRAM[42085] = 8'b0;
    XRAM[42086] = 8'b0;
    XRAM[42087] = 8'b0;
    XRAM[42088] = 8'b0;
    XRAM[42089] = 8'b0;
    XRAM[42090] = 8'b0;
    XRAM[42091] = 8'b0;
    XRAM[42092] = 8'b0;
    XRAM[42093] = 8'b0;
    XRAM[42094] = 8'b0;
    XRAM[42095] = 8'b0;
    XRAM[42096] = 8'b0;
    XRAM[42097] = 8'b0;
    XRAM[42098] = 8'b0;
    XRAM[42099] = 8'b0;
    XRAM[42100] = 8'b0;
    XRAM[42101] = 8'b0;
    XRAM[42102] = 8'b0;
    XRAM[42103] = 8'b0;
    XRAM[42104] = 8'b0;
    XRAM[42105] = 8'b0;
    XRAM[42106] = 8'b0;
    XRAM[42107] = 8'b0;
    XRAM[42108] = 8'b0;
    XRAM[42109] = 8'b0;
    XRAM[42110] = 8'b0;
    XRAM[42111] = 8'b0;
    XRAM[42112] = 8'b0;
    XRAM[42113] = 8'b0;
    XRAM[42114] = 8'b0;
    XRAM[42115] = 8'b0;
    XRAM[42116] = 8'b0;
    XRAM[42117] = 8'b0;
    XRAM[42118] = 8'b0;
    XRAM[42119] = 8'b0;
    XRAM[42120] = 8'b0;
    XRAM[42121] = 8'b0;
    XRAM[42122] = 8'b0;
    XRAM[42123] = 8'b0;
    XRAM[42124] = 8'b0;
    XRAM[42125] = 8'b0;
    XRAM[42126] = 8'b0;
    XRAM[42127] = 8'b0;
    XRAM[42128] = 8'b0;
    XRAM[42129] = 8'b0;
    XRAM[42130] = 8'b0;
    XRAM[42131] = 8'b0;
    XRAM[42132] = 8'b0;
    XRAM[42133] = 8'b0;
    XRAM[42134] = 8'b0;
    XRAM[42135] = 8'b0;
    XRAM[42136] = 8'b0;
    XRAM[42137] = 8'b0;
    XRAM[42138] = 8'b0;
    XRAM[42139] = 8'b0;
    XRAM[42140] = 8'b0;
    XRAM[42141] = 8'b0;
    XRAM[42142] = 8'b0;
    XRAM[42143] = 8'b0;
    XRAM[42144] = 8'b0;
    XRAM[42145] = 8'b0;
    XRAM[42146] = 8'b0;
    XRAM[42147] = 8'b0;
    XRAM[42148] = 8'b0;
    XRAM[42149] = 8'b0;
    XRAM[42150] = 8'b0;
    XRAM[42151] = 8'b0;
    XRAM[42152] = 8'b0;
    XRAM[42153] = 8'b0;
    XRAM[42154] = 8'b0;
    XRAM[42155] = 8'b0;
    XRAM[42156] = 8'b0;
    XRAM[42157] = 8'b0;
    XRAM[42158] = 8'b0;
    XRAM[42159] = 8'b0;
    XRAM[42160] = 8'b0;
    XRAM[42161] = 8'b0;
    XRAM[42162] = 8'b0;
    XRAM[42163] = 8'b0;
    XRAM[42164] = 8'b0;
    XRAM[42165] = 8'b0;
    XRAM[42166] = 8'b0;
    XRAM[42167] = 8'b0;
    XRAM[42168] = 8'b0;
    XRAM[42169] = 8'b0;
    XRAM[42170] = 8'b0;
    XRAM[42171] = 8'b0;
    XRAM[42172] = 8'b0;
    XRAM[42173] = 8'b0;
    XRAM[42174] = 8'b0;
    XRAM[42175] = 8'b0;
    XRAM[42176] = 8'b0;
    XRAM[42177] = 8'b0;
    XRAM[42178] = 8'b0;
    XRAM[42179] = 8'b0;
    XRAM[42180] = 8'b0;
    XRAM[42181] = 8'b0;
    XRAM[42182] = 8'b0;
    XRAM[42183] = 8'b0;
    XRAM[42184] = 8'b0;
    XRAM[42185] = 8'b0;
    XRAM[42186] = 8'b0;
    XRAM[42187] = 8'b0;
    XRAM[42188] = 8'b0;
    XRAM[42189] = 8'b0;
    XRAM[42190] = 8'b0;
    XRAM[42191] = 8'b0;
    XRAM[42192] = 8'b0;
    XRAM[42193] = 8'b0;
    XRAM[42194] = 8'b0;
    XRAM[42195] = 8'b0;
    XRAM[42196] = 8'b0;
    XRAM[42197] = 8'b0;
    XRAM[42198] = 8'b0;
    XRAM[42199] = 8'b0;
    XRAM[42200] = 8'b0;
    XRAM[42201] = 8'b0;
    XRAM[42202] = 8'b0;
    XRAM[42203] = 8'b0;
    XRAM[42204] = 8'b0;
    XRAM[42205] = 8'b0;
    XRAM[42206] = 8'b0;
    XRAM[42207] = 8'b0;
    XRAM[42208] = 8'b0;
    XRAM[42209] = 8'b0;
    XRAM[42210] = 8'b0;
    XRAM[42211] = 8'b0;
    XRAM[42212] = 8'b0;
    XRAM[42213] = 8'b0;
    XRAM[42214] = 8'b0;
    XRAM[42215] = 8'b0;
    XRAM[42216] = 8'b0;
    XRAM[42217] = 8'b0;
    XRAM[42218] = 8'b0;
    XRAM[42219] = 8'b0;
    XRAM[42220] = 8'b0;
    XRAM[42221] = 8'b0;
    XRAM[42222] = 8'b0;
    XRAM[42223] = 8'b0;
    XRAM[42224] = 8'b0;
    XRAM[42225] = 8'b0;
    XRAM[42226] = 8'b0;
    XRAM[42227] = 8'b0;
    XRAM[42228] = 8'b0;
    XRAM[42229] = 8'b0;
    XRAM[42230] = 8'b0;
    XRAM[42231] = 8'b0;
    XRAM[42232] = 8'b0;
    XRAM[42233] = 8'b0;
    XRAM[42234] = 8'b0;
    XRAM[42235] = 8'b0;
    XRAM[42236] = 8'b0;
    XRAM[42237] = 8'b0;
    XRAM[42238] = 8'b0;
    XRAM[42239] = 8'b0;
    XRAM[42240] = 8'b0;
    XRAM[42241] = 8'b0;
    XRAM[42242] = 8'b0;
    XRAM[42243] = 8'b0;
    XRAM[42244] = 8'b0;
    XRAM[42245] = 8'b0;
    XRAM[42246] = 8'b0;
    XRAM[42247] = 8'b0;
    XRAM[42248] = 8'b0;
    XRAM[42249] = 8'b0;
    XRAM[42250] = 8'b0;
    XRAM[42251] = 8'b0;
    XRAM[42252] = 8'b0;
    XRAM[42253] = 8'b0;
    XRAM[42254] = 8'b0;
    XRAM[42255] = 8'b0;
    XRAM[42256] = 8'b0;
    XRAM[42257] = 8'b0;
    XRAM[42258] = 8'b0;
    XRAM[42259] = 8'b0;
    XRAM[42260] = 8'b0;
    XRAM[42261] = 8'b0;
    XRAM[42262] = 8'b0;
    XRAM[42263] = 8'b0;
    XRAM[42264] = 8'b0;
    XRAM[42265] = 8'b0;
    XRAM[42266] = 8'b0;
    XRAM[42267] = 8'b0;
    XRAM[42268] = 8'b0;
    XRAM[42269] = 8'b0;
    XRAM[42270] = 8'b0;
    XRAM[42271] = 8'b0;
    XRAM[42272] = 8'b0;
    XRAM[42273] = 8'b0;
    XRAM[42274] = 8'b0;
    XRAM[42275] = 8'b0;
    XRAM[42276] = 8'b0;
    XRAM[42277] = 8'b0;
    XRAM[42278] = 8'b0;
    XRAM[42279] = 8'b0;
    XRAM[42280] = 8'b0;
    XRAM[42281] = 8'b0;
    XRAM[42282] = 8'b0;
    XRAM[42283] = 8'b0;
    XRAM[42284] = 8'b0;
    XRAM[42285] = 8'b0;
    XRAM[42286] = 8'b0;
    XRAM[42287] = 8'b0;
    XRAM[42288] = 8'b0;
    XRAM[42289] = 8'b0;
    XRAM[42290] = 8'b0;
    XRAM[42291] = 8'b0;
    XRAM[42292] = 8'b0;
    XRAM[42293] = 8'b0;
    XRAM[42294] = 8'b0;
    XRAM[42295] = 8'b0;
    XRAM[42296] = 8'b0;
    XRAM[42297] = 8'b0;
    XRAM[42298] = 8'b0;
    XRAM[42299] = 8'b0;
    XRAM[42300] = 8'b0;
    XRAM[42301] = 8'b0;
    XRAM[42302] = 8'b0;
    XRAM[42303] = 8'b0;
    XRAM[42304] = 8'b0;
    XRAM[42305] = 8'b0;
    XRAM[42306] = 8'b0;
    XRAM[42307] = 8'b0;
    XRAM[42308] = 8'b0;
    XRAM[42309] = 8'b0;
    XRAM[42310] = 8'b0;
    XRAM[42311] = 8'b0;
    XRAM[42312] = 8'b0;
    XRAM[42313] = 8'b0;
    XRAM[42314] = 8'b0;
    XRAM[42315] = 8'b0;
    XRAM[42316] = 8'b0;
    XRAM[42317] = 8'b0;
    XRAM[42318] = 8'b0;
    XRAM[42319] = 8'b0;
    XRAM[42320] = 8'b0;
    XRAM[42321] = 8'b0;
    XRAM[42322] = 8'b0;
    XRAM[42323] = 8'b0;
    XRAM[42324] = 8'b0;
    XRAM[42325] = 8'b0;
    XRAM[42326] = 8'b0;
    XRAM[42327] = 8'b0;
    XRAM[42328] = 8'b0;
    XRAM[42329] = 8'b0;
    XRAM[42330] = 8'b0;
    XRAM[42331] = 8'b0;
    XRAM[42332] = 8'b0;
    XRAM[42333] = 8'b0;
    XRAM[42334] = 8'b0;
    XRAM[42335] = 8'b0;
    XRAM[42336] = 8'b0;
    XRAM[42337] = 8'b0;
    XRAM[42338] = 8'b0;
    XRAM[42339] = 8'b0;
    XRAM[42340] = 8'b0;
    XRAM[42341] = 8'b0;
    XRAM[42342] = 8'b0;
    XRAM[42343] = 8'b0;
    XRAM[42344] = 8'b0;
    XRAM[42345] = 8'b0;
    XRAM[42346] = 8'b0;
    XRAM[42347] = 8'b0;
    XRAM[42348] = 8'b0;
    XRAM[42349] = 8'b0;
    XRAM[42350] = 8'b0;
    XRAM[42351] = 8'b0;
    XRAM[42352] = 8'b0;
    XRAM[42353] = 8'b0;
    XRAM[42354] = 8'b0;
    XRAM[42355] = 8'b0;
    XRAM[42356] = 8'b0;
    XRAM[42357] = 8'b0;
    XRAM[42358] = 8'b0;
    XRAM[42359] = 8'b0;
    XRAM[42360] = 8'b0;
    XRAM[42361] = 8'b0;
    XRAM[42362] = 8'b0;
    XRAM[42363] = 8'b0;
    XRAM[42364] = 8'b0;
    XRAM[42365] = 8'b0;
    XRAM[42366] = 8'b0;
    XRAM[42367] = 8'b0;
    XRAM[42368] = 8'b0;
    XRAM[42369] = 8'b0;
    XRAM[42370] = 8'b0;
    XRAM[42371] = 8'b0;
    XRAM[42372] = 8'b0;
    XRAM[42373] = 8'b0;
    XRAM[42374] = 8'b0;
    XRAM[42375] = 8'b0;
    XRAM[42376] = 8'b0;
    XRAM[42377] = 8'b0;
    XRAM[42378] = 8'b0;
    XRAM[42379] = 8'b0;
    XRAM[42380] = 8'b0;
    XRAM[42381] = 8'b0;
    XRAM[42382] = 8'b0;
    XRAM[42383] = 8'b0;
    XRAM[42384] = 8'b0;
    XRAM[42385] = 8'b0;
    XRAM[42386] = 8'b0;
    XRAM[42387] = 8'b0;
    XRAM[42388] = 8'b0;
    XRAM[42389] = 8'b0;
    XRAM[42390] = 8'b0;
    XRAM[42391] = 8'b0;
    XRAM[42392] = 8'b0;
    XRAM[42393] = 8'b0;
    XRAM[42394] = 8'b0;
    XRAM[42395] = 8'b0;
    XRAM[42396] = 8'b0;
    XRAM[42397] = 8'b0;
    XRAM[42398] = 8'b0;
    XRAM[42399] = 8'b0;
    XRAM[42400] = 8'b0;
    XRAM[42401] = 8'b0;
    XRAM[42402] = 8'b0;
    XRAM[42403] = 8'b0;
    XRAM[42404] = 8'b0;
    XRAM[42405] = 8'b0;
    XRAM[42406] = 8'b0;
    XRAM[42407] = 8'b0;
    XRAM[42408] = 8'b0;
    XRAM[42409] = 8'b0;
    XRAM[42410] = 8'b0;
    XRAM[42411] = 8'b0;
    XRAM[42412] = 8'b0;
    XRAM[42413] = 8'b0;
    XRAM[42414] = 8'b0;
    XRAM[42415] = 8'b0;
    XRAM[42416] = 8'b0;
    XRAM[42417] = 8'b0;
    XRAM[42418] = 8'b0;
    XRAM[42419] = 8'b0;
    XRAM[42420] = 8'b0;
    XRAM[42421] = 8'b0;
    XRAM[42422] = 8'b0;
    XRAM[42423] = 8'b0;
    XRAM[42424] = 8'b0;
    XRAM[42425] = 8'b0;
    XRAM[42426] = 8'b0;
    XRAM[42427] = 8'b0;
    XRAM[42428] = 8'b0;
    XRAM[42429] = 8'b0;
    XRAM[42430] = 8'b0;
    XRAM[42431] = 8'b0;
    XRAM[42432] = 8'b0;
    XRAM[42433] = 8'b0;
    XRAM[42434] = 8'b0;
    XRAM[42435] = 8'b0;
    XRAM[42436] = 8'b0;
    XRAM[42437] = 8'b0;
    XRAM[42438] = 8'b0;
    XRAM[42439] = 8'b0;
    XRAM[42440] = 8'b0;
    XRAM[42441] = 8'b0;
    XRAM[42442] = 8'b0;
    XRAM[42443] = 8'b0;
    XRAM[42444] = 8'b0;
    XRAM[42445] = 8'b0;
    XRAM[42446] = 8'b0;
    XRAM[42447] = 8'b0;
    XRAM[42448] = 8'b0;
    XRAM[42449] = 8'b0;
    XRAM[42450] = 8'b0;
    XRAM[42451] = 8'b0;
    XRAM[42452] = 8'b0;
    XRAM[42453] = 8'b0;
    XRAM[42454] = 8'b0;
    XRAM[42455] = 8'b0;
    XRAM[42456] = 8'b0;
    XRAM[42457] = 8'b0;
    XRAM[42458] = 8'b0;
    XRAM[42459] = 8'b0;
    XRAM[42460] = 8'b0;
    XRAM[42461] = 8'b0;
    XRAM[42462] = 8'b0;
    XRAM[42463] = 8'b0;
    XRAM[42464] = 8'b0;
    XRAM[42465] = 8'b0;
    XRAM[42466] = 8'b0;
    XRAM[42467] = 8'b0;
    XRAM[42468] = 8'b0;
    XRAM[42469] = 8'b0;
    XRAM[42470] = 8'b0;
    XRAM[42471] = 8'b0;
    XRAM[42472] = 8'b0;
    XRAM[42473] = 8'b0;
    XRAM[42474] = 8'b0;
    XRAM[42475] = 8'b0;
    XRAM[42476] = 8'b0;
    XRAM[42477] = 8'b0;
    XRAM[42478] = 8'b0;
    XRAM[42479] = 8'b0;
    XRAM[42480] = 8'b0;
    XRAM[42481] = 8'b0;
    XRAM[42482] = 8'b0;
    XRAM[42483] = 8'b0;
    XRAM[42484] = 8'b0;
    XRAM[42485] = 8'b0;
    XRAM[42486] = 8'b0;
    XRAM[42487] = 8'b0;
    XRAM[42488] = 8'b0;
    XRAM[42489] = 8'b0;
    XRAM[42490] = 8'b0;
    XRAM[42491] = 8'b0;
    XRAM[42492] = 8'b0;
    XRAM[42493] = 8'b0;
    XRAM[42494] = 8'b0;
    XRAM[42495] = 8'b0;
    XRAM[42496] = 8'b0;
    XRAM[42497] = 8'b0;
    XRAM[42498] = 8'b0;
    XRAM[42499] = 8'b0;
    XRAM[42500] = 8'b0;
    XRAM[42501] = 8'b0;
    XRAM[42502] = 8'b0;
    XRAM[42503] = 8'b0;
    XRAM[42504] = 8'b0;
    XRAM[42505] = 8'b0;
    XRAM[42506] = 8'b0;
    XRAM[42507] = 8'b0;
    XRAM[42508] = 8'b0;
    XRAM[42509] = 8'b0;
    XRAM[42510] = 8'b0;
    XRAM[42511] = 8'b0;
    XRAM[42512] = 8'b0;
    XRAM[42513] = 8'b0;
    XRAM[42514] = 8'b0;
    XRAM[42515] = 8'b0;
    XRAM[42516] = 8'b0;
    XRAM[42517] = 8'b0;
    XRAM[42518] = 8'b0;
    XRAM[42519] = 8'b0;
    XRAM[42520] = 8'b0;
    XRAM[42521] = 8'b0;
    XRAM[42522] = 8'b0;
    XRAM[42523] = 8'b0;
    XRAM[42524] = 8'b0;
    XRAM[42525] = 8'b0;
    XRAM[42526] = 8'b0;
    XRAM[42527] = 8'b0;
    XRAM[42528] = 8'b0;
    XRAM[42529] = 8'b0;
    XRAM[42530] = 8'b0;
    XRAM[42531] = 8'b0;
    XRAM[42532] = 8'b0;
    XRAM[42533] = 8'b0;
    XRAM[42534] = 8'b0;
    XRAM[42535] = 8'b0;
    XRAM[42536] = 8'b0;
    XRAM[42537] = 8'b0;
    XRAM[42538] = 8'b0;
    XRAM[42539] = 8'b0;
    XRAM[42540] = 8'b0;
    XRAM[42541] = 8'b0;
    XRAM[42542] = 8'b0;
    XRAM[42543] = 8'b0;
    XRAM[42544] = 8'b0;
    XRAM[42545] = 8'b0;
    XRAM[42546] = 8'b0;
    XRAM[42547] = 8'b0;
    XRAM[42548] = 8'b0;
    XRAM[42549] = 8'b0;
    XRAM[42550] = 8'b0;
    XRAM[42551] = 8'b0;
    XRAM[42552] = 8'b0;
    XRAM[42553] = 8'b0;
    XRAM[42554] = 8'b0;
    XRAM[42555] = 8'b0;
    XRAM[42556] = 8'b0;
    XRAM[42557] = 8'b0;
    XRAM[42558] = 8'b0;
    XRAM[42559] = 8'b0;
    XRAM[42560] = 8'b0;
    XRAM[42561] = 8'b0;
    XRAM[42562] = 8'b0;
    XRAM[42563] = 8'b0;
    XRAM[42564] = 8'b0;
    XRAM[42565] = 8'b0;
    XRAM[42566] = 8'b0;
    XRAM[42567] = 8'b0;
    XRAM[42568] = 8'b0;
    XRAM[42569] = 8'b0;
    XRAM[42570] = 8'b0;
    XRAM[42571] = 8'b0;
    XRAM[42572] = 8'b0;
    XRAM[42573] = 8'b0;
    XRAM[42574] = 8'b0;
    XRAM[42575] = 8'b0;
    XRAM[42576] = 8'b0;
    XRAM[42577] = 8'b0;
    XRAM[42578] = 8'b0;
    XRAM[42579] = 8'b0;
    XRAM[42580] = 8'b0;
    XRAM[42581] = 8'b0;
    XRAM[42582] = 8'b0;
    XRAM[42583] = 8'b0;
    XRAM[42584] = 8'b0;
    XRAM[42585] = 8'b0;
    XRAM[42586] = 8'b0;
    XRAM[42587] = 8'b0;
    XRAM[42588] = 8'b0;
    XRAM[42589] = 8'b0;
    XRAM[42590] = 8'b0;
    XRAM[42591] = 8'b0;
    XRAM[42592] = 8'b0;
    XRAM[42593] = 8'b0;
    XRAM[42594] = 8'b0;
    XRAM[42595] = 8'b0;
    XRAM[42596] = 8'b0;
    XRAM[42597] = 8'b0;
    XRAM[42598] = 8'b0;
    XRAM[42599] = 8'b0;
    XRAM[42600] = 8'b0;
    XRAM[42601] = 8'b0;
    XRAM[42602] = 8'b0;
    XRAM[42603] = 8'b0;
    XRAM[42604] = 8'b0;
    XRAM[42605] = 8'b0;
    XRAM[42606] = 8'b0;
    XRAM[42607] = 8'b0;
    XRAM[42608] = 8'b0;
    XRAM[42609] = 8'b0;
    XRAM[42610] = 8'b0;
    XRAM[42611] = 8'b0;
    XRAM[42612] = 8'b0;
    XRAM[42613] = 8'b0;
    XRAM[42614] = 8'b0;
    XRAM[42615] = 8'b0;
    XRAM[42616] = 8'b0;
    XRAM[42617] = 8'b0;
    XRAM[42618] = 8'b0;
    XRAM[42619] = 8'b0;
    XRAM[42620] = 8'b0;
    XRAM[42621] = 8'b0;
    XRAM[42622] = 8'b0;
    XRAM[42623] = 8'b0;
    XRAM[42624] = 8'b0;
    XRAM[42625] = 8'b0;
    XRAM[42626] = 8'b0;
    XRAM[42627] = 8'b0;
    XRAM[42628] = 8'b0;
    XRAM[42629] = 8'b0;
    XRAM[42630] = 8'b0;
    XRAM[42631] = 8'b0;
    XRAM[42632] = 8'b0;
    XRAM[42633] = 8'b0;
    XRAM[42634] = 8'b0;
    XRAM[42635] = 8'b0;
    XRAM[42636] = 8'b0;
    XRAM[42637] = 8'b0;
    XRAM[42638] = 8'b0;
    XRAM[42639] = 8'b0;
    XRAM[42640] = 8'b0;
    XRAM[42641] = 8'b0;
    XRAM[42642] = 8'b0;
    XRAM[42643] = 8'b0;
    XRAM[42644] = 8'b0;
    XRAM[42645] = 8'b0;
    XRAM[42646] = 8'b0;
    XRAM[42647] = 8'b0;
    XRAM[42648] = 8'b0;
    XRAM[42649] = 8'b0;
    XRAM[42650] = 8'b0;
    XRAM[42651] = 8'b0;
    XRAM[42652] = 8'b0;
    XRAM[42653] = 8'b0;
    XRAM[42654] = 8'b0;
    XRAM[42655] = 8'b0;
    XRAM[42656] = 8'b0;
    XRAM[42657] = 8'b0;
    XRAM[42658] = 8'b0;
    XRAM[42659] = 8'b0;
    XRAM[42660] = 8'b0;
    XRAM[42661] = 8'b0;
    XRAM[42662] = 8'b0;
    XRAM[42663] = 8'b0;
    XRAM[42664] = 8'b0;
    XRAM[42665] = 8'b0;
    XRAM[42666] = 8'b0;
    XRAM[42667] = 8'b0;
    XRAM[42668] = 8'b0;
    XRAM[42669] = 8'b0;
    XRAM[42670] = 8'b0;
    XRAM[42671] = 8'b0;
    XRAM[42672] = 8'b0;
    XRAM[42673] = 8'b0;
    XRAM[42674] = 8'b0;
    XRAM[42675] = 8'b0;
    XRAM[42676] = 8'b0;
    XRAM[42677] = 8'b0;
    XRAM[42678] = 8'b0;
    XRAM[42679] = 8'b0;
    XRAM[42680] = 8'b0;
    XRAM[42681] = 8'b0;
    XRAM[42682] = 8'b0;
    XRAM[42683] = 8'b0;
    XRAM[42684] = 8'b0;
    XRAM[42685] = 8'b0;
    XRAM[42686] = 8'b0;
    XRAM[42687] = 8'b0;
    XRAM[42688] = 8'b0;
    XRAM[42689] = 8'b0;
    XRAM[42690] = 8'b0;
    XRAM[42691] = 8'b0;
    XRAM[42692] = 8'b0;
    XRAM[42693] = 8'b0;
    XRAM[42694] = 8'b0;
    XRAM[42695] = 8'b0;
    XRAM[42696] = 8'b0;
    XRAM[42697] = 8'b0;
    XRAM[42698] = 8'b0;
    XRAM[42699] = 8'b0;
    XRAM[42700] = 8'b0;
    XRAM[42701] = 8'b0;
    XRAM[42702] = 8'b0;
    XRAM[42703] = 8'b0;
    XRAM[42704] = 8'b0;
    XRAM[42705] = 8'b0;
    XRAM[42706] = 8'b0;
    XRAM[42707] = 8'b0;
    XRAM[42708] = 8'b0;
    XRAM[42709] = 8'b0;
    XRAM[42710] = 8'b0;
    XRAM[42711] = 8'b0;
    XRAM[42712] = 8'b0;
    XRAM[42713] = 8'b0;
    XRAM[42714] = 8'b0;
    XRAM[42715] = 8'b0;
    XRAM[42716] = 8'b0;
    XRAM[42717] = 8'b0;
    XRAM[42718] = 8'b0;
    XRAM[42719] = 8'b0;
    XRAM[42720] = 8'b0;
    XRAM[42721] = 8'b0;
    XRAM[42722] = 8'b0;
    XRAM[42723] = 8'b0;
    XRAM[42724] = 8'b0;
    XRAM[42725] = 8'b0;
    XRAM[42726] = 8'b0;
    XRAM[42727] = 8'b0;
    XRAM[42728] = 8'b0;
    XRAM[42729] = 8'b0;
    XRAM[42730] = 8'b0;
    XRAM[42731] = 8'b0;
    XRAM[42732] = 8'b0;
    XRAM[42733] = 8'b0;
    XRAM[42734] = 8'b0;
    XRAM[42735] = 8'b0;
    XRAM[42736] = 8'b0;
    XRAM[42737] = 8'b0;
    XRAM[42738] = 8'b0;
    XRAM[42739] = 8'b0;
    XRAM[42740] = 8'b0;
    XRAM[42741] = 8'b0;
    XRAM[42742] = 8'b0;
    XRAM[42743] = 8'b0;
    XRAM[42744] = 8'b0;
    XRAM[42745] = 8'b0;
    XRAM[42746] = 8'b0;
    XRAM[42747] = 8'b0;
    XRAM[42748] = 8'b0;
    XRAM[42749] = 8'b0;
    XRAM[42750] = 8'b0;
    XRAM[42751] = 8'b0;
    XRAM[42752] = 8'b0;
    XRAM[42753] = 8'b0;
    XRAM[42754] = 8'b0;
    XRAM[42755] = 8'b0;
    XRAM[42756] = 8'b0;
    XRAM[42757] = 8'b0;
    XRAM[42758] = 8'b0;
    XRAM[42759] = 8'b0;
    XRAM[42760] = 8'b0;
    XRAM[42761] = 8'b0;
    XRAM[42762] = 8'b0;
    XRAM[42763] = 8'b0;
    XRAM[42764] = 8'b0;
    XRAM[42765] = 8'b0;
    XRAM[42766] = 8'b0;
    XRAM[42767] = 8'b0;
    XRAM[42768] = 8'b0;
    XRAM[42769] = 8'b0;
    XRAM[42770] = 8'b0;
    XRAM[42771] = 8'b0;
    XRAM[42772] = 8'b0;
    XRAM[42773] = 8'b0;
    XRAM[42774] = 8'b0;
    XRAM[42775] = 8'b0;
    XRAM[42776] = 8'b0;
    XRAM[42777] = 8'b0;
    XRAM[42778] = 8'b0;
    XRAM[42779] = 8'b0;
    XRAM[42780] = 8'b0;
    XRAM[42781] = 8'b0;
    XRAM[42782] = 8'b0;
    XRAM[42783] = 8'b0;
    XRAM[42784] = 8'b0;
    XRAM[42785] = 8'b0;
    XRAM[42786] = 8'b0;
    XRAM[42787] = 8'b0;
    XRAM[42788] = 8'b0;
    XRAM[42789] = 8'b0;
    XRAM[42790] = 8'b0;
    XRAM[42791] = 8'b0;
    XRAM[42792] = 8'b0;
    XRAM[42793] = 8'b0;
    XRAM[42794] = 8'b0;
    XRAM[42795] = 8'b0;
    XRAM[42796] = 8'b0;
    XRAM[42797] = 8'b0;
    XRAM[42798] = 8'b0;
    XRAM[42799] = 8'b0;
    XRAM[42800] = 8'b0;
    XRAM[42801] = 8'b0;
    XRAM[42802] = 8'b0;
    XRAM[42803] = 8'b0;
    XRAM[42804] = 8'b0;
    XRAM[42805] = 8'b0;
    XRAM[42806] = 8'b0;
    XRAM[42807] = 8'b0;
    XRAM[42808] = 8'b0;
    XRAM[42809] = 8'b0;
    XRAM[42810] = 8'b0;
    XRAM[42811] = 8'b0;
    XRAM[42812] = 8'b0;
    XRAM[42813] = 8'b0;
    XRAM[42814] = 8'b0;
    XRAM[42815] = 8'b0;
    XRAM[42816] = 8'b0;
    XRAM[42817] = 8'b0;
    XRAM[42818] = 8'b0;
    XRAM[42819] = 8'b0;
    XRAM[42820] = 8'b0;
    XRAM[42821] = 8'b0;
    XRAM[42822] = 8'b0;
    XRAM[42823] = 8'b0;
    XRAM[42824] = 8'b0;
    XRAM[42825] = 8'b0;
    XRAM[42826] = 8'b0;
    XRAM[42827] = 8'b0;
    XRAM[42828] = 8'b0;
    XRAM[42829] = 8'b0;
    XRAM[42830] = 8'b0;
    XRAM[42831] = 8'b0;
    XRAM[42832] = 8'b0;
    XRAM[42833] = 8'b0;
    XRAM[42834] = 8'b0;
    XRAM[42835] = 8'b0;
    XRAM[42836] = 8'b0;
    XRAM[42837] = 8'b0;
    XRAM[42838] = 8'b0;
    XRAM[42839] = 8'b0;
    XRAM[42840] = 8'b0;
    XRAM[42841] = 8'b0;
    XRAM[42842] = 8'b0;
    XRAM[42843] = 8'b0;
    XRAM[42844] = 8'b0;
    XRAM[42845] = 8'b0;
    XRAM[42846] = 8'b0;
    XRAM[42847] = 8'b0;
    XRAM[42848] = 8'b0;
    XRAM[42849] = 8'b0;
    XRAM[42850] = 8'b0;
    XRAM[42851] = 8'b0;
    XRAM[42852] = 8'b0;
    XRAM[42853] = 8'b0;
    XRAM[42854] = 8'b0;
    XRAM[42855] = 8'b0;
    XRAM[42856] = 8'b0;
    XRAM[42857] = 8'b0;
    XRAM[42858] = 8'b0;
    XRAM[42859] = 8'b0;
    XRAM[42860] = 8'b0;
    XRAM[42861] = 8'b0;
    XRAM[42862] = 8'b0;
    XRAM[42863] = 8'b0;
    XRAM[42864] = 8'b0;
    XRAM[42865] = 8'b0;
    XRAM[42866] = 8'b0;
    XRAM[42867] = 8'b0;
    XRAM[42868] = 8'b0;
    XRAM[42869] = 8'b0;
    XRAM[42870] = 8'b0;
    XRAM[42871] = 8'b0;
    XRAM[42872] = 8'b0;
    XRAM[42873] = 8'b0;
    XRAM[42874] = 8'b0;
    XRAM[42875] = 8'b0;
    XRAM[42876] = 8'b0;
    XRAM[42877] = 8'b0;
    XRAM[42878] = 8'b0;
    XRAM[42879] = 8'b0;
    XRAM[42880] = 8'b0;
    XRAM[42881] = 8'b0;
    XRAM[42882] = 8'b0;
    XRAM[42883] = 8'b0;
    XRAM[42884] = 8'b0;
    XRAM[42885] = 8'b0;
    XRAM[42886] = 8'b0;
    XRAM[42887] = 8'b0;
    XRAM[42888] = 8'b0;
    XRAM[42889] = 8'b0;
    XRAM[42890] = 8'b0;
    XRAM[42891] = 8'b0;
    XRAM[42892] = 8'b0;
    XRAM[42893] = 8'b0;
    XRAM[42894] = 8'b0;
    XRAM[42895] = 8'b0;
    XRAM[42896] = 8'b0;
    XRAM[42897] = 8'b0;
    XRAM[42898] = 8'b0;
    XRAM[42899] = 8'b0;
    XRAM[42900] = 8'b0;
    XRAM[42901] = 8'b0;
    XRAM[42902] = 8'b0;
    XRAM[42903] = 8'b0;
    XRAM[42904] = 8'b0;
    XRAM[42905] = 8'b0;
    XRAM[42906] = 8'b0;
    XRAM[42907] = 8'b0;
    XRAM[42908] = 8'b0;
    XRAM[42909] = 8'b0;
    XRAM[42910] = 8'b0;
    XRAM[42911] = 8'b0;
    XRAM[42912] = 8'b0;
    XRAM[42913] = 8'b0;
    XRAM[42914] = 8'b0;
    XRAM[42915] = 8'b0;
    XRAM[42916] = 8'b0;
    XRAM[42917] = 8'b0;
    XRAM[42918] = 8'b0;
    XRAM[42919] = 8'b0;
    XRAM[42920] = 8'b0;
    XRAM[42921] = 8'b0;
    XRAM[42922] = 8'b0;
    XRAM[42923] = 8'b0;
    XRAM[42924] = 8'b0;
    XRAM[42925] = 8'b0;
    XRAM[42926] = 8'b0;
    XRAM[42927] = 8'b0;
    XRAM[42928] = 8'b0;
    XRAM[42929] = 8'b0;
    XRAM[42930] = 8'b0;
    XRAM[42931] = 8'b0;
    XRAM[42932] = 8'b0;
    XRAM[42933] = 8'b0;
    XRAM[42934] = 8'b0;
    XRAM[42935] = 8'b0;
    XRAM[42936] = 8'b0;
    XRAM[42937] = 8'b0;
    XRAM[42938] = 8'b0;
    XRAM[42939] = 8'b0;
    XRAM[42940] = 8'b0;
    XRAM[42941] = 8'b0;
    XRAM[42942] = 8'b0;
    XRAM[42943] = 8'b0;
    XRAM[42944] = 8'b0;
    XRAM[42945] = 8'b0;
    XRAM[42946] = 8'b0;
    XRAM[42947] = 8'b0;
    XRAM[42948] = 8'b0;
    XRAM[42949] = 8'b0;
    XRAM[42950] = 8'b0;
    XRAM[42951] = 8'b0;
    XRAM[42952] = 8'b0;
    XRAM[42953] = 8'b0;
    XRAM[42954] = 8'b0;
    XRAM[42955] = 8'b0;
    XRAM[42956] = 8'b0;
    XRAM[42957] = 8'b0;
    XRAM[42958] = 8'b0;
    XRAM[42959] = 8'b0;
    XRAM[42960] = 8'b0;
    XRAM[42961] = 8'b0;
    XRAM[42962] = 8'b0;
    XRAM[42963] = 8'b0;
    XRAM[42964] = 8'b0;
    XRAM[42965] = 8'b0;
    XRAM[42966] = 8'b0;
    XRAM[42967] = 8'b0;
    XRAM[42968] = 8'b0;
    XRAM[42969] = 8'b0;
    XRAM[42970] = 8'b0;
    XRAM[42971] = 8'b0;
    XRAM[42972] = 8'b0;
    XRAM[42973] = 8'b0;
    XRAM[42974] = 8'b0;
    XRAM[42975] = 8'b0;
    XRAM[42976] = 8'b0;
    XRAM[42977] = 8'b0;
    XRAM[42978] = 8'b0;
    XRAM[42979] = 8'b0;
    XRAM[42980] = 8'b0;
    XRAM[42981] = 8'b0;
    XRAM[42982] = 8'b0;
    XRAM[42983] = 8'b0;
    XRAM[42984] = 8'b0;
    XRAM[42985] = 8'b0;
    XRAM[42986] = 8'b0;
    XRAM[42987] = 8'b0;
    XRAM[42988] = 8'b0;
    XRAM[42989] = 8'b0;
    XRAM[42990] = 8'b0;
    XRAM[42991] = 8'b0;
    XRAM[42992] = 8'b0;
    XRAM[42993] = 8'b0;
    XRAM[42994] = 8'b0;
    XRAM[42995] = 8'b0;
    XRAM[42996] = 8'b0;
    XRAM[42997] = 8'b0;
    XRAM[42998] = 8'b0;
    XRAM[42999] = 8'b0;
    XRAM[43000] = 8'b0;
    XRAM[43001] = 8'b0;
    XRAM[43002] = 8'b0;
    XRAM[43003] = 8'b0;
    XRAM[43004] = 8'b0;
    XRAM[43005] = 8'b0;
    XRAM[43006] = 8'b0;
    XRAM[43007] = 8'b0;
    XRAM[43008] = 8'b0;
    XRAM[43009] = 8'b0;
    XRAM[43010] = 8'b0;
    XRAM[43011] = 8'b0;
    XRAM[43012] = 8'b0;
    XRAM[43013] = 8'b0;
    XRAM[43014] = 8'b0;
    XRAM[43015] = 8'b0;
    XRAM[43016] = 8'b0;
    XRAM[43017] = 8'b0;
    XRAM[43018] = 8'b0;
    XRAM[43019] = 8'b0;
    XRAM[43020] = 8'b0;
    XRAM[43021] = 8'b0;
    XRAM[43022] = 8'b0;
    XRAM[43023] = 8'b0;
    XRAM[43024] = 8'b0;
    XRAM[43025] = 8'b0;
    XRAM[43026] = 8'b0;
    XRAM[43027] = 8'b0;
    XRAM[43028] = 8'b0;
    XRAM[43029] = 8'b0;
    XRAM[43030] = 8'b0;
    XRAM[43031] = 8'b0;
    XRAM[43032] = 8'b0;
    XRAM[43033] = 8'b0;
    XRAM[43034] = 8'b0;
    XRAM[43035] = 8'b0;
    XRAM[43036] = 8'b0;
    XRAM[43037] = 8'b0;
    XRAM[43038] = 8'b0;
    XRAM[43039] = 8'b0;
    XRAM[43040] = 8'b0;
    XRAM[43041] = 8'b0;
    XRAM[43042] = 8'b0;
    XRAM[43043] = 8'b0;
    XRAM[43044] = 8'b0;
    XRAM[43045] = 8'b0;
    XRAM[43046] = 8'b0;
    XRAM[43047] = 8'b0;
    XRAM[43048] = 8'b0;
    XRAM[43049] = 8'b0;
    XRAM[43050] = 8'b0;
    XRAM[43051] = 8'b0;
    XRAM[43052] = 8'b0;
    XRAM[43053] = 8'b0;
    XRAM[43054] = 8'b0;
    XRAM[43055] = 8'b0;
    XRAM[43056] = 8'b0;
    XRAM[43057] = 8'b0;
    XRAM[43058] = 8'b0;
    XRAM[43059] = 8'b0;
    XRAM[43060] = 8'b0;
    XRAM[43061] = 8'b0;
    XRAM[43062] = 8'b0;
    XRAM[43063] = 8'b0;
    XRAM[43064] = 8'b0;
    XRAM[43065] = 8'b0;
    XRAM[43066] = 8'b0;
    XRAM[43067] = 8'b0;
    XRAM[43068] = 8'b0;
    XRAM[43069] = 8'b0;
    XRAM[43070] = 8'b0;
    XRAM[43071] = 8'b0;
    XRAM[43072] = 8'b0;
    XRAM[43073] = 8'b0;
    XRAM[43074] = 8'b0;
    XRAM[43075] = 8'b0;
    XRAM[43076] = 8'b0;
    XRAM[43077] = 8'b0;
    XRAM[43078] = 8'b0;
    XRAM[43079] = 8'b0;
    XRAM[43080] = 8'b0;
    XRAM[43081] = 8'b0;
    XRAM[43082] = 8'b0;
    XRAM[43083] = 8'b0;
    XRAM[43084] = 8'b0;
    XRAM[43085] = 8'b0;
    XRAM[43086] = 8'b0;
    XRAM[43087] = 8'b0;
    XRAM[43088] = 8'b0;
    XRAM[43089] = 8'b0;
    XRAM[43090] = 8'b0;
    XRAM[43091] = 8'b0;
    XRAM[43092] = 8'b0;
    XRAM[43093] = 8'b0;
    XRAM[43094] = 8'b0;
    XRAM[43095] = 8'b0;
    XRAM[43096] = 8'b0;
    XRAM[43097] = 8'b0;
    XRAM[43098] = 8'b0;
    XRAM[43099] = 8'b0;
    XRAM[43100] = 8'b0;
    XRAM[43101] = 8'b0;
    XRAM[43102] = 8'b0;
    XRAM[43103] = 8'b0;
    XRAM[43104] = 8'b0;
    XRAM[43105] = 8'b0;
    XRAM[43106] = 8'b0;
    XRAM[43107] = 8'b0;
    XRAM[43108] = 8'b0;
    XRAM[43109] = 8'b0;
    XRAM[43110] = 8'b0;
    XRAM[43111] = 8'b0;
    XRAM[43112] = 8'b0;
    XRAM[43113] = 8'b0;
    XRAM[43114] = 8'b0;
    XRAM[43115] = 8'b0;
    XRAM[43116] = 8'b0;
    XRAM[43117] = 8'b0;
    XRAM[43118] = 8'b0;
    XRAM[43119] = 8'b0;
    XRAM[43120] = 8'b0;
    XRAM[43121] = 8'b0;
    XRAM[43122] = 8'b0;
    XRAM[43123] = 8'b0;
    XRAM[43124] = 8'b0;
    XRAM[43125] = 8'b0;
    XRAM[43126] = 8'b0;
    XRAM[43127] = 8'b0;
    XRAM[43128] = 8'b0;
    XRAM[43129] = 8'b0;
    XRAM[43130] = 8'b0;
    XRAM[43131] = 8'b0;
    XRAM[43132] = 8'b0;
    XRAM[43133] = 8'b0;
    XRAM[43134] = 8'b0;
    XRAM[43135] = 8'b0;
    XRAM[43136] = 8'b0;
    XRAM[43137] = 8'b0;
    XRAM[43138] = 8'b0;
    XRAM[43139] = 8'b0;
    XRAM[43140] = 8'b0;
    XRAM[43141] = 8'b0;
    XRAM[43142] = 8'b0;
    XRAM[43143] = 8'b0;
    XRAM[43144] = 8'b0;
    XRAM[43145] = 8'b0;
    XRAM[43146] = 8'b0;
    XRAM[43147] = 8'b0;
    XRAM[43148] = 8'b0;
    XRAM[43149] = 8'b0;
    XRAM[43150] = 8'b0;
    XRAM[43151] = 8'b0;
    XRAM[43152] = 8'b0;
    XRAM[43153] = 8'b0;
    XRAM[43154] = 8'b0;
    XRAM[43155] = 8'b0;
    XRAM[43156] = 8'b0;
    XRAM[43157] = 8'b0;
    XRAM[43158] = 8'b0;
    XRAM[43159] = 8'b0;
    XRAM[43160] = 8'b0;
    XRAM[43161] = 8'b0;
    XRAM[43162] = 8'b0;
    XRAM[43163] = 8'b0;
    XRAM[43164] = 8'b0;
    XRAM[43165] = 8'b0;
    XRAM[43166] = 8'b0;
    XRAM[43167] = 8'b0;
    XRAM[43168] = 8'b0;
    XRAM[43169] = 8'b0;
    XRAM[43170] = 8'b0;
    XRAM[43171] = 8'b0;
    XRAM[43172] = 8'b0;
    XRAM[43173] = 8'b0;
    XRAM[43174] = 8'b0;
    XRAM[43175] = 8'b0;
    XRAM[43176] = 8'b0;
    XRAM[43177] = 8'b0;
    XRAM[43178] = 8'b0;
    XRAM[43179] = 8'b0;
    XRAM[43180] = 8'b0;
    XRAM[43181] = 8'b0;
    XRAM[43182] = 8'b0;
    XRAM[43183] = 8'b0;
    XRAM[43184] = 8'b0;
    XRAM[43185] = 8'b0;
    XRAM[43186] = 8'b0;
    XRAM[43187] = 8'b0;
    XRAM[43188] = 8'b0;
    XRAM[43189] = 8'b0;
    XRAM[43190] = 8'b0;
    XRAM[43191] = 8'b0;
    XRAM[43192] = 8'b0;
    XRAM[43193] = 8'b0;
    XRAM[43194] = 8'b0;
    XRAM[43195] = 8'b0;
    XRAM[43196] = 8'b0;
    XRAM[43197] = 8'b0;
    XRAM[43198] = 8'b0;
    XRAM[43199] = 8'b0;
    XRAM[43200] = 8'b0;
    XRAM[43201] = 8'b0;
    XRAM[43202] = 8'b0;
    XRAM[43203] = 8'b0;
    XRAM[43204] = 8'b0;
    XRAM[43205] = 8'b0;
    XRAM[43206] = 8'b0;
    XRAM[43207] = 8'b0;
    XRAM[43208] = 8'b0;
    XRAM[43209] = 8'b0;
    XRAM[43210] = 8'b0;
    XRAM[43211] = 8'b0;
    XRAM[43212] = 8'b0;
    XRAM[43213] = 8'b0;
    XRAM[43214] = 8'b0;
    XRAM[43215] = 8'b0;
    XRAM[43216] = 8'b0;
    XRAM[43217] = 8'b0;
    XRAM[43218] = 8'b0;
    XRAM[43219] = 8'b0;
    XRAM[43220] = 8'b0;
    XRAM[43221] = 8'b0;
    XRAM[43222] = 8'b0;
    XRAM[43223] = 8'b0;
    XRAM[43224] = 8'b0;
    XRAM[43225] = 8'b0;
    XRAM[43226] = 8'b0;
    XRAM[43227] = 8'b0;
    XRAM[43228] = 8'b0;
    XRAM[43229] = 8'b0;
    XRAM[43230] = 8'b0;
    XRAM[43231] = 8'b0;
    XRAM[43232] = 8'b0;
    XRAM[43233] = 8'b0;
    XRAM[43234] = 8'b0;
    XRAM[43235] = 8'b0;
    XRAM[43236] = 8'b0;
    XRAM[43237] = 8'b0;
    XRAM[43238] = 8'b0;
    XRAM[43239] = 8'b0;
    XRAM[43240] = 8'b0;
    XRAM[43241] = 8'b0;
    XRAM[43242] = 8'b0;
    XRAM[43243] = 8'b0;
    XRAM[43244] = 8'b0;
    XRAM[43245] = 8'b0;
    XRAM[43246] = 8'b0;
    XRAM[43247] = 8'b0;
    XRAM[43248] = 8'b0;
    XRAM[43249] = 8'b0;
    XRAM[43250] = 8'b0;
    XRAM[43251] = 8'b0;
    XRAM[43252] = 8'b0;
    XRAM[43253] = 8'b0;
    XRAM[43254] = 8'b0;
    XRAM[43255] = 8'b0;
    XRAM[43256] = 8'b0;
    XRAM[43257] = 8'b0;
    XRAM[43258] = 8'b0;
    XRAM[43259] = 8'b0;
    XRAM[43260] = 8'b0;
    XRAM[43261] = 8'b0;
    XRAM[43262] = 8'b0;
    XRAM[43263] = 8'b0;
    XRAM[43264] = 8'b0;
    XRAM[43265] = 8'b0;
    XRAM[43266] = 8'b0;
    XRAM[43267] = 8'b0;
    XRAM[43268] = 8'b0;
    XRAM[43269] = 8'b0;
    XRAM[43270] = 8'b0;
    XRAM[43271] = 8'b0;
    XRAM[43272] = 8'b0;
    XRAM[43273] = 8'b0;
    XRAM[43274] = 8'b0;
    XRAM[43275] = 8'b0;
    XRAM[43276] = 8'b0;
    XRAM[43277] = 8'b0;
    XRAM[43278] = 8'b0;
    XRAM[43279] = 8'b0;
    XRAM[43280] = 8'b0;
    XRAM[43281] = 8'b0;
    XRAM[43282] = 8'b0;
    XRAM[43283] = 8'b0;
    XRAM[43284] = 8'b0;
    XRAM[43285] = 8'b0;
    XRAM[43286] = 8'b0;
    XRAM[43287] = 8'b0;
    XRAM[43288] = 8'b0;
    XRAM[43289] = 8'b0;
    XRAM[43290] = 8'b0;
    XRAM[43291] = 8'b0;
    XRAM[43292] = 8'b0;
    XRAM[43293] = 8'b0;
    XRAM[43294] = 8'b0;
    XRAM[43295] = 8'b0;
    XRAM[43296] = 8'b0;
    XRAM[43297] = 8'b0;
    XRAM[43298] = 8'b0;
    XRAM[43299] = 8'b0;
    XRAM[43300] = 8'b0;
    XRAM[43301] = 8'b0;
    XRAM[43302] = 8'b0;
    XRAM[43303] = 8'b0;
    XRAM[43304] = 8'b0;
    XRAM[43305] = 8'b0;
    XRAM[43306] = 8'b0;
    XRAM[43307] = 8'b0;
    XRAM[43308] = 8'b0;
    XRAM[43309] = 8'b0;
    XRAM[43310] = 8'b0;
    XRAM[43311] = 8'b0;
    XRAM[43312] = 8'b0;
    XRAM[43313] = 8'b0;
    XRAM[43314] = 8'b0;
    XRAM[43315] = 8'b0;
    XRAM[43316] = 8'b0;
    XRAM[43317] = 8'b0;
    XRAM[43318] = 8'b0;
    XRAM[43319] = 8'b0;
    XRAM[43320] = 8'b0;
    XRAM[43321] = 8'b0;
    XRAM[43322] = 8'b0;
    XRAM[43323] = 8'b0;
    XRAM[43324] = 8'b0;
    XRAM[43325] = 8'b0;
    XRAM[43326] = 8'b0;
    XRAM[43327] = 8'b0;
    XRAM[43328] = 8'b0;
    XRAM[43329] = 8'b0;
    XRAM[43330] = 8'b0;
    XRAM[43331] = 8'b0;
    XRAM[43332] = 8'b0;
    XRAM[43333] = 8'b0;
    XRAM[43334] = 8'b0;
    XRAM[43335] = 8'b0;
    XRAM[43336] = 8'b0;
    XRAM[43337] = 8'b0;
    XRAM[43338] = 8'b0;
    XRAM[43339] = 8'b0;
    XRAM[43340] = 8'b0;
    XRAM[43341] = 8'b0;
    XRAM[43342] = 8'b0;
    XRAM[43343] = 8'b0;
    XRAM[43344] = 8'b0;
    XRAM[43345] = 8'b0;
    XRAM[43346] = 8'b0;
    XRAM[43347] = 8'b0;
    XRAM[43348] = 8'b0;
    XRAM[43349] = 8'b0;
    XRAM[43350] = 8'b0;
    XRAM[43351] = 8'b0;
    XRAM[43352] = 8'b0;
    XRAM[43353] = 8'b0;
    XRAM[43354] = 8'b0;
    XRAM[43355] = 8'b0;
    XRAM[43356] = 8'b0;
    XRAM[43357] = 8'b0;
    XRAM[43358] = 8'b0;
    XRAM[43359] = 8'b0;
    XRAM[43360] = 8'b0;
    XRAM[43361] = 8'b0;
    XRAM[43362] = 8'b0;
    XRAM[43363] = 8'b0;
    XRAM[43364] = 8'b0;
    XRAM[43365] = 8'b0;
    XRAM[43366] = 8'b0;
    XRAM[43367] = 8'b0;
    XRAM[43368] = 8'b0;
    XRAM[43369] = 8'b0;
    XRAM[43370] = 8'b0;
    XRAM[43371] = 8'b0;
    XRAM[43372] = 8'b0;
    XRAM[43373] = 8'b0;
    XRAM[43374] = 8'b0;
    XRAM[43375] = 8'b0;
    XRAM[43376] = 8'b0;
    XRAM[43377] = 8'b0;
    XRAM[43378] = 8'b0;
    XRAM[43379] = 8'b0;
    XRAM[43380] = 8'b0;
    XRAM[43381] = 8'b0;
    XRAM[43382] = 8'b0;
    XRAM[43383] = 8'b0;
    XRAM[43384] = 8'b0;
    XRAM[43385] = 8'b0;
    XRAM[43386] = 8'b0;
    XRAM[43387] = 8'b0;
    XRAM[43388] = 8'b0;
    XRAM[43389] = 8'b0;
    XRAM[43390] = 8'b0;
    XRAM[43391] = 8'b0;
    XRAM[43392] = 8'b0;
    XRAM[43393] = 8'b0;
    XRAM[43394] = 8'b0;
    XRAM[43395] = 8'b0;
    XRAM[43396] = 8'b0;
    XRAM[43397] = 8'b0;
    XRAM[43398] = 8'b0;
    XRAM[43399] = 8'b0;
    XRAM[43400] = 8'b0;
    XRAM[43401] = 8'b0;
    XRAM[43402] = 8'b0;
    XRAM[43403] = 8'b0;
    XRAM[43404] = 8'b0;
    XRAM[43405] = 8'b0;
    XRAM[43406] = 8'b0;
    XRAM[43407] = 8'b0;
    XRAM[43408] = 8'b0;
    XRAM[43409] = 8'b0;
    XRAM[43410] = 8'b0;
    XRAM[43411] = 8'b0;
    XRAM[43412] = 8'b0;
    XRAM[43413] = 8'b0;
    XRAM[43414] = 8'b0;
    XRAM[43415] = 8'b0;
    XRAM[43416] = 8'b0;
    XRAM[43417] = 8'b0;
    XRAM[43418] = 8'b0;
    XRAM[43419] = 8'b0;
    XRAM[43420] = 8'b0;
    XRAM[43421] = 8'b0;
    XRAM[43422] = 8'b0;
    XRAM[43423] = 8'b0;
    XRAM[43424] = 8'b0;
    XRAM[43425] = 8'b0;
    XRAM[43426] = 8'b0;
    XRAM[43427] = 8'b0;
    XRAM[43428] = 8'b0;
    XRAM[43429] = 8'b0;
    XRAM[43430] = 8'b0;
    XRAM[43431] = 8'b0;
    XRAM[43432] = 8'b0;
    XRAM[43433] = 8'b0;
    XRAM[43434] = 8'b0;
    XRAM[43435] = 8'b0;
    XRAM[43436] = 8'b0;
    XRAM[43437] = 8'b0;
    XRAM[43438] = 8'b0;
    XRAM[43439] = 8'b0;
    XRAM[43440] = 8'b0;
    XRAM[43441] = 8'b0;
    XRAM[43442] = 8'b0;
    XRAM[43443] = 8'b0;
    XRAM[43444] = 8'b0;
    XRAM[43445] = 8'b0;
    XRAM[43446] = 8'b0;
    XRAM[43447] = 8'b0;
    XRAM[43448] = 8'b0;
    XRAM[43449] = 8'b0;
    XRAM[43450] = 8'b0;
    XRAM[43451] = 8'b0;
    XRAM[43452] = 8'b0;
    XRAM[43453] = 8'b0;
    XRAM[43454] = 8'b0;
    XRAM[43455] = 8'b0;
    XRAM[43456] = 8'b0;
    XRAM[43457] = 8'b0;
    XRAM[43458] = 8'b0;
    XRAM[43459] = 8'b0;
    XRAM[43460] = 8'b0;
    XRAM[43461] = 8'b0;
    XRAM[43462] = 8'b0;
    XRAM[43463] = 8'b0;
    XRAM[43464] = 8'b0;
    XRAM[43465] = 8'b0;
    XRAM[43466] = 8'b0;
    XRAM[43467] = 8'b0;
    XRAM[43468] = 8'b0;
    XRAM[43469] = 8'b0;
    XRAM[43470] = 8'b0;
    XRAM[43471] = 8'b0;
    XRAM[43472] = 8'b0;
    XRAM[43473] = 8'b0;
    XRAM[43474] = 8'b0;
    XRAM[43475] = 8'b0;
    XRAM[43476] = 8'b0;
    XRAM[43477] = 8'b0;
    XRAM[43478] = 8'b0;
    XRAM[43479] = 8'b0;
    XRAM[43480] = 8'b0;
    XRAM[43481] = 8'b0;
    XRAM[43482] = 8'b0;
    XRAM[43483] = 8'b0;
    XRAM[43484] = 8'b0;
    XRAM[43485] = 8'b0;
    XRAM[43486] = 8'b0;
    XRAM[43487] = 8'b0;
    XRAM[43488] = 8'b0;
    XRAM[43489] = 8'b0;
    XRAM[43490] = 8'b0;
    XRAM[43491] = 8'b0;
    XRAM[43492] = 8'b0;
    XRAM[43493] = 8'b0;
    XRAM[43494] = 8'b0;
    XRAM[43495] = 8'b0;
    XRAM[43496] = 8'b0;
    XRAM[43497] = 8'b0;
    XRAM[43498] = 8'b0;
    XRAM[43499] = 8'b0;
    XRAM[43500] = 8'b0;
    XRAM[43501] = 8'b0;
    XRAM[43502] = 8'b0;
    XRAM[43503] = 8'b0;
    XRAM[43504] = 8'b0;
    XRAM[43505] = 8'b0;
    XRAM[43506] = 8'b0;
    XRAM[43507] = 8'b0;
    XRAM[43508] = 8'b0;
    XRAM[43509] = 8'b0;
    XRAM[43510] = 8'b0;
    XRAM[43511] = 8'b0;
    XRAM[43512] = 8'b0;
    XRAM[43513] = 8'b0;
    XRAM[43514] = 8'b0;
    XRAM[43515] = 8'b0;
    XRAM[43516] = 8'b0;
    XRAM[43517] = 8'b0;
    XRAM[43518] = 8'b0;
    XRAM[43519] = 8'b0;
    XRAM[43520] = 8'b0;
    XRAM[43521] = 8'b0;
    XRAM[43522] = 8'b0;
    XRAM[43523] = 8'b0;
    XRAM[43524] = 8'b0;
    XRAM[43525] = 8'b0;
    XRAM[43526] = 8'b0;
    XRAM[43527] = 8'b0;
    XRAM[43528] = 8'b0;
    XRAM[43529] = 8'b0;
    XRAM[43530] = 8'b0;
    XRAM[43531] = 8'b0;
    XRAM[43532] = 8'b0;
    XRAM[43533] = 8'b0;
    XRAM[43534] = 8'b0;
    XRAM[43535] = 8'b0;
    XRAM[43536] = 8'b0;
    XRAM[43537] = 8'b0;
    XRAM[43538] = 8'b0;
    XRAM[43539] = 8'b0;
    XRAM[43540] = 8'b0;
    XRAM[43541] = 8'b0;
    XRAM[43542] = 8'b0;
    XRAM[43543] = 8'b0;
    XRAM[43544] = 8'b0;
    XRAM[43545] = 8'b0;
    XRAM[43546] = 8'b0;
    XRAM[43547] = 8'b0;
    XRAM[43548] = 8'b0;
    XRAM[43549] = 8'b0;
    XRAM[43550] = 8'b0;
    XRAM[43551] = 8'b0;
    XRAM[43552] = 8'b0;
    XRAM[43553] = 8'b0;
    XRAM[43554] = 8'b0;
    XRAM[43555] = 8'b0;
    XRAM[43556] = 8'b0;
    XRAM[43557] = 8'b0;
    XRAM[43558] = 8'b0;
    XRAM[43559] = 8'b0;
    XRAM[43560] = 8'b0;
    XRAM[43561] = 8'b0;
    XRAM[43562] = 8'b0;
    XRAM[43563] = 8'b0;
    XRAM[43564] = 8'b0;
    XRAM[43565] = 8'b0;
    XRAM[43566] = 8'b0;
    XRAM[43567] = 8'b0;
    XRAM[43568] = 8'b0;
    XRAM[43569] = 8'b0;
    XRAM[43570] = 8'b0;
    XRAM[43571] = 8'b0;
    XRAM[43572] = 8'b0;
    XRAM[43573] = 8'b0;
    XRAM[43574] = 8'b0;
    XRAM[43575] = 8'b0;
    XRAM[43576] = 8'b0;
    XRAM[43577] = 8'b0;
    XRAM[43578] = 8'b0;
    XRAM[43579] = 8'b0;
    XRAM[43580] = 8'b0;
    XRAM[43581] = 8'b0;
    XRAM[43582] = 8'b0;
    XRAM[43583] = 8'b0;
    XRAM[43584] = 8'b0;
    XRAM[43585] = 8'b0;
    XRAM[43586] = 8'b0;
    XRAM[43587] = 8'b0;
    XRAM[43588] = 8'b0;
    XRAM[43589] = 8'b0;
    XRAM[43590] = 8'b0;
    XRAM[43591] = 8'b0;
    XRAM[43592] = 8'b0;
    XRAM[43593] = 8'b0;
    XRAM[43594] = 8'b0;
    XRAM[43595] = 8'b0;
    XRAM[43596] = 8'b0;
    XRAM[43597] = 8'b0;
    XRAM[43598] = 8'b0;
    XRAM[43599] = 8'b0;
    XRAM[43600] = 8'b0;
    XRAM[43601] = 8'b0;
    XRAM[43602] = 8'b0;
    XRAM[43603] = 8'b0;
    XRAM[43604] = 8'b0;
    XRAM[43605] = 8'b0;
    XRAM[43606] = 8'b0;
    XRAM[43607] = 8'b0;
    XRAM[43608] = 8'b0;
    XRAM[43609] = 8'b0;
    XRAM[43610] = 8'b0;
    XRAM[43611] = 8'b0;
    XRAM[43612] = 8'b0;
    XRAM[43613] = 8'b0;
    XRAM[43614] = 8'b0;
    XRAM[43615] = 8'b0;
    XRAM[43616] = 8'b0;
    XRAM[43617] = 8'b0;
    XRAM[43618] = 8'b0;
    XRAM[43619] = 8'b0;
    XRAM[43620] = 8'b0;
    XRAM[43621] = 8'b0;
    XRAM[43622] = 8'b0;
    XRAM[43623] = 8'b0;
    XRAM[43624] = 8'b0;
    XRAM[43625] = 8'b0;
    XRAM[43626] = 8'b0;
    XRAM[43627] = 8'b0;
    XRAM[43628] = 8'b0;
    XRAM[43629] = 8'b0;
    XRAM[43630] = 8'b0;
    XRAM[43631] = 8'b0;
    XRAM[43632] = 8'b0;
    XRAM[43633] = 8'b0;
    XRAM[43634] = 8'b0;
    XRAM[43635] = 8'b0;
    XRAM[43636] = 8'b0;
    XRAM[43637] = 8'b0;
    XRAM[43638] = 8'b0;
    XRAM[43639] = 8'b0;
    XRAM[43640] = 8'b0;
    XRAM[43641] = 8'b0;
    XRAM[43642] = 8'b0;
    XRAM[43643] = 8'b0;
    XRAM[43644] = 8'b0;
    XRAM[43645] = 8'b0;
    XRAM[43646] = 8'b0;
    XRAM[43647] = 8'b0;
    XRAM[43648] = 8'b0;
    XRAM[43649] = 8'b0;
    XRAM[43650] = 8'b0;
    XRAM[43651] = 8'b0;
    XRAM[43652] = 8'b0;
    XRAM[43653] = 8'b0;
    XRAM[43654] = 8'b0;
    XRAM[43655] = 8'b0;
    XRAM[43656] = 8'b0;
    XRAM[43657] = 8'b0;
    XRAM[43658] = 8'b0;
    XRAM[43659] = 8'b0;
    XRAM[43660] = 8'b0;
    XRAM[43661] = 8'b0;
    XRAM[43662] = 8'b0;
    XRAM[43663] = 8'b0;
    XRAM[43664] = 8'b0;
    XRAM[43665] = 8'b0;
    XRAM[43666] = 8'b0;
    XRAM[43667] = 8'b0;
    XRAM[43668] = 8'b0;
    XRAM[43669] = 8'b0;
    XRAM[43670] = 8'b0;
    XRAM[43671] = 8'b0;
    XRAM[43672] = 8'b0;
    XRAM[43673] = 8'b0;
    XRAM[43674] = 8'b0;
    XRAM[43675] = 8'b0;
    XRAM[43676] = 8'b0;
    XRAM[43677] = 8'b0;
    XRAM[43678] = 8'b0;
    XRAM[43679] = 8'b0;
    XRAM[43680] = 8'b0;
    XRAM[43681] = 8'b0;
    XRAM[43682] = 8'b0;
    XRAM[43683] = 8'b0;
    XRAM[43684] = 8'b0;
    XRAM[43685] = 8'b0;
    XRAM[43686] = 8'b0;
    XRAM[43687] = 8'b0;
    XRAM[43688] = 8'b0;
    XRAM[43689] = 8'b0;
    XRAM[43690] = 8'b0;
    XRAM[43691] = 8'b0;
    XRAM[43692] = 8'b0;
    XRAM[43693] = 8'b0;
    XRAM[43694] = 8'b0;
    XRAM[43695] = 8'b0;
    XRAM[43696] = 8'b0;
    XRAM[43697] = 8'b0;
    XRAM[43698] = 8'b0;
    XRAM[43699] = 8'b0;
    XRAM[43700] = 8'b0;
    XRAM[43701] = 8'b0;
    XRAM[43702] = 8'b0;
    XRAM[43703] = 8'b0;
    XRAM[43704] = 8'b0;
    XRAM[43705] = 8'b0;
    XRAM[43706] = 8'b0;
    XRAM[43707] = 8'b0;
    XRAM[43708] = 8'b0;
    XRAM[43709] = 8'b0;
    XRAM[43710] = 8'b0;
    XRAM[43711] = 8'b0;
    XRAM[43712] = 8'b0;
    XRAM[43713] = 8'b0;
    XRAM[43714] = 8'b0;
    XRAM[43715] = 8'b0;
    XRAM[43716] = 8'b0;
    XRAM[43717] = 8'b0;
    XRAM[43718] = 8'b0;
    XRAM[43719] = 8'b0;
    XRAM[43720] = 8'b0;
    XRAM[43721] = 8'b0;
    XRAM[43722] = 8'b0;
    XRAM[43723] = 8'b0;
    XRAM[43724] = 8'b0;
    XRAM[43725] = 8'b0;
    XRAM[43726] = 8'b0;
    XRAM[43727] = 8'b0;
    XRAM[43728] = 8'b0;
    XRAM[43729] = 8'b0;
    XRAM[43730] = 8'b0;
    XRAM[43731] = 8'b0;
    XRAM[43732] = 8'b0;
    XRAM[43733] = 8'b0;
    XRAM[43734] = 8'b0;
    XRAM[43735] = 8'b0;
    XRAM[43736] = 8'b0;
    XRAM[43737] = 8'b0;
    XRAM[43738] = 8'b0;
    XRAM[43739] = 8'b0;
    XRAM[43740] = 8'b0;
    XRAM[43741] = 8'b0;
    XRAM[43742] = 8'b0;
    XRAM[43743] = 8'b0;
    XRAM[43744] = 8'b0;
    XRAM[43745] = 8'b0;
    XRAM[43746] = 8'b0;
    XRAM[43747] = 8'b0;
    XRAM[43748] = 8'b0;
    XRAM[43749] = 8'b0;
    XRAM[43750] = 8'b0;
    XRAM[43751] = 8'b0;
    XRAM[43752] = 8'b0;
    XRAM[43753] = 8'b0;
    XRAM[43754] = 8'b0;
    XRAM[43755] = 8'b0;
    XRAM[43756] = 8'b0;
    XRAM[43757] = 8'b0;
    XRAM[43758] = 8'b0;
    XRAM[43759] = 8'b0;
    XRAM[43760] = 8'b0;
    XRAM[43761] = 8'b0;
    XRAM[43762] = 8'b0;
    XRAM[43763] = 8'b0;
    XRAM[43764] = 8'b0;
    XRAM[43765] = 8'b0;
    XRAM[43766] = 8'b0;
    XRAM[43767] = 8'b0;
    XRAM[43768] = 8'b0;
    XRAM[43769] = 8'b0;
    XRAM[43770] = 8'b0;
    XRAM[43771] = 8'b0;
    XRAM[43772] = 8'b0;
    XRAM[43773] = 8'b0;
    XRAM[43774] = 8'b0;
    XRAM[43775] = 8'b0;
    XRAM[43776] = 8'b0;
    XRAM[43777] = 8'b0;
    XRAM[43778] = 8'b0;
    XRAM[43779] = 8'b0;
    XRAM[43780] = 8'b0;
    XRAM[43781] = 8'b0;
    XRAM[43782] = 8'b0;
    XRAM[43783] = 8'b0;
    XRAM[43784] = 8'b0;
    XRAM[43785] = 8'b0;
    XRAM[43786] = 8'b0;
    XRAM[43787] = 8'b0;
    XRAM[43788] = 8'b0;
    XRAM[43789] = 8'b0;
    XRAM[43790] = 8'b0;
    XRAM[43791] = 8'b0;
    XRAM[43792] = 8'b0;
    XRAM[43793] = 8'b0;
    XRAM[43794] = 8'b0;
    XRAM[43795] = 8'b0;
    XRAM[43796] = 8'b0;
    XRAM[43797] = 8'b0;
    XRAM[43798] = 8'b0;
    XRAM[43799] = 8'b0;
    XRAM[43800] = 8'b0;
    XRAM[43801] = 8'b0;
    XRAM[43802] = 8'b0;
    XRAM[43803] = 8'b0;
    XRAM[43804] = 8'b0;
    XRAM[43805] = 8'b0;
    XRAM[43806] = 8'b0;
    XRAM[43807] = 8'b0;
    XRAM[43808] = 8'b0;
    XRAM[43809] = 8'b0;
    XRAM[43810] = 8'b0;
    XRAM[43811] = 8'b0;
    XRAM[43812] = 8'b0;
    XRAM[43813] = 8'b0;
    XRAM[43814] = 8'b0;
    XRAM[43815] = 8'b0;
    XRAM[43816] = 8'b0;
    XRAM[43817] = 8'b0;
    XRAM[43818] = 8'b0;
    XRAM[43819] = 8'b0;
    XRAM[43820] = 8'b0;
    XRAM[43821] = 8'b0;
    XRAM[43822] = 8'b0;
    XRAM[43823] = 8'b0;
    XRAM[43824] = 8'b0;
    XRAM[43825] = 8'b0;
    XRAM[43826] = 8'b0;
    XRAM[43827] = 8'b0;
    XRAM[43828] = 8'b0;
    XRAM[43829] = 8'b0;
    XRAM[43830] = 8'b0;
    XRAM[43831] = 8'b0;
    XRAM[43832] = 8'b0;
    XRAM[43833] = 8'b0;
    XRAM[43834] = 8'b0;
    XRAM[43835] = 8'b0;
    XRAM[43836] = 8'b0;
    XRAM[43837] = 8'b0;
    XRAM[43838] = 8'b0;
    XRAM[43839] = 8'b0;
    XRAM[43840] = 8'b0;
    XRAM[43841] = 8'b0;
    XRAM[43842] = 8'b0;
    XRAM[43843] = 8'b0;
    XRAM[43844] = 8'b0;
    XRAM[43845] = 8'b0;
    XRAM[43846] = 8'b0;
    XRAM[43847] = 8'b0;
    XRAM[43848] = 8'b0;
    XRAM[43849] = 8'b0;
    XRAM[43850] = 8'b0;
    XRAM[43851] = 8'b0;
    XRAM[43852] = 8'b0;
    XRAM[43853] = 8'b0;
    XRAM[43854] = 8'b0;
    XRAM[43855] = 8'b0;
    XRAM[43856] = 8'b0;
    XRAM[43857] = 8'b0;
    XRAM[43858] = 8'b0;
    XRAM[43859] = 8'b0;
    XRAM[43860] = 8'b0;
    XRAM[43861] = 8'b0;
    XRAM[43862] = 8'b0;
    XRAM[43863] = 8'b0;
    XRAM[43864] = 8'b0;
    XRAM[43865] = 8'b0;
    XRAM[43866] = 8'b0;
    XRAM[43867] = 8'b0;
    XRAM[43868] = 8'b0;
    XRAM[43869] = 8'b0;
    XRAM[43870] = 8'b0;
    XRAM[43871] = 8'b0;
    XRAM[43872] = 8'b0;
    XRAM[43873] = 8'b0;
    XRAM[43874] = 8'b0;
    XRAM[43875] = 8'b0;
    XRAM[43876] = 8'b0;
    XRAM[43877] = 8'b0;
    XRAM[43878] = 8'b0;
    XRAM[43879] = 8'b0;
    XRAM[43880] = 8'b0;
    XRAM[43881] = 8'b0;
    XRAM[43882] = 8'b0;
    XRAM[43883] = 8'b0;
    XRAM[43884] = 8'b0;
    XRAM[43885] = 8'b0;
    XRAM[43886] = 8'b0;
    XRAM[43887] = 8'b0;
    XRAM[43888] = 8'b0;
    XRAM[43889] = 8'b0;
    XRAM[43890] = 8'b0;
    XRAM[43891] = 8'b0;
    XRAM[43892] = 8'b0;
    XRAM[43893] = 8'b0;
    XRAM[43894] = 8'b0;
    XRAM[43895] = 8'b0;
    XRAM[43896] = 8'b0;
    XRAM[43897] = 8'b0;
    XRAM[43898] = 8'b0;
    XRAM[43899] = 8'b0;
    XRAM[43900] = 8'b0;
    XRAM[43901] = 8'b0;
    XRAM[43902] = 8'b0;
    XRAM[43903] = 8'b0;
    XRAM[43904] = 8'b0;
    XRAM[43905] = 8'b0;
    XRAM[43906] = 8'b0;
    XRAM[43907] = 8'b0;
    XRAM[43908] = 8'b0;
    XRAM[43909] = 8'b0;
    XRAM[43910] = 8'b0;
    XRAM[43911] = 8'b0;
    XRAM[43912] = 8'b0;
    XRAM[43913] = 8'b0;
    XRAM[43914] = 8'b0;
    XRAM[43915] = 8'b0;
    XRAM[43916] = 8'b0;
    XRAM[43917] = 8'b0;
    XRAM[43918] = 8'b0;
    XRAM[43919] = 8'b0;
    XRAM[43920] = 8'b0;
    XRAM[43921] = 8'b0;
    XRAM[43922] = 8'b0;
    XRAM[43923] = 8'b0;
    XRAM[43924] = 8'b0;
    XRAM[43925] = 8'b0;
    XRAM[43926] = 8'b0;
    XRAM[43927] = 8'b0;
    XRAM[43928] = 8'b0;
    XRAM[43929] = 8'b0;
    XRAM[43930] = 8'b0;
    XRAM[43931] = 8'b0;
    XRAM[43932] = 8'b0;
    XRAM[43933] = 8'b0;
    XRAM[43934] = 8'b0;
    XRAM[43935] = 8'b0;
    XRAM[43936] = 8'b0;
    XRAM[43937] = 8'b0;
    XRAM[43938] = 8'b0;
    XRAM[43939] = 8'b0;
    XRAM[43940] = 8'b0;
    XRAM[43941] = 8'b0;
    XRAM[43942] = 8'b0;
    XRAM[43943] = 8'b0;
    XRAM[43944] = 8'b0;
    XRAM[43945] = 8'b0;
    XRAM[43946] = 8'b0;
    XRAM[43947] = 8'b0;
    XRAM[43948] = 8'b0;
    XRAM[43949] = 8'b0;
    XRAM[43950] = 8'b0;
    XRAM[43951] = 8'b0;
    XRAM[43952] = 8'b0;
    XRAM[43953] = 8'b0;
    XRAM[43954] = 8'b0;
    XRAM[43955] = 8'b0;
    XRAM[43956] = 8'b0;
    XRAM[43957] = 8'b0;
    XRAM[43958] = 8'b0;
    XRAM[43959] = 8'b0;
    XRAM[43960] = 8'b0;
    XRAM[43961] = 8'b0;
    XRAM[43962] = 8'b0;
    XRAM[43963] = 8'b0;
    XRAM[43964] = 8'b0;
    XRAM[43965] = 8'b0;
    XRAM[43966] = 8'b0;
    XRAM[43967] = 8'b0;
    XRAM[43968] = 8'b0;
    XRAM[43969] = 8'b0;
    XRAM[43970] = 8'b0;
    XRAM[43971] = 8'b0;
    XRAM[43972] = 8'b0;
    XRAM[43973] = 8'b0;
    XRAM[43974] = 8'b0;
    XRAM[43975] = 8'b0;
    XRAM[43976] = 8'b0;
    XRAM[43977] = 8'b0;
    XRAM[43978] = 8'b0;
    XRAM[43979] = 8'b0;
    XRAM[43980] = 8'b0;
    XRAM[43981] = 8'b0;
    XRAM[43982] = 8'b0;
    XRAM[43983] = 8'b0;
    XRAM[43984] = 8'b0;
    XRAM[43985] = 8'b0;
    XRAM[43986] = 8'b0;
    XRAM[43987] = 8'b0;
    XRAM[43988] = 8'b0;
    XRAM[43989] = 8'b0;
    XRAM[43990] = 8'b0;
    XRAM[43991] = 8'b0;
    XRAM[43992] = 8'b0;
    XRAM[43993] = 8'b0;
    XRAM[43994] = 8'b0;
    XRAM[43995] = 8'b0;
    XRAM[43996] = 8'b0;
    XRAM[43997] = 8'b0;
    XRAM[43998] = 8'b0;
    XRAM[43999] = 8'b0;
    XRAM[44000] = 8'b0;
    XRAM[44001] = 8'b0;
    XRAM[44002] = 8'b0;
    XRAM[44003] = 8'b0;
    XRAM[44004] = 8'b0;
    XRAM[44005] = 8'b0;
    XRAM[44006] = 8'b0;
    XRAM[44007] = 8'b0;
    XRAM[44008] = 8'b0;
    XRAM[44009] = 8'b0;
    XRAM[44010] = 8'b0;
    XRAM[44011] = 8'b0;
    XRAM[44012] = 8'b0;
    XRAM[44013] = 8'b0;
    XRAM[44014] = 8'b0;
    XRAM[44015] = 8'b0;
    XRAM[44016] = 8'b0;
    XRAM[44017] = 8'b0;
    XRAM[44018] = 8'b0;
    XRAM[44019] = 8'b0;
    XRAM[44020] = 8'b0;
    XRAM[44021] = 8'b0;
    XRAM[44022] = 8'b0;
    XRAM[44023] = 8'b0;
    XRAM[44024] = 8'b0;
    XRAM[44025] = 8'b0;
    XRAM[44026] = 8'b0;
    XRAM[44027] = 8'b0;
    XRAM[44028] = 8'b0;
    XRAM[44029] = 8'b0;
    XRAM[44030] = 8'b0;
    XRAM[44031] = 8'b0;
    XRAM[44032] = 8'b0;
    XRAM[44033] = 8'b0;
    XRAM[44034] = 8'b0;
    XRAM[44035] = 8'b0;
    XRAM[44036] = 8'b0;
    XRAM[44037] = 8'b0;
    XRAM[44038] = 8'b0;
    XRAM[44039] = 8'b0;
    XRAM[44040] = 8'b0;
    XRAM[44041] = 8'b0;
    XRAM[44042] = 8'b0;
    XRAM[44043] = 8'b0;
    XRAM[44044] = 8'b0;
    XRAM[44045] = 8'b0;
    XRAM[44046] = 8'b0;
    XRAM[44047] = 8'b0;
    XRAM[44048] = 8'b0;
    XRAM[44049] = 8'b0;
    XRAM[44050] = 8'b0;
    XRAM[44051] = 8'b0;
    XRAM[44052] = 8'b0;
    XRAM[44053] = 8'b0;
    XRAM[44054] = 8'b0;
    XRAM[44055] = 8'b0;
    XRAM[44056] = 8'b0;
    XRAM[44057] = 8'b0;
    XRAM[44058] = 8'b0;
    XRAM[44059] = 8'b0;
    XRAM[44060] = 8'b0;
    XRAM[44061] = 8'b0;
    XRAM[44062] = 8'b0;
    XRAM[44063] = 8'b0;
    XRAM[44064] = 8'b0;
    XRAM[44065] = 8'b0;
    XRAM[44066] = 8'b0;
    XRAM[44067] = 8'b0;
    XRAM[44068] = 8'b0;
    XRAM[44069] = 8'b0;
    XRAM[44070] = 8'b0;
    XRAM[44071] = 8'b0;
    XRAM[44072] = 8'b0;
    XRAM[44073] = 8'b0;
    XRAM[44074] = 8'b0;
    XRAM[44075] = 8'b0;
    XRAM[44076] = 8'b0;
    XRAM[44077] = 8'b0;
    XRAM[44078] = 8'b0;
    XRAM[44079] = 8'b0;
    XRAM[44080] = 8'b0;
    XRAM[44081] = 8'b0;
    XRAM[44082] = 8'b0;
    XRAM[44083] = 8'b0;
    XRAM[44084] = 8'b0;
    XRAM[44085] = 8'b0;
    XRAM[44086] = 8'b0;
    XRAM[44087] = 8'b0;
    XRAM[44088] = 8'b0;
    XRAM[44089] = 8'b0;
    XRAM[44090] = 8'b0;
    XRAM[44091] = 8'b0;
    XRAM[44092] = 8'b0;
    XRAM[44093] = 8'b0;
    XRAM[44094] = 8'b0;
    XRAM[44095] = 8'b0;
    XRAM[44096] = 8'b0;
    XRAM[44097] = 8'b0;
    XRAM[44098] = 8'b0;
    XRAM[44099] = 8'b0;
    XRAM[44100] = 8'b0;
    XRAM[44101] = 8'b0;
    XRAM[44102] = 8'b0;
    XRAM[44103] = 8'b0;
    XRAM[44104] = 8'b0;
    XRAM[44105] = 8'b0;
    XRAM[44106] = 8'b0;
    XRAM[44107] = 8'b0;
    XRAM[44108] = 8'b0;
    XRAM[44109] = 8'b0;
    XRAM[44110] = 8'b0;
    XRAM[44111] = 8'b0;
    XRAM[44112] = 8'b0;
    XRAM[44113] = 8'b0;
    XRAM[44114] = 8'b0;
    XRAM[44115] = 8'b0;
    XRAM[44116] = 8'b0;
    XRAM[44117] = 8'b0;
    XRAM[44118] = 8'b0;
    XRAM[44119] = 8'b0;
    XRAM[44120] = 8'b0;
    XRAM[44121] = 8'b0;
    XRAM[44122] = 8'b0;
    XRAM[44123] = 8'b0;
    XRAM[44124] = 8'b0;
    XRAM[44125] = 8'b0;
    XRAM[44126] = 8'b0;
    XRAM[44127] = 8'b0;
    XRAM[44128] = 8'b0;
    XRAM[44129] = 8'b0;
    XRAM[44130] = 8'b0;
    XRAM[44131] = 8'b0;
    XRAM[44132] = 8'b0;
    XRAM[44133] = 8'b0;
    XRAM[44134] = 8'b0;
    XRAM[44135] = 8'b0;
    XRAM[44136] = 8'b0;
    XRAM[44137] = 8'b0;
    XRAM[44138] = 8'b0;
    XRAM[44139] = 8'b0;
    XRAM[44140] = 8'b0;
    XRAM[44141] = 8'b0;
    XRAM[44142] = 8'b0;
    XRAM[44143] = 8'b0;
    XRAM[44144] = 8'b0;
    XRAM[44145] = 8'b0;
    XRAM[44146] = 8'b0;
    XRAM[44147] = 8'b0;
    XRAM[44148] = 8'b0;
    XRAM[44149] = 8'b0;
    XRAM[44150] = 8'b0;
    XRAM[44151] = 8'b0;
    XRAM[44152] = 8'b0;
    XRAM[44153] = 8'b0;
    XRAM[44154] = 8'b0;
    XRAM[44155] = 8'b0;
    XRAM[44156] = 8'b0;
    XRAM[44157] = 8'b0;
    XRAM[44158] = 8'b0;
    XRAM[44159] = 8'b0;
    XRAM[44160] = 8'b0;
    XRAM[44161] = 8'b0;
    XRAM[44162] = 8'b0;
    XRAM[44163] = 8'b0;
    XRAM[44164] = 8'b0;
    XRAM[44165] = 8'b0;
    XRAM[44166] = 8'b0;
    XRAM[44167] = 8'b0;
    XRAM[44168] = 8'b0;
    XRAM[44169] = 8'b0;
    XRAM[44170] = 8'b0;
    XRAM[44171] = 8'b0;
    XRAM[44172] = 8'b0;
    XRAM[44173] = 8'b0;
    XRAM[44174] = 8'b0;
    XRAM[44175] = 8'b0;
    XRAM[44176] = 8'b0;
    XRAM[44177] = 8'b0;
    XRAM[44178] = 8'b0;
    XRAM[44179] = 8'b0;
    XRAM[44180] = 8'b0;
    XRAM[44181] = 8'b0;
    XRAM[44182] = 8'b0;
    XRAM[44183] = 8'b0;
    XRAM[44184] = 8'b0;
    XRAM[44185] = 8'b0;
    XRAM[44186] = 8'b0;
    XRAM[44187] = 8'b0;
    XRAM[44188] = 8'b0;
    XRAM[44189] = 8'b0;
    XRAM[44190] = 8'b0;
    XRAM[44191] = 8'b0;
    XRAM[44192] = 8'b0;
    XRAM[44193] = 8'b0;
    XRAM[44194] = 8'b0;
    XRAM[44195] = 8'b0;
    XRAM[44196] = 8'b0;
    XRAM[44197] = 8'b0;
    XRAM[44198] = 8'b0;
    XRAM[44199] = 8'b0;
    XRAM[44200] = 8'b0;
    XRAM[44201] = 8'b0;
    XRAM[44202] = 8'b0;
    XRAM[44203] = 8'b0;
    XRAM[44204] = 8'b0;
    XRAM[44205] = 8'b0;
    XRAM[44206] = 8'b0;
    XRAM[44207] = 8'b0;
    XRAM[44208] = 8'b0;
    XRAM[44209] = 8'b0;
    XRAM[44210] = 8'b0;
    XRAM[44211] = 8'b0;
    XRAM[44212] = 8'b0;
    XRAM[44213] = 8'b0;
    XRAM[44214] = 8'b0;
    XRAM[44215] = 8'b0;
    XRAM[44216] = 8'b0;
    XRAM[44217] = 8'b0;
    XRAM[44218] = 8'b0;
    XRAM[44219] = 8'b0;
    XRAM[44220] = 8'b0;
    XRAM[44221] = 8'b0;
    XRAM[44222] = 8'b0;
    XRAM[44223] = 8'b0;
    XRAM[44224] = 8'b0;
    XRAM[44225] = 8'b0;
    XRAM[44226] = 8'b0;
    XRAM[44227] = 8'b0;
    XRAM[44228] = 8'b0;
    XRAM[44229] = 8'b0;
    XRAM[44230] = 8'b0;
    XRAM[44231] = 8'b0;
    XRAM[44232] = 8'b0;
    XRAM[44233] = 8'b0;
    XRAM[44234] = 8'b0;
    XRAM[44235] = 8'b0;
    XRAM[44236] = 8'b0;
    XRAM[44237] = 8'b0;
    XRAM[44238] = 8'b0;
    XRAM[44239] = 8'b0;
    XRAM[44240] = 8'b0;
    XRAM[44241] = 8'b0;
    XRAM[44242] = 8'b0;
    XRAM[44243] = 8'b0;
    XRAM[44244] = 8'b0;
    XRAM[44245] = 8'b0;
    XRAM[44246] = 8'b0;
    XRAM[44247] = 8'b0;
    XRAM[44248] = 8'b0;
    XRAM[44249] = 8'b0;
    XRAM[44250] = 8'b0;
    XRAM[44251] = 8'b0;
    XRAM[44252] = 8'b0;
    XRAM[44253] = 8'b0;
    XRAM[44254] = 8'b0;
    XRAM[44255] = 8'b0;
    XRAM[44256] = 8'b0;
    XRAM[44257] = 8'b0;
    XRAM[44258] = 8'b0;
    XRAM[44259] = 8'b0;
    XRAM[44260] = 8'b0;
    XRAM[44261] = 8'b0;
    XRAM[44262] = 8'b0;
    XRAM[44263] = 8'b0;
    XRAM[44264] = 8'b0;
    XRAM[44265] = 8'b0;
    XRAM[44266] = 8'b0;
    XRAM[44267] = 8'b0;
    XRAM[44268] = 8'b0;
    XRAM[44269] = 8'b0;
    XRAM[44270] = 8'b0;
    XRAM[44271] = 8'b0;
    XRAM[44272] = 8'b0;
    XRAM[44273] = 8'b0;
    XRAM[44274] = 8'b0;
    XRAM[44275] = 8'b0;
    XRAM[44276] = 8'b0;
    XRAM[44277] = 8'b0;
    XRAM[44278] = 8'b0;
    XRAM[44279] = 8'b0;
    XRAM[44280] = 8'b0;
    XRAM[44281] = 8'b0;
    XRAM[44282] = 8'b0;
    XRAM[44283] = 8'b0;
    XRAM[44284] = 8'b0;
    XRAM[44285] = 8'b0;
    XRAM[44286] = 8'b0;
    XRAM[44287] = 8'b0;
    XRAM[44288] = 8'b0;
    XRAM[44289] = 8'b0;
    XRAM[44290] = 8'b0;
    XRAM[44291] = 8'b0;
    XRAM[44292] = 8'b0;
    XRAM[44293] = 8'b0;
    XRAM[44294] = 8'b0;
    XRAM[44295] = 8'b0;
    XRAM[44296] = 8'b0;
    XRAM[44297] = 8'b0;
    XRAM[44298] = 8'b0;
    XRAM[44299] = 8'b0;
    XRAM[44300] = 8'b0;
    XRAM[44301] = 8'b0;
    XRAM[44302] = 8'b0;
    XRAM[44303] = 8'b0;
    XRAM[44304] = 8'b0;
    XRAM[44305] = 8'b0;
    XRAM[44306] = 8'b0;
    XRAM[44307] = 8'b0;
    XRAM[44308] = 8'b0;
    XRAM[44309] = 8'b0;
    XRAM[44310] = 8'b0;
    XRAM[44311] = 8'b0;
    XRAM[44312] = 8'b0;
    XRAM[44313] = 8'b0;
    XRAM[44314] = 8'b0;
    XRAM[44315] = 8'b0;
    XRAM[44316] = 8'b0;
    XRAM[44317] = 8'b0;
    XRAM[44318] = 8'b0;
    XRAM[44319] = 8'b0;
    XRAM[44320] = 8'b0;
    XRAM[44321] = 8'b0;
    XRAM[44322] = 8'b0;
    XRAM[44323] = 8'b0;
    XRAM[44324] = 8'b0;
    XRAM[44325] = 8'b0;
    XRAM[44326] = 8'b0;
    XRAM[44327] = 8'b0;
    XRAM[44328] = 8'b0;
    XRAM[44329] = 8'b0;
    XRAM[44330] = 8'b0;
    XRAM[44331] = 8'b0;
    XRAM[44332] = 8'b0;
    XRAM[44333] = 8'b0;
    XRAM[44334] = 8'b0;
    XRAM[44335] = 8'b0;
    XRAM[44336] = 8'b0;
    XRAM[44337] = 8'b0;
    XRAM[44338] = 8'b0;
    XRAM[44339] = 8'b0;
    XRAM[44340] = 8'b0;
    XRAM[44341] = 8'b0;
    XRAM[44342] = 8'b0;
    XRAM[44343] = 8'b0;
    XRAM[44344] = 8'b0;
    XRAM[44345] = 8'b0;
    XRAM[44346] = 8'b0;
    XRAM[44347] = 8'b0;
    XRAM[44348] = 8'b0;
    XRAM[44349] = 8'b0;
    XRAM[44350] = 8'b0;
    XRAM[44351] = 8'b0;
    XRAM[44352] = 8'b0;
    XRAM[44353] = 8'b0;
    XRAM[44354] = 8'b0;
    XRAM[44355] = 8'b0;
    XRAM[44356] = 8'b0;
    XRAM[44357] = 8'b0;
    XRAM[44358] = 8'b0;
    XRAM[44359] = 8'b0;
    XRAM[44360] = 8'b0;
    XRAM[44361] = 8'b0;
    XRAM[44362] = 8'b0;
    XRAM[44363] = 8'b0;
    XRAM[44364] = 8'b0;
    XRAM[44365] = 8'b0;
    XRAM[44366] = 8'b0;
    XRAM[44367] = 8'b0;
    XRAM[44368] = 8'b0;
    XRAM[44369] = 8'b0;
    XRAM[44370] = 8'b0;
    XRAM[44371] = 8'b0;
    XRAM[44372] = 8'b0;
    XRAM[44373] = 8'b0;
    XRAM[44374] = 8'b0;
    XRAM[44375] = 8'b0;
    XRAM[44376] = 8'b0;
    XRAM[44377] = 8'b0;
    XRAM[44378] = 8'b0;
    XRAM[44379] = 8'b0;
    XRAM[44380] = 8'b0;
    XRAM[44381] = 8'b0;
    XRAM[44382] = 8'b0;
    XRAM[44383] = 8'b0;
    XRAM[44384] = 8'b0;
    XRAM[44385] = 8'b0;
    XRAM[44386] = 8'b0;
    XRAM[44387] = 8'b0;
    XRAM[44388] = 8'b0;
    XRAM[44389] = 8'b0;
    XRAM[44390] = 8'b0;
    XRAM[44391] = 8'b0;
    XRAM[44392] = 8'b0;
    XRAM[44393] = 8'b0;
    XRAM[44394] = 8'b0;
    XRAM[44395] = 8'b0;
    XRAM[44396] = 8'b0;
    XRAM[44397] = 8'b0;
    XRAM[44398] = 8'b0;
    XRAM[44399] = 8'b0;
    XRAM[44400] = 8'b0;
    XRAM[44401] = 8'b0;
    XRAM[44402] = 8'b0;
    XRAM[44403] = 8'b0;
    XRAM[44404] = 8'b0;
    XRAM[44405] = 8'b0;
    XRAM[44406] = 8'b0;
    XRAM[44407] = 8'b0;
    XRAM[44408] = 8'b0;
    XRAM[44409] = 8'b0;
    XRAM[44410] = 8'b0;
    XRAM[44411] = 8'b0;
    XRAM[44412] = 8'b0;
    XRAM[44413] = 8'b0;
    XRAM[44414] = 8'b0;
    XRAM[44415] = 8'b0;
    XRAM[44416] = 8'b0;
    XRAM[44417] = 8'b0;
    XRAM[44418] = 8'b0;
    XRAM[44419] = 8'b0;
    XRAM[44420] = 8'b0;
    XRAM[44421] = 8'b0;
    XRAM[44422] = 8'b0;
    XRAM[44423] = 8'b0;
    XRAM[44424] = 8'b0;
    XRAM[44425] = 8'b0;
    XRAM[44426] = 8'b0;
    XRAM[44427] = 8'b0;
    XRAM[44428] = 8'b0;
    XRAM[44429] = 8'b0;
    XRAM[44430] = 8'b0;
    XRAM[44431] = 8'b0;
    XRAM[44432] = 8'b0;
    XRAM[44433] = 8'b0;
    XRAM[44434] = 8'b0;
    XRAM[44435] = 8'b0;
    XRAM[44436] = 8'b0;
    XRAM[44437] = 8'b0;
    XRAM[44438] = 8'b0;
    XRAM[44439] = 8'b0;
    XRAM[44440] = 8'b0;
    XRAM[44441] = 8'b0;
    XRAM[44442] = 8'b0;
    XRAM[44443] = 8'b0;
    XRAM[44444] = 8'b0;
    XRAM[44445] = 8'b0;
    XRAM[44446] = 8'b0;
    XRAM[44447] = 8'b0;
    XRAM[44448] = 8'b0;
    XRAM[44449] = 8'b0;
    XRAM[44450] = 8'b0;
    XRAM[44451] = 8'b0;
    XRAM[44452] = 8'b0;
    XRAM[44453] = 8'b0;
    XRAM[44454] = 8'b0;
    XRAM[44455] = 8'b0;
    XRAM[44456] = 8'b0;
    XRAM[44457] = 8'b0;
    XRAM[44458] = 8'b0;
    XRAM[44459] = 8'b0;
    XRAM[44460] = 8'b0;
    XRAM[44461] = 8'b0;
    XRAM[44462] = 8'b0;
    XRAM[44463] = 8'b0;
    XRAM[44464] = 8'b0;
    XRAM[44465] = 8'b0;
    XRAM[44466] = 8'b0;
    XRAM[44467] = 8'b0;
    XRAM[44468] = 8'b0;
    XRAM[44469] = 8'b0;
    XRAM[44470] = 8'b0;
    XRAM[44471] = 8'b0;
    XRAM[44472] = 8'b0;
    XRAM[44473] = 8'b0;
    XRAM[44474] = 8'b0;
    XRAM[44475] = 8'b0;
    XRAM[44476] = 8'b0;
    XRAM[44477] = 8'b0;
    XRAM[44478] = 8'b0;
    XRAM[44479] = 8'b0;
    XRAM[44480] = 8'b0;
    XRAM[44481] = 8'b0;
    XRAM[44482] = 8'b0;
    XRAM[44483] = 8'b0;
    XRAM[44484] = 8'b0;
    XRAM[44485] = 8'b0;
    XRAM[44486] = 8'b0;
    XRAM[44487] = 8'b0;
    XRAM[44488] = 8'b0;
    XRAM[44489] = 8'b0;
    XRAM[44490] = 8'b0;
    XRAM[44491] = 8'b0;
    XRAM[44492] = 8'b0;
    XRAM[44493] = 8'b0;
    XRAM[44494] = 8'b0;
    XRAM[44495] = 8'b0;
    XRAM[44496] = 8'b0;
    XRAM[44497] = 8'b0;
    XRAM[44498] = 8'b0;
    XRAM[44499] = 8'b0;
    XRAM[44500] = 8'b0;
    XRAM[44501] = 8'b0;
    XRAM[44502] = 8'b0;
    XRAM[44503] = 8'b0;
    XRAM[44504] = 8'b0;
    XRAM[44505] = 8'b0;
    XRAM[44506] = 8'b0;
    XRAM[44507] = 8'b0;
    XRAM[44508] = 8'b0;
    XRAM[44509] = 8'b0;
    XRAM[44510] = 8'b0;
    XRAM[44511] = 8'b0;
    XRAM[44512] = 8'b0;
    XRAM[44513] = 8'b0;
    XRAM[44514] = 8'b0;
    XRAM[44515] = 8'b0;
    XRAM[44516] = 8'b0;
    XRAM[44517] = 8'b0;
    XRAM[44518] = 8'b0;
    XRAM[44519] = 8'b0;
    XRAM[44520] = 8'b0;
    XRAM[44521] = 8'b0;
    XRAM[44522] = 8'b0;
    XRAM[44523] = 8'b0;
    XRAM[44524] = 8'b0;
    XRAM[44525] = 8'b0;
    XRAM[44526] = 8'b0;
    XRAM[44527] = 8'b0;
    XRAM[44528] = 8'b0;
    XRAM[44529] = 8'b0;
    XRAM[44530] = 8'b0;
    XRAM[44531] = 8'b0;
    XRAM[44532] = 8'b0;
    XRAM[44533] = 8'b0;
    XRAM[44534] = 8'b0;
    XRAM[44535] = 8'b0;
    XRAM[44536] = 8'b0;
    XRAM[44537] = 8'b0;
    XRAM[44538] = 8'b0;
    XRAM[44539] = 8'b0;
    XRAM[44540] = 8'b0;
    XRAM[44541] = 8'b0;
    XRAM[44542] = 8'b0;
    XRAM[44543] = 8'b0;
    XRAM[44544] = 8'b0;
    XRAM[44545] = 8'b0;
    XRAM[44546] = 8'b0;
    XRAM[44547] = 8'b0;
    XRAM[44548] = 8'b0;
    XRAM[44549] = 8'b0;
    XRAM[44550] = 8'b0;
    XRAM[44551] = 8'b0;
    XRAM[44552] = 8'b0;
    XRAM[44553] = 8'b0;
    XRAM[44554] = 8'b0;
    XRAM[44555] = 8'b0;
    XRAM[44556] = 8'b0;
    XRAM[44557] = 8'b0;
    XRAM[44558] = 8'b0;
    XRAM[44559] = 8'b0;
    XRAM[44560] = 8'b0;
    XRAM[44561] = 8'b0;
    XRAM[44562] = 8'b0;
    XRAM[44563] = 8'b0;
    XRAM[44564] = 8'b0;
    XRAM[44565] = 8'b0;
    XRAM[44566] = 8'b0;
    XRAM[44567] = 8'b0;
    XRAM[44568] = 8'b0;
    XRAM[44569] = 8'b0;
    XRAM[44570] = 8'b0;
    XRAM[44571] = 8'b0;
    XRAM[44572] = 8'b0;
    XRAM[44573] = 8'b0;
    XRAM[44574] = 8'b0;
    XRAM[44575] = 8'b0;
    XRAM[44576] = 8'b0;
    XRAM[44577] = 8'b0;
    XRAM[44578] = 8'b0;
    XRAM[44579] = 8'b0;
    XRAM[44580] = 8'b0;
    XRAM[44581] = 8'b0;
    XRAM[44582] = 8'b0;
    XRAM[44583] = 8'b0;
    XRAM[44584] = 8'b0;
    XRAM[44585] = 8'b0;
    XRAM[44586] = 8'b0;
    XRAM[44587] = 8'b0;
    XRAM[44588] = 8'b0;
    XRAM[44589] = 8'b0;
    XRAM[44590] = 8'b0;
    XRAM[44591] = 8'b0;
    XRAM[44592] = 8'b0;
    XRAM[44593] = 8'b0;
    XRAM[44594] = 8'b0;
    XRAM[44595] = 8'b0;
    XRAM[44596] = 8'b0;
    XRAM[44597] = 8'b0;
    XRAM[44598] = 8'b0;
    XRAM[44599] = 8'b0;
    XRAM[44600] = 8'b0;
    XRAM[44601] = 8'b0;
    XRAM[44602] = 8'b0;
    XRAM[44603] = 8'b0;
    XRAM[44604] = 8'b0;
    XRAM[44605] = 8'b0;
    XRAM[44606] = 8'b0;
    XRAM[44607] = 8'b0;
    XRAM[44608] = 8'b0;
    XRAM[44609] = 8'b0;
    XRAM[44610] = 8'b0;
    XRAM[44611] = 8'b0;
    XRAM[44612] = 8'b0;
    XRAM[44613] = 8'b0;
    XRAM[44614] = 8'b0;
    XRAM[44615] = 8'b0;
    XRAM[44616] = 8'b0;
    XRAM[44617] = 8'b0;
    XRAM[44618] = 8'b0;
    XRAM[44619] = 8'b0;
    XRAM[44620] = 8'b0;
    XRAM[44621] = 8'b0;
    XRAM[44622] = 8'b0;
    XRAM[44623] = 8'b0;
    XRAM[44624] = 8'b0;
    XRAM[44625] = 8'b0;
    XRAM[44626] = 8'b0;
    XRAM[44627] = 8'b0;
    XRAM[44628] = 8'b0;
    XRAM[44629] = 8'b0;
    XRAM[44630] = 8'b0;
    XRAM[44631] = 8'b0;
    XRAM[44632] = 8'b0;
    XRAM[44633] = 8'b0;
    XRAM[44634] = 8'b0;
    XRAM[44635] = 8'b0;
    XRAM[44636] = 8'b0;
    XRAM[44637] = 8'b0;
    XRAM[44638] = 8'b0;
    XRAM[44639] = 8'b0;
    XRAM[44640] = 8'b0;
    XRAM[44641] = 8'b0;
    XRAM[44642] = 8'b0;
    XRAM[44643] = 8'b0;
    XRAM[44644] = 8'b0;
    XRAM[44645] = 8'b0;
    XRAM[44646] = 8'b0;
    XRAM[44647] = 8'b0;
    XRAM[44648] = 8'b0;
    XRAM[44649] = 8'b0;
    XRAM[44650] = 8'b0;
    XRAM[44651] = 8'b0;
    XRAM[44652] = 8'b0;
    XRAM[44653] = 8'b0;
    XRAM[44654] = 8'b0;
    XRAM[44655] = 8'b0;
    XRAM[44656] = 8'b0;
    XRAM[44657] = 8'b0;
    XRAM[44658] = 8'b0;
    XRAM[44659] = 8'b0;
    XRAM[44660] = 8'b0;
    XRAM[44661] = 8'b0;
    XRAM[44662] = 8'b0;
    XRAM[44663] = 8'b0;
    XRAM[44664] = 8'b0;
    XRAM[44665] = 8'b0;
    XRAM[44666] = 8'b0;
    XRAM[44667] = 8'b0;
    XRAM[44668] = 8'b0;
    XRAM[44669] = 8'b0;
    XRAM[44670] = 8'b0;
    XRAM[44671] = 8'b0;
    XRAM[44672] = 8'b0;
    XRAM[44673] = 8'b0;
    XRAM[44674] = 8'b0;
    XRAM[44675] = 8'b0;
    XRAM[44676] = 8'b0;
    XRAM[44677] = 8'b0;
    XRAM[44678] = 8'b0;
    XRAM[44679] = 8'b0;
    XRAM[44680] = 8'b0;
    XRAM[44681] = 8'b0;
    XRAM[44682] = 8'b0;
    XRAM[44683] = 8'b0;
    XRAM[44684] = 8'b0;
    XRAM[44685] = 8'b0;
    XRAM[44686] = 8'b0;
    XRAM[44687] = 8'b0;
    XRAM[44688] = 8'b0;
    XRAM[44689] = 8'b0;
    XRAM[44690] = 8'b0;
    XRAM[44691] = 8'b0;
    XRAM[44692] = 8'b0;
    XRAM[44693] = 8'b0;
    XRAM[44694] = 8'b0;
    XRAM[44695] = 8'b0;
    XRAM[44696] = 8'b0;
    XRAM[44697] = 8'b0;
    XRAM[44698] = 8'b0;
    XRAM[44699] = 8'b0;
    XRAM[44700] = 8'b0;
    XRAM[44701] = 8'b0;
    XRAM[44702] = 8'b0;
    XRAM[44703] = 8'b0;
    XRAM[44704] = 8'b0;
    XRAM[44705] = 8'b0;
    XRAM[44706] = 8'b0;
    XRAM[44707] = 8'b0;
    XRAM[44708] = 8'b0;
    XRAM[44709] = 8'b0;
    XRAM[44710] = 8'b0;
    XRAM[44711] = 8'b0;
    XRAM[44712] = 8'b0;
    XRAM[44713] = 8'b0;
    XRAM[44714] = 8'b0;
    XRAM[44715] = 8'b0;
    XRAM[44716] = 8'b0;
    XRAM[44717] = 8'b0;
    XRAM[44718] = 8'b0;
    XRAM[44719] = 8'b0;
    XRAM[44720] = 8'b0;
    XRAM[44721] = 8'b0;
    XRAM[44722] = 8'b0;
    XRAM[44723] = 8'b0;
    XRAM[44724] = 8'b0;
    XRAM[44725] = 8'b0;
    XRAM[44726] = 8'b0;
    XRAM[44727] = 8'b0;
    XRAM[44728] = 8'b0;
    XRAM[44729] = 8'b0;
    XRAM[44730] = 8'b0;
    XRAM[44731] = 8'b0;
    XRAM[44732] = 8'b0;
    XRAM[44733] = 8'b0;
    XRAM[44734] = 8'b0;
    XRAM[44735] = 8'b0;
    XRAM[44736] = 8'b0;
    XRAM[44737] = 8'b0;
    XRAM[44738] = 8'b0;
    XRAM[44739] = 8'b0;
    XRAM[44740] = 8'b0;
    XRAM[44741] = 8'b0;
    XRAM[44742] = 8'b0;
    XRAM[44743] = 8'b0;
    XRAM[44744] = 8'b0;
    XRAM[44745] = 8'b0;
    XRAM[44746] = 8'b0;
    XRAM[44747] = 8'b0;
    XRAM[44748] = 8'b0;
    XRAM[44749] = 8'b0;
    XRAM[44750] = 8'b0;
    XRAM[44751] = 8'b0;
    XRAM[44752] = 8'b0;
    XRAM[44753] = 8'b0;
    XRAM[44754] = 8'b0;
    XRAM[44755] = 8'b0;
    XRAM[44756] = 8'b0;
    XRAM[44757] = 8'b0;
    XRAM[44758] = 8'b0;
    XRAM[44759] = 8'b0;
    XRAM[44760] = 8'b0;
    XRAM[44761] = 8'b0;
    XRAM[44762] = 8'b0;
    XRAM[44763] = 8'b0;
    XRAM[44764] = 8'b0;
    XRAM[44765] = 8'b0;
    XRAM[44766] = 8'b0;
    XRAM[44767] = 8'b0;
    XRAM[44768] = 8'b0;
    XRAM[44769] = 8'b0;
    XRAM[44770] = 8'b0;
    XRAM[44771] = 8'b0;
    XRAM[44772] = 8'b0;
    XRAM[44773] = 8'b0;
    XRAM[44774] = 8'b0;
    XRAM[44775] = 8'b0;
    XRAM[44776] = 8'b0;
    XRAM[44777] = 8'b0;
    XRAM[44778] = 8'b0;
    XRAM[44779] = 8'b0;
    XRAM[44780] = 8'b0;
    XRAM[44781] = 8'b0;
    XRAM[44782] = 8'b0;
    XRAM[44783] = 8'b0;
    XRAM[44784] = 8'b0;
    XRAM[44785] = 8'b0;
    XRAM[44786] = 8'b0;
    XRAM[44787] = 8'b0;
    XRAM[44788] = 8'b0;
    XRAM[44789] = 8'b0;
    XRAM[44790] = 8'b0;
    XRAM[44791] = 8'b0;
    XRAM[44792] = 8'b0;
    XRAM[44793] = 8'b0;
    XRAM[44794] = 8'b0;
    XRAM[44795] = 8'b0;
    XRAM[44796] = 8'b0;
    XRAM[44797] = 8'b0;
    XRAM[44798] = 8'b0;
    XRAM[44799] = 8'b0;
    XRAM[44800] = 8'b0;
    XRAM[44801] = 8'b0;
    XRAM[44802] = 8'b0;
    XRAM[44803] = 8'b0;
    XRAM[44804] = 8'b0;
    XRAM[44805] = 8'b0;
    XRAM[44806] = 8'b0;
    XRAM[44807] = 8'b0;
    XRAM[44808] = 8'b0;
    XRAM[44809] = 8'b0;
    XRAM[44810] = 8'b0;
    XRAM[44811] = 8'b0;
    XRAM[44812] = 8'b0;
    XRAM[44813] = 8'b0;
    XRAM[44814] = 8'b0;
    XRAM[44815] = 8'b0;
    XRAM[44816] = 8'b0;
    XRAM[44817] = 8'b0;
    XRAM[44818] = 8'b0;
    XRAM[44819] = 8'b0;
    XRAM[44820] = 8'b0;
    XRAM[44821] = 8'b0;
    XRAM[44822] = 8'b0;
    XRAM[44823] = 8'b0;
    XRAM[44824] = 8'b0;
    XRAM[44825] = 8'b0;
    XRAM[44826] = 8'b0;
    XRAM[44827] = 8'b0;
    XRAM[44828] = 8'b0;
    XRAM[44829] = 8'b0;
    XRAM[44830] = 8'b0;
    XRAM[44831] = 8'b0;
    XRAM[44832] = 8'b0;
    XRAM[44833] = 8'b0;
    XRAM[44834] = 8'b0;
    XRAM[44835] = 8'b0;
    XRAM[44836] = 8'b0;
    XRAM[44837] = 8'b0;
    XRAM[44838] = 8'b0;
    XRAM[44839] = 8'b0;
    XRAM[44840] = 8'b0;
    XRAM[44841] = 8'b0;
    XRAM[44842] = 8'b0;
    XRAM[44843] = 8'b0;
    XRAM[44844] = 8'b0;
    XRAM[44845] = 8'b0;
    XRAM[44846] = 8'b0;
    XRAM[44847] = 8'b0;
    XRAM[44848] = 8'b0;
    XRAM[44849] = 8'b0;
    XRAM[44850] = 8'b0;
    XRAM[44851] = 8'b0;
    XRAM[44852] = 8'b0;
    XRAM[44853] = 8'b0;
    XRAM[44854] = 8'b0;
    XRAM[44855] = 8'b0;
    XRAM[44856] = 8'b0;
    XRAM[44857] = 8'b0;
    XRAM[44858] = 8'b0;
    XRAM[44859] = 8'b0;
    XRAM[44860] = 8'b0;
    XRAM[44861] = 8'b0;
    XRAM[44862] = 8'b0;
    XRAM[44863] = 8'b0;
    XRAM[44864] = 8'b0;
    XRAM[44865] = 8'b0;
    XRAM[44866] = 8'b0;
    XRAM[44867] = 8'b0;
    XRAM[44868] = 8'b0;
    XRAM[44869] = 8'b0;
    XRAM[44870] = 8'b0;
    XRAM[44871] = 8'b0;
    XRAM[44872] = 8'b0;
    XRAM[44873] = 8'b0;
    XRAM[44874] = 8'b0;
    XRAM[44875] = 8'b0;
    XRAM[44876] = 8'b0;
    XRAM[44877] = 8'b0;
    XRAM[44878] = 8'b0;
    XRAM[44879] = 8'b0;
    XRAM[44880] = 8'b0;
    XRAM[44881] = 8'b0;
    XRAM[44882] = 8'b0;
    XRAM[44883] = 8'b0;
    XRAM[44884] = 8'b0;
    XRAM[44885] = 8'b0;
    XRAM[44886] = 8'b0;
    XRAM[44887] = 8'b0;
    XRAM[44888] = 8'b0;
    XRAM[44889] = 8'b0;
    XRAM[44890] = 8'b0;
    XRAM[44891] = 8'b0;
    XRAM[44892] = 8'b0;
    XRAM[44893] = 8'b0;
    XRAM[44894] = 8'b0;
    XRAM[44895] = 8'b0;
    XRAM[44896] = 8'b0;
    XRAM[44897] = 8'b0;
    XRAM[44898] = 8'b0;
    XRAM[44899] = 8'b0;
    XRAM[44900] = 8'b0;
    XRAM[44901] = 8'b0;
    XRAM[44902] = 8'b0;
    XRAM[44903] = 8'b0;
    XRAM[44904] = 8'b0;
    XRAM[44905] = 8'b0;
    XRAM[44906] = 8'b0;
    XRAM[44907] = 8'b0;
    XRAM[44908] = 8'b0;
    XRAM[44909] = 8'b0;
    XRAM[44910] = 8'b0;
    XRAM[44911] = 8'b0;
    XRAM[44912] = 8'b0;
    XRAM[44913] = 8'b0;
    XRAM[44914] = 8'b0;
    XRAM[44915] = 8'b0;
    XRAM[44916] = 8'b0;
    XRAM[44917] = 8'b0;
    XRAM[44918] = 8'b0;
    XRAM[44919] = 8'b0;
    XRAM[44920] = 8'b0;
    XRAM[44921] = 8'b0;
    XRAM[44922] = 8'b0;
    XRAM[44923] = 8'b0;
    XRAM[44924] = 8'b0;
    XRAM[44925] = 8'b0;
    XRAM[44926] = 8'b0;
    XRAM[44927] = 8'b0;
    XRAM[44928] = 8'b0;
    XRAM[44929] = 8'b0;
    XRAM[44930] = 8'b0;
    XRAM[44931] = 8'b0;
    XRAM[44932] = 8'b0;
    XRAM[44933] = 8'b0;
    XRAM[44934] = 8'b0;
    XRAM[44935] = 8'b0;
    XRAM[44936] = 8'b0;
    XRAM[44937] = 8'b0;
    XRAM[44938] = 8'b0;
    XRAM[44939] = 8'b0;
    XRAM[44940] = 8'b0;
    XRAM[44941] = 8'b0;
    XRAM[44942] = 8'b0;
    XRAM[44943] = 8'b0;
    XRAM[44944] = 8'b0;
    XRAM[44945] = 8'b0;
    XRAM[44946] = 8'b0;
    XRAM[44947] = 8'b0;
    XRAM[44948] = 8'b0;
    XRAM[44949] = 8'b0;
    XRAM[44950] = 8'b0;
    XRAM[44951] = 8'b0;
    XRAM[44952] = 8'b0;
    XRAM[44953] = 8'b0;
    XRAM[44954] = 8'b0;
    XRAM[44955] = 8'b0;
    XRAM[44956] = 8'b0;
    XRAM[44957] = 8'b0;
    XRAM[44958] = 8'b0;
    XRAM[44959] = 8'b0;
    XRAM[44960] = 8'b0;
    XRAM[44961] = 8'b0;
    XRAM[44962] = 8'b0;
    XRAM[44963] = 8'b0;
    XRAM[44964] = 8'b0;
    XRAM[44965] = 8'b0;
    XRAM[44966] = 8'b0;
    XRAM[44967] = 8'b0;
    XRAM[44968] = 8'b0;
    XRAM[44969] = 8'b0;
    XRAM[44970] = 8'b0;
    XRAM[44971] = 8'b0;
    XRAM[44972] = 8'b0;
    XRAM[44973] = 8'b0;
    XRAM[44974] = 8'b0;
    XRAM[44975] = 8'b0;
    XRAM[44976] = 8'b0;
    XRAM[44977] = 8'b0;
    XRAM[44978] = 8'b0;
    XRAM[44979] = 8'b0;
    XRAM[44980] = 8'b0;
    XRAM[44981] = 8'b0;
    XRAM[44982] = 8'b0;
    XRAM[44983] = 8'b0;
    XRAM[44984] = 8'b0;
    XRAM[44985] = 8'b0;
    XRAM[44986] = 8'b0;
    XRAM[44987] = 8'b0;
    XRAM[44988] = 8'b0;
    XRAM[44989] = 8'b0;
    XRAM[44990] = 8'b0;
    XRAM[44991] = 8'b0;
    XRAM[44992] = 8'b0;
    XRAM[44993] = 8'b0;
    XRAM[44994] = 8'b0;
    XRAM[44995] = 8'b0;
    XRAM[44996] = 8'b0;
    XRAM[44997] = 8'b0;
    XRAM[44998] = 8'b0;
    XRAM[44999] = 8'b0;
    XRAM[45000] = 8'b0;
    XRAM[45001] = 8'b0;
    XRAM[45002] = 8'b0;
    XRAM[45003] = 8'b0;
    XRAM[45004] = 8'b0;
    XRAM[45005] = 8'b0;
    XRAM[45006] = 8'b0;
    XRAM[45007] = 8'b0;
    XRAM[45008] = 8'b0;
    XRAM[45009] = 8'b0;
    XRAM[45010] = 8'b0;
    XRAM[45011] = 8'b0;
    XRAM[45012] = 8'b0;
    XRAM[45013] = 8'b0;
    XRAM[45014] = 8'b0;
    XRAM[45015] = 8'b0;
    XRAM[45016] = 8'b0;
    XRAM[45017] = 8'b0;
    XRAM[45018] = 8'b0;
    XRAM[45019] = 8'b0;
    XRAM[45020] = 8'b0;
    XRAM[45021] = 8'b0;
    XRAM[45022] = 8'b0;
    XRAM[45023] = 8'b0;
    XRAM[45024] = 8'b0;
    XRAM[45025] = 8'b0;
    XRAM[45026] = 8'b0;
    XRAM[45027] = 8'b0;
    XRAM[45028] = 8'b0;
    XRAM[45029] = 8'b0;
    XRAM[45030] = 8'b0;
    XRAM[45031] = 8'b0;
    XRAM[45032] = 8'b0;
    XRAM[45033] = 8'b0;
    XRAM[45034] = 8'b0;
    XRAM[45035] = 8'b0;
    XRAM[45036] = 8'b0;
    XRAM[45037] = 8'b0;
    XRAM[45038] = 8'b0;
    XRAM[45039] = 8'b0;
    XRAM[45040] = 8'b0;
    XRAM[45041] = 8'b0;
    XRAM[45042] = 8'b0;
    XRAM[45043] = 8'b0;
    XRAM[45044] = 8'b0;
    XRAM[45045] = 8'b0;
    XRAM[45046] = 8'b0;
    XRAM[45047] = 8'b0;
    XRAM[45048] = 8'b0;
    XRAM[45049] = 8'b0;
    XRAM[45050] = 8'b0;
    XRAM[45051] = 8'b0;
    XRAM[45052] = 8'b0;
    XRAM[45053] = 8'b0;
    XRAM[45054] = 8'b0;
    XRAM[45055] = 8'b0;
    XRAM[45056] = 8'b0;
    XRAM[45057] = 8'b0;
    XRAM[45058] = 8'b0;
    XRAM[45059] = 8'b0;
    XRAM[45060] = 8'b0;
    XRAM[45061] = 8'b0;
    XRAM[45062] = 8'b0;
    XRAM[45063] = 8'b0;
    XRAM[45064] = 8'b0;
    XRAM[45065] = 8'b0;
    XRAM[45066] = 8'b0;
    XRAM[45067] = 8'b0;
    XRAM[45068] = 8'b0;
    XRAM[45069] = 8'b0;
    XRAM[45070] = 8'b0;
    XRAM[45071] = 8'b0;
    XRAM[45072] = 8'b0;
    XRAM[45073] = 8'b0;
    XRAM[45074] = 8'b0;
    XRAM[45075] = 8'b0;
    XRAM[45076] = 8'b0;
    XRAM[45077] = 8'b0;
    XRAM[45078] = 8'b0;
    XRAM[45079] = 8'b0;
    XRAM[45080] = 8'b0;
    XRAM[45081] = 8'b0;
    XRAM[45082] = 8'b0;
    XRAM[45083] = 8'b0;
    XRAM[45084] = 8'b0;
    XRAM[45085] = 8'b0;
    XRAM[45086] = 8'b0;
    XRAM[45087] = 8'b0;
    XRAM[45088] = 8'b0;
    XRAM[45089] = 8'b0;
    XRAM[45090] = 8'b0;
    XRAM[45091] = 8'b0;
    XRAM[45092] = 8'b0;
    XRAM[45093] = 8'b0;
    XRAM[45094] = 8'b0;
    XRAM[45095] = 8'b0;
    XRAM[45096] = 8'b0;
    XRAM[45097] = 8'b0;
    XRAM[45098] = 8'b0;
    XRAM[45099] = 8'b0;
    XRAM[45100] = 8'b0;
    XRAM[45101] = 8'b0;
    XRAM[45102] = 8'b0;
    XRAM[45103] = 8'b0;
    XRAM[45104] = 8'b0;
    XRAM[45105] = 8'b0;
    XRAM[45106] = 8'b0;
    XRAM[45107] = 8'b0;
    XRAM[45108] = 8'b0;
    XRAM[45109] = 8'b0;
    XRAM[45110] = 8'b0;
    XRAM[45111] = 8'b0;
    XRAM[45112] = 8'b0;
    XRAM[45113] = 8'b0;
    XRAM[45114] = 8'b0;
    XRAM[45115] = 8'b0;
    XRAM[45116] = 8'b0;
    XRAM[45117] = 8'b0;
    XRAM[45118] = 8'b0;
    XRAM[45119] = 8'b0;
    XRAM[45120] = 8'b0;
    XRAM[45121] = 8'b0;
    XRAM[45122] = 8'b0;
    XRAM[45123] = 8'b0;
    XRAM[45124] = 8'b0;
    XRAM[45125] = 8'b0;
    XRAM[45126] = 8'b0;
    XRAM[45127] = 8'b0;
    XRAM[45128] = 8'b0;
    XRAM[45129] = 8'b0;
    XRAM[45130] = 8'b0;
    XRAM[45131] = 8'b0;
    XRAM[45132] = 8'b0;
    XRAM[45133] = 8'b0;
    XRAM[45134] = 8'b0;
    XRAM[45135] = 8'b0;
    XRAM[45136] = 8'b0;
    XRAM[45137] = 8'b0;
    XRAM[45138] = 8'b0;
    XRAM[45139] = 8'b0;
    XRAM[45140] = 8'b0;
    XRAM[45141] = 8'b0;
    XRAM[45142] = 8'b0;
    XRAM[45143] = 8'b0;
    XRAM[45144] = 8'b0;
    XRAM[45145] = 8'b0;
    XRAM[45146] = 8'b0;
    XRAM[45147] = 8'b0;
    XRAM[45148] = 8'b0;
    XRAM[45149] = 8'b0;
    XRAM[45150] = 8'b0;
    XRAM[45151] = 8'b0;
    XRAM[45152] = 8'b0;
    XRAM[45153] = 8'b0;
    XRAM[45154] = 8'b0;
    XRAM[45155] = 8'b0;
    XRAM[45156] = 8'b0;
    XRAM[45157] = 8'b0;
    XRAM[45158] = 8'b0;
    XRAM[45159] = 8'b0;
    XRAM[45160] = 8'b0;
    XRAM[45161] = 8'b0;
    XRAM[45162] = 8'b0;
    XRAM[45163] = 8'b0;
    XRAM[45164] = 8'b0;
    XRAM[45165] = 8'b0;
    XRAM[45166] = 8'b0;
    XRAM[45167] = 8'b0;
    XRAM[45168] = 8'b0;
    XRAM[45169] = 8'b0;
    XRAM[45170] = 8'b0;
    XRAM[45171] = 8'b0;
    XRAM[45172] = 8'b0;
    XRAM[45173] = 8'b0;
    XRAM[45174] = 8'b0;
    XRAM[45175] = 8'b0;
    XRAM[45176] = 8'b0;
    XRAM[45177] = 8'b0;
    XRAM[45178] = 8'b0;
    XRAM[45179] = 8'b0;
    XRAM[45180] = 8'b0;
    XRAM[45181] = 8'b0;
    XRAM[45182] = 8'b0;
    XRAM[45183] = 8'b0;
    XRAM[45184] = 8'b0;
    XRAM[45185] = 8'b0;
    XRAM[45186] = 8'b0;
    XRAM[45187] = 8'b0;
    XRAM[45188] = 8'b0;
    XRAM[45189] = 8'b0;
    XRAM[45190] = 8'b0;
    XRAM[45191] = 8'b0;
    XRAM[45192] = 8'b0;
    XRAM[45193] = 8'b0;
    XRAM[45194] = 8'b0;
    XRAM[45195] = 8'b0;
    XRAM[45196] = 8'b0;
    XRAM[45197] = 8'b0;
    XRAM[45198] = 8'b0;
    XRAM[45199] = 8'b0;
    XRAM[45200] = 8'b0;
    XRAM[45201] = 8'b0;
    XRAM[45202] = 8'b0;
    XRAM[45203] = 8'b0;
    XRAM[45204] = 8'b0;
    XRAM[45205] = 8'b0;
    XRAM[45206] = 8'b0;
    XRAM[45207] = 8'b0;
    XRAM[45208] = 8'b0;
    XRAM[45209] = 8'b0;
    XRAM[45210] = 8'b0;
    XRAM[45211] = 8'b0;
    XRAM[45212] = 8'b0;
    XRAM[45213] = 8'b0;
    XRAM[45214] = 8'b0;
    XRAM[45215] = 8'b0;
    XRAM[45216] = 8'b0;
    XRAM[45217] = 8'b0;
    XRAM[45218] = 8'b0;
    XRAM[45219] = 8'b0;
    XRAM[45220] = 8'b0;
    XRAM[45221] = 8'b0;
    XRAM[45222] = 8'b0;
    XRAM[45223] = 8'b0;
    XRAM[45224] = 8'b0;
    XRAM[45225] = 8'b0;
    XRAM[45226] = 8'b0;
    XRAM[45227] = 8'b0;
    XRAM[45228] = 8'b0;
    XRAM[45229] = 8'b0;
    XRAM[45230] = 8'b0;
    XRAM[45231] = 8'b0;
    XRAM[45232] = 8'b0;
    XRAM[45233] = 8'b0;
    XRAM[45234] = 8'b0;
    XRAM[45235] = 8'b0;
    XRAM[45236] = 8'b0;
    XRAM[45237] = 8'b0;
    XRAM[45238] = 8'b0;
    XRAM[45239] = 8'b0;
    XRAM[45240] = 8'b0;
    XRAM[45241] = 8'b0;
    XRAM[45242] = 8'b0;
    XRAM[45243] = 8'b0;
    XRAM[45244] = 8'b0;
    XRAM[45245] = 8'b0;
    XRAM[45246] = 8'b0;
    XRAM[45247] = 8'b0;
    XRAM[45248] = 8'b0;
    XRAM[45249] = 8'b0;
    XRAM[45250] = 8'b0;
    XRAM[45251] = 8'b0;
    XRAM[45252] = 8'b0;
    XRAM[45253] = 8'b0;
    XRAM[45254] = 8'b0;
    XRAM[45255] = 8'b0;
    XRAM[45256] = 8'b0;
    XRAM[45257] = 8'b0;
    XRAM[45258] = 8'b0;
    XRAM[45259] = 8'b0;
    XRAM[45260] = 8'b0;
    XRAM[45261] = 8'b0;
    XRAM[45262] = 8'b0;
    XRAM[45263] = 8'b0;
    XRAM[45264] = 8'b0;
    XRAM[45265] = 8'b0;
    XRAM[45266] = 8'b0;
    XRAM[45267] = 8'b0;
    XRAM[45268] = 8'b0;
    XRAM[45269] = 8'b0;
    XRAM[45270] = 8'b0;
    XRAM[45271] = 8'b0;
    XRAM[45272] = 8'b0;
    XRAM[45273] = 8'b0;
    XRAM[45274] = 8'b0;
    XRAM[45275] = 8'b0;
    XRAM[45276] = 8'b0;
    XRAM[45277] = 8'b0;
    XRAM[45278] = 8'b0;
    XRAM[45279] = 8'b0;
    XRAM[45280] = 8'b0;
    XRAM[45281] = 8'b0;
    XRAM[45282] = 8'b0;
    XRAM[45283] = 8'b0;
    XRAM[45284] = 8'b0;
    XRAM[45285] = 8'b0;
    XRAM[45286] = 8'b0;
    XRAM[45287] = 8'b0;
    XRAM[45288] = 8'b0;
    XRAM[45289] = 8'b0;
    XRAM[45290] = 8'b0;
    XRAM[45291] = 8'b0;
    XRAM[45292] = 8'b0;
    XRAM[45293] = 8'b0;
    XRAM[45294] = 8'b0;
    XRAM[45295] = 8'b0;
    XRAM[45296] = 8'b0;
    XRAM[45297] = 8'b0;
    XRAM[45298] = 8'b0;
    XRAM[45299] = 8'b0;
    XRAM[45300] = 8'b0;
    XRAM[45301] = 8'b0;
    XRAM[45302] = 8'b0;
    XRAM[45303] = 8'b0;
    XRAM[45304] = 8'b0;
    XRAM[45305] = 8'b0;
    XRAM[45306] = 8'b0;
    XRAM[45307] = 8'b0;
    XRAM[45308] = 8'b0;
    XRAM[45309] = 8'b0;
    XRAM[45310] = 8'b0;
    XRAM[45311] = 8'b0;
    XRAM[45312] = 8'b0;
    XRAM[45313] = 8'b0;
    XRAM[45314] = 8'b0;
    XRAM[45315] = 8'b0;
    XRAM[45316] = 8'b0;
    XRAM[45317] = 8'b0;
    XRAM[45318] = 8'b0;
    XRAM[45319] = 8'b0;
    XRAM[45320] = 8'b0;
    XRAM[45321] = 8'b0;
    XRAM[45322] = 8'b0;
    XRAM[45323] = 8'b0;
    XRAM[45324] = 8'b0;
    XRAM[45325] = 8'b0;
    XRAM[45326] = 8'b0;
    XRAM[45327] = 8'b0;
    XRAM[45328] = 8'b0;
    XRAM[45329] = 8'b0;
    XRAM[45330] = 8'b0;
    XRAM[45331] = 8'b0;
    XRAM[45332] = 8'b0;
    XRAM[45333] = 8'b0;
    XRAM[45334] = 8'b0;
    XRAM[45335] = 8'b0;
    XRAM[45336] = 8'b0;
    XRAM[45337] = 8'b0;
    XRAM[45338] = 8'b0;
    XRAM[45339] = 8'b0;
    XRAM[45340] = 8'b0;
    XRAM[45341] = 8'b0;
    XRAM[45342] = 8'b0;
    XRAM[45343] = 8'b0;
    XRAM[45344] = 8'b0;
    XRAM[45345] = 8'b0;
    XRAM[45346] = 8'b0;
    XRAM[45347] = 8'b0;
    XRAM[45348] = 8'b0;
    XRAM[45349] = 8'b0;
    XRAM[45350] = 8'b0;
    XRAM[45351] = 8'b0;
    XRAM[45352] = 8'b0;
    XRAM[45353] = 8'b0;
    XRAM[45354] = 8'b0;
    XRAM[45355] = 8'b0;
    XRAM[45356] = 8'b0;
    XRAM[45357] = 8'b0;
    XRAM[45358] = 8'b0;
    XRAM[45359] = 8'b0;
    XRAM[45360] = 8'b0;
    XRAM[45361] = 8'b0;
    XRAM[45362] = 8'b0;
    XRAM[45363] = 8'b0;
    XRAM[45364] = 8'b0;
    XRAM[45365] = 8'b0;
    XRAM[45366] = 8'b0;
    XRAM[45367] = 8'b0;
    XRAM[45368] = 8'b0;
    XRAM[45369] = 8'b0;
    XRAM[45370] = 8'b0;
    XRAM[45371] = 8'b0;
    XRAM[45372] = 8'b0;
    XRAM[45373] = 8'b0;
    XRAM[45374] = 8'b0;
    XRAM[45375] = 8'b0;
    XRAM[45376] = 8'b0;
    XRAM[45377] = 8'b0;
    XRAM[45378] = 8'b0;
    XRAM[45379] = 8'b0;
    XRAM[45380] = 8'b0;
    XRAM[45381] = 8'b0;
    XRAM[45382] = 8'b0;
    XRAM[45383] = 8'b0;
    XRAM[45384] = 8'b0;
    XRAM[45385] = 8'b0;
    XRAM[45386] = 8'b0;
    XRAM[45387] = 8'b0;
    XRAM[45388] = 8'b0;
    XRAM[45389] = 8'b0;
    XRAM[45390] = 8'b0;
    XRAM[45391] = 8'b0;
    XRAM[45392] = 8'b0;
    XRAM[45393] = 8'b0;
    XRAM[45394] = 8'b0;
    XRAM[45395] = 8'b0;
    XRAM[45396] = 8'b0;
    XRAM[45397] = 8'b0;
    XRAM[45398] = 8'b0;
    XRAM[45399] = 8'b0;
    XRAM[45400] = 8'b0;
    XRAM[45401] = 8'b0;
    XRAM[45402] = 8'b0;
    XRAM[45403] = 8'b0;
    XRAM[45404] = 8'b0;
    XRAM[45405] = 8'b0;
    XRAM[45406] = 8'b0;
    XRAM[45407] = 8'b0;
    XRAM[45408] = 8'b0;
    XRAM[45409] = 8'b0;
    XRAM[45410] = 8'b0;
    XRAM[45411] = 8'b0;
    XRAM[45412] = 8'b0;
    XRAM[45413] = 8'b0;
    XRAM[45414] = 8'b0;
    XRAM[45415] = 8'b0;
    XRAM[45416] = 8'b0;
    XRAM[45417] = 8'b0;
    XRAM[45418] = 8'b0;
    XRAM[45419] = 8'b0;
    XRAM[45420] = 8'b0;
    XRAM[45421] = 8'b0;
    XRAM[45422] = 8'b0;
    XRAM[45423] = 8'b0;
    XRAM[45424] = 8'b0;
    XRAM[45425] = 8'b0;
    XRAM[45426] = 8'b0;
    XRAM[45427] = 8'b0;
    XRAM[45428] = 8'b0;
    XRAM[45429] = 8'b0;
    XRAM[45430] = 8'b0;
    XRAM[45431] = 8'b0;
    XRAM[45432] = 8'b0;
    XRAM[45433] = 8'b0;
    XRAM[45434] = 8'b0;
    XRAM[45435] = 8'b0;
    XRAM[45436] = 8'b0;
    XRAM[45437] = 8'b0;
    XRAM[45438] = 8'b0;
    XRAM[45439] = 8'b0;
    XRAM[45440] = 8'b0;
    XRAM[45441] = 8'b0;
    XRAM[45442] = 8'b0;
    XRAM[45443] = 8'b0;
    XRAM[45444] = 8'b0;
    XRAM[45445] = 8'b0;
    XRAM[45446] = 8'b0;
    XRAM[45447] = 8'b0;
    XRAM[45448] = 8'b0;
    XRAM[45449] = 8'b0;
    XRAM[45450] = 8'b0;
    XRAM[45451] = 8'b0;
    XRAM[45452] = 8'b0;
    XRAM[45453] = 8'b0;
    XRAM[45454] = 8'b0;
    XRAM[45455] = 8'b0;
    XRAM[45456] = 8'b0;
    XRAM[45457] = 8'b0;
    XRAM[45458] = 8'b0;
    XRAM[45459] = 8'b0;
    XRAM[45460] = 8'b0;
    XRAM[45461] = 8'b0;
    XRAM[45462] = 8'b0;
    XRAM[45463] = 8'b0;
    XRAM[45464] = 8'b0;
    XRAM[45465] = 8'b0;
    XRAM[45466] = 8'b0;
    XRAM[45467] = 8'b0;
    XRAM[45468] = 8'b0;
    XRAM[45469] = 8'b0;
    XRAM[45470] = 8'b0;
    XRAM[45471] = 8'b0;
    XRAM[45472] = 8'b0;
    XRAM[45473] = 8'b0;
    XRAM[45474] = 8'b0;
    XRAM[45475] = 8'b0;
    XRAM[45476] = 8'b0;
    XRAM[45477] = 8'b0;
    XRAM[45478] = 8'b0;
    XRAM[45479] = 8'b0;
    XRAM[45480] = 8'b0;
    XRAM[45481] = 8'b0;
    XRAM[45482] = 8'b0;
    XRAM[45483] = 8'b0;
    XRAM[45484] = 8'b0;
    XRAM[45485] = 8'b0;
    XRAM[45486] = 8'b0;
    XRAM[45487] = 8'b0;
    XRAM[45488] = 8'b0;
    XRAM[45489] = 8'b0;
    XRAM[45490] = 8'b0;
    XRAM[45491] = 8'b0;
    XRAM[45492] = 8'b0;
    XRAM[45493] = 8'b0;
    XRAM[45494] = 8'b0;
    XRAM[45495] = 8'b0;
    XRAM[45496] = 8'b0;
    XRAM[45497] = 8'b0;
    XRAM[45498] = 8'b0;
    XRAM[45499] = 8'b0;
    XRAM[45500] = 8'b0;
    XRAM[45501] = 8'b0;
    XRAM[45502] = 8'b0;
    XRAM[45503] = 8'b0;
    XRAM[45504] = 8'b0;
    XRAM[45505] = 8'b0;
    XRAM[45506] = 8'b0;
    XRAM[45507] = 8'b0;
    XRAM[45508] = 8'b0;
    XRAM[45509] = 8'b0;
    XRAM[45510] = 8'b0;
    XRAM[45511] = 8'b0;
    XRAM[45512] = 8'b0;
    XRAM[45513] = 8'b0;
    XRAM[45514] = 8'b0;
    XRAM[45515] = 8'b0;
    XRAM[45516] = 8'b0;
    XRAM[45517] = 8'b0;
    XRAM[45518] = 8'b0;
    XRAM[45519] = 8'b0;
    XRAM[45520] = 8'b0;
    XRAM[45521] = 8'b0;
    XRAM[45522] = 8'b0;
    XRAM[45523] = 8'b0;
    XRAM[45524] = 8'b0;
    XRAM[45525] = 8'b0;
    XRAM[45526] = 8'b0;
    XRAM[45527] = 8'b0;
    XRAM[45528] = 8'b0;
    XRAM[45529] = 8'b0;
    XRAM[45530] = 8'b0;
    XRAM[45531] = 8'b0;
    XRAM[45532] = 8'b0;
    XRAM[45533] = 8'b0;
    XRAM[45534] = 8'b0;
    XRAM[45535] = 8'b0;
    XRAM[45536] = 8'b0;
    XRAM[45537] = 8'b0;
    XRAM[45538] = 8'b0;
    XRAM[45539] = 8'b0;
    XRAM[45540] = 8'b0;
    XRAM[45541] = 8'b0;
    XRAM[45542] = 8'b0;
    XRAM[45543] = 8'b0;
    XRAM[45544] = 8'b0;
    XRAM[45545] = 8'b0;
    XRAM[45546] = 8'b0;
    XRAM[45547] = 8'b0;
    XRAM[45548] = 8'b0;
    XRAM[45549] = 8'b0;
    XRAM[45550] = 8'b0;
    XRAM[45551] = 8'b0;
    XRAM[45552] = 8'b0;
    XRAM[45553] = 8'b0;
    XRAM[45554] = 8'b0;
    XRAM[45555] = 8'b0;
    XRAM[45556] = 8'b0;
    XRAM[45557] = 8'b0;
    XRAM[45558] = 8'b0;
    XRAM[45559] = 8'b0;
    XRAM[45560] = 8'b0;
    XRAM[45561] = 8'b0;
    XRAM[45562] = 8'b0;
    XRAM[45563] = 8'b0;
    XRAM[45564] = 8'b0;
    XRAM[45565] = 8'b0;
    XRAM[45566] = 8'b0;
    XRAM[45567] = 8'b0;
    XRAM[45568] = 8'b0;
    XRAM[45569] = 8'b0;
    XRAM[45570] = 8'b0;
    XRAM[45571] = 8'b0;
    XRAM[45572] = 8'b0;
    XRAM[45573] = 8'b0;
    XRAM[45574] = 8'b0;
    XRAM[45575] = 8'b0;
    XRAM[45576] = 8'b0;
    XRAM[45577] = 8'b0;
    XRAM[45578] = 8'b0;
    XRAM[45579] = 8'b0;
    XRAM[45580] = 8'b0;
    XRAM[45581] = 8'b0;
    XRAM[45582] = 8'b0;
    XRAM[45583] = 8'b0;
    XRAM[45584] = 8'b0;
    XRAM[45585] = 8'b0;
    XRAM[45586] = 8'b0;
    XRAM[45587] = 8'b0;
    XRAM[45588] = 8'b0;
    XRAM[45589] = 8'b0;
    XRAM[45590] = 8'b0;
    XRAM[45591] = 8'b0;
    XRAM[45592] = 8'b0;
    XRAM[45593] = 8'b0;
    XRAM[45594] = 8'b0;
    XRAM[45595] = 8'b0;
    XRAM[45596] = 8'b0;
    XRAM[45597] = 8'b0;
    XRAM[45598] = 8'b0;
    XRAM[45599] = 8'b0;
    XRAM[45600] = 8'b0;
    XRAM[45601] = 8'b0;
    XRAM[45602] = 8'b0;
    XRAM[45603] = 8'b0;
    XRAM[45604] = 8'b0;
    XRAM[45605] = 8'b0;
    XRAM[45606] = 8'b0;
    XRAM[45607] = 8'b0;
    XRAM[45608] = 8'b0;
    XRAM[45609] = 8'b0;
    XRAM[45610] = 8'b0;
    XRAM[45611] = 8'b0;
    XRAM[45612] = 8'b0;
    XRAM[45613] = 8'b0;
    XRAM[45614] = 8'b0;
    XRAM[45615] = 8'b0;
    XRAM[45616] = 8'b0;
    XRAM[45617] = 8'b0;
    XRAM[45618] = 8'b0;
    XRAM[45619] = 8'b0;
    XRAM[45620] = 8'b0;
    XRAM[45621] = 8'b0;
    XRAM[45622] = 8'b0;
    XRAM[45623] = 8'b0;
    XRAM[45624] = 8'b0;
    XRAM[45625] = 8'b0;
    XRAM[45626] = 8'b0;
    XRAM[45627] = 8'b0;
    XRAM[45628] = 8'b0;
    XRAM[45629] = 8'b0;
    XRAM[45630] = 8'b0;
    XRAM[45631] = 8'b0;
    XRAM[45632] = 8'b0;
    XRAM[45633] = 8'b0;
    XRAM[45634] = 8'b0;
    XRAM[45635] = 8'b0;
    XRAM[45636] = 8'b0;
    XRAM[45637] = 8'b0;
    XRAM[45638] = 8'b0;
    XRAM[45639] = 8'b0;
    XRAM[45640] = 8'b0;
    XRAM[45641] = 8'b0;
    XRAM[45642] = 8'b0;
    XRAM[45643] = 8'b0;
    XRAM[45644] = 8'b0;
    XRAM[45645] = 8'b0;
    XRAM[45646] = 8'b0;
    XRAM[45647] = 8'b0;
    XRAM[45648] = 8'b0;
    XRAM[45649] = 8'b0;
    XRAM[45650] = 8'b0;
    XRAM[45651] = 8'b0;
    XRAM[45652] = 8'b0;
    XRAM[45653] = 8'b0;
    XRAM[45654] = 8'b0;
    XRAM[45655] = 8'b0;
    XRAM[45656] = 8'b0;
    XRAM[45657] = 8'b0;
    XRAM[45658] = 8'b0;
    XRAM[45659] = 8'b0;
    XRAM[45660] = 8'b0;
    XRAM[45661] = 8'b0;
    XRAM[45662] = 8'b0;
    XRAM[45663] = 8'b0;
    XRAM[45664] = 8'b0;
    XRAM[45665] = 8'b0;
    XRAM[45666] = 8'b0;
    XRAM[45667] = 8'b0;
    XRAM[45668] = 8'b0;
    XRAM[45669] = 8'b0;
    XRAM[45670] = 8'b0;
    XRAM[45671] = 8'b0;
    XRAM[45672] = 8'b0;
    XRAM[45673] = 8'b0;
    XRAM[45674] = 8'b0;
    XRAM[45675] = 8'b0;
    XRAM[45676] = 8'b0;
    XRAM[45677] = 8'b0;
    XRAM[45678] = 8'b0;
    XRAM[45679] = 8'b0;
    XRAM[45680] = 8'b0;
    XRAM[45681] = 8'b0;
    XRAM[45682] = 8'b0;
    XRAM[45683] = 8'b0;
    XRAM[45684] = 8'b0;
    XRAM[45685] = 8'b0;
    XRAM[45686] = 8'b0;
    XRAM[45687] = 8'b0;
    XRAM[45688] = 8'b0;
    XRAM[45689] = 8'b0;
    XRAM[45690] = 8'b0;
    XRAM[45691] = 8'b0;
    XRAM[45692] = 8'b0;
    XRAM[45693] = 8'b0;
    XRAM[45694] = 8'b0;
    XRAM[45695] = 8'b0;
    XRAM[45696] = 8'b0;
    XRAM[45697] = 8'b0;
    XRAM[45698] = 8'b0;
    XRAM[45699] = 8'b0;
    XRAM[45700] = 8'b0;
    XRAM[45701] = 8'b0;
    XRAM[45702] = 8'b0;
    XRAM[45703] = 8'b0;
    XRAM[45704] = 8'b0;
    XRAM[45705] = 8'b0;
    XRAM[45706] = 8'b0;
    XRAM[45707] = 8'b0;
    XRAM[45708] = 8'b0;
    XRAM[45709] = 8'b0;
    XRAM[45710] = 8'b0;
    XRAM[45711] = 8'b0;
    XRAM[45712] = 8'b0;
    XRAM[45713] = 8'b0;
    XRAM[45714] = 8'b0;
    XRAM[45715] = 8'b0;
    XRAM[45716] = 8'b0;
    XRAM[45717] = 8'b0;
    XRAM[45718] = 8'b0;
    XRAM[45719] = 8'b0;
    XRAM[45720] = 8'b0;
    XRAM[45721] = 8'b0;
    XRAM[45722] = 8'b0;
    XRAM[45723] = 8'b0;
    XRAM[45724] = 8'b0;
    XRAM[45725] = 8'b0;
    XRAM[45726] = 8'b0;
    XRAM[45727] = 8'b0;
    XRAM[45728] = 8'b0;
    XRAM[45729] = 8'b0;
    XRAM[45730] = 8'b0;
    XRAM[45731] = 8'b0;
    XRAM[45732] = 8'b0;
    XRAM[45733] = 8'b0;
    XRAM[45734] = 8'b0;
    XRAM[45735] = 8'b0;
    XRAM[45736] = 8'b0;
    XRAM[45737] = 8'b0;
    XRAM[45738] = 8'b0;
    XRAM[45739] = 8'b0;
    XRAM[45740] = 8'b0;
    XRAM[45741] = 8'b0;
    XRAM[45742] = 8'b0;
    XRAM[45743] = 8'b0;
    XRAM[45744] = 8'b0;
    XRAM[45745] = 8'b0;
    XRAM[45746] = 8'b0;
    XRAM[45747] = 8'b0;
    XRAM[45748] = 8'b0;
    XRAM[45749] = 8'b0;
    XRAM[45750] = 8'b0;
    XRAM[45751] = 8'b0;
    XRAM[45752] = 8'b0;
    XRAM[45753] = 8'b0;
    XRAM[45754] = 8'b0;
    XRAM[45755] = 8'b0;
    XRAM[45756] = 8'b0;
    XRAM[45757] = 8'b0;
    XRAM[45758] = 8'b0;
    XRAM[45759] = 8'b0;
    XRAM[45760] = 8'b0;
    XRAM[45761] = 8'b0;
    XRAM[45762] = 8'b0;
    XRAM[45763] = 8'b0;
    XRAM[45764] = 8'b0;
    XRAM[45765] = 8'b0;
    XRAM[45766] = 8'b0;
    XRAM[45767] = 8'b0;
    XRAM[45768] = 8'b0;
    XRAM[45769] = 8'b0;
    XRAM[45770] = 8'b0;
    XRAM[45771] = 8'b0;
    XRAM[45772] = 8'b0;
    XRAM[45773] = 8'b0;
    XRAM[45774] = 8'b0;
    XRAM[45775] = 8'b0;
    XRAM[45776] = 8'b0;
    XRAM[45777] = 8'b0;
    XRAM[45778] = 8'b0;
    XRAM[45779] = 8'b0;
    XRAM[45780] = 8'b0;
    XRAM[45781] = 8'b0;
    XRAM[45782] = 8'b0;
    XRAM[45783] = 8'b0;
    XRAM[45784] = 8'b0;
    XRAM[45785] = 8'b0;
    XRAM[45786] = 8'b0;
    XRAM[45787] = 8'b0;
    XRAM[45788] = 8'b0;
    XRAM[45789] = 8'b0;
    XRAM[45790] = 8'b0;
    XRAM[45791] = 8'b0;
    XRAM[45792] = 8'b0;
    XRAM[45793] = 8'b0;
    XRAM[45794] = 8'b0;
    XRAM[45795] = 8'b0;
    XRAM[45796] = 8'b0;
    XRAM[45797] = 8'b0;
    XRAM[45798] = 8'b0;
    XRAM[45799] = 8'b0;
    XRAM[45800] = 8'b0;
    XRAM[45801] = 8'b0;
    XRAM[45802] = 8'b0;
    XRAM[45803] = 8'b0;
    XRAM[45804] = 8'b0;
    XRAM[45805] = 8'b0;
    XRAM[45806] = 8'b0;
    XRAM[45807] = 8'b0;
    XRAM[45808] = 8'b0;
    XRAM[45809] = 8'b0;
    XRAM[45810] = 8'b0;
    XRAM[45811] = 8'b0;
    XRAM[45812] = 8'b0;
    XRAM[45813] = 8'b0;
    XRAM[45814] = 8'b0;
    XRAM[45815] = 8'b0;
    XRAM[45816] = 8'b0;
    XRAM[45817] = 8'b0;
    XRAM[45818] = 8'b0;
    XRAM[45819] = 8'b0;
    XRAM[45820] = 8'b0;
    XRAM[45821] = 8'b0;
    XRAM[45822] = 8'b0;
    XRAM[45823] = 8'b0;
    XRAM[45824] = 8'b0;
    XRAM[45825] = 8'b0;
    XRAM[45826] = 8'b0;
    XRAM[45827] = 8'b0;
    XRAM[45828] = 8'b0;
    XRAM[45829] = 8'b0;
    XRAM[45830] = 8'b0;
    XRAM[45831] = 8'b0;
    XRAM[45832] = 8'b0;
    XRAM[45833] = 8'b0;
    XRAM[45834] = 8'b0;
    XRAM[45835] = 8'b0;
    XRAM[45836] = 8'b0;
    XRAM[45837] = 8'b0;
    XRAM[45838] = 8'b0;
    XRAM[45839] = 8'b0;
    XRAM[45840] = 8'b0;
    XRAM[45841] = 8'b0;
    XRAM[45842] = 8'b0;
    XRAM[45843] = 8'b0;
    XRAM[45844] = 8'b0;
    XRAM[45845] = 8'b0;
    XRAM[45846] = 8'b0;
    XRAM[45847] = 8'b0;
    XRAM[45848] = 8'b0;
    XRAM[45849] = 8'b0;
    XRAM[45850] = 8'b0;
    XRAM[45851] = 8'b0;
    XRAM[45852] = 8'b0;
    XRAM[45853] = 8'b0;
    XRAM[45854] = 8'b0;
    XRAM[45855] = 8'b0;
    XRAM[45856] = 8'b0;
    XRAM[45857] = 8'b0;
    XRAM[45858] = 8'b0;
    XRAM[45859] = 8'b0;
    XRAM[45860] = 8'b0;
    XRAM[45861] = 8'b0;
    XRAM[45862] = 8'b0;
    XRAM[45863] = 8'b0;
    XRAM[45864] = 8'b0;
    XRAM[45865] = 8'b0;
    XRAM[45866] = 8'b0;
    XRAM[45867] = 8'b0;
    XRAM[45868] = 8'b0;
    XRAM[45869] = 8'b0;
    XRAM[45870] = 8'b0;
    XRAM[45871] = 8'b0;
    XRAM[45872] = 8'b0;
    XRAM[45873] = 8'b0;
    XRAM[45874] = 8'b0;
    XRAM[45875] = 8'b0;
    XRAM[45876] = 8'b0;
    XRAM[45877] = 8'b0;
    XRAM[45878] = 8'b0;
    XRAM[45879] = 8'b0;
    XRAM[45880] = 8'b0;
    XRAM[45881] = 8'b0;
    XRAM[45882] = 8'b0;
    XRAM[45883] = 8'b0;
    XRAM[45884] = 8'b0;
    XRAM[45885] = 8'b0;
    XRAM[45886] = 8'b0;
    XRAM[45887] = 8'b0;
    XRAM[45888] = 8'b0;
    XRAM[45889] = 8'b0;
    XRAM[45890] = 8'b0;
    XRAM[45891] = 8'b0;
    XRAM[45892] = 8'b0;
    XRAM[45893] = 8'b0;
    XRAM[45894] = 8'b0;
    XRAM[45895] = 8'b0;
    XRAM[45896] = 8'b0;
    XRAM[45897] = 8'b0;
    XRAM[45898] = 8'b0;
    XRAM[45899] = 8'b0;
    XRAM[45900] = 8'b0;
    XRAM[45901] = 8'b0;
    XRAM[45902] = 8'b0;
    XRAM[45903] = 8'b0;
    XRAM[45904] = 8'b0;
    XRAM[45905] = 8'b0;
    XRAM[45906] = 8'b0;
    XRAM[45907] = 8'b0;
    XRAM[45908] = 8'b0;
    XRAM[45909] = 8'b0;
    XRAM[45910] = 8'b0;
    XRAM[45911] = 8'b0;
    XRAM[45912] = 8'b0;
    XRAM[45913] = 8'b0;
    XRAM[45914] = 8'b0;
    XRAM[45915] = 8'b0;
    XRAM[45916] = 8'b0;
    XRAM[45917] = 8'b0;
    XRAM[45918] = 8'b0;
    XRAM[45919] = 8'b0;
    XRAM[45920] = 8'b0;
    XRAM[45921] = 8'b0;
    XRAM[45922] = 8'b0;
    XRAM[45923] = 8'b0;
    XRAM[45924] = 8'b0;
    XRAM[45925] = 8'b0;
    XRAM[45926] = 8'b0;
    XRAM[45927] = 8'b0;
    XRAM[45928] = 8'b0;
    XRAM[45929] = 8'b0;
    XRAM[45930] = 8'b0;
    XRAM[45931] = 8'b0;
    XRAM[45932] = 8'b0;
    XRAM[45933] = 8'b0;
    XRAM[45934] = 8'b0;
    XRAM[45935] = 8'b0;
    XRAM[45936] = 8'b0;
    XRAM[45937] = 8'b0;
    XRAM[45938] = 8'b0;
    XRAM[45939] = 8'b0;
    XRAM[45940] = 8'b0;
    XRAM[45941] = 8'b0;
    XRAM[45942] = 8'b0;
    XRAM[45943] = 8'b0;
    XRAM[45944] = 8'b0;
    XRAM[45945] = 8'b0;
    XRAM[45946] = 8'b0;
    XRAM[45947] = 8'b0;
    XRAM[45948] = 8'b0;
    XRAM[45949] = 8'b0;
    XRAM[45950] = 8'b0;
    XRAM[45951] = 8'b0;
    XRAM[45952] = 8'b0;
    XRAM[45953] = 8'b0;
    XRAM[45954] = 8'b0;
    XRAM[45955] = 8'b0;
    XRAM[45956] = 8'b0;
    XRAM[45957] = 8'b0;
    XRAM[45958] = 8'b0;
    XRAM[45959] = 8'b0;
    XRAM[45960] = 8'b0;
    XRAM[45961] = 8'b0;
    XRAM[45962] = 8'b0;
    XRAM[45963] = 8'b0;
    XRAM[45964] = 8'b0;
    XRAM[45965] = 8'b0;
    XRAM[45966] = 8'b0;
    XRAM[45967] = 8'b0;
    XRAM[45968] = 8'b0;
    XRAM[45969] = 8'b0;
    XRAM[45970] = 8'b0;
    XRAM[45971] = 8'b0;
    XRAM[45972] = 8'b0;
    XRAM[45973] = 8'b0;
    XRAM[45974] = 8'b0;
    XRAM[45975] = 8'b0;
    XRAM[45976] = 8'b0;
    XRAM[45977] = 8'b0;
    XRAM[45978] = 8'b0;
    XRAM[45979] = 8'b0;
    XRAM[45980] = 8'b0;
    XRAM[45981] = 8'b0;
    XRAM[45982] = 8'b0;
    XRAM[45983] = 8'b0;
    XRAM[45984] = 8'b0;
    XRAM[45985] = 8'b0;
    XRAM[45986] = 8'b0;
    XRAM[45987] = 8'b0;
    XRAM[45988] = 8'b0;
    XRAM[45989] = 8'b0;
    XRAM[45990] = 8'b0;
    XRAM[45991] = 8'b0;
    XRAM[45992] = 8'b0;
    XRAM[45993] = 8'b0;
    XRAM[45994] = 8'b0;
    XRAM[45995] = 8'b0;
    XRAM[45996] = 8'b0;
    XRAM[45997] = 8'b0;
    XRAM[45998] = 8'b0;
    XRAM[45999] = 8'b0;
    XRAM[46000] = 8'b0;
    XRAM[46001] = 8'b0;
    XRAM[46002] = 8'b0;
    XRAM[46003] = 8'b0;
    XRAM[46004] = 8'b0;
    XRAM[46005] = 8'b0;
    XRAM[46006] = 8'b0;
    XRAM[46007] = 8'b0;
    XRAM[46008] = 8'b0;
    XRAM[46009] = 8'b0;
    XRAM[46010] = 8'b0;
    XRAM[46011] = 8'b0;
    XRAM[46012] = 8'b0;
    XRAM[46013] = 8'b0;
    XRAM[46014] = 8'b0;
    XRAM[46015] = 8'b0;
    XRAM[46016] = 8'b0;
    XRAM[46017] = 8'b0;
    XRAM[46018] = 8'b0;
    XRAM[46019] = 8'b0;
    XRAM[46020] = 8'b0;
    XRAM[46021] = 8'b0;
    XRAM[46022] = 8'b0;
    XRAM[46023] = 8'b0;
    XRAM[46024] = 8'b0;
    XRAM[46025] = 8'b0;
    XRAM[46026] = 8'b0;
    XRAM[46027] = 8'b0;
    XRAM[46028] = 8'b0;
    XRAM[46029] = 8'b0;
    XRAM[46030] = 8'b0;
    XRAM[46031] = 8'b0;
    XRAM[46032] = 8'b0;
    XRAM[46033] = 8'b0;
    XRAM[46034] = 8'b0;
    XRAM[46035] = 8'b0;
    XRAM[46036] = 8'b0;
    XRAM[46037] = 8'b0;
    XRAM[46038] = 8'b0;
    XRAM[46039] = 8'b0;
    XRAM[46040] = 8'b0;
    XRAM[46041] = 8'b0;
    XRAM[46042] = 8'b0;
    XRAM[46043] = 8'b0;
    XRAM[46044] = 8'b0;
    XRAM[46045] = 8'b0;
    XRAM[46046] = 8'b0;
    XRAM[46047] = 8'b0;
    XRAM[46048] = 8'b0;
    XRAM[46049] = 8'b0;
    XRAM[46050] = 8'b0;
    XRAM[46051] = 8'b0;
    XRAM[46052] = 8'b0;
    XRAM[46053] = 8'b0;
    XRAM[46054] = 8'b0;
    XRAM[46055] = 8'b0;
    XRAM[46056] = 8'b0;
    XRAM[46057] = 8'b0;
    XRAM[46058] = 8'b0;
    XRAM[46059] = 8'b0;
    XRAM[46060] = 8'b0;
    XRAM[46061] = 8'b0;
    XRAM[46062] = 8'b0;
    XRAM[46063] = 8'b0;
    XRAM[46064] = 8'b0;
    XRAM[46065] = 8'b0;
    XRAM[46066] = 8'b0;
    XRAM[46067] = 8'b0;
    XRAM[46068] = 8'b0;
    XRAM[46069] = 8'b0;
    XRAM[46070] = 8'b0;
    XRAM[46071] = 8'b0;
    XRAM[46072] = 8'b0;
    XRAM[46073] = 8'b0;
    XRAM[46074] = 8'b0;
    XRAM[46075] = 8'b0;
    XRAM[46076] = 8'b0;
    XRAM[46077] = 8'b0;
    XRAM[46078] = 8'b0;
    XRAM[46079] = 8'b0;
    XRAM[46080] = 8'b0;
    XRAM[46081] = 8'b0;
    XRAM[46082] = 8'b0;
    XRAM[46083] = 8'b0;
    XRAM[46084] = 8'b0;
    XRAM[46085] = 8'b0;
    XRAM[46086] = 8'b0;
    XRAM[46087] = 8'b0;
    XRAM[46088] = 8'b0;
    XRAM[46089] = 8'b0;
    XRAM[46090] = 8'b0;
    XRAM[46091] = 8'b0;
    XRAM[46092] = 8'b0;
    XRAM[46093] = 8'b0;
    XRAM[46094] = 8'b0;
    XRAM[46095] = 8'b0;
    XRAM[46096] = 8'b0;
    XRAM[46097] = 8'b0;
    XRAM[46098] = 8'b0;
    XRAM[46099] = 8'b0;
    XRAM[46100] = 8'b0;
    XRAM[46101] = 8'b0;
    XRAM[46102] = 8'b0;
    XRAM[46103] = 8'b0;
    XRAM[46104] = 8'b0;
    XRAM[46105] = 8'b0;
    XRAM[46106] = 8'b0;
    XRAM[46107] = 8'b0;
    XRAM[46108] = 8'b0;
    XRAM[46109] = 8'b0;
    XRAM[46110] = 8'b0;
    XRAM[46111] = 8'b0;
    XRAM[46112] = 8'b0;
    XRAM[46113] = 8'b0;
    XRAM[46114] = 8'b0;
    XRAM[46115] = 8'b0;
    XRAM[46116] = 8'b0;
    XRAM[46117] = 8'b0;
    XRAM[46118] = 8'b0;
    XRAM[46119] = 8'b0;
    XRAM[46120] = 8'b0;
    XRAM[46121] = 8'b0;
    XRAM[46122] = 8'b0;
    XRAM[46123] = 8'b0;
    XRAM[46124] = 8'b0;
    XRAM[46125] = 8'b0;
    XRAM[46126] = 8'b0;
    XRAM[46127] = 8'b0;
    XRAM[46128] = 8'b0;
    XRAM[46129] = 8'b0;
    XRAM[46130] = 8'b0;
    XRAM[46131] = 8'b0;
    XRAM[46132] = 8'b0;
    XRAM[46133] = 8'b0;
    XRAM[46134] = 8'b0;
    XRAM[46135] = 8'b0;
    XRAM[46136] = 8'b0;
    XRAM[46137] = 8'b0;
    XRAM[46138] = 8'b0;
    XRAM[46139] = 8'b0;
    XRAM[46140] = 8'b0;
    XRAM[46141] = 8'b0;
    XRAM[46142] = 8'b0;
    XRAM[46143] = 8'b0;
    XRAM[46144] = 8'b0;
    XRAM[46145] = 8'b0;
    XRAM[46146] = 8'b0;
    XRAM[46147] = 8'b0;
    XRAM[46148] = 8'b0;
    XRAM[46149] = 8'b0;
    XRAM[46150] = 8'b0;
    XRAM[46151] = 8'b0;
    XRAM[46152] = 8'b0;
    XRAM[46153] = 8'b0;
    XRAM[46154] = 8'b0;
    XRAM[46155] = 8'b0;
    XRAM[46156] = 8'b0;
    XRAM[46157] = 8'b0;
    XRAM[46158] = 8'b0;
    XRAM[46159] = 8'b0;
    XRAM[46160] = 8'b0;
    XRAM[46161] = 8'b0;
    XRAM[46162] = 8'b0;
    XRAM[46163] = 8'b0;
    XRAM[46164] = 8'b0;
    XRAM[46165] = 8'b0;
    XRAM[46166] = 8'b0;
    XRAM[46167] = 8'b0;
    XRAM[46168] = 8'b0;
    XRAM[46169] = 8'b0;
    XRAM[46170] = 8'b0;
    XRAM[46171] = 8'b0;
    XRAM[46172] = 8'b0;
    XRAM[46173] = 8'b0;
    XRAM[46174] = 8'b0;
    XRAM[46175] = 8'b0;
    XRAM[46176] = 8'b0;
    XRAM[46177] = 8'b0;
    XRAM[46178] = 8'b0;
    XRAM[46179] = 8'b0;
    XRAM[46180] = 8'b0;
    XRAM[46181] = 8'b0;
    XRAM[46182] = 8'b0;
    XRAM[46183] = 8'b0;
    XRAM[46184] = 8'b0;
    XRAM[46185] = 8'b0;
    XRAM[46186] = 8'b0;
    XRAM[46187] = 8'b0;
    XRAM[46188] = 8'b0;
    XRAM[46189] = 8'b0;
    XRAM[46190] = 8'b0;
    XRAM[46191] = 8'b0;
    XRAM[46192] = 8'b0;
    XRAM[46193] = 8'b0;
    XRAM[46194] = 8'b0;
    XRAM[46195] = 8'b0;
    XRAM[46196] = 8'b0;
    XRAM[46197] = 8'b0;
    XRAM[46198] = 8'b0;
    XRAM[46199] = 8'b0;
    XRAM[46200] = 8'b0;
    XRAM[46201] = 8'b0;
    XRAM[46202] = 8'b0;
    XRAM[46203] = 8'b0;
    XRAM[46204] = 8'b0;
    XRAM[46205] = 8'b0;
    XRAM[46206] = 8'b0;
    XRAM[46207] = 8'b0;
    XRAM[46208] = 8'b0;
    XRAM[46209] = 8'b0;
    XRAM[46210] = 8'b0;
    XRAM[46211] = 8'b0;
    XRAM[46212] = 8'b0;
    XRAM[46213] = 8'b0;
    XRAM[46214] = 8'b0;
    XRAM[46215] = 8'b0;
    XRAM[46216] = 8'b0;
    XRAM[46217] = 8'b0;
    XRAM[46218] = 8'b0;
    XRAM[46219] = 8'b0;
    XRAM[46220] = 8'b0;
    XRAM[46221] = 8'b0;
    XRAM[46222] = 8'b0;
    XRAM[46223] = 8'b0;
    XRAM[46224] = 8'b0;
    XRAM[46225] = 8'b0;
    XRAM[46226] = 8'b0;
    XRAM[46227] = 8'b0;
    XRAM[46228] = 8'b0;
    XRAM[46229] = 8'b0;
    XRAM[46230] = 8'b0;
    XRAM[46231] = 8'b0;
    XRAM[46232] = 8'b0;
    XRAM[46233] = 8'b0;
    XRAM[46234] = 8'b0;
    XRAM[46235] = 8'b0;
    XRAM[46236] = 8'b0;
    XRAM[46237] = 8'b0;
    XRAM[46238] = 8'b0;
    XRAM[46239] = 8'b0;
    XRAM[46240] = 8'b0;
    XRAM[46241] = 8'b0;
    XRAM[46242] = 8'b0;
    XRAM[46243] = 8'b0;
    XRAM[46244] = 8'b0;
    XRAM[46245] = 8'b0;
    XRAM[46246] = 8'b0;
    XRAM[46247] = 8'b0;
    XRAM[46248] = 8'b0;
    XRAM[46249] = 8'b0;
    XRAM[46250] = 8'b0;
    XRAM[46251] = 8'b0;
    XRAM[46252] = 8'b0;
    XRAM[46253] = 8'b0;
    XRAM[46254] = 8'b0;
    XRAM[46255] = 8'b0;
    XRAM[46256] = 8'b0;
    XRAM[46257] = 8'b0;
    XRAM[46258] = 8'b0;
    XRAM[46259] = 8'b0;
    XRAM[46260] = 8'b0;
    XRAM[46261] = 8'b0;
    XRAM[46262] = 8'b0;
    XRAM[46263] = 8'b0;
    XRAM[46264] = 8'b0;
    XRAM[46265] = 8'b0;
    XRAM[46266] = 8'b0;
    XRAM[46267] = 8'b0;
    XRAM[46268] = 8'b0;
    XRAM[46269] = 8'b0;
    XRAM[46270] = 8'b0;
    XRAM[46271] = 8'b0;
    XRAM[46272] = 8'b0;
    XRAM[46273] = 8'b0;
    XRAM[46274] = 8'b0;
    XRAM[46275] = 8'b0;
    XRAM[46276] = 8'b0;
    XRAM[46277] = 8'b0;
    XRAM[46278] = 8'b0;
    XRAM[46279] = 8'b0;
    XRAM[46280] = 8'b0;
    XRAM[46281] = 8'b0;
    XRAM[46282] = 8'b0;
    XRAM[46283] = 8'b0;
    XRAM[46284] = 8'b0;
    XRAM[46285] = 8'b0;
    XRAM[46286] = 8'b0;
    XRAM[46287] = 8'b0;
    XRAM[46288] = 8'b0;
    XRAM[46289] = 8'b0;
    XRAM[46290] = 8'b0;
    XRAM[46291] = 8'b0;
    XRAM[46292] = 8'b0;
    XRAM[46293] = 8'b0;
    XRAM[46294] = 8'b0;
    XRAM[46295] = 8'b0;
    XRAM[46296] = 8'b0;
    XRAM[46297] = 8'b0;
    XRAM[46298] = 8'b0;
    XRAM[46299] = 8'b0;
    XRAM[46300] = 8'b0;
    XRAM[46301] = 8'b0;
    XRAM[46302] = 8'b0;
    XRAM[46303] = 8'b0;
    XRAM[46304] = 8'b0;
    XRAM[46305] = 8'b0;
    XRAM[46306] = 8'b0;
    XRAM[46307] = 8'b0;
    XRAM[46308] = 8'b0;
    XRAM[46309] = 8'b0;
    XRAM[46310] = 8'b0;
    XRAM[46311] = 8'b0;
    XRAM[46312] = 8'b0;
    XRAM[46313] = 8'b0;
    XRAM[46314] = 8'b0;
    XRAM[46315] = 8'b0;
    XRAM[46316] = 8'b0;
    XRAM[46317] = 8'b0;
    XRAM[46318] = 8'b0;
    XRAM[46319] = 8'b0;
    XRAM[46320] = 8'b0;
    XRAM[46321] = 8'b0;
    XRAM[46322] = 8'b0;
    XRAM[46323] = 8'b0;
    XRAM[46324] = 8'b0;
    XRAM[46325] = 8'b0;
    XRAM[46326] = 8'b0;
    XRAM[46327] = 8'b0;
    XRAM[46328] = 8'b0;
    XRAM[46329] = 8'b0;
    XRAM[46330] = 8'b0;
    XRAM[46331] = 8'b0;
    XRAM[46332] = 8'b0;
    XRAM[46333] = 8'b0;
    XRAM[46334] = 8'b0;
    XRAM[46335] = 8'b0;
    XRAM[46336] = 8'b0;
    XRAM[46337] = 8'b0;
    XRAM[46338] = 8'b0;
    XRAM[46339] = 8'b0;
    XRAM[46340] = 8'b0;
    XRAM[46341] = 8'b0;
    XRAM[46342] = 8'b0;
    XRAM[46343] = 8'b0;
    XRAM[46344] = 8'b0;
    XRAM[46345] = 8'b0;
    XRAM[46346] = 8'b0;
    XRAM[46347] = 8'b0;
    XRAM[46348] = 8'b0;
    XRAM[46349] = 8'b0;
    XRAM[46350] = 8'b0;
    XRAM[46351] = 8'b0;
    XRAM[46352] = 8'b0;
    XRAM[46353] = 8'b0;
    XRAM[46354] = 8'b0;
    XRAM[46355] = 8'b0;
    XRAM[46356] = 8'b0;
    XRAM[46357] = 8'b0;
    XRAM[46358] = 8'b0;
    XRAM[46359] = 8'b0;
    XRAM[46360] = 8'b0;
    XRAM[46361] = 8'b0;
    XRAM[46362] = 8'b0;
    XRAM[46363] = 8'b0;
    XRAM[46364] = 8'b0;
    XRAM[46365] = 8'b0;
    XRAM[46366] = 8'b0;
    XRAM[46367] = 8'b0;
    XRAM[46368] = 8'b0;
    XRAM[46369] = 8'b0;
    XRAM[46370] = 8'b0;
    XRAM[46371] = 8'b0;
    XRAM[46372] = 8'b0;
    XRAM[46373] = 8'b0;
    XRAM[46374] = 8'b0;
    XRAM[46375] = 8'b0;
    XRAM[46376] = 8'b0;
    XRAM[46377] = 8'b0;
    XRAM[46378] = 8'b0;
    XRAM[46379] = 8'b0;
    XRAM[46380] = 8'b0;
    XRAM[46381] = 8'b0;
    XRAM[46382] = 8'b0;
    XRAM[46383] = 8'b0;
    XRAM[46384] = 8'b0;
    XRAM[46385] = 8'b0;
    XRAM[46386] = 8'b0;
    XRAM[46387] = 8'b0;
    XRAM[46388] = 8'b0;
    XRAM[46389] = 8'b0;
    XRAM[46390] = 8'b0;
    XRAM[46391] = 8'b0;
    XRAM[46392] = 8'b0;
    XRAM[46393] = 8'b0;
    XRAM[46394] = 8'b0;
    XRAM[46395] = 8'b0;
    XRAM[46396] = 8'b0;
    XRAM[46397] = 8'b0;
    XRAM[46398] = 8'b0;
    XRAM[46399] = 8'b0;
    XRAM[46400] = 8'b0;
    XRAM[46401] = 8'b0;
    XRAM[46402] = 8'b0;
    XRAM[46403] = 8'b0;
    XRAM[46404] = 8'b0;
    XRAM[46405] = 8'b0;
    XRAM[46406] = 8'b0;
    XRAM[46407] = 8'b0;
    XRAM[46408] = 8'b0;
    XRAM[46409] = 8'b0;
    XRAM[46410] = 8'b0;
    XRAM[46411] = 8'b0;
    XRAM[46412] = 8'b0;
    XRAM[46413] = 8'b0;
    XRAM[46414] = 8'b0;
    XRAM[46415] = 8'b0;
    XRAM[46416] = 8'b0;
    XRAM[46417] = 8'b0;
    XRAM[46418] = 8'b0;
    XRAM[46419] = 8'b0;
    XRAM[46420] = 8'b0;
    XRAM[46421] = 8'b0;
    XRAM[46422] = 8'b0;
    XRAM[46423] = 8'b0;
    XRAM[46424] = 8'b0;
    XRAM[46425] = 8'b0;
    XRAM[46426] = 8'b0;
    XRAM[46427] = 8'b0;
    XRAM[46428] = 8'b0;
    XRAM[46429] = 8'b0;
    XRAM[46430] = 8'b0;
    XRAM[46431] = 8'b0;
    XRAM[46432] = 8'b0;
    XRAM[46433] = 8'b0;
    XRAM[46434] = 8'b0;
    XRAM[46435] = 8'b0;
    XRAM[46436] = 8'b0;
    XRAM[46437] = 8'b0;
    XRAM[46438] = 8'b0;
    XRAM[46439] = 8'b0;
    XRAM[46440] = 8'b0;
    XRAM[46441] = 8'b0;
    XRAM[46442] = 8'b0;
    XRAM[46443] = 8'b0;
    XRAM[46444] = 8'b0;
    XRAM[46445] = 8'b0;
    XRAM[46446] = 8'b0;
    XRAM[46447] = 8'b0;
    XRAM[46448] = 8'b0;
    XRAM[46449] = 8'b0;
    XRAM[46450] = 8'b0;
    XRAM[46451] = 8'b0;
    XRAM[46452] = 8'b0;
    XRAM[46453] = 8'b0;
    XRAM[46454] = 8'b0;
    XRAM[46455] = 8'b0;
    XRAM[46456] = 8'b0;
    XRAM[46457] = 8'b0;
    XRAM[46458] = 8'b0;
    XRAM[46459] = 8'b0;
    XRAM[46460] = 8'b0;
    XRAM[46461] = 8'b0;
    XRAM[46462] = 8'b0;
    XRAM[46463] = 8'b0;
    XRAM[46464] = 8'b0;
    XRAM[46465] = 8'b0;
    XRAM[46466] = 8'b0;
    XRAM[46467] = 8'b0;
    XRAM[46468] = 8'b0;
    XRAM[46469] = 8'b0;
    XRAM[46470] = 8'b0;
    XRAM[46471] = 8'b0;
    XRAM[46472] = 8'b0;
    XRAM[46473] = 8'b0;
    XRAM[46474] = 8'b0;
    XRAM[46475] = 8'b0;
    XRAM[46476] = 8'b0;
    XRAM[46477] = 8'b0;
    XRAM[46478] = 8'b0;
    XRAM[46479] = 8'b0;
    XRAM[46480] = 8'b0;
    XRAM[46481] = 8'b0;
    XRAM[46482] = 8'b0;
    XRAM[46483] = 8'b0;
    XRAM[46484] = 8'b0;
    XRAM[46485] = 8'b0;
    XRAM[46486] = 8'b0;
    XRAM[46487] = 8'b0;
    XRAM[46488] = 8'b0;
    XRAM[46489] = 8'b0;
    XRAM[46490] = 8'b0;
    XRAM[46491] = 8'b0;
    XRAM[46492] = 8'b0;
    XRAM[46493] = 8'b0;
    XRAM[46494] = 8'b0;
    XRAM[46495] = 8'b0;
    XRAM[46496] = 8'b0;
    XRAM[46497] = 8'b0;
    XRAM[46498] = 8'b0;
    XRAM[46499] = 8'b0;
    XRAM[46500] = 8'b0;
    XRAM[46501] = 8'b0;
    XRAM[46502] = 8'b0;
    XRAM[46503] = 8'b0;
    XRAM[46504] = 8'b0;
    XRAM[46505] = 8'b0;
    XRAM[46506] = 8'b0;
    XRAM[46507] = 8'b0;
    XRAM[46508] = 8'b0;
    XRAM[46509] = 8'b0;
    XRAM[46510] = 8'b0;
    XRAM[46511] = 8'b0;
    XRAM[46512] = 8'b0;
    XRAM[46513] = 8'b0;
    XRAM[46514] = 8'b0;
    XRAM[46515] = 8'b0;
    XRAM[46516] = 8'b0;
    XRAM[46517] = 8'b0;
    XRAM[46518] = 8'b0;
    XRAM[46519] = 8'b0;
    XRAM[46520] = 8'b0;
    XRAM[46521] = 8'b0;
    XRAM[46522] = 8'b0;
    XRAM[46523] = 8'b0;
    XRAM[46524] = 8'b0;
    XRAM[46525] = 8'b0;
    XRAM[46526] = 8'b0;
    XRAM[46527] = 8'b0;
    XRAM[46528] = 8'b0;
    XRAM[46529] = 8'b0;
    XRAM[46530] = 8'b0;
    XRAM[46531] = 8'b0;
    XRAM[46532] = 8'b0;
    XRAM[46533] = 8'b0;
    XRAM[46534] = 8'b0;
    XRAM[46535] = 8'b0;
    XRAM[46536] = 8'b0;
    XRAM[46537] = 8'b0;
    XRAM[46538] = 8'b0;
    XRAM[46539] = 8'b0;
    XRAM[46540] = 8'b0;
    XRAM[46541] = 8'b0;
    XRAM[46542] = 8'b0;
    XRAM[46543] = 8'b0;
    XRAM[46544] = 8'b0;
    XRAM[46545] = 8'b0;
    XRAM[46546] = 8'b0;
    XRAM[46547] = 8'b0;
    XRAM[46548] = 8'b0;
    XRAM[46549] = 8'b0;
    XRAM[46550] = 8'b0;
    XRAM[46551] = 8'b0;
    XRAM[46552] = 8'b0;
    XRAM[46553] = 8'b0;
    XRAM[46554] = 8'b0;
    XRAM[46555] = 8'b0;
    XRAM[46556] = 8'b0;
    XRAM[46557] = 8'b0;
    XRAM[46558] = 8'b0;
    XRAM[46559] = 8'b0;
    XRAM[46560] = 8'b0;
    XRAM[46561] = 8'b0;
    XRAM[46562] = 8'b0;
    XRAM[46563] = 8'b0;
    XRAM[46564] = 8'b0;
    XRAM[46565] = 8'b0;
    XRAM[46566] = 8'b0;
    XRAM[46567] = 8'b0;
    XRAM[46568] = 8'b0;
    XRAM[46569] = 8'b0;
    XRAM[46570] = 8'b0;
    XRAM[46571] = 8'b0;
    XRAM[46572] = 8'b0;
    XRAM[46573] = 8'b0;
    XRAM[46574] = 8'b0;
    XRAM[46575] = 8'b0;
    XRAM[46576] = 8'b0;
    XRAM[46577] = 8'b0;
    XRAM[46578] = 8'b0;
    XRAM[46579] = 8'b0;
    XRAM[46580] = 8'b0;
    XRAM[46581] = 8'b0;
    XRAM[46582] = 8'b0;
    XRAM[46583] = 8'b0;
    XRAM[46584] = 8'b0;
    XRAM[46585] = 8'b0;
    XRAM[46586] = 8'b0;
    XRAM[46587] = 8'b0;
    XRAM[46588] = 8'b0;
    XRAM[46589] = 8'b0;
    XRAM[46590] = 8'b0;
    XRAM[46591] = 8'b0;
    XRAM[46592] = 8'b0;
    XRAM[46593] = 8'b0;
    XRAM[46594] = 8'b0;
    XRAM[46595] = 8'b0;
    XRAM[46596] = 8'b0;
    XRAM[46597] = 8'b0;
    XRAM[46598] = 8'b0;
    XRAM[46599] = 8'b0;
    XRAM[46600] = 8'b0;
    XRAM[46601] = 8'b0;
    XRAM[46602] = 8'b0;
    XRAM[46603] = 8'b0;
    XRAM[46604] = 8'b0;
    XRAM[46605] = 8'b0;
    XRAM[46606] = 8'b0;
    XRAM[46607] = 8'b0;
    XRAM[46608] = 8'b0;
    XRAM[46609] = 8'b0;
    XRAM[46610] = 8'b0;
    XRAM[46611] = 8'b0;
    XRAM[46612] = 8'b0;
    XRAM[46613] = 8'b0;
    XRAM[46614] = 8'b0;
    XRAM[46615] = 8'b0;
    XRAM[46616] = 8'b0;
    XRAM[46617] = 8'b0;
    XRAM[46618] = 8'b0;
    XRAM[46619] = 8'b0;
    XRAM[46620] = 8'b0;
    XRAM[46621] = 8'b0;
    XRAM[46622] = 8'b0;
    XRAM[46623] = 8'b0;
    XRAM[46624] = 8'b0;
    XRAM[46625] = 8'b0;
    XRAM[46626] = 8'b0;
    XRAM[46627] = 8'b0;
    XRAM[46628] = 8'b0;
    XRAM[46629] = 8'b0;
    XRAM[46630] = 8'b0;
    XRAM[46631] = 8'b0;
    XRAM[46632] = 8'b0;
    XRAM[46633] = 8'b0;
    XRAM[46634] = 8'b0;
    XRAM[46635] = 8'b0;
    XRAM[46636] = 8'b0;
    XRAM[46637] = 8'b0;
    XRAM[46638] = 8'b0;
    XRAM[46639] = 8'b0;
    XRAM[46640] = 8'b0;
    XRAM[46641] = 8'b0;
    XRAM[46642] = 8'b0;
    XRAM[46643] = 8'b0;
    XRAM[46644] = 8'b0;
    XRAM[46645] = 8'b0;
    XRAM[46646] = 8'b0;
    XRAM[46647] = 8'b0;
    XRAM[46648] = 8'b0;
    XRAM[46649] = 8'b0;
    XRAM[46650] = 8'b0;
    XRAM[46651] = 8'b0;
    XRAM[46652] = 8'b0;
    XRAM[46653] = 8'b0;
    XRAM[46654] = 8'b0;
    XRAM[46655] = 8'b0;
    XRAM[46656] = 8'b0;
    XRAM[46657] = 8'b0;
    XRAM[46658] = 8'b0;
    XRAM[46659] = 8'b0;
    XRAM[46660] = 8'b0;
    XRAM[46661] = 8'b0;
    XRAM[46662] = 8'b0;
    XRAM[46663] = 8'b0;
    XRAM[46664] = 8'b0;
    XRAM[46665] = 8'b0;
    XRAM[46666] = 8'b0;
    XRAM[46667] = 8'b0;
    XRAM[46668] = 8'b0;
    XRAM[46669] = 8'b0;
    XRAM[46670] = 8'b0;
    XRAM[46671] = 8'b0;
    XRAM[46672] = 8'b0;
    XRAM[46673] = 8'b0;
    XRAM[46674] = 8'b0;
    XRAM[46675] = 8'b0;
    XRAM[46676] = 8'b0;
    XRAM[46677] = 8'b0;
    XRAM[46678] = 8'b0;
    XRAM[46679] = 8'b0;
    XRAM[46680] = 8'b0;
    XRAM[46681] = 8'b0;
    XRAM[46682] = 8'b0;
    XRAM[46683] = 8'b0;
    XRAM[46684] = 8'b0;
    XRAM[46685] = 8'b0;
    XRAM[46686] = 8'b0;
    XRAM[46687] = 8'b0;
    XRAM[46688] = 8'b0;
    XRAM[46689] = 8'b0;
    XRAM[46690] = 8'b0;
    XRAM[46691] = 8'b0;
    XRAM[46692] = 8'b0;
    XRAM[46693] = 8'b0;
    XRAM[46694] = 8'b0;
    XRAM[46695] = 8'b0;
    XRAM[46696] = 8'b0;
    XRAM[46697] = 8'b0;
    XRAM[46698] = 8'b0;
    XRAM[46699] = 8'b0;
    XRAM[46700] = 8'b0;
    XRAM[46701] = 8'b0;
    XRAM[46702] = 8'b0;
    XRAM[46703] = 8'b0;
    XRAM[46704] = 8'b0;
    XRAM[46705] = 8'b0;
    XRAM[46706] = 8'b0;
    XRAM[46707] = 8'b0;
    XRAM[46708] = 8'b0;
    XRAM[46709] = 8'b0;
    XRAM[46710] = 8'b0;
    XRAM[46711] = 8'b0;
    XRAM[46712] = 8'b0;
    XRAM[46713] = 8'b0;
    XRAM[46714] = 8'b0;
    XRAM[46715] = 8'b0;
    XRAM[46716] = 8'b0;
    XRAM[46717] = 8'b0;
    XRAM[46718] = 8'b0;
    XRAM[46719] = 8'b0;
    XRAM[46720] = 8'b0;
    XRAM[46721] = 8'b0;
    XRAM[46722] = 8'b0;
    XRAM[46723] = 8'b0;
    XRAM[46724] = 8'b0;
    XRAM[46725] = 8'b0;
    XRAM[46726] = 8'b0;
    XRAM[46727] = 8'b0;
    XRAM[46728] = 8'b0;
    XRAM[46729] = 8'b0;
    XRAM[46730] = 8'b0;
    XRAM[46731] = 8'b0;
    XRAM[46732] = 8'b0;
    XRAM[46733] = 8'b0;
    XRAM[46734] = 8'b0;
    XRAM[46735] = 8'b0;
    XRAM[46736] = 8'b0;
    XRAM[46737] = 8'b0;
    XRAM[46738] = 8'b0;
    XRAM[46739] = 8'b0;
    XRAM[46740] = 8'b0;
    XRAM[46741] = 8'b0;
    XRAM[46742] = 8'b0;
    XRAM[46743] = 8'b0;
    XRAM[46744] = 8'b0;
    XRAM[46745] = 8'b0;
    XRAM[46746] = 8'b0;
    XRAM[46747] = 8'b0;
    XRAM[46748] = 8'b0;
    XRAM[46749] = 8'b0;
    XRAM[46750] = 8'b0;
    XRAM[46751] = 8'b0;
    XRAM[46752] = 8'b0;
    XRAM[46753] = 8'b0;
    XRAM[46754] = 8'b0;
    XRAM[46755] = 8'b0;
    XRAM[46756] = 8'b0;
    XRAM[46757] = 8'b0;
    XRAM[46758] = 8'b0;
    XRAM[46759] = 8'b0;
    XRAM[46760] = 8'b0;
    XRAM[46761] = 8'b0;
    XRAM[46762] = 8'b0;
    XRAM[46763] = 8'b0;
    XRAM[46764] = 8'b0;
    XRAM[46765] = 8'b0;
    XRAM[46766] = 8'b0;
    XRAM[46767] = 8'b0;
    XRAM[46768] = 8'b0;
    XRAM[46769] = 8'b0;
    XRAM[46770] = 8'b0;
    XRAM[46771] = 8'b0;
    XRAM[46772] = 8'b0;
    XRAM[46773] = 8'b0;
    XRAM[46774] = 8'b0;
    XRAM[46775] = 8'b0;
    XRAM[46776] = 8'b0;
    XRAM[46777] = 8'b0;
    XRAM[46778] = 8'b0;
    XRAM[46779] = 8'b0;
    XRAM[46780] = 8'b0;
    XRAM[46781] = 8'b0;
    XRAM[46782] = 8'b0;
    XRAM[46783] = 8'b0;
    XRAM[46784] = 8'b0;
    XRAM[46785] = 8'b0;
    XRAM[46786] = 8'b0;
    XRAM[46787] = 8'b0;
    XRAM[46788] = 8'b0;
    XRAM[46789] = 8'b0;
    XRAM[46790] = 8'b0;
    XRAM[46791] = 8'b0;
    XRAM[46792] = 8'b0;
    XRAM[46793] = 8'b0;
    XRAM[46794] = 8'b0;
    XRAM[46795] = 8'b0;
    XRAM[46796] = 8'b0;
    XRAM[46797] = 8'b0;
    XRAM[46798] = 8'b0;
    XRAM[46799] = 8'b0;
    XRAM[46800] = 8'b0;
    XRAM[46801] = 8'b0;
    XRAM[46802] = 8'b0;
    XRAM[46803] = 8'b0;
    XRAM[46804] = 8'b0;
    XRAM[46805] = 8'b0;
    XRAM[46806] = 8'b0;
    XRAM[46807] = 8'b0;
    XRAM[46808] = 8'b0;
    XRAM[46809] = 8'b0;
    XRAM[46810] = 8'b0;
    XRAM[46811] = 8'b0;
    XRAM[46812] = 8'b0;
    XRAM[46813] = 8'b0;
    XRAM[46814] = 8'b0;
    XRAM[46815] = 8'b0;
    XRAM[46816] = 8'b0;
    XRAM[46817] = 8'b0;
    XRAM[46818] = 8'b0;
    XRAM[46819] = 8'b0;
    XRAM[46820] = 8'b0;
    XRAM[46821] = 8'b0;
    XRAM[46822] = 8'b0;
    XRAM[46823] = 8'b0;
    XRAM[46824] = 8'b0;
    XRAM[46825] = 8'b0;
    XRAM[46826] = 8'b0;
    XRAM[46827] = 8'b0;
    XRAM[46828] = 8'b0;
    XRAM[46829] = 8'b0;
    XRAM[46830] = 8'b0;
    XRAM[46831] = 8'b0;
    XRAM[46832] = 8'b0;
    XRAM[46833] = 8'b0;
    XRAM[46834] = 8'b0;
    XRAM[46835] = 8'b0;
    XRAM[46836] = 8'b0;
    XRAM[46837] = 8'b0;
    XRAM[46838] = 8'b0;
    XRAM[46839] = 8'b0;
    XRAM[46840] = 8'b0;
    XRAM[46841] = 8'b0;
    XRAM[46842] = 8'b0;
    XRAM[46843] = 8'b0;
    XRAM[46844] = 8'b0;
    XRAM[46845] = 8'b0;
    XRAM[46846] = 8'b0;
    XRAM[46847] = 8'b0;
    XRAM[46848] = 8'b0;
    XRAM[46849] = 8'b0;
    XRAM[46850] = 8'b0;
    XRAM[46851] = 8'b0;
    XRAM[46852] = 8'b0;
    XRAM[46853] = 8'b0;
    XRAM[46854] = 8'b0;
    XRAM[46855] = 8'b0;
    XRAM[46856] = 8'b0;
    XRAM[46857] = 8'b0;
    XRAM[46858] = 8'b0;
    XRAM[46859] = 8'b0;
    XRAM[46860] = 8'b0;
    XRAM[46861] = 8'b0;
    XRAM[46862] = 8'b0;
    XRAM[46863] = 8'b0;
    XRAM[46864] = 8'b0;
    XRAM[46865] = 8'b0;
    XRAM[46866] = 8'b0;
    XRAM[46867] = 8'b0;
    XRAM[46868] = 8'b0;
    XRAM[46869] = 8'b0;
    XRAM[46870] = 8'b0;
    XRAM[46871] = 8'b0;
    XRAM[46872] = 8'b0;
    XRAM[46873] = 8'b0;
    XRAM[46874] = 8'b0;
    XRAM[46875] = 8'b0;
    XRAM[46876] = 8'b0;
    XRAM[46877] = 8'b0;
    XRAM[46878] = 8'b0;
    XRAM[46879] = 8'b0;
    XRAM[46880] = 8'b0;
    XRAM[46881] = 8'b0;
    XRAM[46882] = 8'b0;
    XRAM[46883] = 8'b0;
    XRAM[46884] = 8'b0;
    XRAM[46885] = 8'b0;
    XRAM[46886] = 8'b0;
    XRAM[46887] = 8'b0;
    XRAM[46888] = 8'b0;
    XRAM[46889] = 8'b0;
    XRAM[46890] = 8'b0;
    XRAM[46891] = 8'b0;
    XRAM[46892] = 8'b0;
    XRAM[46893] = 8'b0;
    XRAM[46894] = 8'b0;
    XRAM[46895] = 8'b0;
    XRAM[46896] = 8'b0;
    XRAM[46897] = 8'b0;
    XRAM[46898] = 8'b0;
    XRAM[46899] = 8'b0;
    XRAM[46900] = 8'b0;
    XRAM[46901] = 8'b0;
    XRAM[46902] = 8'b0;
    XRAM[46903] = 8'b0;
    XRAM[46904] = 8'b0;
    XRAM[46905] = 8'b0;
    XRAM[46906] = 8'b0;
    XRAM[46907] = 8'b0;
    XRAM[46908] = 8'b0;
    XRAM[46909] = 8'b0;
    XRAM[46910] = 8'b0;
    XRAM[46911] = 8'b0;
    XRAM[46912] = 8'b0;
    XRAM[46913] = 8'b0;
    XRAM[46914] = 8'b0;
    XRAM[46915] = 8'b0;
    XRAM[46916] = 8'b0;
    XRAM[46917] = 8'b0;
    XRAM[46918] = 8'b0;
    XRAM[46919] = 8'b0;
    XRAM[46920] = 8'b0;
    XRAM[46921] = 8'b0;
    XRAM[46922] = 8'b0;
    XRAM[46923] = 8'b0;
    XRAM[46924] = 8'b0;
    XRAM[46925] = 8'b0;
    XRAM[46926] = 8'b0;
    XRAM[46927] = 8'b0;
    XRAM[46928] = 8'b0;
    XRAM[46929] = 8'b0;
    XRAM[46930] = 8'b0;
    XRAM[46931] = 8'b0;
    XRAM[46932] = 8'b0;
    XRAM[46933] = 8'b0;
    XRAM[46934] = 8'b0;
    XRAM[46935] = 8'b0;
    XRAM[46936] = 8'b0;
    XRAM[46937] = 8'b0;
    XRAM[46938] = 8'b0;
    XRAM[46939] = 8'b0;
    XRAM[46940] = 8'b0;
    XRAM[46941] = 8'b0;
    XRAM[46942] = 8'b0;
    XRAM[46943] = 8'b0;
    XRAM[46944] = 8'b0;
    XRAM[46945] = 8'b0;
    XRAM[46946] = 8'b0;
    XRAM[46947] = 8'b0;
    XRAM[46948] = 8'b0;
    XRAM[46949] = 8'b0;
    XRAM[46950] = 8'b0;
    XRAM[46951] = 8'b0;
    XRAM[46952] = 8'b0;
    XRAM[46953] = 8'b0;
    XRAM[46954] = 8'b0;
    XRAM[46955] = 8'b0;
    XRAM[46956] = 8'b0;
    XRAM[46957] = 8'b0;
    XRAM[46958] = 8'b0;
    XRAM[46959] = 8'b0;
    XRAM[46960] = 8'b0;
    XRAM[46961] = 8'b0;
    XRAM[46962] = 8'b0;
    XRAM[46963] = 8'b0;
    XRAM[46964] = 8'b0;
    XRAM[46965] = 8'b0;
    XRAM[46966] = 8'b0;
    XRAM[46967] = 8'b0;
    XRAM[46968] = 8'b0;
    XRAM[46969] = 8'b0;
    XRAM[46970] = 8'b0;
    XRAM[46971] = 8'b0;
    XRAM[46972] = 8'b0;
    XRAM[46973] = 8'b0;
    XRAM[46974] = 8'b0;
    XRAM[46975] = 8'b0;
    XRAM[46976] = 8'b0;
    XRAM[46977] = 8'b0;
    XRAM[46978] = 8'b0;
    XRAM[46979] = 8'b0;
    XRAM[46980] = 8'b0;
    XRAM[46981] = 8'b0;
    XRAM[46982] = 8'b0;
    XRAM[46983] = 8'b0;
    XRAM[46984] = 8'b0;
    XRAM[46985] = 8'b0;
    XRAM[46986] = 8'b0;
    XRAM[46987] = 8'b0;
    XRAM[46988] = 8'b0;
    XRAM[46989] = 8'b0;
    XRAM[46990] = 8'b0;
    XRAM[46991] = 8'b0;
    XRAM[46992] = 8'b0;
    XRAM[46993] = 8'b0;
    XRAM[46994] = 8'b0;
    XRAM[46995] = 8'b0;
    XRAM[46996] = 8'b0;
    XRAM[46997] = 8'b0;
    XRAM[46998] = 8'b0;
    XRAM[46999] = 8'b0;
    XRAM[47000] = 8'b0;
    XRAM[47001] = 8'b0;
    XRAM[47002] = 8'b0;
    XRAM[47003] = 8'b0;
    XRAM[47004] = 8'b0;
    XRAM[47005] = 8'b0;
    XRAM[47006] = 8'b0;
    XRAM[47007] = 8'b0;
    XRAM[47008] = 8'b0;
    XRAM[47009] = 8'b0;
    XRAM[47010] = 8'b0;
    XRAM[47011] = 8'b0;
    XRAM[47012] = 8'b0;
    XRAM[47013] = 8'b0;
    XRAM[47014] = 8'b0;
    XRAM[47015] = 8'b0;
    XRAM[47016] = 8'b0;
    XRAM[47017] = 8'b0;
    XRAM[47018] = 8'b0;
    XRAM[47019] = 8'b0;
    XRAM[47020] = 8'b0;
    XRAM[47021] = 8'b0;
    XRAM[47022] = 8'b0;
    XRAM[47023] = 8'b0;
    XRAM[47024] = 8'b0;
    XRAM[47025] = 8'b0;
    XRAM[47026] = 8'b0;
    XRAM[47027] = 8'b0;
    XRAM[47028] = 8'b0;
    XRAM[47029] = 8'b0;
    XRAM[47030] = 8'b0;
    XRAM[47031] = 8'b0;
    XRAM[47032] = 8'b0;
    XRAM[47033] = 8'b0;
    XRAM[47034] = 8'b0;
    XRAM[47035] = 8'b0;
    XRAM[47036] = 8'b0;
    XRAM[47037] = 8'b0;
    XRAM[47038] = 8'b0;
    XRAM[47039] = 8'b0;
    XRAM[47040] = 8'b0;
    XRAM[47041] = 8'b0;
    XRAM[47042] = 8'b0;
    XRAM[47043] = 8'b0;
    XRAM[47044] = 8'b0;
    XRAM[47045] = 8'b0;
    XRAM[47046] = 8'b0;
    XRAM[47047] = 8'b0;
    XRAM[47048] = 8'b0;
    XRAM[47049] = 8'b0;
    XRAM[47050] = 8'b0;
    XRAM[47051] = 8'b0;
    XRAM[47052] = 8'b0;
    XRAM[47053] = 8'b0;
    XRAM[47054] = 8'b0;
    XRAM[47055] = 8'b0;
    XRAM[47056] = 8'b0;
    XRAM[47057] = 8'b0;
    XRAM[47058] = 8'b0;
    XRAM[47059] = 8'b0;
    XRAM[47060] = 8'b0;
    XRAM[47061] = 8'b0;
    XRAM[47062] = 8'b0;
    XRAM[47063] = 8'b0;
    XRAM[47064] = 8'b0;
    XRAM[47065] = 8'b0;
    XRAM[47066] = 8'b0;
    XRAM[47067] = 8'b0;
    XRAM[47068] = 8'b0;
    XRAM[47069] = 8'b0;
    XRAM[47070] = 8'b0;
    XRAM[47071] = 8'b0;
    XRAM[47072] = 8'b0;
    XRAM[47073] = 8'b0;
    XRAM[47074] = 8'b0;
    XRAM[47075] = 8'b0;
    XRAM[47076] = 8'b0;
    XRAM[47077] = 8'b0;
    XRAM[47078] = 8'b0;
    XRAM[47079] = 8'b0;
    XRAM[47080] = 8'b0;
    XRAM[47081] = 8'b0;
    XRAM[47082] = 8'b0;
    XRAM[47083] = 8'b0;
    XRAM[47084] = 8'b0;
    XRAM[47085] = 8'b0;
    XRAM[47086] = 8'b0;
    XRAM[47087] = 8'b0;
    XRAM[47088] = 8'b0;
    XRAM[47089] = 8'b0;
    XRAM[47090] = 8'b0;
    XRAM[47091] = 8'b0;
    XRAM[47092] = 8'b0;
    XRAM[47093] = 8'b0;
    XRAM[47094] = 8'b0;
    XRAM[47095] = 8'b0;
    XRAM[47096] = 8'b0;
    XRAM[47097] = 8'b0;
    XRAM[47098] = 8'b0;
    XRAM[47099] = 8'b0;
    XRAM[47100] = 8'b0;
    XRAM[47101] = 8'b0;
    XRAM[47102] = 8'b0;
    XRAM[47103] = 8'b0;
    XRAM[47104] = 8'b0;
    XRAM[47105] = 8'b0;
    XRAM[47106] = 8'b0;
    XRAM[47107] = 8'b0;
    XRAM[47108] = 8'b0;
    XRAM[47109] = 8'b0;
    XRAM[47110] = 8'b0;
    XRAM[47111] = 8'b0;
    XRAM[47112] = 8'b0;
    XRAM[47113] = 8'b0;
    XRAM[47114] = 8'b0;
    XRAM[47115] = 8'b0;
    XRAM[47116] = 8'b0;
    XRAM[47117] = 8'b0;
    XRAM[47118] = 8'b0;
    XRAM[47119] = 8'b0;
    XRAM[47120] = 8'b0;
    XRAM[47121] = 8'b0;
    XRAM[47122] = 8'b0;
    XRAM[47123] = 8'b0;
    XRAM[47124] = 8'b0;
    XRAM[47125] = 8'b0;
    XRAM[47126] = 8'b0;
    XRAM[47127] = 8'b0;
    XRAM[47128] = 8'b0;
    XRAM[47129] = 8'b0;
    XRAM[47130] = 8'b0;
    XRAM[47131] = 8'b0;
    XRAM[47132] = 8'b0;
    XRAM[47133] = 8'b0;
    XRAM[47134] = 8'b0;
    XRAM[47135] = 8'b0;
    XRAM[47136] = 8'b0;
    XRAM[47137] = 8'b0;
    XRAM[47138] = 8'b0;
    XRAM[47139] = 8'b0;
    XRAM[47140] = 8'b0;
    XRAM[47141] = 8'b0;
    XRAM[47142] = 8'b0;
    XRAM[47143] = 8'b0;
    XRAM[47144] = 8'b0;
    XRAM[47145] = 8'b0;
    XRAM[47146] = 8'b0;
    XRAM[47147] = 8'b0;
    XRAM[47148] = 8'b0;
    XRAM[47149] = 8'b0;
    XRAM[47150] = 8'b0;
    XRAM[47151] = 8'b0;
    XRAM[47152] = 8'b0;
    XRAM[47153] = 8'b0;
    XRAM[47154] = 8'b0;
    XRAM[47155] = 8'b0;
    XRAM[47156] = 8'b0;
    XRAM[47157] = 8'b0;
    XRAM[47158] = 8'b0;
    XRAM[47159] = 8'b0;
    XRAM[47160] = 8'b0;
    XRAM[47161] = 8'b0;
    XRAM[47162] = 8'b0;
    XRAM[47163] = 8'b0;
    XRAM[47164] = 8'b0;
    XRAM[47165] = 8'b0;
    XRAM[47166] = 8'b0;
    XRAM[47167] = 8'b0;
    XRAM[47168] = 8'b0;
    XRAM[47169] = 8'b0;
    XRAM[47170] = 8'b0;
    XRAM[47171] = 8'b0;
    XRAM[47172] = 8'b0;
    XRAM[47173] = 8'b0;
    XRAM[47174] = 8'b0;
    XRAM[47175] = 8'b0;
    XRAM[47176] = 8'b0;
    XRAM[47177] = 8'b0;
    XRAM[47178] = 8'b0;
    XRAM[47179] = 8'b0;
    XRAM[47180] = 8'b0;
    XRAM[47181] = 8'b0;
    XRAM[47182] = 8'b0;
    XRAM[47183] = 8'b0;
    XRAM[47184] = 8'b0;
    XRAM[47185] = 8'b0;
    XRAM[47186] = 8'b0;
    XRAM[47187] = 8'b0;
    XRAM[47188] = 8'b0;
    XRAM[47189] = 8'b0;
    XRAM[47190] = 8'b0;
    XRAM[47191] = 8'b0;
    XRAM[47192] = 8'b0;
    XRAM[47193] = 8'b0;
    XRAM[47194] = 8'b0;
    XRAM[47195] = 8'b0;
    XRAM[47196] = 8'b0;
    XRAM[47197] = 8'b0;
    XRAM[47198] = 8'b0;
    XRAM[47199] = 8'b0;
    XRAM[47200] = 8'b0;
    XRAM[47201] = 8'b0;
    XRAM[47202] = 8'b0;
    XRAM[47203] = 8'b0;
    XRAM[47204] = 8'b0;
    XRAM[47205] = 8'b0;
    XRAM[47206] = 8'b0;
    XRAM[47207] = 8'b0;
    XRAM[47208] = 8'b0;
    XRAM[47209] = 8'b0;
    XRAM[47210] = 8'b0;
    XRAM[47211] = 8'b0;
    XRAM[47212] = 8'b0;
    XRAM[47213] = 8'b0;
    XRAM[47214] = 8'b0;
    XRAM[47215] = 8'b0;
    XRAM[47216] = 8'b0;
    XRAM[47217] = 8'b0;
    XRAM[47218] = 8'b0;
    XRAM[47219] = 8'b0;
    XRAM[47220] = 8'b0;
    XRAM[47221] = 8'b0;
    XRAM[47222] = 8'b0;
    XRAM[47223] = 8'b0;
    XRAM[47224] = 8'b0;
    XRAM[47225] = 8'b0;
    XRAM[47226] = 8'b0;
    XRAM[47227] = 8'b0;
    XRAM[47228] = 8'b0;
    XRAM[47229] = 8'b0;
    XRAM[47230] = 8'b0;
    XRAM[47231] = 8'b0;
    XRAM[47232] = 8'b0;
    XRAM[47233] = 8'b0;
    XRAM[47234] = 8'b0;
    XRAM[47235] = 8'b0;
    XRAM[47236] = 8'b0;
    XRAM[47237] = 8'b0;
    XRAM[47238] = 8'b0;
    XRAM[47239] = 8'b0;
    XRAM[47240] = 8'b0;
    XRAM[47241] = 8'b0;
    XRAM[47242] = 8'b0;
    XRAM[47243] = 8'b0;
    XRAM[47244] = 8'b0;
    XRAM[47245] = 8'b0;
    XRAM[47246] = 8'b0;
    XRAM[47247] = 8'b0;
    XRAM[47248] = 8'b0;
    XRAM[47249] = 8'b0;
    XRAM[47250] = 8'b0;
    XRAM[47251] = 8'b0;
    XRAM[47252] = 8'b0;
    XRAM[47253] = 8'b0;
    XRAM[47254] = 8'b0;
    XRAM[47255] = 8'b0;
    XRAM[47256] = 8'b0;
    XRAM[47257] = 8'b0;
    XRAM[47258] = 8'b0;
    XRAM[47259] = 8'b0;
    XRAM[47260] = 8'b0;
    XRAM[47261] = 8'b0;
    XRAM[47262] = 8'b0;
    XRAM[47263] = 8'b0;
    XRAM[47264] = 8'b0;
    XRAM[47265] = 8'b0;
    XRAM[47266] = 8'b0;
    XRAM[47267] = 8'b0;
    XRAM[47268] = 8'b0;
    XRAM[47269] = 8'b0;
    XRAM[47270] = 8'b0;
    XRAM[47271] = 8'b0;
    XRAM[47272] = 8'b0;
    XRAM[47273] = 8'b0;
    XRAM[47274] = 8'b0;
    XRAM[47275] = 8'b0;
    XRAM[47276] = 8'b0;
    XRAM[47277] = 8'b0;
    XRAM[47278] = 8'b0;
    XRAM[47279] = 8'b0;
    XRAM[47280] = 8'b0;
    XRAM[47281] = 8'b0;
    XRAM[47282] = 8'b0;
    XRAM[47283] = 8'b0;
    XRAM[47284] = 8'b0;
    XRAM[47285] = 8'b0;
    XRAM[47286] = 8'b0;
    XRAM[47287] = 8'b0;
    XRAM[47288] = 8'b0;
    XRAM[47289] = 8'b0;
    XRAM[47290] = 8'b0;
    XRAM[47291] = 8'b0;
    XRAM[47292] = 8'b0;
    XRAM[47293] = 8'b0;
    XRAM[47294] = 8'b0;
    XRAM[47295] = 8'b0;
    XRAM[47296] = 8'b0;
    XRAM[47297] = 8'b0;
    XRAM[47298] = 8'b0;
    XRAM[47299] = 8'b0;
    XRAM[47300] = 8'b0;
    XRAM[47301] = 8'b0;
    XRAM[47302] = 8'b0;
    XRAM[47303] = 8'b0;
    XRAM[47304] = 8'b0;
    XRAM[47305] = 8'b0;
    XRAM[47306] = 8'b0;
    XRAM[47307] = 8'b0;
    XRAM[47308] = 8'b0;
    XRAM[47309] = 8'b0;
    XRAM[47310] = 8'b0;
    XRAM[47311] = 8'b0;
    XRAM[47312] = 8'b0;
    XRAM[47313] = 8'b0;
    XRAM[47314] = 8'b0;
    XRAM[47315] = 8'b0;
    XRAM[47316] = 8'b0;
    XRAM[47317] = 8'b0;
    XRAM[47318] = 8'b0;
    XRAM[47319] = 8'b0;
    XRAM[47320] = 8'b0;
    XRAM[47321] = 8'b0;
    XRAM[47322] = 8'b0;
    XRAM[47323] = 8'b0;
    XRAM[47324] = 8'b0;
    XRAM[47325] = 8'b0;
    XRAM[47326] = 8'b0;
    XRAM[47327] = 8'b0;
    XRAM[47328] = 8'b0;
    XRAM[47329] = 8'b0;
    XRAM[47330] = 8'b0;
    XRAM[47331] = 8'b0;
    XRAM[47332] = 8'b0;
    XRAM[47333] = 8'b0;
    XRAM[47334] = 8'b0;
    XRAM[47335] = 8'b0;
    XRAM[47336] = 8'b0;
    XRAM[47337] = 8'b0;
    XRAM[47338] = 8'b0;
    XRAM[47339] = 8'b0;
    XRAM[47340] = 8'b0;
    XRAM[47341] = 8'b0;
    XRAM[47342] = 8'b0;
    XRAM[47343] = 8'b0;
    XRAM[47344] = 8'b0;
    XRAM[47345] = 8'b0;
    XRAM[47346] = 8'b0;
    XRAM[47347] = 8'b0;
    XRAM[47348] = 8'b0;
    XRAM[47349] = 8'b0;
    XRAM[47350] = 8'b0;
    XRAM[47351] = 8'b0;
    XRAM[47352] = 8'b0;
    XRAM[47353] = 8'b0;
    XRAM[47354] = 8'b0;
    XRAM[47355] = 8'b0;
    XRAM[47356] = 8'b0;
    XRAM[47357] = 8'b0;
    XRAM[47358] = 8'b0;
    XRAM[47359] = 8'b0;
    XRAM[47360] = 8'b0;
    XRAM[47361] = 8'b0;
    XRAM[47362] = 8'b0;
    XRAM[47363] = 8'b0;
    XRAM[47364] = 8'b0;
    XRAM[47365] = 8'b0;
    XRAM[47366] = 8'b0;
    XRAM[47367] = 8'b0;
    XRAM[47368] = 8'b0;
    XRAM[47369] = 8'b0;
    XRAM[47370] = 8'b0;
    XRAM[47371] = 8'b0;
    XRAM[47372] = 8'b0;
    XRAM[47373] = 8'b0;
    XRAM[47374] = 8'b0;
    XRAM[47375] = 8'b0;
    XRAM[47376] = 8'b0;
    XRAM[47377] = 8'b0;
    XRAM[47378] = 8'b0;
    XRAM[47379] = 8'b0;
    XRAM[47380] = 8'b0;
    XRAM[47381] = 8'b0;
    XRAM[47382] = 8'b0;
    XRAM[47383] = 8'b0;
    XRAM[47384] = 8'b0;
    XRAM[47385] = 8'b0;
    XRAM[47386] = 8'b0;
    XRAM[47387] = 8'b0;
    XRAM[47388] = 8'b0;
    XRAM[47389] = 8'b0;
    XRAM[47390] = 8'b0;
    XRAM[47391] = 8'b0;
    XRAM[47392] = 8'b0;
    XRAM[47393] = 8'b0;
    XRAM[47394] = 8'b0;
    XRAM[47395] = 8'b0;
    XRAM[47396] = 8'b0;
    XRAM[47397] = 8'b0;
    XRAM[47398] = 8'b0;
    XRAM[47399] = 8'b0;
    XRAM[47400] = 8'b0;
    XRAM[47401] = 8'b0;
    XRAM[47402] = 8'b0;
    XRAM[47403] = 8'b0;
    XRAM[47404] = 8'b0;
    XRAM[47405] = 8'b0;
    XRAM[47406] = 8'b0;
    XRAM[47407] = 8'b0;
    XRAM[47408] = 8'b0;
    XRAM[47409] = 8'b0;
    XRAM[47410] = 8'b0;
    XRAM[47411] = 8'b0;
    XRAM[47412] = 8'b0;
    XRAM[47413] = 8'b0;
    XRAM[47414] = 8'b0;
    XRAM[47415] = 8'b0;
    XRAM[47416] = 8'b0;
    XRAM[47417] = 8'b0;
    XRAM[47418] = 8'b0;
    XRAM[47419] = 8'b0;
    XRAM[47420] = 8'b0;
    XRAM[47421] = 8'b0;
    XRAM[47422] = 8'b0;
    XRAM[47423] = 8'b0;
    XRAM[47424] = 8'b0;
    XRAM[47425] = 8'b0;
    XRAM[47426] = 8'b0;
    XRAM[47427] = 8'b0;
    XRAM[47428] = 8'b0;
    XRAM[47429] = 8'b0;
    XRAM[47430] = 8'b0;
    XRAM[47431] = 8'b0;
    XRAM[47432] = 8'b0;
    XRAM[47433] = 8'b0;
    XRAM[47434] = 8'b0;
    XRAM[47435] = 8'b0;
    XRAM[47436] = 8'b0;
    XRAM[47437] = 8'b0;
    XRAM[47438] = 8'b0;
    XRAM[47439] = 8'b0;
    XRAM[47440] = 8'b0;
    XRAM[47441] = 8'b0;
    XRAM[47442] = 8'b0;
    XRAM[47443] = 8'b0;
    XRAM[47444] = 8'b0;
    XRAM[47445] = 8'b0;
    XRAM[47446] = 8'b0;
    XRAM[47447] = 8'b0;
    XRAM[47448] = 8'b0;
    XRAM[47449] = 8'b0;
    XRAM[47450] = 8'b0;
    XRAM[47451] = 8'b0;
    XRAM[47452] = 8'b0;
    XRAM[47453] = 8'b0;
    XRAM[47454] = 8'b0;
    XRAM[47455] = 8'b0;
    XRAM[47456] = 8'b0;
    XRAM[47457] = 8'b0;
    XRAM[47458] = 8'b0;
    XRAM[47459] = 8'b0;
    XRAM[47460] = 8'b0;
    XRAM[47461] = 8'b0;
    XRAM[47462] = 8'b0;
    XRAM[47463] = 8'b0;
    XRAM[47464] = 8'b0;
    XRAM[47465] = 8'b0;
    XRAM[47466] = 8'b0;
    XRAM[47467] = 8'b0;
    XRAM[47468] = 8'b0;
    XRAM[47469] = 8'b0;
    XRAM[47470] = 8'b0;
    XRAM[47471] = 8'b0;
    XRAM[47472] = 8'b0;
    XRAM[47473] = 8'b0;
    XRAM[47474] = 8'b0;
    XRAM[47475] = 8'b0;
    XRAM[47476] = 8'b0;
    XRAM[47477] = 8'b0;
    XRAM[47478] = 8'b0;
    XRAM[47479] = 8'b0;
    XRAM[47480] = 8'b0;
    XRAM[47481] = 8'b0;
    XRAM[47482] = 8'b0;
    XRAM[47483] = 8'b0;
    XRAM[47484] = 8'b0;
    XRAM[47485] = 8'b0;
    XRAM[47486] = 8'b0;
    XRAM[47487] = 8'b0;
    XRAM[47488] = 8'b0;
    XRAM[47489] = 8'b0;
    XRAM[47490] = 8'b0;
    XRAM[47491] = 8'b0;
    XRAM[47492] = 8'b0;
    XRAM[47493] = 8'b0;
    XRAM[47494] = 8'b0;
    XRAM[47495] = 8'b0;
    XRAM[47496] = 8'b0;
    XRAM[47497] = 8'b0;
    XRAM[47498] = 8'b0;
    XRAM[47499] = 8'b0;
    XRAM[47500] = 8'b0;
    XRAM[47501] = 8'b0;
    XRAM[47502] = 8'b0;
    XRAM[47503] = 8'b0;
    XRAM[47504] = 8'b0;
    XRAM[47505] = 8'b0;
    XRAM[47506] = 8'b0;
    XRAM[47507] = 8'b0;
    XRAM[47508] = 8'b0;
    XRAM[47509] = 8'b0;
    XRAM[47510] = 8'b0;
    XRAM[47511] = 8'b0;
    XRAM[47512] = 8'b0;
    XRAM[47513] = 8'b0;
    XRAM[47514] = 8'b0;
    XRAM[47515] = 8'b0;
    XRAM[47516] = 8'b0;
    XRAM[47517] = 8'b0;
    XRAM[47518] = 8'b0;
    XRAM[47519] = 8'b0;
    XRAM[47520] = 8'b0;
    XRAM[47521] = 8'b0;
    XRAM[47522] = 8'b0;
    XRAM[47523] = 8'b0;
    XRAM[47524] = 8'b0;
    XRAM[47525] = 8'b0;
    XRAM[47526] = 8'b0;
    XRAM[47527] = 8'b0;
    XRAM[47528] = 8'b0;
    XRAM[47529] = 8'b0;
    XRAM[47530] = 8'b0;
    XRAM[47531] = 8'b0;
    XRAM[47532] = 8'b0;
    XRAM[47533] = 8'b0;
    XRAM[47534] = 8'b0;
    XRAM[47535] = 8'b0;
    XRAM[47536] = 8'b0;
    XRAM[47537] = 8'b0;
    XRAM[47538] = 8'b0;
    XRAM[47539] = 8'b0;
    XRAM[47540] = 8'b0;
    XRAM[47541] = 8'b0;
    XRAM[47542] = 8'b0;
    XRAM[47543] = 8'b0;
    XRAM[47544] = 8'b0;
    XRAM[47545] = 8'b0;
    XRAM[47546] = 8'b0;
    XRAM[47547] = 8'b0;
    XRAM[47548] = 8'b0;
    XRAM[47549] = 8'b0;
    XRAM[47550] = 8'b0;
    XRAM[47551] = 8'b0;
    XRAM[47552] = 8'b0;
    XRAM[47553] = 8'b0;
    XRAM[47554] = 8'b0;
    XRAM[47555] = 8'b0;
    XRAM[47556] = 8'b0;
    XRAM[47557] = 8'b0;
    XRAM[47558] = 8'b0;
    XRAM[47559] = 8'b0;
    XRAM[47560] = 8'b0;
    XRAM[47561] = 8'b0;
    XRAM[47562] = 8'b0;
    XRAM[47563] = 8'b0;
    XRAM[47564] = 8'b0;
    XRAM[47565] = 8'b0;
    XRAM[47566] = 8'b0;
    XRAM[47567] = 8'b0;
    XRAM[47568] = 8'b0;
    XRAM[47569] = 8'b0;
    XRAM[47570] = 8'b0;
    XRAM[47571] = 8'b0;
    XRAM[47572] = 8'b0;
    XRAM[47573] = 8'b0;
    XRAM[47574] = 8'b0;
    XRAM[47575] = 8'b0;
    XRAM[47576] = 8'b0;
    XRAM[47577] = 8'b0;
    XRAM[47578] = 8'b0;
    XRAM[47579] = 8'b0;
    XRAM[47580] = 8'b0;
    XRAM[47581] = 8'b0;
    XRAM[47582] = 8'b0;
    XRAM[47583] = 8'b0;
    XRAM[47584] = 8'b0;
    XRAM[47585] = 8'b0;
    XRAM[47586] = 8'b0;
    XRAM[47587] = 8'b0;
    XRAM[47588] = 8'b0;
    XRAM[47589] = 8'b0;
    XRAM[47590] = 8'b0;
    XRAM[47591] = 8'b0;
    XRAM[47592] = 8'b0;
    XRAM[47593] = 8'b0;
    XRAM[47594] = 8'b0;
    XRAM[47595] = 8'b0;
    XRAM[47596] = 8'b0;
    XRAM[47597] = 8'b0;
    XRAM[47598] = 8'b0;
    XRAM[47599] = 8'b0;
    XRAM[47600] = 8'b0;
    XRAM[47601] = 8'b0;
    XRAM[47602] = 8'b0;
    XRAM[47603] = 8'b0;
    XRAM[47604] = 8'b0;
    XRAM[47605] = 8'b0;
    XRAM[47606] = 8'b0;
    XRAM[47607] = 8'b0;
    XRAM[47608] = 8'b0;
    XRAM[47609] = 8'b0;
    XRAM[47610] = 8'b0;
    XRAM[47611] = 8'b0;
    XRAM[47612] = 8'b0;
    XRAM[47613] = 8'b0;
    XRAM[47614] = 8'b0;
    XRAM[47615] = 8'b0;
    XRAM[47616] = 8'b0;
    XRAM[47617] = 8'b0;
    XRAM[47618] = 8'b0;
    XRAM[47619] = 8'b0;
    XRAM[47620] = 8'b0;
    XRAM[47621] = 8'b0;
    XRAM[47622] = 8'b0;
    XRAM[47623] = 8'b0;
    XRAM[47624] = 8'b0;
    XRAM[47625] = 8'b0;
    XRAM[47626] = 8'b0;
    XRAM[47627] = 8'b0;
    XRAM[47628] = 8'b0;
    XRAM[47629] = 8'b0;
    XRAM[47630] = 8'b0;
    XRAM[47631] = 8'b0;
    XRAM[47632] = 8'b0;
    XRAM[47633] = 8'b0;
    XRAM[47634] = 8'b0;
    XRAM[47635] = 8'b0;
    XRAM[47636] = 8'b0;
    XRAM[47637] = 8'b0;
    XRAM[47638] = 8'b0;
    XRAM[47639] = 8'b0;
    XRAM[47640] = 8'b0;
    XRAM[47641] = 8'b0;
    XRAM[47642] = 8'b0;
    XRAM[47643] = 8'b0;
    XRAM[47644] = 8'b0;
    XRAM[47645] = 8'b0;
    XRAM[47646] = 8'b0;
    XRAM[47647] = 8'b0;
    XRAM[47648] = 8'b0;
    XRAM[47649] = 8'b0;
    XRAM[47650] = 8'b0;
    XRAM[47651] = 8'b0;
    XRAM[47652] = 8'b0;
    XRAM[47653] = 8'b0;
    XRAM[47654] = 8'b0;
    XRAM[47655] = 8'b0;
    XRAM[47656] = 8'b0;
    XRAM[47657] = 8'b0;
    XRAM[47658] = 8'b0;
    XRAM[47659] = 8'b0;
    XRAM[47660] = 8'b0;
    XRAM[47661] = 8'b0;
    XRAM[47662] = 8'b0;
    XRAM[47663] = 8'b0;
    XRAM[47664] = 8'b0;
    XRAM[47665] = 8'b0;
    XRAM[47666] = 8'b0;
    XRAM[47667] = 8'b0;
    XRAM[47668] = 8'b0;
    XRAM[47669] = 8'b0;
    XRAM[47670] = 8'b0;
    XRAM[47671] = 8'b0;
    XRAM[47672] = 8'b0;
    XRAM[47673] = 8'b0;
    XRAM[47674] = 8'b0;
    XRAM[47675] = 8'b0;
    XRAM[47676] = 8'b0;
    XRAM[47677] = 8'b0;
    XRAM[47678] = 8'b0;
    XRAM[47679] = 8'b0;
    XRAM[47680] = 8'b0;
    XRAM[47681] = 8'b0;
    XRAM[47682] = 8'b0;
    XRAM[47683] = 8'b0;
    XRAM[47684] = 8'b0;
    XRAM[47685] = 8'b0;
    XRAM[47686] = 8'b0;
    XRAM[47687] = 8'b0;
    XRAM[47688] = 8'b0;
    XRAM[47689] = 8'b0;
    XRAM[47690] = 8'b0;
    XRAM[47691] = 8'b0;
    XRAM[47692] = 8'b0;
    XRAM[47693] = 8'b0;
    XRAM[47694] = 8'b0;
    XRAM[47695] = 8'b0;
    XRAM[47696] = 8'b0;
    XRAM[47697] = 8'b0;
    XRAM[47698] = 8'b0;
    XRAM[47699] = 8'b0;
    XRAM[47700] = 8'b0;
    XRAM[47701] = 8'b0;
    XRAM[47702] = 8'b0;
    XRAM[47703] = 8'b0;
    XRAM[47704] = 8'b0;
    XRAM[47705] = 8'b0;
    XRAM[47706] = 8'b0;
    XRAM[47707] = 8'b0;
    XRAM[47708] = 8'b0;
    XRAM[47709] = 8'b0;
    XRAM[47710] = 8'b0;
    XRAM[47711] = 8'b0;
    XRAM[47712] = 8'b0;
    XRAM[47713] = 8'b0;
    XRAM[47714] = 8'b0;
    XRAM[47715] = 8'b0;
    XRAM[47716] = 8'b0;
    XRAM[47717] = 8'b0;
    XRAM[47718] = 8'b0;
    XRAM[47719] = 8'b0;
    XRAM[47720] = 8'b0;
    XRAM[47721] = 8'b0;
    XRAM[47722] = 8'b0;
    XRAM[47723] = 8'b0;
    XRAM[47724] = 8'b0;
    XRAM[47725] = 8'b0;
    XRAM[47726] = 8'b0;
    XRAM[47727] = 8'b0;
    XRAM[47728] = 8'b0;
    XRAM[47729] = 8'b0;
    XRAM[47730] = 8'b0;
    XRAM[47731] = 8'b0;
    XRAM[47732] = 8'b0;
    XRAM[47733] = 8'b0;
    XRAM[47734] = 8'b0;
    XRAM[47735] = 8'b0;
    XRAM[47736] = 8'b0;
    XRAM[47737] = 8'b0;
    XRAM[47738] = 8'b0;
    XRAM[47739] = 8'b0;
    XRAM[47740] = 8'b0;
    XRAM[47741] = 8'b0;
    XRAM[47742] = 8'b0;
    XRAM[47743] = 8'b0;
    XRAM[47744] = 8'b0;
    XRAM[47745] = 8'b0;
    XRAM[47746] = 8'b0;
    XRAM[47747] = 8'b0;
    XRAM[47748] = 8'b0;
    XRAM[47749] = 8'b0;
    XRAM[47750] = 8'b0;
    XRAM[47751] = 8'b0;
    XRAM[47752] = 8'b0;
    XRAM[47753] = 8'b0;
    XRAM[47754] = 8'b0;
    XRAM[47755] = 8'b0;
    XRAM[47756] = 8'b0;
    XRAM[47757] = 8'b0;
    XRAM[47758] = 8'b0;
    XRAM[47759] = 8'b0;
    XRAM[47760] = 8'b0;
    XRAM[47761] = 8'b0;
    XRAM[47762] = 8'b0;
    XRAM[47763] = 8'b0;
    XRAM[47764] = 8'b0;
    XRAM[47765] = 8'b0;
    XRAM[47766] = 8'b0;
    XRAM[47767] = 8'b0;
    XRAM[47768] = 8'b0;
    XRAM[47769] = 8'b0;
    XRAM[47770] = 8'b0;
    XRAM[47771] = 8'b0;
    XRAM[47772] = 8'b0;
    XRAM[47773] = 8'b0;
    XRAM[47774] = 8'b0;
    XRAM[47775] = 8'b0;
    XRAM[47776] = 8'b0;
    XRAM[47777] = 8'b0;
    XRAM[47778] = 8'b0;
    XRAM[47779] = 8'b0;
    XRAM[47780] = 8'b0;
    XRAM[47781] = 8'b0;
    XRAM[47782] = 8'b0;
    XRAM[47783] = 8'b0;
    XRAM[47784] = 8'b0;
    XRAM[47785] = 8'b0;
    XRAM[47786] = 8'b0;
    XRAM[47787] = 8'b0;
    XRAM[47788] = 8'b0;
    XRAM[47789] = 8'b0;
    XRAM[47790] = 8'b0;
    XRAM[47791] = 8'b0;
    XRAM[47792] = 8'b0;
    XRAM[47793] = 8'b0;
    XRAM[47794] = 8'b0;
    XRAM[47795] = 8'b0;
    XRAM[47796] = 8'b0;
    XRAM[47797] = 8'b0;
    XRAM[47798] = 8'b0;
    XRAM[47799] = 8'b0;
    XRAM[47800] = 8'b0;
    XRAM[47801] = 8'b0;
    XRAM[47802] = 8'b0;
    XRAM[47803] = 8'b0;
    XRAM[47804] = 8'b0;
    XRAM[47805] = 8'b0;
    XRAM[47806] = 8'b0;
    XRAM[47807] = 8'b0;
    XRAM[47808] = 8'b0;
    XRAM[47809] = 8'b0;
    XRAM[47810] = 8'b0;
    XRAM[47811] = 8'b0;
    XRAM[47812] = 8'b0;
    XRAM[47813] = 8'b0;
    XRAM[47814] = 8'b0;
    XRAM[47815] = 8'b0;
    XRAM[47816] = 8'b0;
    XRAM[47817] = 8'b0;
    XRAM[47818] = 8'b0;
    XRAM[47819] = 8'b0;
    XRAM[47820] = 8'b0;
    XRAM[47821] = 8'b0;
    XRAM[47822] = 8'b0;
    XRAM[47823] = 8'b0;
    XRAM[47824] = 8'b0;
    XRAM[47825] = 8'b0;
    XRAM[47826] = 8'b0;
    XRAM[47827] = 8'b0;
    XRAM[47828] = 8'b0;
    XRAM[47829] = 8'b0;
    XRAM[47830] = 8'b0;
    XRAM[47831] = 8'b0;
    XRAM[47832] = 8'b0;
    XRAM[47833] = 8'b0;
    XRAM[47834] = 8'b0;
    XRAM[47835] = 8'b0;
    XRAM[47836] = 8'b0;
    XRAM[47837] = 8'b0;
    XRAM[47838] = 8'b0;
    XRAM[47839] = 8'b0;
    XRAM[47840] = 8'b0;
    XRAM[47841] = 8'b0;
    XRAM[47842] = 8'b0;
    XRAM[47843] = 8'b0;
    XRAM[47844] = 8'b0;
    XRAM[47845] = 8'b0;
    XRAM[47846] = 8'b0;
    XRAM[47847] = 8'b0;
    XRAM[47848] = 8'b0;
    XRAM[47849] = 8'b0;
    XRAM[47850] = 8'b0;
    XRAM[47851] = 8'b0;
    XRAM[47852] = 8'b0;
    XRAM[47853] = 8'b0;
    XRAM[47854] = 8'b0;
    XRAM[47855] = 8'b0;
    XRAM[47856] = 8'b0;
    XRAM[47857] = 8'b0;
    XRAM[47858] = 8'b0;
    XRAM[47859] = 8'b0;
    XRAM[47860] = 8'b0;
    XRAM[47861] = 8'b0;
    XRAM[47862] = 8'b0;
    XRAM[47863] = 8'b0;
    XRAM[47864] = 8'b0;
    XRAM[47865] = 8'b0;
    XRAM[47866] = 8'b0;
    XRAM[47867] = 8'b0;
    XRAM[47868] = 8'b0;
    XRAM[47869] = 8'b0;
    XRAM[47870] = 8'b0;
    XRAM[47871] = 8'b0;
    XRAM[47872] = 8'b0;
    XRAM[47873] = 8'b0;
    XRAM[47874] = 8'b0;
    XRAM[47875] = 8'b0;
    XRAM[47876] = 8'b0;
    XRAM[47877] = 8'b0;
    XRAM[47878] = 8'b0;
    XRAM[47879] = 8'b0;
    XRAM[47880] = 8'b0;
    XRAM[47881] = 8'b0;
    XRAM[47882] = 8'b0;
    XRAM[47883] = 8'b0;
    XRAM[47884] = 8'b0;
    XRAM[47885] = 8'b0;
    XRAM[47886] = 8'b0;
    XRAM[47887] = 8'b0;
    XRAM[47888] = 8'b0;
    XRAM[47889] = 8'b0;
    XRAM[47890] = 8'b0;
    XRAM[47891] = 8'b0;
    XRAM[47892] = 8'b0;
    XRAM[47893] = 8'b0;
    XRAM[47894] = 8'b0;
    XRAM[47895] = 8'b0;
    XRAM[47896] = 8'b0;
    XRAM[47897] = 8'b0;
    XRAM[47898] = 8'b0;
    XRAM[47899] = 8'b0;
    XRAM[47900] = 8'b0;
    XRAM[47901] = 8'b0;
    XRAM[47902] = 8'b0;
    XRAM[47903] = 8'b0;
    XRAM[47904] = 8'b0;
    XRAM[47905] = 8'b0;
    XRAM[47906] = 8'b0;
    XRAM[47907] = 8'b0;
    XRAM[47908] = 8'b0;
    XRAM[47909] = 8'b0;
    XRAM[47910] = 8'b0;
    XRAM[47911] = 8'b0;
    XRAM[47912] = 8'b0;
    XRAM[47913] = 8'b0;
    XRAM[47914] = 8'b0;
    XRAM[47915] = 8'b0;
    XRAM[47916] = 8'b0;
    XRAM[47917] = 8'b0;
    XRAM[47918] = 8'b0;
    XRAM[47919] = 8'b0;
    XRAM[47920] = 8'b0;
    XRAM[47921] = 8'b0;
    XRAM[47922] = 8'b0;
    XRAM[47923] = 8'b0;
    XRAM[47924] = 8'b0;
    XRAM[47925] = 8'b0;
    XRAM[47926] = 8'b0;
    XRAM[47927] = 8'b0;
    XRAM[47928] = 8'b0;
    XRAM[47929] = 8'b0;
    XRAM[47930] = 8'b0;
    XRAM[47931] = 8'b0;
    XRAM[47932] = 8'b0;
    XRAM[47933] = 8'b0;
    XRAM[47934] = 8'b0;
    XRAM[47935] = 8'b0;
    XRAM[47936] = 8'b0;
    XRAM[47937] = 8'b0;
    XRAM[47938] = 8'b0;
    XRAM[47939] = 8'b0;
    XRAM[47940] = 8'b0;
    XRAM[47941] = 8'b0;
    XRAM[47942] = 8'b0;
    XRAM[47943] = 8'b0;
    XRAM[47944] = 8'b0;
    XRAM[47945] = 8'b0;
    XRAM[47946] = 8'b0;
    XRAM[47947] = 8'b0;
    XRAM[47948] = 8'b0;
    XRAM[47949] = 8'b0;
    XRAM[47950] = 8'b0;
    XRAM[47951] = 8'b0;
    XRAM[47952] = 8'b0;
    XRAM[47953] = 8'b0;
    XRAM[47954] = 8'b0;
    XRAM[47955] = 8'b0;
    XRAM[47956] = 8'b0;
    XRAM[47957] = 8'b0;
    XRAM[47958] = 8'b0;
    XRAM[47959] = 8'b0;
    XRAM[47960] = 8'b0;
    XRAM[47961] = 8'b0;
    XRAM[47962] = 8'b0;
    XRAM[47963] = 8'b0;
    XRAM[47964] = 8'b0;
    XRAM[47965] = 8'b0;
    XRAM[47966] = 8'b0;
    XRAM[47967] = 8'b0;
    XRAM[47968] = 8'b0;
    XRAM[47969] = 8'b0;
    XRAM[47970] = 8'b0;
    XRAM[47971] = 8'b0;
    XRAM[47972] = 8'b0;
    XRAM[47973] = 8'b0;
    XRAM[47974] = 8'b0;
    XRAM[47975] = 8'b0;
    XRAM[47976] = 8'b0;
    XRAM[47977] = 8'b0;
    XRAM[47978] = 8'b0;
    XRAM[47979] = 8'b0;
    XRAM[47980] = 8'b0;
    XRAM[47981] = 8'b0;
    XRAM[47982] = 8'b0;
    XRAM[47983] = 8'b0;
    XRAM[47984] = 8'b0;
    XRAM[47985] = 8'b0;
    XRAM[47986] = 8'b0;
    XRAM[47987] = 8'b0;
    XRAM[47988] = 8'b0;
    XRAM[47989] = 8'b0;
    XRAM[47990] = 8'b0;
    XRAM[47991] = 8'b0;
    XRAM[47992] = 8'b0;
    XRAM[47993] = 8'b0;
    XRAM[47994] = 8'b0;
    XRAM[47995] = 8'b0;
    XRAM[47996] = 8'b0;
    XRAM[47997] = 8'b0;
    XRAM[47998] = 8'b0;
    XRAM[47999] = 8'b0;
    XRAM[48000] = 8'b0;
    XRAM[48001] = 8'b0;
    XRAM[48002] = 8'b0;
    XRAM[48003] = 8'b0;
    XRAM[48004] = 8'b0;
    XRAM[48005] = 8'b0;
    XRAM[48006] = 8'b0;
    XRAM[48007] = 8'b0;
    XRAM[48008] = 8'b0;
    XRAM[48009] = 8'b0;
    XRAM[48010] = 8'b0;
    XRAM[48011] = 8'b0;
    XRAM[48012] = 8'b0;
    XRAM[48013] = 8'b0;
    XRAM[48014] = 8'b0;
    XRAM[48015] = 8'b0;
    XRAM[48016] = 8'b0;
    XRAM[48017] = 8'b0;
    XRAM[48018] = 8'b0;
    XRAM[48019] = 8'b0;
    XRAM[48020] = 8'b0;
    XRAM[48021] = 8'b0;
    XRAM[48022] = 8'b0;
    XRAM[48023] = 8'b0;
    XRAM[48024] = 8'b0;
    XRAM[48025] = 8'b0;
    XRAM[48026] = 8'b0;
    XRAM[48027] = 8'b0;
    XRAM[48028] = 8'b0;
    XRAM[48029] = 8'b0;
    XRAM[48030] = 8'b0;
    XRAM[48031] = 8'b0;
    XRAM[48032] = 8'b0;
    XRAM[48033] = 8'b0;
    XRAM[48034] = 8'b0;
    XRAM[48035] = 8'b0;
    XRAM[48036] = 8'b0;
    XRAM[48037] = 8'b0;
    XRAM[48038] = 8'b0;
    XRAM[48039] = 8'b0;
    XRAM[48040] = 8'b0;
    XRAM[48041] = 8'b0;
    XRAM[48042] = 8'b0;
    XRAM[48043] = 8'b0;
    XRAM[48044] = 8'b0;
    XRAM[48045] = 8'b0;
    XRAM[48046] = 8'b0;
    XRAM[48047] = 8'b0;
    XRAM[48048] = 8'b0;
    XRAM[48049] = 8'b0;
    XRAM[48050] = 8'b0;
    XRAM[48051] = 8'b0;
    XRAM[48052] = 8'b0;
    XRAM[48053] = 8'b0;
    XRAM[48054] = 8'b0;
    XRAM[48055] = 8'b0;
    XRAM[48056] = 8'b0;
    XRAM[48057] = 8'b0;
    XRAM[48058] = 8'b0;
    XRAM[48059] = 8'b0;
    XRAM[48060] = 8'b0;
    XRAM[48061] = 8'b0;
    XRAM[48062] = 8'b0;
    XRAM[48063] = 8'b0;
    XRAM[48064] = 8'b0;
    XRAM[48065] = 8'b0;
    XRAM[48066] = 8'b0;
    XRAM[48067] = 8'b0;
    XRAM[48068] = 8'b0;
    XRAM[48069] = 8'b0;
    XRAM[48070] = 8'b0;
    XRAM[48071] = 8'b0;
    XRAM[48072] = 8'b0;
    XRAM[48073] = 8'b0;
    XRAM[48074] = 8'b0;
    XRAM[48075] = 8'b0;
    XRAM[48076] = 8'b0;
    XRAM[48077] = 8'b0;
    XRAM[48078] = 8'b0;
    XRAM[48079] = 8'b0;
    XRAM[48080] = 8'b0;
    XRAM[48081] = 8'b0;
    XRAM[48082] = 8'b0;
    XRAM[48083] = 8'b0;
    XRAM[48084] = 8'b0;
    XRAM[48085] = 8'b0;
    XRAM[48086] = 8'b0;
    XRAM[48087] = 8'b0;
    XRAM[48088] = 8'b0;
    XRAM[48089] = 8'b0;
    XRAM[48090] = 8'b0;
    XRAM[48091] = 8'b0;
    XRAM[48092] = 8'b0;
    XRAM[48093] = 8'b0;
    XRAM[48094] = 8'b0;
    XRAM[48095] = 8'b0;
    XRAM[48096] = 8'b0;
    XRAM[48097] = 8'b0;
    XRAM[48098] = 8'b0;
    XRAM[48099] = 8'b0;
    XRAM[48100] = 8'b0;
    XRAM[48101] = 8'b0;
    XRAM[48102] = 8'b0;
    XRAM[48103] = 8'b0;
    XRAM[48104] = 8'b0;
    XRAM[48105] = 8'b0;
    XRAM[48106] = 8'b0;
    XRAM[48107] = 8'b0;
    XRAM[48108] = 8'b0;
    XRAM[48109] = 8'b0;
    XRAM[48110] = 8'b0;
    XRAM[48111] = 8'b0;
    XRAM[48112] = 8'b0;
    XRAM[48113] = 8'b0;
    XRAM[48114] = 8'b0;
    XRAM[48115] = 8'b0;
    XRAM[48116] = 8'b0;
    XRAM[48117] = 8'b0;
    XRAM[48118] = 8'b0;
    XRAM[48119] = 8'b0;
    XRAM[48120] = 8'b0;
    XRAM[48121] = 8'b0;
    XRAM[48122] = 8'b0;
    XRAM[48123] = 8'b0;
    XRAM[48124] = 8'b0;
    XRAM[48125] = 8'b0;
    XRAM[48126] = 8'b0;
    XRAM[48127] = 8'b0;
    XRAM[48128] = 8'b0;
    XRAM[48129] = 8'b0;
    XRAM[48130] = 8'b0;
    XRAM[48131] = 8'b0;
    XRAM[48132] = 8'b0;
    XRAM[48133] = 8'b0;
    XRAM[48134] = 8'b0;
    XRAM[48135] = 8'b0;
    XRAM[48136] = 8'b0;
    XRAM[48137] = 8'b0;
    XRAM[48138] = 8'b0;
    XRAM[48139] = 8'b0;
    XRAM[48140] = 8'b0;
    XRAM[48141] = 8'b0;
    XRAM[48142] = 8'b0;
    XRAM[48143] = 8'b0;
    XRAM[48144] = 8'b0;
    XRAM[48145] = 8'b0;
    XRAM[48146] = 8'b0;
    XRAM[48147] = 8'b0;
    XRAM[48148] = 8'b0;
    XRAM[48149] = 8'b0;
    XRAM[48150] = 8'b0;
    XRAM[48151] = 8'b0;
    XRAM[48152] = 8'b0;
    XRAM[48153] = 8'b0;
    XRAM[48154] = 8'b0;
    XRAM[48155] = 8'b0;
    XRAM[48156] = 8'b0;
    XRAM[48157] = 8'b0;
    XRAM[48158] = 8'b0;
    XRAM[48159] = 8'b0;
    XRAM[48160] = 8'b0;
    XRAM[48161] = 8'b0;
    XRAM[48162] = 8'b0;
    XRAM[48163] = 8'b0;
    XRAM[48164] = 8'b0;
    XRAM[48165] = 8'b0;
    XRAM[48166] = 8'b0;
    XRAM[48167] = 8'b0;
    XRAM[48168] = 8'b0;
    XRAM[48169] = 8'b0;
    XRAM[48170] = 8'b0;
    XRAM[48171] = 8'b0;
    XRAM[48172] = 8'b0;
    XRAM[48173] = 8'b0;
    XRAM[48174] = 8'b0;
    XRAM[48175] = 8'b0;
    XRAM[48176] = 8'b0;
    XRAM[48177] = 8'b0;
    XRAM[48178] = 8'b0;
    XRAM[48179] = 8'b0;
    XRAM[48180] = 8'b0;
    XRAM[48181] = 8'b0;
    XRAM[48182] = 8'b0;
    XRAM[48183] = 8'b0;
    XRAM[48184] = 8'b0;
    XRAM[48185] = 8'b0;
    XRAM[48186] = 8'b0;
    XRAM[48187] = 8'b0;
    XRAM[48188] = 8'b0;
    XRAM[48189] = 8'b0;
    XRAM[48190] = 8'b0;
    XRAM[48191] = 8'b0;
    XRAM[48192] = 8'b0;
    XRAM[48193] = 8'b0;
    XRAM[48194] = 8'b0;
    XRAM[48195] = 8'b0;
    XRAM[48196] = 8'b0;
    XRAM[48197] = 8'b0;
    XRAM[48198] = 8'b0;
    XRAM[48199] = 8'b0;
    XRAM[48200] = 8'b0;
    XRAM[48201] = 8'b0;
    XRAM[48202] = 8'b0;
    XRAM[48203] = 8'b0;
    XRAM[48204] = 8'b0;
    XRAM[48205] = 8'b0;
    XRAM[48206] = 8'b0;
    XRAM[48207] = 8'b0;
    XRAM[48208] = 8'b0;
    XRAM[48209] = 8'b0;
    XRAM[48210] = 8'b0;
    XRAM[48211] = 8'b0;
    XRAM[48212] = 8'b0;
    XRAM[48213] = 8'b0;
    XRAM[48214] = 8'b0;
    XRAM[48215] = 8'b0;
    XRAM[48216] = 8'b0;
    XRAM[48217] = 8'b0;
    XRAM[48218] = 8'b0;
    XRAM[48219] = 8'b0;
    XRAM[48220] = 8'b0;
    XRAM[48221] = 8'b0;
    XRAM[48222] = 8'b0;
    XRAM[48223] = 8'b0;
    XRAM[48224] = 8'b0;
    XRAM[48225] = 8'b0;
    XRAM[48226] = 8'b0;
    XRAM[48227] = 8'b0;
    XRAM[48228] = 8'b0;
    XRAM[48229] = 8'b0;
    XRAM[48230] = 8'b0;
    XRAM[48231] = 8'b0;
    XRAM[48232] = 8'b0;
    XRAM[48233] = 8'b0;
    XRAM[48234] = 8'b0;
    XRAM[48235] = 8'b0;
    XRAM[48236] = 8'b0;
    XRAM[48237] = 8'b0;
    XRAM[48238] = 8'b0;
    XRAM[48239] = 8'b0;
    XRAM[48240] = 8'b0;
    XRAM[48241] = 8'b0;
    XRAM[48242] = 8'b0;
    XRAM[48243] = 8'b0;
    XRAM[48244] = 8'b0;
    XRAM[48245] = 8'b0;
    XRAM[48246] = 8'b0;
    XRAM[48247] = 8'b0;
    XRAM[48248] = 8'b0;
    XRAM[48249] = 8'b0;
    XRAM[48250] = 8'b0;
    XRAM[48251] = 8'b0;
    XRAM[48252] = 8'b0;
    XRAM[48253] = 8'b0;
    XRAM[48254] = 8'b0;
    XRAM[48255] = 8'b0;
    XRAM[48256] = 8'b0;
    XRAM[48257] = 8'b0;
    XRAM[48258] = 8'b0;
    XRAM[48259] = 8'b0;
    XRAM[48260] = 8'b0;
    XRAM[48261] = 8'b0;
    XRAM[48262] = 8'b0;
    XRAM[48263] = 8'b0;
    XRAM[48264] = 8'b0;
    XRAM[48265] = 8'b0;
    XRAM[48266] = 8'b0;
    XRAM[48267] = 8'b0;
    XRAM[48268] = 8'b0;
    XRAM[48269] = 8'b0;
    XRAM[48270] = 8'b0;
    XRAM[48271] = 8'b0;
    XRAM[48272] = 8'b0;
    XRAM[48273] = 8'b0;
    XRAM[48274] = 8'b0;
    XRAM[48275] = 8'b0;
    XRAM[48276] = 8'b0;
    XRAM[48277] = 8'b0;
    XRAM[48278] = 8'b0;
    XRAM[48279] = 8'b0;
    XRAM[48280] = 8'b0;
    XRAM[48281] = 8'b0;
    XRAM[48282] = 8'b0;
    XRAM[48283] = 8'b0;
    XRAM[48284] = 8'b0;
    XRAM[48285] = 8'b0;
    XRAM[48286] = 8'b0;
    XRAM[48287] = 8'b0;
    XRAM[48288] = 8'b0;
    XRAM[48289] = 8'b0;
    XRAM[48290] = 8'b0;
    XRAM[48291] = 8'b0;
    XRAM[48292] = 8'b0;
    XRAM[48293] = 8'b0;
    XRAM[48294] = 8'b0;
    XRAM[48295] = 8'b0;
    XRAM[48296] = 8'b0;
    XRAM[48297] = 8'b0;
    XRAM[48298] = 8'b0;
    XRAM[48299] = 8'b0;
    XRAM[48300] = 8'b0;
    XRAM[48301] = 8'b0;
    XRAM[48302] = 8'b0;
    XRAM[48303] = 8'b0;
    XRAM[48304] = 8'b0;
    XRAM[48305] = 8'b0;
    XRAM[48306] = 8'b0;
    XRAM[48307] = 8'b0;
    XRAM[48308] = 8'b0;
    XRAM[48309] = 8'b0;
    XRAM[48310] = 8'b0;
    XRAM[48311] = 8'b0;
    XRAM[48312] = 8'b0;
    XRAM[48313] = 8'b0;
    XRAM[48314] = 8'b0;
    XRAM[48315] = 8'b0;
    XRAM[48316] = 8'b0;
    XRAM[48317] = 8'b0;
    XRAM[48318] = 8'b0;
    XRAM[48319] = 8'b0;
    XRAM[48320] = 8'b0;
    XRAM[48321] = 8'b0;
    XRAM[48322] = 8'b0;
    XRAM[48323] = 8'b0;
    XRAM[48324] = 8'b0;
    XRAM[48325] = 8'b0;
    XRAM[48326] = 8'b0;
    XRAM[48327] = 8'b0;
    XRAM[48328] = 8'b0;
    XRAM[48329] = 8'b0;
    XRAM[48330] = 8'b0;
    XRAM[48331] = 8'b0;
    XRAM[48332] = 8'b0;
    XRAM[48333] = 8'b0;
    XRAM[48334] = 8'b0;
    XRAM[48335] = 8'b0;
    XRAM[48336] = 8'b0;
    XRAM[48337] = 8'b0;
    XRAM[48338] = 8'b0;
    XRAM[48339] = 8'b0;
    XRAM[48340] = 8'b0;
    XRAM[48341] = 8'b0;
    XRAM[48342] = 8'b0;
    XRAM[48343] = 8'b0;
    XRAM[48344] = 8'b0;
    XRAM[48345] = 8'b0;
    XRAM[48346] = 8'b0;
    XRAM[48347] = 8'b0;
    XRAM[48348] = 8'b0;
    XRAM[48349] = 8'b0;
    XRAM[48350] = 8'b0;
    XRAM[48351] = 8'b0;
    XRAM[48352] = 8'b0;
    XRAM[48353] = 8'b0;
    XRAM[48354] = 8'b0;
    XRAM[48355] = 8'b0;
    XRAM[48356] = 8'b0;
    XRAM[48357] = 8'b0;
    XRAM[48358] = 8'b0;
    XRAM[48359] = 8'b0;
    XRAM[48360] = 8'b0;
    XRAM[48361] = 8'b0;
    XRAM[48362] = 8'b0;
    XRAM[48363] = 8'b0;
    XRAM[48364] = 8'b0;
    XRAM[48365] = 8'b0;
    XRAM[48366] = 8'b0;
    XRAM[48367] = 8'b0;
    XRAM[48368] = 8'b0;
    XRAM[48369] = 8'b0;
    XRAM[48370] = 8'b0;
    XRAM[48371] = 8'b0;
    XRAM[48372] = 8'b0;
    XRAM[48373] = 8'b0;
    XRAM[48374] = 8'b0;
    XRAM[48375] = 8'b0;
    XRAM[48376] = 8'b0;
    XRAM[48377] = 8'b0;
    XRAM[48378] = 8'b0;
    XRAM[48379] = 8'b0;
    XRAM[48380] = 8'b0;
    XRAM[48381] = 8'b0;
    XRAM[48382] = 8'b0;
    XRAM[48383] = 8'b0;
    XRAM[48384] = 8'b0;
    XRAM[48385] = 8'b0;
    XRAM[48386] = 8'b0;
    XRAM[48387] = 8'b0;
    XRAM[48388] = 8'b0;
    XRAM[48389] = 8'b0;
    XRAM[48390] = 8'b0;
    XRAM[48391] = 8'b0;
    XRAM[48392] = 8'b0;
    XRAM[48393] = 8'b0;
    XRAM[48394] = 8'b0;
    XRAM[48395] = 8'b0;
    XRAM[48396] = 8'b0;
    XRAM[48397] = 8'b0;
    XRAM[48398] = 8'b0;
    XRAM[48399] = 8'b0;
    XRAM[48400] = 8'b0;
    XRAM[48401] = 8'b0;
    XRAM[48402] = 8'b0;
    XRAM[48403] = 8'b0;
    XRAM[48404] = 8'b0;
    XRAM[48405] = 8'b0;
    XRAM[48406] = 8'b0;
    XRAM[48407] = 8'b0;
    XRAM[48408] = 8'b0;
    XRAM[48409] = 8'b0;
    XRAM[48410] = 8'b0;
    XRAM[48411] = 8'b0;
    XRAM[48412] = 8'b0;
    XRAM[48413] = 8'b0;
    XRAM[48414] = 8'b0;
    XRAM[48415] = 8'b0;
    XRAM[48416] = 8'b0;
    XRAM[48417] = 8'b0;
    XRAM[48418] = 8'b0;
    XRAM[48419] = 8'b0;
    XRAM[48420] = 8'b0;
    XRAM[48421] = 8'b0;
    XRAM[48422] = 8'b0;
    XRAM[48423] = 8'b0;
    XRAM[48424] = 8'b0;
    XRAM[48425] = 8'b0;
    XRAM[48426] = 8'b0;
    XRAM[48427] = 8'b0;
    XRAM[48428] = 8'b0;
    XRAM[48429] = 8'b0;
    XRAM[48430] = 8'b0;
    XRAM[48431] = 8'b0;
    XRAM[48432] = 8'b0;
    XRAM[48433] = 8'b0;
    XRAM[48434] = 8'b0;
    XRAM[48435] = 8'b0;
    XRAM[48436] = 8'b0;
    XRAM[48437] = 8'b0;
    XRAM[48438] = 8'b0;
    XRAM[48439] = 8'b0;
    XRAM[48440] = 8'b0;
    XRAM[48441] = 8'b0;
    XRAM[48442] = 8'b0;
    XRAM[48443] = 8'b0;
    XRAM[48444] = 8'b0;
    XRAM[48445] = 8'b0;
    XRAM[48446] = 8'b0;
    XRAM[48447] = 8'b0;
    XRAM[48448] = 8'b0;
    XRAM[48449] = 8'b0;
    XRAM[48450] = 8'b0;
    XRAM[48451] = 8'b0;
    XRAM[48452] = 8'b0;
    XRAM[48453] = 8'b0;
    XRAM[48454] = 8'b0;
    XRAM[48455] = 8'b0;
    XRAM[48456] = 8'b0;
    XRAM[48457] = 8'b0;
    XRAM[48458] = 8'b0;
    XRAM[48459] = 8'b0;
    XRAM[48460] = 8'b0;
    XRAM[48461] = 8'b0;
    XRAM[48462] = 8'b0;
    XRAM[48463] = 8'b0;
    XRAM[48464] = 8'b0;
    XRAM[48465] = 8'b0;
    XRAM[48466] = 8'b0;
    XRAM[48467] = 8'b0;
    XRAM[48468] = 8'b0;
    XRAM[48469] = 8'b0;
    XRAM[48470] = 8'b0;
    XRAM[48471] = 8'b0;
    XRAM[48472] = 8'b0;
    XRAM[48473] = 8'b0;
    XRAM[48474] = 8'b0;
    XRAM[48475] = 8'b0;
    XRAM[48476] = 8'b0;
    XRAM[48477] = 8'b0;
    XRAM[48478] = 8'b0;
    XRAM[48479] = 8'b0;
    XRAM[48480] = 8'b0;
    XRAM[48481] = 8'b0;
    XRAM[48482] = 8'b0;
    XRAM[48483] = 8'b0;
    XRAM[48484] = 8'b0;
    XRAM[48485] = 8'b0;
    XRAM[48486] = 8'b0;
    XRAM[48487] = 8'b0;
    XRAM[48488] = 8'b0;
    XRAM[48489] = 8'b0;
    XRAM[48490] = 8'b0;
    XRAM[48491] = 8'b0;
    XRAM[48492] = 8'b0;
    XRAM[48493] = 8'b0;
    XRAM[48494] = 8'b0;
    XRAM[48495] = 8'b0;
    XRAM[48496] = 8'b0;
    XRAM[48497] = 8'b0;
    XRAM[48498] = 8'b0;
    XRAM[48499] = 8'b0;
    XRAM[48500] = 8'b0;
    XRAM[48501] = 8'b0;
    XRAM[48502] = 8'b0;
    XRAM[48503] = 8'b0;
    XRAM[48504] = 8'b0;
    XRAM[48505] = 8'b0;
    XRAM[48506] = 8'b0;
    XRAM[48507] = 8'b0;
    XRAM[48508] = 8'b0;
    XRAM[48509] = 8'b0;
    XRAM[48510] = 8'b0;
    XRAM[48511] = 8'b0;
    XRAM[48512] = 8'b0;
    XRAM[48513] = 8'b0;
    XRAM[48514] = 8'b0;
    XRAM[48515] = 8'b0;
    XRAM[48516] = 8'b0;
    XRAM[48517] = 8'b0;
    XRAM[48518] = 8'b0;
    XRAM[48519] = 8'b0;
    XRAM[48520] = 8'b0;
    XRAM[48521] = 8'b0;
    XRAM[48522] = 8'b0;
    XRAM[48523] = 8'b0;
    XRAM[48524] = 8'b0;
    XRAM[48525] = 8'b0;
    XRAM[48526] = 8'b0;
    XRAM[48527] = 8'b0;
    XRAM[48528] = 8'b0;
    XRAM[48529] = 8'b0;
    XRAM[48530] = 8'b0;
    XRAM[48531] = 8'b0;
    XRAM[48532] = 8'b0;
    XRAM[48533] = 8'b0;
    XRAM[48534] = 8'b0;
    XRAM[48535] = 8'b0;
    XRAM[48536] = 8'b0;
    XRAM[48537] = 8'b0;
    XRAM[48538] = 8'b0;
    XRAM[48539] = 8'b0;
    XRAM[48540] = 8'b0;
    XRAM[48541] = 8'b0;
    XRAM[48542] = 8'b0;
    XRAM[48543] = 8'b0;
    XRAM[48544] = 8'b0;
    XRAM[48545] = 8'b0;
    XRAM[48546] = 8'b0;
    XRAM[48547] = 8'b0;
    XRAM[48548] = 8'b0;
    XRAM[48549] = 8'b0;
    XRAM[48550] = 8'b0;
    XRAM[48551] = 8'b0;
    XRAM[48552] = 8'b0;
    XRAM[48553] = 8'b0;
    XRAM[48554] = 8'b0;
    XRAM[48555] = 8'b0;
    XRAM[48556] = 8'b0;
    XRAM[48557] = 8'b0;
    XRAM[48558] = 8'b0;
    XRAM[48559] = 8'b0;
    XRAM[48560] = 8'b0;
    XRAM[48561] = 8'b0;
    XRAM[48562] = 8'b0;
    XRAM[48563] = 8'b0;
    XRAM[48564] = 8'b0;
    XRAM[48565] = 8'b0;
    XRAM[48566] = 8'b0;
    XRAM[48567] = 8'b0;
    XRAM[48568] = 8'b0;
    XRAM[48569] = 8'b0;
    XRAM[48570] = 8'b0;
    XRAM[48571] = 8'b0;
    XRAM[48572] = 8'b0;
    XRAM[48573] = 8'b0;
    XRAM[48574] = 8'b0;
    XRAM[48575] = 8'b0;
    XRAM[48576] = 8'b0;
    XRAM[48577] = 8'b0;
    XRAM[48578] = 8'b0;
    XRAM[48579] = 8'b0;
    XRAM[48580] = 8'b0;
    XRAM[48581] = 8'b0;
    XRAM[48582] = 8'b0;
    XRAM[48583] = 8'b0;
    XRAM[48584] = 8'b0;
    XRAM[48585] = 8'b0;
    XRAM[48586] = 8'b0;
    XRAM[48587] = 8'b0;
    XRAM[48588] = 8'b0;
    XRAM[48589] = 8'b0;
    XRAM[48590] = 8'b0;
    XRAM[48591] = 8'b0;
    XRAM[48592] = 8'b0;
    XRAM[48593] = 8'b0;
    XRAM[48594] = 8'b0;
    XRAM[48595] = 8'b0;
    XRAM[48596] = 8'b0;
    XRAM[48597] = 8'b0;
    XRAM[48598] = 8'b0;
    XRAM[48599] = 8'b0;
    XRAM[48600] = 8'b0;
    XRAM[48601] = 8'b0;
    XRAM[48602] = 8'b0;
    XRAM[48603] = 8'b0;
    XRAM[48604] = 8'b0;
    XRAM[48605] = 8'b0;
    XRAM[48606] = 8'b0;
    XRAM[48607] = 8'b0;
    XRAM[48608] = 8'b0;
    XRAM[48609] = 8'b0;
    XRAM[48610] = 8'b0;
    XRAM[48611] = 8'b0;
    XRAM[48612] = 8'b0;
    XRAM[48613] = 8'b0;
    XRAM[48614] = 8'b0;
    XRAM[48615] = 8'b0;
    XRAM[48616] = 8'b0;
    XRAM[48617] = 8'b0;
    XRAM[48618] = 8'b0;
    XRAM[48619] = 8'b0;
    XRAM[48620] = 8'b0;
    XRAM[48621] = 8'b0;
    XRAM[48622] = 8'b0;
    XRAM[48623] = 8'b0;
    XRAM[48624] = 8'b0;
    XRAM[48625] = 8'b0;
    XRAM[48626] = 8'b0;
    XRAM[48627] = 8'b0;
    XRAM[48628] = 8'b0;
    XRAM[48629] = 8'b0;
    XRAM[48630] = 8'b0;
    XRAM[48631] = 8'b0;
    XRAM[48632] = 8'b0;
    XRAM[48633] = 8'b0;
    XRAM[48634] = 8'b0;
    XRAM[48635] = 8'b0;
    XRAM[48636] = 8'b0;
    XRAM[48637] = 8'b0;
    XRAM[48638] = 8'b0;
    XRAM[48639] = 8'b0;
    XRAM[48640] = 8'b0;
    XRAM[48641] = 8'b0;
    XRAM[48642] = 8'b0;
    XRAM[48643] = 8'b0;
    XRAM[48644] = 8'b0;
    XRAM[48645] = 8'b0;
    XRAM[48646] = 8'b0;
    XRAM[48647] = 8'b0;
    XRAM[48648] = 8'b0;
    XRAM[48649] = 8'b0;
    XRAM[48650] = 8'b0;
    XRAM[48651] = 8'b0;
    XRAM[48652] = 8'b0;
    XRAM[48653] = 8'b0;
    XRAM[48654] = 8'b0;
    XRAM[48655] = 8'b0;
    XRAM[48656] = 8'b0;
    XRAM[48657] = 8'b0;
    XRAM[48658] = 8'b0;
    XRAM[48659] = 8'b0;
    XRAM[48660] = 8'b0;
    XRAM[48661] = 8'b0;
    XRAM[48662] = 8'b0;
    XRAM[48663] = 8'b0;
    XRAM[48664] = 8'b0;
    XRAM[48665] = 8'b0;
    XRAM[48666] = 8'b0;
    XRAM[48667] = 8'b0;
    XRAM[48668] = 8'b0;
    XRAM[48669] = 8'b0;
    XRAM[48670] = 8'b0;
    XRAM[48671] = 8'b0;
    XRAM[48672] = 8'b0;
    XRAM[48673] = 8'b0;
    XRAM[48674] = 8'b0;
    XRAM[48675] = 8'b0;
    XRAM[48676] = 8'b0;
    XRAM[48677] = 8'b0;
    XRAM[48678] = 8'b0;
    XRAM[48679] = 8'b0;
    XRAM[48680] = 8'b0;
    XRAM[48681] = 8'b0;
    XRAM[48682] = 8'b0;
    XRAM[48683] = 8'b0;
    XRAM[48684] = 8'b0;
    XRAM[48685] = 8'b0;
    XRAM[48686] = 8'b0;
    XRAM[48687] = 8'b0;
    XRAM[48688] = 8'b0;
    XRAM[48689] = 8'b0;
    XRAM[48690] = 8'b0;
    XRAM[48691] = 8'b0;
    XRAM[48692] = 8'b0;
    XRAM[48693] = 8'b0;
    XRAM[48694] = 8'b0;
    XRAM[48695] = 8'b0;
    XRAM[48696] = 8'b0;
    XRAM[48697] = 8'b0;
    XRAM[48698] = 8'b0;
    XRAM[48699] = 8'b0;
    XRAM[48700] = 8'b0;
    XRAM[48701] = 8'b0;
    XRAM[48702] = 8'b0;
    XRAM[48703] = 8'b0;
    XRAM[48704] = 8'b0;
    XRAM[48705] = 8'b0;
    XRAM[48706] = 8'b0;
    XRAM[48707] = 8'b0;
    XRAM[48708] = 8'b0;
    XRAM[48709] = 8'b0;
    XRAM[48710] = 8'b0;
    XRAM[48711] = 8'b0;
    XRAM[48712] = 8'b0;
    XRAM[48713] = 8'b0;
    XRAM[48714] = 8'b0;
    XRAM[48715] = 8'b0;
    XRAM[48716] = 8'b0;
    XRAM[48717] = 8'b0;
    XRAM[48718] = 8'b0;
    XRAM[48719] = 8'b0;
    XRAM[48720] = 8'b0;
    XRAM[48721] = 8'b0;
    XRAM[48722] = 8'b0;
    XRAM[48723] = 8'b0;
    XRAM[48724] = 8'b0;
    XRAM[48725] = 8'b0;
    XRAM[48726] = 8'b0;
    XRAM[48727] = 8'b0;
    XRAM[48728] = 8'b0;
    XRAM[48729] = 8'b0;
    XRAM[48730] = 8'b0;
    XRAM[48731] = 8'b0;
    XRAM[48732] = 8'b0;
    XRAM[48733] = 8'b0;
    XRAM[48734] = 8'b0;
    XRAM[48735] = 8'b0;
    XRAM[48736] = 8'b0;
    XRAM[48737] = 8'b0;
    XRAM[48738] = 8'b0;
    XRAM[48739] = 8'b0;
    XRAM[48740] = 8'b0;
    XRAM[48741] = 8'b0;
    XRAM[48742] = 8'b0;
    XRAM[48743] = 8'b0;
    XRAM[48744] = 8'b0;
    XRAM[48745] = 8'b0;
    XRAM[48746] = 8'b0;
    XRAM[48747] = 8'b0;
    XRAM[48748] = 8'b0;
    XRAM[48749] = 8'b0;
    XRAM[48750] = 8'b0;
    XRAM[48751] = 8'b0;
    XRAM[48752] = 8'b0;
    XRAM[48753] = 8'b0;
    XRAM[48754] = 8'b0;
    XRAM[48755] = 8'b0;
    XRAM[48756] = 8'b0;
    XRAM[48757] = 8'b0;
    XRAM[48758] = 8'b0;
    XRAM[48759] = 8'b0;
    XRAM[48760] = 8'b0;
    XRAM[48761] = 8'b0;
    XRAM[48762] = 8'b0;
    XRAM[48763] = 8'b0;
    XRAM[48764] = 8'b0;
    XRAM[48765] = 8'b0;
    XRAM[48766] = 8'b0;
    XRAM[48767] = 8'b0;
    XRAM[48768] = 8'b0;
    XRAM[48769] = 8'b0;
    XRAM[48770] = 8'b0;
    XRAM[48771] = 8'b0;
    XRAM[48772] = 8'b0;
    XRAM[48773] = 8'b0;
    XRAM[48774] = 8'b0;
    XRAM[48775] = 8'b0;
    XRAM[48776] = 8'b0;
    XRAM[48777] = 8'b0;
    XRAM[48778] = 8'b0;
    XRAM[48779] = 8'b0;
    XRAM[48780] = 8'b0;
    XRAM[48781] = 8'b0;
    XRAM[48782] = 8'b0;
    XRAM[48783] = 8'b0;
    XRAM[48784] = 8'b0;
    XRAM[48785] = 8'b0;
    XRAM[48786] = 8'b0;
    XRAM[48787] = 8'b0;
    XRAM[48788] = 8'b0;
    XRAM[48789] = 8'b0;
    XRAM[48790] = 8'b0;
    XRAM[48791] = 8'b0;
    XRAM[48792] = 8'b0;
    XRAM[48793] = 8'b0;
    XRAM[48794] = 8'b0;
    XRAM[48795] = 8'b0;
    XRAM[48796] = 8'b0;
    XRAM[48797] = 8'b0;
    XRAM[48798] = 8'b0;
    XRAM[48799] = 8'b0;
    XRAM[48800] = 8'b0;
    XRAM[48801] = 8'b0;
    XRAM[48802] = 8'b0;
    XRAM[48803] = 8'b0;
    XRAM[48804] = 8'b0;
    XRAM[48805] = 8'b0;
    XRAM[48806] = 8'b0;
    XRAM[48807] = 8'b0;
    XRAM[48808] = 8'b0;
    XRAM[48809] = 8'b0;
    XRAM[48810] = 8'b0;
    XRAM[48811] = 8'b0;
    XRAM[48812] = 8'b0;
    XRAM[48813] = 8'b0;
    XRAM[48814] = 8'b0;
    XRAM[48815] = 8'b0;
    XRAM[48816] = 8'b0;
    XRAM[48817] = 8'b0;
    XRAM[48818] = 8'b0;
    XRAM[48819] = 8'b0;
    XRAM[48820] = 8'b0;
    XRAM[48821] = 8'b0;
    XRAM[48822] = 8'b0;
    XRAM[48823] = 8'b0;
    XRAM[48824] = 8'b0;
    XRAM[48825] = 8'b0;
    XRAM[48826] = 8'b0;
    XRAM[48827] = 8'b0;
    XRAM[48828] = 8'b0;
    XRAM[48829] = 8'b0;
    XRAM[48830] = 8'b0;
    XRAM[48831] = 8'b0;
    XRAM[48832] = 8'b0;
    XRAM[48833] = 8'b0;
    XRAM[48834] = 8'b0;
    XRAM[48835] = 8'b0;
    XRAM[48836] = 8'b0;
    XRAM[48837] = 8'b0;
    XRAM[48838] = 8'b0;
    XRAM[48839] = 8'b0;
    XRAM[48840] = 8'b0;
    XRAM[48841] = 8'b0;
    XRAM[48842] = 8'b0;
    XRAM[48843] = 8'b0;
    XRAM[48844] = 8'b0;
    XRAM[48845] = 8'b0;
    XRAM[48846] = 8'b0;
    XRAM[48847] = 8'b0;
    XRAM[48848] = 8'b0;
    XRAM[48849] = 8'b0;
    XRAM[48850] = 8'b0;
    XRAM[48851] = 8'b0;
    XRAM[48852] = 8'b0;
    XRAM[48853] = 8'b0;
    XRAM[48854] = 8'b0;
    XRAM[48855] = 8'b0;
    XRAM[48856] = 8'b0;
    XRAM[48857] = 8'b0;
    XRAM[48858] = 8'b0;
    XRAM[48859] = 8'b0;
    XRAM[48860] = 8'b0;
    XRAM[48861] = 8'b0;
    XRAM[48862] = 8'b0;
    XRAM[48863] = 8'b0;
    XRAM[48864] = 8'b0;
    XRAM[48865] = 8'b0;
    XRAM[48866] = 8'b0;
    XRAM[48867] = 8'b0;
    XRAM[48868] = 8'b0;
    XRAM[48869] = 8'b0;
    XRAM[48870] = 8'b0;
    XRAM[48871] = 8'b0;
    XRAM[48872] = 8'b0;
    XRAM[48873] = 8'b0;
    XRAM[48874] = 8'b0;
    XRAM[48875] = 8'b0;
    XRAM[48876] = 8'b0;
    XRAM[48877] = 8'b0;
    XRAM[48878] = 8'b0;
    XRAM[48879] = 8'b0;
    XRAM[48880] = 8'b0;
    XRAM[48881] = 8'b0;
    XRAM[48882] = 8'b0;
    XRAM[48883] = 8'b0;
    XRAM[48884] = 8'b0;
    XRAM[48885] = 8'b0;
    XRAM[48886] = 8'b0;
    XRAM[48887] = 8'b0;
    XRAM[48888] = 8'b0;
    XRAM[48889] = 8'b0;
    XRAM[48890] = 8'b0;
    XRAM[48891] = 8'b0;
    XRAM[48892] = 8'b0;
    XRAM[48893] = 8'b0;
    XRAM[48894] = 8'b0;
    XRAM[48895] = 8'b0;
    XRAM[48896] = 8'b0;
    XRAM[48897] = 8'b0;
    XRAM[48898] = 8'b0;
    XRAM[48899] = 8'b0;
    XRAM[48900] = 8'b0;
    XRAM[48901] = 8'b0;
    XRAM[48902] = 8'b0;
    XRAM[48903] = 8'b0;
    XRAM[48904] = 8'b0;
    XRAM[48905] = 8'b0;
    XRAM[48906] = 8'b0;
    XRAM[48907] = 8'b0;
    XRAM[48908] = 8'b0;
    XRAM[48909] = 8'b0;
    XRAM[48910] = 8'b0;
    XRAM[48911] = 8'b0;
    XRAM[48912] = 8'b0;
    XRAM[48913] = 8'b0;
    XRAM[48914] = 8'b0;
    XRAM[48915] = 8'b0;
    XRAM[48916] = 8'b0;
    XRAM[48917] = 8'b0;
    XRAM[48918] = 8'b0;
    XRAM[48919] = 8'b0;
    XRAM[48920] = 8'b0;
    XRAM[48921] = 8'b0;
    XRAM[48922] = 8'b0;
    XRAM[48923] = 8'b0;
    XRAM[48924] = 8'b0;
    XRAM[48925] = 8'b0;
    XRAM[48926] = 8'b0;
    XRAM[48927] = 8'b0;
    XRAM[48928] = 8'b0;
    XRAM[48929] = 8'b0;
    XRAM[48930] = 8'b0;
    XRAM[48931] = 8'b0;
    XRAM[48932] = 8'b0;
    XRAM[48933] = 8'b0;
    XRAM[48934] = 8'b0;
    XRAM[48935] = 8'b0;
    XRAM[48936] = 8'b0;
    XRAM[48937] = 8'b0;
    XRAM[48938] = 8'b0;
    XRAM[48939] = 8'b0;
    XRAM[48940] = 8'b0;
    XRAM[48941] = 8'b0;
    XRAM[48942] = 8'b0;
    XRAM[48943] = 8'b0;
    XRAM[48944] = 8'b0;
    XRAM[48945] = 8'b0;
    XRAM[48946] = 8'b0;
    XRAM[48947] = 8'b0;
    XRAM[48948] = 8'b0;
    XRAM[48949] = 8'b0;
    XRAM[48950] = 8'b0;
    XRAM[48951] = 8'b0;
    XRAM[48952] = 8'b0;
    XRAM[48953] = 8'b0;
    XRAM[48954] = 8'b0;
    XRAM[48955] = 8'b0;
    XRAM[48956] = 8'b0;
    XRAM[48957] = 8'b0;
    XRAM[48958] = 8'b0;
    XRAM[48959] = 8'b0;
    XRAM[48960] = 8'b0;
    XRAM[48961] = 8'b0;
    XRAM[48962] = 8'b0;
    XRAM[48963] = 8'b0;
    XRAM[48964] = 8'b0;
    XRAM[48965] = 8'b0;
    XRAM[48966] = 8'b0;
    XRAM[48967] = 8'b0;
    XRAM[48968] = 8'b0;
    XRAM[48969] = 8'b0;
    XRAM[48970] = 8'b0;
    XRAM[48971] = 8'b0;
    XRAM[48972] = 8'b0;
    XRAM[48973] = 8'b0;
    XRAM[48974] = 8'b0;
    XRAM[48975] = 8'b0;
    XRAM[48976] = 8'b0;
    XRAM[48977] = 8'b0;
    XRAM[48978] = 8'b0;
    XRAM[48979] = 8'b0;
    XRAM[48980] = 8'b0;
    XRAM[48981] = 8'b0;
    XRAM[48982] = 8'b0;
    XRAM[48983] = 8'b0;
    XRAM[48984] = 8'b0;
    XRAM[48985] = 8'b0;
    XRAM[48986] = 8'b0;
    XRAM[48987] = 8'b0;
    XRAM[48988] = 8'b0;
    XRAM[48989] = 8'b0;
    XRAM[48990] = 8'b0;
    XRAM[48991] = 8'b0;
    XRAM[48992] = 8'b0;
    XRAM[48993] = 8'b0;
    XRAM[48994] = 8'b0;
    XRAM[48995] = 8'b0;
    XRAM[48996] = 8'b0;
    XRAM[48997] = 8'b0;
    XRAM[48998] = 8'b0;
    XRAM[48999] = 8'b0;
    XRAM[49000] = 8'b0;
    XRAM[49001] = 8'b0;
    XRAM[49002] = 8'b0;
    XRAM[49003] = 8'b0;
    XRAM[49004] = 8'b0;
    XRAM[49005] = 8'b0;
    XRAM[49006] = 8'b0;
    XRAM[49007] = 8'b0;
    XRAM[49008] = 8'b0;
    XRAM[49009] = 8'b0;
    XRAM[49010] = 8'b0;
    XRAM[49011] = 8'b0;
    XRAM[49012] = 8'b0;
    XRAM[49013] = 8'b0;
    XRAM[49014] = 8'b0;
    XRAM[49015] = 8'b0;
    XRAM[49016] = 8'b0;
    XRAM[49017] = 8'b0;
    XRAM[49018] = 8'b0;
    XRAM[49019] = 8'b0;
    XRAM[49020] = 8'b0;
    XRAM[49021] = 8'b0;
    XRAM[49022] = 8'b0;
    XRAM[49023] = 8'b0;
    XRAM[49024] = 8'b0;
    XRAM[49025] = 8'b0;
    XRAM[49026] = 8'b0;
    XRAM[49027] = 8'b0;
    XRAM[49028] = 8'b0;
    XRAM[49029] = 8'b0;
    XRAM[49030] = 8'b0;
    XRAM[49031] = 8'b0;
    XRAM[49032] = 8'b0;
    XRAM[49033] = 8'b0;
    XRAM[49034] = 8'b0;
    XRAM[49035] = 8'b0;
    XRAM[49036] = 8'b0;
    XRAM[49037] = 8'b0;
    XRAM[49038] = 8'b0;
    XRAM[49039] = 8'b0;
    XRAM[49040] = 8'b0;
    XRAM[49041] = 8'b0;
    XRAM[49042] = 8'b0;
    XRAM[49043] = 8'b0;
    XRAM[49044] = 8'b0;
    XRAM[49045] = 8'b0;
    XRAM[49046] = 8'b0;
    XRAM[49047] = 8'b0;
    XRAM[49048] = 8'b0;
    XRAM[49049] = 8'b0;
    XRAM[49050] = 8'b0;
    XRAM[49051] = 8'b0;
    XRAM[49052] = 8'b0;
    XRAM[49053] = 8'b0;
    XRAM[49054] = 8'b0;
    XRAM[49055] = 8'b0;
    XRAM[49056] = 8'b0;
    XRAM[49057] = 8'b0;
    XRAM[49058] = 8'b0;
    XRAM[49059] = 8'b0;
    XRAM[49060] = 8'b0;
    XRAM[49061] = 8'b0;
    XRAM[49062] = 8'b0;
    XRAM[49063] = 8'b0;
    XRAM[49064] = 8'b0;
    XRAM[49065] = 8'b0;
    XRAM[49066] = 8'b0;
    XRAM[49067] = 8'b0;
    XRAM[49068] = 8'b0;
    XRAM[49069] = 8'b0;
    XRAM[49070] = 8'b0;
    XRAM[49071] = 8'b0;
    XRAM[49072] = 8'b0;
    XRAM[49073] = 8'b0;
    XRAM[49074] = 8'b0;
    XRAM[49075] = 8'b0;
    XRAM[49076] = 8'b0;
    XRAM[49077] = 8'b0;
    XRAM[49078] = 8'b0;
    XRAM[49079] = 8'b0;
    XRAM[49080] = 8'b0;
    XRAM[49081] = 8'b0;
    XRAM[49082] = 8'b0;
    XRAM[49083] = 8'b0;
    XRAM[49084] = 8'b0;
    XRAM[49085] = 8'b0;
    XRAM[49086] = 8'b0;
    XRAM[49087] = 8'b0;
    XRAM[49088] = 8'b0;
    XRAM[49089] = 8'b0;
    XRAM[49090] = 8'b0;
    XRAM[49091] = 8'b0;
    XRAM[49092] = 8'b0;
    XRAM[49093] = 8'b0;
    XRAM[49094] = 8'b0;
    XRAM[49095] = 8'b0;
    XRAM[49096] = 8'b0;
    XRAM[49097] = 8'b0;
    XRAM[49098] = 8'b0;
    XRAM[49099] = 8'b0;
    XRAM[49100] = 8'b0;
    XRAM[49101] = 8'b0;
    XRAM[49102] = 8'b0;
    XRAM[49103] = 8'b0;
    XRAM[49104] = 8'b0;
    XRAM[49105] = 8'b0;
    XRAM[49106] = 8'b0;
    XRAM[49107] = 8'b0;
    XRAM[49108] = 8'b0;
    XRAM[49109] = 8'b0;
    XRAM[49110] = 8'b0;
    XRAM[49111] = 8'b0;
    XRAM[49112] = 8'b0;
    XRAM[49113] = 8'b0;
    XRAM[49114] = 8'b0;
    XRAM[49115] = 8'b0;
    XRAM[49116] = 8'b0;
    XRAM[49117] = 8'b0;
    XRAM[49118] = 8'b0;
    XRAM[49119] = 8'b0;
    XRAM[49120] = 8'b0;
    XRAM[49121] = 8'b0;
    XRAM[49122] = 8'b0;
    XRAM[49123] = 8'b0;
    XRAM[49124] = 8'b0;
    XRAM[49125] = 8'b0;
    XRAM[49126] = 8'b0;
    XRAM[49127] = 8'b0;
    XRAM[49128] = 8'b0;
    XRAM[49129] = 8'b0;
    XRAM[49130] = 8'b0;
    XRAM[49131] = 8'b0;
    XRAM[49132] = 8'b0;
    XRAM[49133] = 8'b0;
    XRAM[49134] = 8'b0;
    XRAM[49135] = 8'b0;
    XRAM[49136] = 8'b0;
    XRAM[49137] = 8'b0;
    XRAM[49138] = 8'b0;
    XRAM[49139] = 8'b0;
    XRAM[49140] = 8'b0;
    XRAM[49141] = 8'b0;
    XRAM[49142] = 8'b0;
    XRAM[49143] = 8'b0;
    XRAM[49144] = 8'b0;
    XRAM[49145] = 8'b0;
    XRAM[49146] = 8'b0;
    XRAM[49147] = 8'b0;
    XRAM[49148] = 8'b0;
    XRAM[49149] = 8'b0;
    XRAM[49150] = 8'b0;
    XRAM[49151] = 8'b0;
    XRAM[49152] = 8'b0;
    XRAM[49153] = 8'b0;
    XRAM[49154] = 8'b0;
    XRAM[49155] = 8'b0;
    XRAM[49156] = 8'b0;
    XRAM[49157] = 8'b0;
    XRAM[49158] = 8'b0;
    XRAM[49159] = 8'b0;
    XRAM[49160] = 8'b0;
    XRAM[49161] = 8'b0;
    XRAM[49162] = 8'b0;
    XRAM[49163] = 8'b0;
    XRAM[49164] = 8'b0;
    XRAM[49165] = 8'b0;
    XRAM[49166] = 8'b0;
    XRAM[49167] = 8'b0;
    XRAM[49168] = 8'b0;
    XRAM[49169] = 8'b0;
    XRAM[49170] = 8'b0;
    XRAM[49171] = 8'b0;
    XRAM[49172] = 8'b0;
    XRAM[49173] = 8'b0;
    XRAM[49174] = 8'b0;
    XRAM[49175] = 8'b0;
    XRAM[49176] = 8'b0;
    XRAM[49177] = 8'b0;
    XRAM[49178] = 8'b0;
    XRAM[49179] = 8'b0;
    XRAM[49180] = 8'b0;
    XRAM[49181] = 8'b0;
    XRAM[49182] = 8'b0;
    XRAM[49183] = 8'b0;
    XRAM[49184] = 8'b0;
    XRAM[49185] = 8'b0;
    XRAM[49186] = 8'b0;
    XRAM[49187] = 8'b0;
    XRAM[49188] = 8'b0;
    XRAM[49189] = 8'b0;
    XRAM[49190] = 8'b0;
    XRAM[49191] = 8'b0;
    XRAM[49192] = 8'b0;
    XRAM[49193] = 8'b0;
    XRAM[49194] = 8'b0;
    XRAM[49195] = 8'b0;
    XRAM[49196] = 8'b0;
    XRAM[49197] = 8'b0;
    XRAM[49198] = 8'b0;
    XRAM[49199] = 8'b0;
    XRAM[49200] = 8'b0;
    XRAM[49201] = 8'b0;
    XRAM[49202] = 8'b0;
    XRAM[49203] = 8'b0;
    XRAM[49204] = 8'b0;
    XRAM[49205] = 8'b0;
    XRAM[49206] = 8'b0;
    XRAM[49207] = 8'b0;
    XRAM[49208] = 8'b0;
    XRAM[49209] = 8'b0;
    XRAM[49210] = 8'b0;
    XRAM[49211] = 8'b0;
    XRAM[49212] = 8'b0;
    XRAM[49213] = 8'b0;
    XRAM[49214] = 8'b0;
    XRAM[49215] = 8'b0;
    XRAM[49216] = 8'b0;
    XRAM[49217] = 8'b0;
    XRAM[49218] = 8'b0;
    XRAM[49219] = 8'b0;
    XRAM[49220] = 8'b0;
    XRAM[49221] = 8'b0;
    XRAM[49222] = 8'b0;
    XRAM[49223] = 8'b0;
    XRAM[49224] = 8'b0;
    XRAM[49225] = 8'b0;
    XRAM[49226] = 8'b0;
    XRAM[49227] = 8'b0;
    XRAM[49228] = 8'b0;
    XRAM[49229] = 8'b0;
    XRAM[49230] = 8'b0;
    XRAM[49231] = 8'b0;
    XRAM[49232] = 8'b0;
    XRAM[49233] = 8'b0;
    XRAM[49234] = 8'b0;
    XRAM[49235] = 8'b0;
    XRAM[49236] = 8'b0;
    XRAM[49237] = 8'b0;
    XRAM[49238] = 8'b0;
    XRAM[49239] = 8'b0;
    XRAM[49240] = 8'b0;
    XRAM[49241] = 8'b0;
    XRAM[49242] = 8'b0;
    XRAM[49243] = 8'b0;
    XRAM[49244] = 8'b0;
    XRAM[49245] = 8'b0;
    XRAM[49246] = 8'b0;
    XRAM[49247] = 8'b0;
    XRAM[49248] = 8'b0;
    XRAM[49249] = 8'b0;
    XRAM[49250] = 8'b0;
    XRAM[49251] = 8'b0;
    XRAM[49252] = 8'b0;
    XRAM[49253] = 8'b0;
    XRAM[49254] = 8'b0;
    XRAM[49255] = 8'b0;
    XRAM[49256] = 8'b0;
    XRAM[49257] = 8'b0;
    XRAM[49258] = 8'b0;
    XRAM[49259] = 8'b0;
    XRAM[49260] = 8'b0;
    XRAM[49261] = 8'b0;
    XRAM[49262] = 8'b0;
    XRAM[49263] = 8'b0;
    XRAM[49264] = 8'b0;
    XRAM[49265] = 8'b0;
    XRAM[49266] = 8'b0;
    XRAM[49267] = 8'b0;
    XRAM[49268] = 8'b0;
    XRAM[49269] = 8'b0;
    XRAM[49270] = 8'b0;
    XRAM[49271] = 8'b0;
    XRAM[49272] = 8'b0;
    XRAM[49273] = 8'b0;
    XRAM[49274] = 8'b0;
    XRAM[49275] = 8'b0;
    XRAM[49276] = 8'b0;
    XRAM[49277] = 8'b0;
    XRAM[49278] = 8'b0;
    XRAM[49279] = 8'b0;
    XRAM[49280] = 8'b0;
    XRAM[49281] = 8'b0;
    XRAM[49282] = 8'b0;
    XRAM[49283] = 8'b0;
    XRAM[49284] = 8'b0;
    XRAM[49285] = 8'b0;
    XRAM[49286] = 8'b0;
    XRAM[49287] = 8'b0;
    XRAM[49288] = 8'b0;
    XRAM[49289] = 8'b0;
    XRAM[49290] = 8'b0;
    XRAM[49291] = 8'b0;
    XRAM[49292] = 8'b0;
    XRAM[49293] = 8'b0;
    XRAM[49294] = 8'b0;
    XRAM[49295] = 8'b0;
    XRAM[49296] = 8'b0;
    XRAM[49297] = 8'b0;
    XRAM[49298] = 8'b0;
    XRAM[49299] = 8'b0;
    XRAM[49300] = 8'b0;
    XRAM[49301] = 8'b0;
    XRAM[49302] = 8'b0;
    XRAM[49303] = 8'b0;
    XRAM[49304] = 8'b0;
    XRAM[49305] = 8'b0;
    XRAM[49306] = 8'b0;
    XRAM[49307] = 8'b0;
    XRAM[49308] = 8'b0;
    XRAM[49309] = 8'b0;
    XRAM[49310] = 8'b0;
    XRAM[49311] = 8'b0;
    XRAM[49312] = 8'b0;
    XRAM[49313] = 8'b0;
    XRAM[49314] = 8'b0;
    XRAM[49315] = 8'b0;
    XRAM[49316] = 8'b0;
    XRAM[49317] = 8'b0;
    XRAM[49318] = 8'b0;
    XRAM[49319] = 8'b0;
    XRAM[49320] = 8'b0;
    XRAM[49321] = 8'b0;
    XRAM[49322] = 8'b0;
    XRAM[49323] = 8'b0;
    XRAM[49324] = 8'b0;
    XRAM[49325] = 8'b0;
    XRAM[49326] = 8'b0;
    XRAM[49327] = 8'b0;
    XRAM[49328] = 8'b0;
    XRAM[49329] = 8'b0;
    XRAM[49330] = 8'b0;
    XRAM[49331] = 8'b0;
    XRAM[49332] = 8'b0;
    XRAM[49333] = 8'b0;
    XRAM[49334] = 8'b0;
    XRAM[49335] = 8'b0;
    XRAM[49336] = 8'b0;
    XRAM[49337] = 8'b0;
    XRAM[49338] = 8'b0;
    XRAM[49339] = 8'b0;
    XRAM[49340] = 8'b0;
    XRAM[49341] = 8'b0;
    XRAM[49342] = 8'b0;
    XRAM[49343] = 8'b0;
    XRAM[49344] = 8'b0;
    XRAM[49345] = 8'b0;
    XRAM[49346] = 8'b0;
    XRAM[49347] = 8'b0;
    XRAM[49348] = 8'b0;
    XRAM[49349] = 8'b0;
    XRAM[49350] = 8'b0;
    XRAM[49351] = 8'b0;
    XRAM[49352] = 8'b0;
    XRAM[49353] = 8'b0;
    XRAM[49354] = 8'b0;
    XRAM[49355] = 8'b0;
    XRAM[49356] = 8'b0;
    XRAM[49357] = 8'b0;
    XRAM[49358] = 8'b0;
    XRAM[49359] = 8'b0;
    XRAM[49360] = 8'b0;
    XRAM[49361] = 8'b0;
    XRAM[49362] = 8'b0;
    XRAM[49363] = 8'b0;
    XRAM[49364] = 8'b0;
    XRAM[49365] = 8'b0;
    XRAM[49366] = 8'b0;
    XRAM[49367] = 8'b0;
    XRAM[49368] = 8'b0;
    XRAM[49369] = 8'b0;
    XRAM[49370] = 8'b0;
    XRAM[49371] = 8'b0;
    XRAM[49372] = 8'b0;
    XRAM[49373] = 8'b0;
    XRAM[49374] = 8'b0;
    XRAM[49375] = 8'b0;
    XRAM[49376] = 8'b0;
    XRAM[49377] = 8'b0;
    XRAM[49378] = 8'b0;
    XRAM[49379] = 8'b0;
    XRAM[49380] = 8'b0;
    XRAM[49381] = 8'b0;
    XRAM[49382] = 8'b0;
    XRAM[49383] = 8'b0;
    XRAM[49384] = 8'b0;
    XRAM[49385] = 8'b0;
    XRAM[49386] = 8'b0;
    XRAM[49387] = 8'b0;
    XRAM[49388] = 8'b0;
    XRAM[49389] = 8'b0;
    XRAM[49390] = 8'b0;
    XRAM[49391] = 8'b0;
    XRAM[49392] = 8'b0;
    XRAM[49393] = 8'b0;
    XRAM[49394] = 8'b0;
    XRAM[49395] = 8'b0;
    XRAM[49396] = 8'b0;
    XRAM[49397] = 8'b0;
    XRAM[49398] = 8'b0;
    XRAM[49399] = 8'b0;
    XRAM[49400] = 8'b0;
    XRAM[49401] = 8'b0;
    XRAM[49402] = 8'b0;
    XRAM[49403] = 8'b0;
    XRAM[49404] = 8'b0;
    XRAM[49405] = 8'b0;
    XRAM[49406] = 8'b0;
    XRAM[49407] = 8'b0;
    XRAM[49408] = 8'b0;
    XRAM[49409] = 8'b0;
    XRAM[49410] = 8'b0;
    XRAM[49411] = 8'b0;
    XRAM[49412] = 8'b0;
    XRAM[49413] = 8'b0;
    XRAM[49414] = 8'b0;
    XRAM[49415] = 8'b0;
    XRAM[49416] = 8'b0;
    XRAM[49417] = 8'b0;
    XRAM[49418] = 8'b0;
    XRAM[49419] = 8'b0;
    XRAM[49420] = 8'b0;
    XRAM[49421] = 8'b0;
    XRAM[49422] = 8'b0;
    XRAM[49423] = 8'b0;
    XRAM[49424] = 8'b0;
    XRAM[49425] = 8'b0;
    XRAM[49426] = 8'b0;
    XRAM[49427] = 8'b0;
    XRAM[49428] = 8'b0;
    XRAM[49429] = 8'b0;
    XRAM[49430] = 8'b0;
    XRAM[49431] = 8'b0;
    XRAM[49432] = 8'b0;
    XRAM[49433] = 8'b0;
    XRAM[49434] = 8'b0;
    XRAM[49435] = 8'b0;
    XRAM[49436] = 8'b0;
    XRAM[49437] = 8'b0;
    XRAM[49438] = 8'b0;
    XRAM[49439] = 8'b0;
    XRAM[49440] = 8'b0;
    XRAM[49441] = 8'b0;
    XRAM[49442] = 8'b0;
    XRAM[49443] = 8'b0;
    XRAM[49444] = 8'b0;
    XRAM[49445] = 8'b0;
    XRAM[49446] = 8'b0;
    XRAM[49447] = 8'b0;
    XRAM[49448] = 8'b0;
    XRAM[49449] = 8'b0;
    XRAM[49450] = 8'b0;
    XRAM[49451] = 8'b0;
    XRAM[49452] = 8'b0;
    XRAM[49453] = 8'b0;
    XRAM[49454] = 8'b0;
    XRAM[49455] = 8'b0;
    XRAM[49456] = 8'b0;
    XRAM[49457] = 8'b0;
    XRAM[49458] = 8'b0;
    XRAM[49459] = 8'b0;
    XRAM[49460] = 8'b0;
    XRAM[49461] = 8'b0;
    XRAM[49462] = 8'b0;
    XRAM[49463] = 8'b0;
    XRAM[49464] = 8'b0;
    XRAM[49465] = 8'b0;
    XRAM[49466] = 8'b0;
    XRAM[49467] = 8'b0;
    XRAM[49468] = 8'b0;
    XRAM[49469] = 8'b0;
    XRAM[49470] = 8'b0;
    XRAM[49471] = 8'b0;
    XRAM[49472] = 8'b0;
    XRAM[49473] = 8'b0;
    XRAM[49474] = 8'b0;
    XRAM[49475] = 8'b0;
    XRAM[49476] = 8'b0;
    XRAM[49477] = 8'b0;
    XRAM[49478] = 8'b0;
    XRAM[49479] = 8'b0;
    XRAM[49480] = 8'b0;
    XRAM[49481] = 8'b0;
    XRAM[49482] = 8'b0;
    XRAM[49483] = 8'b0;
    XRAM[49484] = 8'b0;
    XRAM[49485] = 8'b0;
    XRAM[49486] = 8'b0;
    XRAM[49487] = 8'b0;
    XRAM[49488] = 8'b0;
    XRAM[49489] = 8'b0;
    XRAM[49490] = 8'b0;
    XRAM[49491] = 8'b0;
    XRAM[49492] = 8'b0;
    XRAM[49493] = 8'b0;
    XRAM[49494] = 8'b0;
    XRAM[49495] = 8'b0;
    XRAM[49496] = 8'b0;
    XRAM[49497] = 8'b0;
    XRAM[49498] = 8'b0;
    XRAM[49499] = 8'b0;
    XRAM[49500] = 8'b0;
    XRAM[49501] = 8'b0;
    XRAM[49502] = 8'b0;
    XRAM[49503] = 8'b0;
    XRAM[49504] = 8'b0;
    XRAM[49505] = 8'b0;
    XRAM[49506] = 8'b0;
    XRAM[49507] = 8'b0;
    XRAM[49508] = 8'b0;
    XRAM[49509] = 8'b0;
    XRAM[49510] = 8'b0;
    XRAM[49511] = 8'b0;
    XRAM[49512] = 8'b0;
    XRAM[49513] = 8'b0;
    XRAM[49514] = 8'b0;
    XRAM[49515] = 8'b0;
    XRAM[49516] = 8'b0;
    XRAM[49517] = 8'b0;
    XRAM[49518] = 8'b0;
    XRAM[49519] = 8'b0;
    XRAM[49520] = 8'b0;
    XRAM[49521] = 8'b0;
    XRAM[49522] = 8'b0;
    XRAM[49523] = 8'b0;
    XRAM[49524] = 8'b0;
    XRAM[49525] = 8'b0;
    XRAM[49526] = 8'b0;
    XRAM[49527] = 8'b0;
    XRAM[49528] = 8'b0;
    XRAM[49529] = 8'b0;
    XRAM[49530] = 8'b0;
    XRAM[49531] = 8'b0;
    XRAM[49532] = 8'b0;
    XRAM[49533] = 8'b0;
    XRAM[49534] = 8'b0;
    XRAM[49535] = 8'b0;
    XRAM[49536] = 8'b0;
    XRAM[49537] = 8'b0;
    XRAM[49538] = 8'b0;
    XRAM[49539] = 8'b0;
    XRAM[49540] = 8'b0;
    XRAM[49541] = 8'b0;
    XRAM[49542] = 8'b0;
    XRAM[49543] = 8'b0;
    XRAM[49544] = 8'b0;
    XRAM[49545] = 8'b0;
    XRAM[49546] = 8'b0;
    XRAM[49547] = 8'b0;
    XRAM[49548] = 8'b0;
    XRAM[49549] = 8'b0;
    XRAM[49550] = 8'b0;
    XRAM[49551] = 8'b0;
    XRAM[49552] = 8'b0;
    XRAM[49553] = 8'b0;
    XRAM[49554] = 8'b0;
    XRAM[49555] = 8'b0;
    XRAM[49556] = 8'b0;
    XRAM[49557] = 8'b0;
    XRAM[49558] = 8'b0;
    XRAM[49559] = 8'b0;
    XRAM[49560] = 8'b0;
    XRAM[49561] = 8'b0;
    XRAM[49562] = 8'b0;
    XRAM[49563] = 8'b0;
    XRAM[49564] = 8'b0;
    XRAM[49565] = 8'b0;
    XRAM[49566] = 8'b0;
    XRAM[49567] = 8'b0;
    XRAM[49568] = 8'b0;
    XRAM[49569] = 8'b0;
    XRAM[49570] = 8'b0;
    XRAM[49571] = 8'b0;
    XRAM[49572] = 8'b0;
    XRAM[49573] = 8'b0;
    XRAM[49574] = 8'b0;
    XRAM[49575] = 8'b0;
    XRAM[49576] = 8'b0;
    XRAM[49577] = 8'b0;
    XRAM[49578] = 8'b0;
    XRAM[49579] = 8'b0;
    XRAM[49580] = 8'b0;
    XRAM[49581] = 8'b0;
    XRAM[49582] = 8'b0;
    XRAM[49583] = 8'b0;
    XRAM[49584] = 8'b0;
    XRAM[49585] = 8'b0;
    XRAM[49586] = 8'b0;
    XRAM[49587] = 8'b0;
    XRAM[49588] = 8'b0;
    XRAM[49589] = 8'b0;
    XRAM[49590] = 8'b0;
    XRAM[49591] = 8'b0;
    XRAM[49592] = 8'b0;
    XRAM[49593] = 8'b0;
    XRAM[49594] = 8'b0;
    XRAM[49595] = 8'b0;
    XRAM[49596] = 8'b0;
    XRAM[49597] = 8'b0;
    XRAM[49598] = 8'b0;
    XRAM[49599] = 8'b0;
    XRAM[49600] = 8'b0;
    XRAM[49601] = 8'b0;
    XRAM[49602] = 8'b0;
    XRAM[49603] = 8'b0;
    XRAM[49604] = 8'b0;
    XRAM[49605] = 8'b0;
    XRAM[49606] = 8'b0;
    XRAM[49607] = 8'b0;
    XRAM[49608] = 8'b0;
    XRAM[49609] = 8'b0;
    XRAM[49610] = 8'b0;
    XRAM[49611] = 8'b0;
    XRAM[49612] = 8'b0;
    XRAM[49613] = 8'b0;
    XRAM[49614] = 8'b0;
    XRAM[49615] = 8'b0;
    XRAM[49616] = 8'b0;
    XRAM[49617] = 8'b0;
    XRAM[49618] = 8'b0;
    XRAM[49619] = 8'b0;
    XRAM[49620] = 8'b0;
    XRAM[49621] = 8'b0;
    XRAM[49622] = 8'b0;
    XRAM[49623] = 8'b0;
    XRAM[49624] = 8'b0;
    XRAM[49625] = 8'b0;
    XRAM[49626] = 8'b0;
    XRAM[49627] = 8'b0;
    XRAM[49628] = 8'b0;
    XRAM[49629] = 8'b0;
    XRAM[49630] = 8'b0;
    XRAM[49631] = 8'b0;
    XRAM[49632] = 8'b0;
    XRAM[49633] = 8'b0;
    XRAM[49634] = 8'b0;
    XRAM[49635] = 8'b0;
    XRAM[49636] = 8'b0;
    XRAM[49637] = 8'b0;
    XRAM[49638] = 8'b0;
    XRAM[49639] = 8'b0;
    XRAM[49640] = 8'b0;
    XRAM[49641] = 8'b0;
    XRAM[49642] = 8'b0;
    XRAM[49643] = 8'b0;
    XRAM[49644] = 8'b0;
    XRAM[49645] = 8'b0;
    XRAM[49646] = 8'b0;
    XRAM[49647] = 8'b0;
    XRAM[49648] = 8'b0;
    XRAM[49649] = 8'b0;
    XRAM[49650] = 8'b0;
    XRAM[49651] = 8'b0;
    XRAM[49652] = 8'b0;
    XRAM[49653] = 8'b0;
    XRAM[49654] = 8'b0;
    XRAM[49655] = 8'b0;
    XRAM[49656] = 8'b0;
    XRAM[49657] = 8'b0;
    XRAM[49658] = 8'b0;
    XRAM[49659] = 8'b0;
    XRAM[49660] = 8'b0;
    XRAM[49661] = 8'b0;
    XRAM[49662] = 8'b0;
    XRAM[49663] = 8'b0;
    XRAM[49664] = 8'b0;
    XRAM[49665] = 8'b0;
    XRAM[49666] = 8'b0;
    XRAM[49667] = 8'b0;
    XRAM[49668] = 8'b0;
    XRAM[49669] = 8'b0;
    XRAM[49670] = 8'b0;
    XRAM[49671] = 8'b0;
    XRAM[49672] = 8'b0;
    XRAM[49673] = 8'b0;
    XRAM[49674] = 8'b0;
    XRAM[49675] = 8'b0;
    XRAM[49676] = 8'b0;
    XRAM[49677] = 8'b0;
    XRAM[49678] = 8'b0;
    XRAM[49679] = 8'b0;
    XRAM[49680] = 8'b0;
    XRAM[49681] = 8'b0;
    XRAM[49682] = 8'b0;
    XRAM[49683] = 8'b0;
    XRAM[49684] = 8'b0;
    XRAM[49685] = 8'b0;
    XRAM[49686] = 8'b0;
    XRAM[49687] = 8'b0;
    XRAM[49688] = 8'b0;
    XRAM[49689] = 8'b0;
    XRAM[49690] = 8'b0;
    XRAM[49691] = 8'b0;
    XRAM[49692] = 8'b0;
    XRAM[49693] = 8'b0;
    XRAM[49694] = 8'b0;
    XRAM[49695] = 8'b0;
    XRAM[49696] = 8'b0;
    XRAM[49697] = 8'b0;
    XRAM[49698] = 8'b0;
    XRAM[49699] = 8'b0;
    XRAM[49700] = 8'b0;
    XRAM[49701] = 8'b0;
    XRAM[49702] = 8'b0;
    XRAM[49703] = 8'b0;
    XRAM[49704] = 8'b0;
    XRAM[49705] = 8'b0;
    XRAM[49706] = 8'b0;
    XRAM[49707] = 8'b0;
    XRAM[49708] = 8'b0;
    XRAM[49709] = 8'b0;
    XRAM[49710] = 8'b0;
    XRAM[49711] = 8'b0;
    XRAM[49712] = 8'b0;
    XRAM[49713] = 8'b0;
    XRAM[49714] = 8'b0;
    XRAM[49715] = 8'b0;
    XRAM[49716] = 8'b0;
    XRAM[49717] = 8'b0;
    XRAM[49718] = 8'b0;
    XRAM[49719] = 8'b0;
    XRAM[49720] = 8'b0;
    XRAM[49721] = 8'b0;
    XRAM[49722] = 8'b0;
    XRAM[49723] = 8'b0;
    XRAM[49724] = 8'b0;
    XRAM[49725] = 8'b0;
    XRAM[49726] = 8'b0;
    XRAM[49727] = 8'b0;
    XRAM[49728] = 8'b0;
    XRAM[49729] = 8'b0;
    XRAM[49730] = 8'b0;
    XRAM[49731] = 8'b0;
    XRAM[49732] = 8'b0;
    XRAM[49733] = 8'b0;
    XRAM[49734] = 8'b0;
    XRAM[49735] = 8'b0;
    XRAM[49736] = 8'b0;
    XRAM[49737] = 8'b0;
    XRAM[49738] = 8'b0;
    XRAM[49739] = 8'b0;
    XRAM[49740] = 8'b0;
    XRAM[49741] = 8'b0;
    XRAM[49742] = 8'b0;
    XRAM[49743] = 8'b0;
    XRAM[49744] = 8'b0;
    XRAM[49745] = 8'b0;
    XRAM[49746] = 8'b0;
    XRAM[49747] = 8'b0;
    XRAM[49748] = 8'b0;
    XRAM[49749] = 8'b0;
    XRAM[49750] = 8'b0;
    XRAM[49751] = 8'b0;
    XRAM[49752] = 8'b0;
    XRAM[49753] = 8'b0;
    XRAM[49754] = 8'b0;
    XRAM[49755] = 8'b0;
    XRAM[49756] = 8'b0;
    XRAM[49757] = 8'b0;
    XRAM[49758] = 8'b0;
    XRAM[49759] = 8'b0;
    XRAM[49760] = 8'b0;
    XRAM[49761] = 8'b0;
    XRAM[49762] = 8'b0;
    XRAM[49763] = 8'b0;
    XRAM[49764] = 8'b0;
    XRAM[49765] = 8'b0;
    XRAM[49766] = 8'b0;
    XRAM[49767] = 8'b0;
    XRAM[49768] = 8'b0;
    XRAM[49769] = 8'b0;
    XRAM[49770] = 8'b0;
    XRAM[49771] = 8'b0;
    XRAM[49772] = 8'b0;
    XRAM[49773] = 8'b0;
    XRAM[49774] = 8'b0;
    XRAM[49775] = 8'b0;
    XRAM[49776] = 8'b0;
    XRAM[49777] = 8'b0;
    XRAM[49778] = 8'b0;
    XRAM[49779] = 8'b0;
    XRAM[49780] = 8'b0;
    XRAM[49781] = 8'b0;
    XRAM[49782] = 8'b0;
    XRAM[49783] = 8'b0;
    XRAM[49784] = 8'b0;
    XRAM[49785] = 8'b0;
    XRAM[49786] = 8'b0;
    XRAM[49787] = 8'b0;
    XRAM[49788] = 8'b0;
    XRAM[49789] = 8'b0;
    XRAM[49790] = 8'b0;
    XRAM[49791] = 8'b0;
    XRAM[49792] = 8'b0;
    XRAM[49793] = 8'b0;
    XRAM[49794] = 8'b0;
    XRAM[49795] = 8'b0;
    XRAM[49796] = 8'b0;
    XRAM[49797] = 8'b0;
    XRAM[49798] = 8'b0;
    XRAM[49799] = 8'b0;
    XRAM[49800] = 8'b0;
    XRAM[49801] = 8'b0;
    XRAM[49802] = 8'b0;
    XRAM[49803] = 8'b0;
    XRAM[49804] = 8'b0;
    XRAM[49805] = 8'b0;
    XRAM[49806] = 8'b0;
    XRAM[49807] = 8'b0;
    XRAM[49808] = 8'b0;
    XRAM[49809] = 8'b0;
    XRAM[49810] = 8'b0;
    XRAM[49811] = 8'b0;
    XRAM[49812] = 8'b0;
    XRAM[49813] = 8'b0;
    XRAM[49814] = 8'b0;
    XRAM[49815] = 8'b0;
    XRAM[49816] = 8'b0;
    XRAM[49817] = 8'b0;
    XRAM[49818] = 8'b0;
    XRAM[49819] = 8'b0;
    XRAM[49820] = 8'b0;
    XRAM[49821] = 8'b0;
    XRAM[49822] = 8'b0;
    XRAM[49823] = 8'b0;
    XRAM[49824] = 8'b0;
    XRAM[49825] = 8'b0;
    XRAM[49826] = 8'b0;
    XRAM[49827] = 8'b0;
    XRAM[49828] = 8'b0;
    XRAM[49829] = 8'b0;
    XRAM[49830] = 8'b0;
    XRAM[49831] = 8'b0;
    XRAM[49832] = 8'b0;
    XRAM[49833] = 8'b0;
    XRAM[49834] = 8'b0;
    XRAM[49835] = 8'b0;
    XRAM[49836] = 8'b0;
    XRAM[49837] = 8'b0;
    XRAM[49838] = 8'b0;
    XRAM[49839] = 8'b0;
    XRAM[49840] = 8'b0;
    XRAM[49841] = 8'b0;
    XRAM[49842] = 8'b0;
    XRAM[49843] = 8'b0;
    XRAM[49844] = 8'b0;
    XRAM[49845] = 8'b0;
    XRAM[49846] = 8'b0;
    XRAM[49847] = 8'b0;
    XRAM[49848] = 8'b0;
    XRAM[49849] = 8'b0;
    XRAM[49850] = 8'b0;
    XRAM[49851] = 8'b0;
    XRAM[49852] = 8'b0;
    XRAM[49853] = 8'b0;
    XRAM[49854] = 8'b0;
    XRAM[49855] = 8'b0;
    XRAM[49856] = 8'b0;
    XRAM[49857] = 8'b0;
    XRAM[49858] = 8'b0;
    XRAM[49859] = 8'b0;
    XRAM[49860] = 8'b0;
    XRAM[49861] = 8'b0;
    XRAM[49862] = 8'b0;
    XRAM[49863] = 8'b0;
    XRAM[49864] = 8'b0;
    XRAM[49865] = 8'b0;
    XRAM[49866] = 8'b0;
    XRAM[49867] = 8'b0;
    XRAM[49868] = 8'b0;
    XRAM[49869] = 8'b0;
    XRAM[49870] = 8'b0;
    XRAM[49871] = 8'b0;
    XRAM[49872] = 8'b0;
    XRAM[49873] = 8'b0;
    XRAM[49874] = 8'b0;
    XRAM[49875] = 8'b0;
    XRAM[49876] = 8'b0;
    XRAM[49877] = 8'b0;
    XRAM[49878] = 8'b0;
    XRAM[49879] = 8'b0;
    XRAM[49880] = 8'b0;
    XRAM[49881] = 8'b0;
    XRAM[49882] = 8'b0;
    XRAM[49883] = 8'b0;
    XRAM[49884] = 8'b0;
    XRAM[49885] = 8'b0;
    XRAM[49886] = 8'b0;
    XRAM[49887] = 8'b0;
    XRAM[49888] = 8'b0;
    XRAM[49889] = 8'b0;
    XRAM[49890] = 8'b0;
    XRAM[49891] = 8'b0;
    XRAM[49892] = 8'b0;
    XRAM[49893] = 8'b0;
    XRAM[49894] = 8'b0;
    XRAM[49895] = 8'b0;
    XRAM[49896] = 8'b0;
    XRAM[49897] = 8'b0;
    XRAM[49898] = 8'b0;
    XRAM[49899] = 8'b0;
    XRAM[49900] = 8'b0;
    XRAM[49901] = 8'b0;
    XRAM[49902] = 8'b0;
    XRAM[49903] = 8'b0;
    XRAM[49904] = 8'b0;
    XRAM[49905] = 8'b0;
    XRAM[49906] = 8'b0;
    XRAM[49907] = 8'b0;
    XRAM[49908] = 8'b0;
    XRAM[49909] = 8'b0;
    XRAM[49910] = 8'b0;
    XRAM[49911] = 8'b0;
    XRAM[49912] = 8'b0;
    XRAM[49913] = 8'b0;
    XRAM[49914] = 8'b0;
    XRAM[49915] = 8'b0;
    XRAM[49916] = 8'b0;
    XRAM[49917] = 8'b0;
    XRAM[49918] = 8'b0;
    XRAM[49919] = 8'b0;
    XRAM[49920] = 8'b0;
    XRAM[49921] = 8'b0;
    XRAM[49922] = 8'b0;
    XRAM[49923] = 8'b0;
    XRAM[49924] = 8'b0;
    XRAM[49925] = 8'b0;
    XRAM[49926] = 8'b0;
    XRAM[49927] = 8'b0;
    XRAM[49928] = 8'b0;
    XRAM[49929] = 8'b0;
    XRAM[49930] = 8'b0;
    XRAM[49931] = 8'b0;
    XRAM[49932] = 8'b0;
    XRAM[49933] = 8'b0;
    XRAM[49934] = 8'b0;
    XRAM[49935] = 8'b0;
    XRAM[49936] = 8'b0;
    XRAM[49937] = 8'b0;
    XRAM[49938] = 8'b0;
    XRAM[49939] = 8'b0;
    XRAM[49940] = 8'b0;
    XRAM[49941] = 8'b0;
    XRAM[49942] = 8'b0;
    XRAM[49943] = 8'b0;
    XRAM[49944] = 8'b0;
    XRAM[49945] = 8'b0;
    XRAM[49946] = 8'b0;
    XRAM[49947] = 8'b0;
    XRAM[49948] = 8'b0;
    XRAM[49949] = 8'b0;
    XRAM[49950] = 8'b0;
    XRAM[49951] = 8'b0;
    XRAM[49952] = 8'b0;
    XRAM[49953] = 8'b0;
    XRAM[49954] = 8'b0;
    XRAM[49955] = 8'b0;
    XRAM[49956] = 8'b0;
    XRAM[49957] = 8'b0;
    XRAM[49958] = 8'b0;
    XRAM[49959] = 8'b0;
    XRAM[49960] = 8'b0;
    XRAM[49961] = 8'b0;
    XRAM[49962] = 8'b0;
    XRAM[49963] = 8'b0;
    XRAM[49964] = 8'b0;
    XRAM[49965] = 8'b0;
    XRAM[49966] = 8'b0;
    XRAM[49967] = 8'b0;
    XRAM[49968] = 8'b0;
    XRAM[49969] = 8'b0;
    XRAM[49970] = 8'b0;
    XRAM[49971] = 8'b0;
    XRAM[49972] = 8'b0;
    XRAM[49973] = 8'b0;
    XRAM[49974] = 8'b0;
    XRAM[49975] = 8'b0;
    XRAM[49976] = 8'b0;
    XRAM[49977] = 8'b0;
    XRAM[49978] = 8'b0;
    XRAM[49979] = 8'b0;
    XRAM[49980] = 8'b0;
    XRAM[49981] = 8'b0;
    XRAM[49982] = 8'b0;
    XRAM[49983] = 8'b0;
    XRAM[49984] = 8'b0;
    XRAM[49985] = 8'b0;
    XRAM[49986] = 8'b0;
    XRAM[49987] = 8'b0;
    XRAM[49988] = 8'b0;
    XRAM[49989] = 8'b0;
    XRAM[49990] = 8'b0;
    XRAM[49991] = 8'b0;
    XRAM[49992] = 8'b0;
    XRAM[49993] = 8'b0;
    XRAM[49994] = 8'b0;
    XRAM[49995] = 8'b0;
    XRAM[49996] = 8'b0;
    XRAM[49997] = 8'b0;
    XRAM[49998] = 8'b0;
    XRAM[49999] = 8'b0;
    XRAM[50000] = 8'b0;
    XRAM[50001] = 8'b0;
    XRAM[50002] = 8'b0;
    XRAM[50003] = 8'b0;
    XRAM[50004] = 8'b0;
    XRAM[50005] = 8'b0;
    XRAM[50006] = 8'b0;
    XRAM[50007] = 8'b0;
    XRAM[50008] = 8'b0;
    XRAM[50009] = 8'b0;
    XRAM[50010] = 8'b0;
    XRAM[50011] = 8'b0;
    XRAM[50012] = 8'b0;
    XRAM[50013] = 8'b0;
    XRAM[50014] = 8'b0;
    XRAM[50015] = 8'b0;
    XRAM[50016] = 8'b0;
    XRAM[50017] = 8'b0;
    XRAM[50018] = 8'b0;
    XRAM[50019] = 8'b0;
    XRAM[50020] = 8'b0;
    XRAM[50021] = 8'b0;
    XRAM[50022] = 8'b0;
    XRAM[50023] = 8'b0;
    XRAM[50024] = 8'b0;
    XRAM[50025] = 8'b0;
    XRAM[50026] = 8'b0;
    XRAM[50027] = 8'b0;
    XRAM[50028] = 8'b0;
    XRAM[50029] = 8'b0;
    XRAM[50030] = 8'b0;
    XRAM[50031] = 8'b0;
    XRAM[50032] = 8'b0;
    XRAM[50033] = 8'b0;
    XRAM[50034] = 8'b0;
    XRAM[50035] = 8'b0;
    XRAM[50036] = 8'b0;
    XRAM[50037] = 8'b0;
    XRAM[50038] = 8'b0;
    XRAM[50039] = 8'b0;
    XRAM[50040] = 8'b0;
    XRAM[50041] = 8'b0;
    XRAM[50042] = 8'b0;
    XRAM[50043] = 8'b0;
    XRAM[50044] = 8'b0;
    XRAM[50045] = 8'b0;
    XRAM[50046] = 8'b0;
    XRAM[50047] = 8'b0;
    XRAM[50048] = 8'b0;
    XRAM[50049] = 8'b0;
    XRAM[50050] = 8'b0;
    XRAM[50051] = 8'b0;
    XRAM[50052] = 8'b0;
    XRAM[50053] = 8'b0;
    XRAM[50054] = 8'b0;
    XRAM[50055] = 8'b0;
    XRAM[50056] = 8'b0;
    XRAM[50057] = 8'b0;
    XRAM[50058] = 8'b0;
    XRAM[50059] = 8'b0;
    XRAM[50060] = 8'b0;
    XRAM[50061] = 8'b0;
    XRAM[50062] = 8'b0;
    XRAM[50063] = 8'b0;
    XRAM[50064] = 8'b0;
    XRAM[50065] = 8'b0;
    XRAM[50066] = 8'b0;
    XRAM[50067] = 8'b0;
    XRAM[50068] = 8'b0;
    XRAM[50069] = 8'b0;
    XRAM[50070] = 8'b0;
    XRAM[50071] = 8'b0;
    XRAM[50072] = 8'b0;
    XRAM[50073] = 8'b0;
    XRAM[50074] = 8'b0;
    XRAM[50075] = 8'b0;
    XRAM[50076] = 8'b0;
    XRAM[50077] = 8'b0;
    XRAM[50078] = 8'b0;
    XRAM[50079] = 8'b0;
    XRAM[50080] = 8'b0;
    XRAM[50081] = 8'b0;
    XRAM[50082] = 8'b0;
    XRAM[50083] = 8'b0;
    XRAM[50084] = 8'b0;
    XRAM[50085] = 8'b0;
    XRAM[50086] = 8'b0;
    XRAM[50087] = 8'b0;
    XRAM[50088] = 8'b0;
    XRAM[50089] = 8'b0;
    XRAM[50090] = 8'b0;
    XRAM[50091] = 8'b0;
    XRAM[50092] = 8'b0;
    XRAM[50093] = 8'b0;
    XRAM[50094] = 8'b0;
    XRAM[50095] = 8'b0;
    XRAM[50096] = 8'b0;
    XRAM[50097] = 8'b0;
    XRAM[50098] = 8'b0;
    XRAM[50099] = 8'b0;
    XRAM[50100] = 8'b0;
    XRAM[50101] = 8'b0;
    XRAM[50102] = 8'b0;
    XRAM[50103] = 8'b0;
    XRAM[50104] = 8'b0;
    XRAM[50105] = 8'b0;
    XRAM[50106] = 8'b0;
    XRAM[50107] = 8'b0;
    XRAM[50108] = 8'b0;
    XRAM[50109] = 8'b0;
    XRAM[50110] = 8'b0;
    XRAM[50111] = 8'b0;
    XRAM[50112] = 8'b0;
    XRAM[50113] = 8'b0;
    XRAM[50114] = 8'b0;
    XRAM[50115] = 8'b0;
    XRAM[50116] = 8'b0;
    XRAM[50117] = 8'b0;
    XRAM[50118] = 8'b0;
    XRAM[50119] = 8'b0;
    XRAM[50120] = 8'b0;
    XRAM[50121] = 8'b0;
    XRAM[50122] = 8'b0;
    XRAM[50123] = 8'b0;
    XRAM[50124] = 8'b0;
    XRAM[50125] = 8'b0;
    XRAM[50126] = 8'b0;
    XRAM[50127] = 8'b0;
    XRAM[50128] = 8'b0;
    XRAM[50129] = 8'b0;
    XRAM[50130] = 8'b0;
    XRAM[50131] = 8'b0;
    XRAM[50132] = 8'b0;
    XRAM[50133] = 8'b0;
    XRAM[50134] = 8'b0;
    XRAM[50135] = 8'b0;
    XRAM[50136] = 8'b0;
    XRAM[50137] = 8'b0;
    XRAM[50138] = 8'b0;
    XRAM[50139] = 8'b0;
    XRAM[50140] = 8'b0;
    XRAM[50141] = 8'b0;
    XRAM[50142] = 8'b0;
    XRAM[50143] = 8'b0;
    XRAM[50144] = 8'b0;
    XRAM[50145] = 8'b0;
    XRAM[50146] = 8'b0;
    XRAM[50147] = 8'b0;
    XRAM[50148] = 8'b0;
    XRAM[50149] = 8'b0;
    XRAM[50150] = 8'b0;
    XRAM[50151] = 8'b0;
    XRAM[50152] = 8'b0;
    XRAM[50153] = 8'b0;
    XRAM[50154] = 8'b0;
    XRAM[50155] = 8'b0;
    XRAM[50156] = 8'b0;
    XRAM[50157] = 8'b0;
    XRAM[50158] = 8'b0;
    XRAM[50159] = 8'b0;
    XRAM[50160] = 8'b0;
    XRAM[50161] = 8'b0;
    XRAM[50162] = 8'b0;
    XRAM[50163] = 8'b0;
    XRAM[50164] = 8'b0;
    XRAM[50165] = 8'b0;
    XRAM[50166] = 8'b0;
    XRAM[50167] = 8'b0;
    XRAM[50168] = 8'b0;
    XRAM[50169] = 8'b0;
    XRAM[50170] = 8'b0;
    XRAM[50171] = 8'b0;
    XRAM[50172] = 8'b0;
    XRAM[50173] = 8'b0;
    XRAM[50174] = 8'b0;
    XRAM[50175] = 8'b0;
    XRAM[50176] = 8'b0;
    XRAM[50177] = 8'b0;
    XRAM[50178] = 8'b0;
    XRAM[50179] = 8'b0;
    XRAM[50180] = 8'b0;
    XRAM[50181] = 8'b0;
    XRAM[50182] = 8'b0;
    XRAM[50183] = 8'b0;
    XRAM[50184] = 8'b0;
    XRAM[50185] = 8'b0;
    XRAM[50186] = 8'b0;
    XRAM[50187] = 8'b0;
    XRAM[50188] = 8'b0;
    XRAM[50189] = 8'b0;
    XRAM[50190] = 8'b0;
    XRAM[50191] = 8'b0;
    XRAM[50192] = 8'b0;
    XRAM[50193] = 8'b0;
    XRAM[50194] = 8'b0;
    XRAM[50195] = 8'b0;
    XRAM[50196] = 8'b0;
    XRAM[50197] = 8'b0;
    XRAM[50198] = 8'b0;
    XRAM[50199] = 8'b0;
    XRAM[50200] = 8'b0;
    XRAM[50201] = 8'b0;
    XRAM[50202] = 8'b0;
    XRAM[50203] = 8'b0;
    XRAM[50204] = 8'b0;
    XRAM[50205] = 8'b0;
    XRAM[50206] = 8'b0;
    XRAM[50207] = 8'b0;
    XRAM[50208] = 8'b0;
    XRAM[50209] = 8'b0;
    XRAM[50210] = 8'b0;
    XRAM[50211] = 8'b0;
    XRAM[50212] = 8'b0;
    XRAM[50213] = 8'b0;
    XRAM[50214] = 8'b0;
    XRAM[50215] = 8'b0;
    XRAM[50216] = 8'b0;
    XRAM[50217] = 8'b0;
    XRAM[50218] = 8'b0;
    XRAM[50219] = 8'b0;
    XRAM[50220] = 8'b0;
    XRAM[50221] = 8'b0;
    XRAM[50222] = 8'b0;
    XRAM[50223] = 8'b0;
    XRAM[50224] = 8'b0;
    XRAM[50225] = 8'b0;
    XRAM[50226] = 8'b0;
    XRAM[50227] = 8'b0;
    XRAM[50228] = 8'b0;
    XRAM[50229] = 8'b0;
    XRAM[50230] = 8'b0;
    XRAM[50231] = 8'b0;
    XRAM[50232] = 8'b0;
    XRAM[50233] = 8'b0;
    XRAM[50234] = 8'b0;
    XRAM[50235] = 8'b0;
    XRAM[50236] = 8'b0;
    XRAM[50237] = 8'b0;
    XRAM[50238] = 8'b0;
    XRAM[50239] = 8'b0;
    XRAM[50240] = 8'b0;
    XRAM[50241] = 8'b0;
    XRAM[50242] = 8'b0;
    XRAM[50243] = 8'b0;
    XRAM[50244] = 8'b0;
    XRAM[50245] = 8'b0;
    XRAM[50246] = 8'b0;
    XRAM[50247] = 8'b0;
    XRAM[50248] = 8'b0;
    XRAM[50249] = 8'b0;
    XRAM[50250] = 8'b0;
    XRAM[50251] = 8'b0;
    XRAM[50252] = 8'b0;
    XRAM[50253] = 8'b0;
    XRAM[50254] = 8'b0;
    XRAM[50255] = 8'b0;
    XRAM[50256] = 8'b0;
    XRAM[50257] = 8'b0;
    XRAM[50258] = 8'b0;
    XRAM[50259] = 8'b0;
    XRAM[50260] = 8'b0;
    XRAM[50261] = 8'b0;
    XRAM[50262] = 8'b0;
    XRAM[50263] = 8'b0;
    XRAM[50264] = 8'b0;
    XRAM[50265] = 8'b0;
    XRAM[50266] = 8'b0;
    XRAM[50267] = 8'b0;
    XRAM[50268] = 8'b0;
    XRAM[50269] = 8'b0;
    XRAM[50270] = 8'b0;
    XRAM[50271] = 8'b0;
    XRAM[50272] = 8'b0;
    XRAM[50273] = 8'b0;
    XRAM[50274] = 8'b0;
    XRAM[50275] = 8'b0;
    XRAM[50276] = 8'b0;
    XRAM[50277] = 8'b0;
    XRAM[50278] = 8'b0;
    XRAM[50279] = 8'b0;
    XRAM[50280] = 8'b0;
    XRAM[50281] = 8'b0;
    XRAM[50282] = 8'b0;
    XRAM[50283] = 8'b0;
    XRAM[50284] = 8'b0;
    XRAM[50285] = 8'b0;
    XRAM[50286] = 8'b0;
    XRAM[50287] = 8'b0;
    XRAM[50288] = 8'b0;
    XRAM[50289] = 8'b0;
    XRAM[50290] = 8'b0;
    XRAM[50291] = 8'b0;
    XRAM[50292] = 8'b0;
    XRAM[50293] = 8'b0;
    XRAM[50294] = 8'b0;
    XRAM[50295] = 8'b0;
    XRAM[50296] = 8'b0;
    XRAM[50297] = 8'b0;
    XRAM[50298] = 8'b0;
    XRAM[50299] = 8'b0;
    XRAM[50300] = 8'b0;
    XRAM[50301] = 8'b0;
    XRAM[50302] = 8'b0;
    XRAM[50303] = 8'b0;
    XRAM[50304] = 8'b0;
    XRAM[50305] = 8'b0;
    XRAM[50306] = 8'b0;
    XRAM[50307] = 8'b0;
    XRAM[50308] = 8'b0;
    XRAM[50309] = 8'b0;
    XRAM[50310] = 8'b0;
    XRAM[50311] = 8'b0;
    XRAM[50312] = 8'b0;
    XRAM[50313] = 8'b0;
    XRAM[50314] = 8'b0;
    XRAM[50315] = 8'b0;
    XRAM[50316] = 8'b0;
    XRAM[50317] = 8'b0;
    XRAM[50318] = 8'b0;
    XRAM[50319] = 8'b0;
    XRAM[50320] = 8'b0;
    XRAM[50321] = 8'b0;
    XRAM[50322] = 8'b0;
    XRAM[50323] = 8'b0;
    XRAM[50324] = 8'b0;
    XRAM[50325] = 8'b0;
    XRAM[50326] = 8'b0;
    XRAM[50327] = 8'b0;
    XRAM[50328] = 8'b0;
    XRAM[50329] = 8'b0;
    XRAM[50330] = 8'b0;
    XRAM[50331] = 8'b0;
    XRAM[50332] = 8'b0;
    XRAM[50333] = 8'b0;
    XRAM[50334] = 8'b0;
    XRAM[50335] = 8'b0;
    XRAM[50336] = 8'b0;
    XRAM[50337] = 8'b0;
    XRAM[50338] = 8'b0;
    XRAM[50339] = 8'b0;
    XRAM[50340] = 8'b0;
    XRAM[50341] = 8'b0;
    XRAM[50342] = 8'b0;
    XRAM[50343] = 8'b0;
    XRAM[50344] = 8'b0;
    XRAM[50345] = 8'b0;
    XRAM[50346] = 8'b0;
    XRAM[50347] = 8'b0;
    XRAM[50348] = 8'b0;
    XRAM[50349] = 8'b0;
    XRAM[50350] = 8'b0;
    XRAM[50351] = 8'b0;
    XRAM[50352] = 8'b0;
    XRAM[50353] = 8'b0;
    XRAM[50354] = 8'b0;
    XRAM[50355] = 8'b0;
    XRAM[50356] = 8'b0;
    XRAM[50357] = 8'b0;
    XRAM[50358] = 8'b0;
    XRAM[50359] = 8'b0;
    XRAM[50360] = 8'b0;
    XRAM[50361] = 8'b0;
    XRAM[50362] = 8'b0;
    XRAM[50363] = 8'b0;
    XRAM[50364] = 8'b0;
    XRAM[50365] = 8'b0;
    XRAM[50366] = 8'b0;
    XRAM[50367] = 8'b0;
    XRAM[50368] = 8'b0;
    XRAM[50369] = 8'b0;
    XRAM[50370] = 8'b0;
    XRAM[50371] = 8'b0;
    XRAM[50372] = 8'b0;
    XRAM[50373] = 8'b0;
    XRAM[50374] = 8'b0;
    XRAM[50375] = 8'b0;
    XRAM[50376] = 8'b0;
    XRAM[50377] = 8'b0;
    XRAM[50378] = 8'b0;
    XRAM[50379] = 8'b0;
    XRAM[50380] = 8'b0;
    XRAM[50381] = 8'b0;
    XRAM[50382] = 8'b0;
    XRAM[50383] = 8'b0;
    XRAM[50384] = 8'b0;
    XRAM[50385] = 8'b0;
    XRAM[50386] = 8'b0;
    XRAM[50387] = 8'b0;
    XRAM[50388] = 8'b0;
    XRAM[50389] = 8'b0;
    XRAM[50390] = 8'b0;
    XRAM[50391] = 8'b0;
    XRAM[50392] = 8'b0;
    XRAM[50393] = 8'b0;
    XRAM[50394] = 8'b0;
    XRAM[50395] = 8'b0;
    XRAM[50396] = 8'b0;
    XRAM[50397] = 8'b0;
    XRAM[50398] = 8'b0;
    XRAM[50399] = 8'b0;
    XRAM[50400] = 8'b0;
    XRAM[50401] = 8'b0;
    XRAM[50402] = 8'b0;
    XRAM[50403] = 8'b0;
    XRAM[50404] = 8'b0;
    XRAM[50405] = 8'b0;
    XRAM[50406] = 8'b0;
    XRAM[50407] = 8'b0;
    XRAM[50408] = 8'b0;
    XRAM[50409] = 8'b0;
    XRAM[50410] = 8'b0;
    XRAM[50411] = 8'b0;
    XRAM[50412] = 8'b0;
    XRAM[50413] = 8'b0;
    XRAM[50414] = 8'b0;
    XRAM[50415] = 8'b0;
    XRAM[50416] = 8'b0;
    XRAM[50417] = 8'b0;
    XRAM[50418] = 8'b0;
    XRAM[50419] = 8'b0;
    XRAM[50420] = 8'b0;
    XRAM[50421] = 8'b0;
    XRAM[50422] = 8'b0;
    XRAM[50423] = 8'b0;
    XRAM[50424] = 8'b0;
    XRAM[50425] = 8'b0;
    XRAM[50426] = 8'b0;
    XRAM[50427] = 8'b0;
    XRAM[50428] = 8'b0;
    XRAM[50429] = 8'b0;
    XRAM[50430] = 8'b0;
    XRAM[50431] = 8'b0;
    XRAM[50432] = 8'b0;
    XRAM[50433] = 8'b0;
    XRAM[50434] = 8'b0;
    XRAM[50435] = 8'b0;
    XRAM[50436] = 8'b0;
    XRAM[50437] = 8'b0;
    XRAM[50438] = 8'b0;
    XRAM[50439] = 8'b0;
    XRAM[50440] = 8'b0;
    XRAM[50441] = 8'b0;
    XRAM[50442] = 8'b0;
    XRAM[50443] = 8'b0;
    XRAM[50444] = 8'b0;
    XRAM[50445] = 8'b0;
    XRAM[50446] = 8'b0;
    XRAM[50447] = 8'b0;
    XRAM[50448] = 8'b0;
    XRAM[50449] = 8'b0;
    XRAM[50450] = 8'b0;
    XRAM[50451] = 8'b0;
    XRAM[50452] = 8'b0;
    XRAM[50453] = 8'b0;
    XRAM[50454] = 8'b0;
    XRAM[50455] = 8'b0;
    XRAM[50456] = 8'b0;
    XRAM[50457] = 8'b0;
    XRAM[50458] = 8'b0;
    XRAM[50459] = 8'b0;
    XRAM[50460] = 8'b0;
    XRAM[50461] = 8'b0;
    XRAM[50462] = 8'b0;
    XRAM[50463] = 8'b0;
    XRAM[50464] = 8'b0;
    XRAM[50465] = 8'b0;
    XRAM[50466] = 8'b0;
    XRAM[50467] = 8'b0;
    XRAM[50468] = 8'b0;
    XRAM[50469] = 8'b0;
    XRAM[50470] = 8'b0;
    XRAM[50471] = 8'b0;
    XRAM[50472] = 8'b0;
    XRAM[50473] = 8'b0;
    XRAM[50474] = 8'b0;
    XRAM[50475] = 8'b0;
    XRAM[50476] = 8'b0;
    XRAM[50477] = 8'b0;
    XRAM[50478] = 8'b0;
    XRAM[50479] = 8'b0;
    XRAM[50480] = 8'b0;
    XRAM[50481] = 8'b0;
    XRAM[50482] = 8'b0;
    XRAM[50483] = 8'b0;
    XRAM[50484] = 8'b0;
    XRAM[50485] = 8'b0;
    XRAM[50486] = 8'b0;
    XRAM[50487] = 8'b0;
    XRAM[50488] = 8'b0;
    XRAM[50489] = 8'b0;
    XRAM[50490] = 8'b0;
    XRAM[50491] = 8'b0;
    XRAM[50492] = 8'b0;
    XRAM[50493] = 8'b0;
    XRAM[50494] = 8'b0;
    XRAM[50495] = 8'b0;
    XRAM[50496] = 8'b0;
    XRAM[50497] = 8'b0;
    XRAM[50498] = 8'b0;
    XRAM[50499] = 8'b0;
    XRAM[50500] = 8'b0;
    XRAM[50501] = 8'b0;
    XRAM[50502] = 8'b0;
    XRAM[50503] = 8'b0;
    XRAM[50504] = 8'b0;
    XRAM[50505] = 8'b0;
    XRAM[50506] = 8'b0;
    XRAM[50507] = 8'b0;
    XRAM[50508] = 8'b0;
    XRAM[50509] = 8'b0;
    XRAM[50510] = 8'b0;
    XRAM[50511] = 8'b0;
    XRAM[50512] = 8'b0;
    XRAM[50513] = 8'b0;
    XRAM[50514] = 8'b0;
    XRAM[50515] = 8'b0;
    XRAM[50516] = 8'b0;
    XRAM[50517] = 8'b0;
    XRAM[50518] = 8'b0;
    XRAM[50519] = 8'b0;
    XRAM[50520] = 8'b0;
    XRAM[50521] = 8'b0;
    XRAM[50522] = 8'b0;
    XRAM[50523] = 8'b0;
    XRAM[50524] = 8'b0;
    XRAM[50525] = 8'b0;
    XRAM[50526] = 8'b0;
    XRAM[50527] = 8'b0;
    XRAM[50528] = 8'b0;
    XRAM[50529] = 8'b0;
    XRAM[50530] = 8'b0;
    XRAM[50531] = 8'b0;
    XRAM[50532] = 8'b0;
    XRAM[50533] = 8'b0;
    XRAM[50534] = 8'b0;
    XRAM[50535] = 8'b0;
    XRAM[50536] = 8'b0;
    XRAM[50537] = 8'b0;
    XRAM[50538] = 8'b0;
    XRAM[50539] = 8'b0;
    XRAM[50540] = 8'b0;
    XRAM[50541] = 8'b0;
    XRAM[50542] = 8'b0;
    XRAM[50543] = 8'b0;
    XRAM[50544] = 8'b0;
    XRAM[50545] = 8'b0;
    XRAM[50546] = 8'b0;
    XRAM[50547] = 8'b0;
    XRAM[50548] = 8'b0;
    XRAM[50549] = 8'b0;
    XRAM[50550] = 8'b0;
    XRAM[50551] = 8'b0;
    XRAM[50552] = 8'b0;
    XRAM[50553] = 8'b0;
    XRAM[50554] = 8'b0;
    XRAM[50555] = 8'b0;
    XRAM[50556] = 8'b0;
    XRAM[50557] = 8'b0;
    XRAM[50558] = 8'b0;
    XRAM[50559] = 8'b0;
    XRAM[50560] = 8'b0;
    XRAM[50561] = 8'b0;
    XRAM[50562] = 8'b0;
    XRAM[50563] = 8'b0;
    XRAM[50564] = 8'b0;
    XRAM[50565] = 8'b0;
    XRAM[50566] = 8'b0;
    XRAM[50567] = 8'b0;
    XRAM[50568] = 8'b0;
    XRAM[50569] = 8'b0;
    XRAM[50570] = 8'b0;
    XRAM[50571] = 8'b0;
    XRAM[50572] = 8'b0;
    XRAM[50573] = 8'b0;
    XRAM[50574] = 8'b0;
    XRAM[50575] = 8'b0;
    XRAM[50576] = 8'b0;
    XRAM[50577] = 8'b0;
    XRAM[50578] = 8'b0;
    XRAM[50579] = 8'b0;
    XRAM[50580] = 8'b0;
    XRAM[50581] = 8'b0;
    XRAM[50582] = 8'b0;
    XRAM[50583] = 8'b0;
    XRAM[50584] = 8'b0;
    XRAM[50585] = 8'b0;
    XRAM[50586] = 8'b0;
    XRAM[50587] = 8'b0;
    XRAM[50588] = 8'b0;
    XRAM[50589] = 8'b0;
    XRAM[50590] = 8'b0;
    XRAM[50591] = 8'b0;
    XRAM[50592] = 8'b0;
    XRAM[50593] = 8'b0;
    XRAM[50594] = 8'b0;
    XRAM[50595] = 8'b0;
    XRAM[50596] = 8'b0;
    XRAM[50597] = 8'b0;
    XRAM[50598] = 8'b0;
    XRAM[50599] = 8'b0;
    XRAM[50600] = 8'b0;
    XRAM[50601] = 8'b0;
    XRAM[50602] = 8'b0;
    XRAM[50603] = 8'b0;
    XRAM[50604] = 8'b0;
    XRAM[50605] = 8'b0;
    XRAM[50606] = 8'b0;
    XRAM[50607] = 8'b0;
    XRAM[50608] = 8'b0;
    XRAM[50609] = 8'b0;
    XRAM[50610] = 8'b0;
    XRAM[50611] = 8'b0;
    XRAM[50612] = 8'b0;
    XRAM[50613] = 8'b0;
    XRAM[50614] = 8'b0;
    XRAM[50615] = 8'b0;
    XRAM[50616] = 8'b0;
    XRAM[50617] = 8'b0;
    XRAM[50618] = 8'b0;
    XRAM[50619] = 8'b0;
    XRAM[50620] = 8'b0;
    XRAM[50621] = 8'b0;
    XRAM[50622] = 8'b0;
    XRAM[50623] = 8'b0;
    XRAM[50624] = 8'b0;
    XRAM[50625] = 8'b0;
    XRAM[50626] = 8'b0;
    XRAM[50627] = 8'b0;
    XRAM[50628] = 8'b0;
    XRAM[50629] = 8'b0;
    XRAM[50630] = 8'b0;
    XRAM[50631] = 8'b0;
    XRAM[50632] = 8'b0;
    XRAM[50633] = 8'b0;
    XRAM[50634] = 8'b0;
    XRAM[50635] = 8'b0;
    XRAM[50636] = 8'b0;
    XRAM[50637] = 8'b0;
    XRAM[50638] = 8'b0;
    XRAM[50639] = 8'b0;
    XRAM[50640] = 8'b0;
    XRAM[50641] = 8'b0;
    XRAM[50642] = 8'b0;
    XRAM[50643] = 8'b0;
    XRAM[50644] = 8'b0;
    XRAM[50645] = 8'b0;
    XRAM[50646] = 8'b0;
    XRAM[50647] = 8'b0;
    XRAM[50648] = 8'b0;
    XRAM[50649] = 8'b0;
    XRAM[50650] = 8'b0;
    XRAM[50651] = 8'b0;
    XRAM[50652] = 8'b0;
    XRAM[50653] = 8'b0;
    XRAM[50654] = 8'b0;
    XRAM[50655] = 8'b0;
    XRAM[50656] = 8'b0;
    XRAM[50657] = 8'b0;
    XRAM[50658] = 8'b0;
    XRAM[50659] = 8'b0;
    XRAM[50660] = 8'b0;
    XRAM[50661] = 8'b0;
    XRAM[50662] = 8'b0;
    XRAM[50663] = 8'b0;
    XRAM[50664] = 8'b0;
    XRAM[50665] = 8'b0;
    XRAM[50666] = 8'b0;
    XRAM[50667] = 8'b0;
    XRAM[50668] = 8'b0;
    XRAM[50669] = 8'b0;
    XRAM[50670] = 8'b0;
    XRAM[50671] = 8'b0;
    XRAM[50672] = 8'b0;
    XRAM[50673] = 8'b0;
    XRAM[50674] = 8'b0;
    XRAM[50675] = 8'b0;
    XRAM[50676] = 8'b0;
    XRAM[50677] = 8'b0;
    XRAM[50678] = 8'b0;
    XRAM[50679] = 8'b0;
    XRAM[50680] = 8'b0;
    XRAM[50681] = 8'b0;
    XRAM[50682] = 8'b0;
    XRAM[50683] = 8'b0;
    XRAM[50684] = 8'b0;
    XRAM[50685] = 8'b0;
    XRAM[50686] = 8'b0;
    XRAM[50687] = 8'b0;
    XRAM[50688] = 8'b0;
    XRAM[50689] = 8'b0;
    XRAM[50690] = 8'b0;
    XRAM[50691] = 8'b0;
    XRAM[50692] = 8'b0;
    XRAM[50693] = 8'b0;
    XRAM[50694] = 8'b0;
    XRAM[50695] = 8'b0;
    XRAM[50696] = 8'b0;
    XRAM[50697] = 8'b0;
    XRAM[50698] = 8'b0;
    XRAM[50699] = 8'b0;
    XRAM[50700] = 8'b0;
    XRAM[50701] = 8'b0;
    XRAM[50702] = 8'b0;
    XRAM[50703] = 8'b0;
    XRAM[50704] = 8'b0;
    XRAM[50705] = 8'b0;
    XRAM[50706] = 8'b0;
    XRAM[50707] = 8'b0;
    XRAM[50708] = 8'b0;
    XRAM[50709] = 8'b0;
    XRAM[50710] = 8'b0;
    XRAM[50711] = 8'b0;
    XRAM[50712] = 8'b0;
    XRAM[50713] = 8'b0;
    XRAM[50714] = 8'b0;
    XRAM[50715] = 8'b0;
    XRAM[50716] = 8'b0;
    XRAM[50717] = 8'b0;
    XRAM[50718] = 8'b0;
    XRAM[50719] = 8'b0;
    XRAM[50720] = 8'b0;
    XRAM[50721] = 8'b0;
    XRAM[50722] = 8'b0;
    XRAM[50723] = 8'b0;
    XRAM[50724] = 8'b0;
    XRAM[50725] = 8'b0;
    XRAM[50726] = 8'b0;
    XRAM[50727] = 8'b0;
    XRAM[50728] = 8'b0;
    XRAM[50729] = 8'b0;
    XRAM[50730] = 8'b0;
    XRAM[50731] = 8'b0;
    XRAM[50732] = 8'b0;
    XRAM[50733] = 8'b0;
    XRAM[50734] = 8'b0;
    XRAM[50735] = 8'b0;
    XRAM[50736] = 8'b0;
    XRAM[50737] = 8'b0;
    XRAM[50738] = 8'b0;
    XRAM[50739] = 8'b0;
    XRAM[50740] = 8'b0;
    XRAM[50741] = 8'b0;
    XRAM[50742] = 8'b0;
    XRAM[50743] = 8'b0;
    XRAM[50744] = 8'b0;
    XRAM[50745] = 8'b0;
    XRAM[50746] = 8'b0;
    XRAM[50747] = 8'b0;
    XRAM[50748] = 8'b0;
    XRAM[50749] = 8'b0;
    XRAM[50750] = 8'b0;
    XRAM[50751] = 8'b0;
    XRAM[50752] = 8'b0;
    XRAM[50753] = 8'b0;
    XRAM[50754] = 8'b0;
    XRAM[50755] = 8'b0;
    XRAM[50756] = 8'b0;
    XRAM[50757] = 8'b0;
    XRAM[50758] = 8'b0;
    XRAM[50759] = 8'b0;
    XRAM[50760] = 8'b0;
    XRAM[50761] = 8'b0;
    XRAM[50762] = 8'b0;
    XRAM[50763] = 8'b0;
    XRAM[50764] = 8'b0;
    XRAM[50765] = 8'b0;
    XRAM[50766] = 8'b0;
    XRAM[50767] = 8'b0;
    XRAM[50768] = 8'b0;
    XRAM[50769] = 8'b0;
    XRAM[50770] = 8'b0;
    XRAM[50771] = 8'b0;
    XRAM[50772] = 8'b0;
    XRAM[50773] = 8'b0;
    XRAM[50774] = 8'b0;
    XRAM[50775] = 8'b0;
    XRAM[50776] = 8'b0;
    XRAM[50777] = 8'b0;
    XRAM[50778] = 8'b0;
    XRAM[50779] = 8'b0;
    XRAM[50780] = 8'b0;
    XRAM[50781] = 8'b0;
    XRAM[50782] = 8'b0;
    XRAM[50783] = 8'b0;
    XRAM[50784] = 8'b0;
    XRAM[50785] = 8'b0;
    XRAM[50786] = 8'b0;
    XRAM[50787] = 8'b0;
    XRAM[50788] = 8'b0;
    XRAM[50789] = 8'b0;
    XRAM[50790] = 8'b0;
    XRAM[50791] = 8'b0;
    XRAM[50792] = 8'b0;
    XRAM[50793] = 8'b0;
    XRAM[50794] = 8'b0;
    XRAM[50795] = 8'b0;
    XRAM[50796] = 8'b0;
    XRAM[50797] = 8'b0;
    XRAM[50798] = 8'b0;
    XRAM[50799] = 8'b0;
    XRAM[50800] = 8'b0;
    XRAM[50801] = 8'b0;
    XRAM[50802] = 8'b0;
    XRAM[50803] = 8'b0;
    XRAM[50804] = 8'b0;
    XRAM[50805] = 8'b0;
    XRAM[50806] = 8'b0;
    XRAM[50807] = 8'b0;
    XRAM[50808] = 8'b0;
    XRAM[50809] = 8'b0;
    XRAM[50810] = 8'b0;
    XRAM[50811] = 8'b0;
    XRAM[50812] = 8'b0;
    XRAM[50813] = 8'b0;
    XRAM[50814] = 8'b0;
    XRAM[50815] = 8'b0;
    XRAM[50816] = 8'b0;
    XRAM[50817] = 8'b0;
    XRAM[50818] = 8'b0;
    XRAM[50819] = 8'b0;
    XRAM[50820] = 8'b0;
    XRAM[50821] = 8'b0;
    XRAM[50822] = 8'b0;
    XRAM[50823] = 8'b0;
    XRAM[50824] = 8'b0;
    XRAM[50825] = 8'b0;
    XRAM[50826] = 8'b0;
    XRAM[50827] = 8'b0;
    XRAM[50828] = 8'b0;
    XRAM[50829] = 8'b0;
    XRAM[50830] = 8'b0;
    XRAM[50831] = 8'b0;
    XRAM[50832] = 8'b0;
    XRAM[50833] = 8'b0;
    XRAM[50834] = 8'b0;
    XRAM[50835] = 8'b0;
    XRAM[50836] = 8'b0;
    XRAM[50837] = 8'b0;
    XRAM[50838] = 8'b0;
    XRAM[50839] = 8'b0;
    XRAM[50840] = 8'b0;
    XRAM[50841] = 8'b0;
    XRAM[50842] = 8'b0;
    XRAM[50843] = 8'b0;
    XRAM[50844] = 8'b0;
    XRAM[50845] = 8'b0;
    XRAM[50846] = 8'b0;
    XRAM[50847] = 8'b0;
    XRAM[50848] = 8'b0;
    XRAM[50849] = 8'b0;
    XRAM[50850] = 8'b0;
    XRAM[50851] = 8'b0;
    XRAM[50852] = 8'b0;
    XRAM[50853] = 8'b0;
    XRAM[50854] = 8'b0;
    XRAM[50855] = 8'b0;
    XRAM[50856] = 8'b0;
    XRAM[50857] = 8'b0;
    XRAM[50858] = 8'b0;
    XRAM[50859] = 8'b0;
    XRAM[50860] = 8'b0;
    XRAM[50861] = 8'b0;
    XRAM[50862] = 8'b0;
    XRAM[50863] = 8'b0;
    XRAM[50864] = 8'b0;
    XRAM[50865] = 8'b0;
    XRAM[50866] = 8'b0;
    XRAM[50867] = 8'b0;
    XRAM[50868] = 8'b0;
    XRAM[50869] = 8'b0;
    XRAM[50870] = 8'b0;
    XRAM[50871] = 8'b0;
    XRAM[50872] = 8'b0;
    XRAM[50873] = 8'b0;
    XRAM[50874] = 8'b0;
    XRAM[50875] = 8'b0;
    XRAM[50876] = 8'b0;
    XRAM[50877] = 8'b0;
    XRAM[50878] = 8'b0;
    XRAM[50879] = 8'b0;
    XRAM[50880] = 8'b0;
    XRAM[50881] = 8'b0;
    XRAM[50882] = 8'b0;
    XRAM[50883] = 8'b0;
    XRAM[50884] = 8'b0;
    XRAM[50885] = 8'b0;
    XRAM[50886] = 8'b0;
    XRAM[50887] = 8'b0;
    XRAM[50888] = 8'b0;
    XRAM[50889] = 8'b0;
    XRAM[50890] = 8'b0;
    XRAM[50891] = 8'b0;
    XRAM[50892] = 8'b0;
    XRAM[50893] = 8'b0;
    XRAM[50894] = 8'b0;
    XRAM[50895] = 8'b0;
    XRAM[50896] = 8'b0;
    XRAM[50897] = 8'b0;
    XRAM[50898] = 8'b0;
    XRAM[50899] = 8'b0;
    XRAM[50900] = 8'b0;
    XRAM[50901] = 8'b0;
    XRAM[50902] = 8'b0;
    XRAM[50903] = 8'b0;
    XRAM[50904] = 8'b0;
    XRAM[50905] = 8'b0;
    XRAM[50906] = 8'b0;
    XRAM[50907] = 8'b0;
    XRAM[50908] = 8'b0;
    XRAM[50909] = 8'b0;
    XRAM[50910] = 8'b0;
    XRAM[50911] = 8'b0;
    XRAM[50912] = 8'b0;
    XRAM[50913] = 8'b0;
    XRAM[50914] = 8'b0;
    XRAM[50915] = 8'b0;
    XRAM[50916] = 8'b0;
    XRAM[50917] = 8'b0;
    XRAM[50918] = 8'b0;
    XRAM[50919] = 8'b0;
    XRAM[50920] = 8'b0;
    XRAM[50921] = 8'b0;
    XRAM[50922] = 8'b0;
    XRAM[50923] = 8'b0;
    XRAM[50924] = 8'b0;
    XRAM[50925] = 8'b0;
    XRAM[50926] = 8'b0;
    XRAM[50927] = 8'b0;
    XRAM[50928] = 8'b0;
    XRAM[50929] = 8'b0;
    XRAM[50930] = 8'b0;
    XRAM[50931] = 8'b0;
    XRAM[50932] = 8'b0;
    XRAM[50933] = 8'b0;
    XRAM[50934] = 8'b0;
    XRAM[50935] = 8'b0;
    XRAM[50936] = 8'b0;
    XRAM[50937] = 8'b0;
    XRAM[50938] = 8'b0;
    XRAM[50939] = 8'b0;
    XRAM[50940] = 8'b0;
    XRAM[50941] = 8'b0;
    XRAM[50942] = 8'b0;
    XRAM[50943] = 8'b0;
    XRAM[50944] = 8'b0;
    XRAM[50945] = 8'b0;
    XRAM[50946] = 8'b0;
    XRAM[50947] = 8'b0;
    XRAM[50948] = 8'b0;
    XRAM[50949] = 8'b0;
    XRAM[50950] = 8'b0;
    XRAM[50951] = 8'b0;
    XRAM[50952] = 8'b0;
    XRAM[50953] = 8'b0;
    XRAM[50954] = 8'b0;
    XRAM[50955] = 8'b0;
    XRAM[50956] = 8'b0;
    XRAM[50957] = 8'b0;
    XRAM[50958] = 8'b0;
    XRAM[50959] = 8'b0;
    XRAM[50960] = 8'b0;
    XRAM[50961] = 8'b0;
    XRAM[50962] = 8'b0;
    XRAM[50963] = 8'b0;
    XRAM[50964] = 8'b0;
    XRAM[50965] = 8'b0;
    XRAM[50966] = 8'b0;
    XRAM[50967] = 8'b0;
    XRAM[50968] = 8'b0;
    XRAM[50969] = 8'b0;
    XRAM[50970] = 8'b0;
    XRAM[50971] = 8'b0;
    XRAM[50972] = 8'b0;
    XRAM[50973] = 8'b0;
    XRAM[50974] = 8'b0;
    XRAM[50975] = 8'b0;
    XRAM[50976] = 8'b0;
    XRAM[50977] = 8'b0;
    XRAM[50978] = 8'b0;
    XRAM[50979] = 8'b0;
    XRAM[50980] = 8'b0;
    XRAM[50981] = 8'b0;
    XRAM[50982] = 8'b0;
    XRAM[50983] = 8'b0;
    XRAM[50984] = 8'b0;
    XRAM[50985] = 8'b0;
    XRAM[50986] = 8'b0;
    XRAM[50987] = 8'b0;
    XRAM[50988] = 8'b0;
    XRAM[50989] = 8'b0;
    XRAM[50990] = 8'b0;
    XRAM[50991] = 8'b0;
    XRAM[50992] = 8'b0;
    XRAM[50993] = 8'b0;
    XRAM[50994] = 8'b0;
    XRAM[50995] = 8'b0;
    XRAM[50996] = 8'b0;
    XRAM[50997] = 8'b0;
    XRAM[50998] = 8'b0;
    XRAM[50999] = 8'b0;
    XRAM[51000] = 8'b0;
    XRAM[51001] = 8'b0;
    XRAM[51002] = 8'b0;
    XRAM[51003] = 8'b0;
    XRAM[51004] = 8'b0;
    XRAM[51005] = 8'b0;
    XRAM[51006] = 8'b0;
    XRAM[51007] = 8'b0;
    XRAM[51008] = 8'b0;
    XRAM[51009] = 8'b0;
    XRAM[51010] = 8'b0;
    XRAM[51011] = 8'b0;
    XRAM[51012] = 8'b0;
    XRAM[51013] = 8'b0;
    XRAM[51014] = 8'b0;
    XRAM[51015] = 8'b0;
    XRAM[51016] = 8'b0;
    XRAM[51017] = 8'b0;
    XRAM[51018] = 8'b0;
    XRAM[51019] = 8'b0;
    XRAM[51020] = 8'b0;
    XRAM[51021] = 8'b0;
    XRAM[51022] = 8'b0;
    XRAM[51023] = 8'b0;
    XRAM[51024] = 8'b0;
    XRAM[51025] = 8'b0;
    XRAM[51026] = 8'b0;
    XRAM[51027] = 8'b0;
    XRAM[51028] = 8'b0;
    XRAM[51029] = 8'b0;
    XRAM[51030] = 8'b0;
    XRAM[51031] = 8'b0;
    XRAM[51032] = 8'b0;
    XRAM[51033] = 8'b0;
    XRAM[51034] = 8'b0;
    XRAM[51035] = 8'b0;
    XRAM[51036] = 8'b0;
    XRAM[51037] = 8'b0;
    XRAM[51038] = 8'b0;
    XRAM[51039] = 8'b0;
    XRAM[51040] = 8'b0;
    XRAM[51041] = 8'b0;
    XRAM[51042] = 8'b0;
    XRAM[51043] = 8'b0;
    XRAM[51044] = 8'b0;
    XRAM[51045] = 8'b0;
    XRAM[51046] = 8'b0;
    XRAM[51047] = 8'b0;
    XRAM[51048] = 8'b0;
    XRAM[51049] = 8'b0;
    XRAM[51050] = 8'b0;
    XRAM[51051] = 8'b0;
    XRAM[51052] = 8'b0;
    XRAM[51053] = 8'b0;
    XRAM[51054] = 8'b0;
    XRAM[51055] = 8'b0;
    XRAM[51056] = 8'b0;
    XRAM[51057] = 8'b0;
    XRAM[51058] = 8'b0;
    XRAM[51059] = 8'b0;
    XRAM[51060] = 8'b0;
    XRAM[51061] = 8'b0;
    XRAM[51062] = 8'b0;
    XRAM[51063] = 8'b0;
    XRAM[51064] = 8'b0;
    XRAM[51065] = 8'b0;
    XRAM[51066] = 8'b0;
    XRAM[51067] = 8'b0;
    XRAM[51068] = 8'b0;
    XRAM[51069] = 8'b0;
    XRAM[51070] = 8'b0;
    XRAM[51071] = 8'b0;
    XRAM[51072] = 8'b0;
    XRAM[51073] = 8'b0;
    XRAM[51074] = 8'b0;
    XRAM[51075] = 8'b0;
    XRAM[51076] = 8'b0;
    XRAM[51077] = 8'b0;
    XRAM[51078] = 8'b0;
    XRAM[51079] = 8'b0;
    XRAM[51080] = 8'b0;
    XRAM[51081] = 8'b0;
    XRAM[51082] = 8'b0;
    XRAM[51083] = 8'b0;
    XRAM[51084] = 8'b0;
    XRAM[51085] = 8'b0;
    XRAM[51086] = 8'b0;
    XRAM[51087] = 8'b0;
    XRAM[51088] = 8'b0;
    XRAM[51089] = 8'b0;
    XRAM[51090] = 8'b0;
    XRAM[51091] = 8'b0;
    XRAM[51092] = 8'b0;
    XRAM[51093] = 8'b0;
    XRAM[51094] = 8'b0;
    XRAM[51095] = 8'b0;
    XRAM[51096] = 8'b0;
    XRAM[51097] = 8'b0;
    XRAM[51098] = 8'b0;
    XRAM[51099] = 8'b0;
    XRAM[51100] = 8'b0;
    XRAM[51101] = 8'b0;
    XRAM[51102] = 8'b0;
    XRAM[51103] = 8'b0;
    XRAM[51104] = 8'b0;
    XRAM[51105] = 8'b0;
    XRAM[51106] = 8'b0;
    XRAM[51107] = 8'b0;
    XRAM[51108] = 8'b0;
    XRAM[51109] = 8'b0;
    XRAM[51110] = 8'b0;
    XRAM[51111] = 8'b0;
    XRAM[51112] = 8'b0;
    XRAM[51113] = 8'b0;
    XRAM[51114] = 8'b0;
    XRAM[51115] = 8'b0;
    XRAM[51116] = 8'b0;
    XRAM[51117] = 8'b0;
    XRAM[51118] = 8'b0;
    XRAM[51119] = 8'b0;
    XRAM[51120] = 8'b0;
    XRAM[51121] = 8'b0;
    XRAM[51122] = 8'b0;
    XRAM[51123] = 8'b0;
    XRAM[51124] = 8'b0;
    XRAM[51125] = 8'b0;
    XRAM[51126] = 8'b0;
    XRAM[51127] = 8'b0;
    XRAM[51128] = 8'b0;
    XRAM[51129] = 8'b0;
    XRAM[51130] = 8'b0;
    XRAM[51131] = 8'b0;
    XRAM[51132] = 8'b0;
    XRAM[51133] = 8'b0;
    XRAM[51134] = 8'b0;
    XRAM[51135] = 8'b0;
    XRAM[51136] = 8'b0;
    XRAM[51137] = 8'b0;
    XRAM[51138] = 8'b0;
    XRAM[51139] = 8'b0;
    XRAM[51140] = 8'b0;
    XRAM[51141] = 8'b0;
    XRAM[51142] = 8'b0;
    XRAM[51143] = 8'b0;
    XRAM[51144] = 8'b0;
    XRAM[51145] = 8'b0;
    XRAM[51146] = 8'b0;
    XRAM[51147] = 8'b0;
    XRAM[51148] = 8'b0;
    XRAM[51149] = 8'b0;
    XRAM[51150] = 8'b0;
    XRAM[51151] = 8'b0;
    XRAM[51152] = 8'b0;
    XRAM[51153] = 8'b0;
    XRAM[51154] = 8'b0;
    XRAM[51155] = 8'b0;
    XRAM[51156] = 8'b0;
    XRAM[51157] = 8'b0;
    XRAM[51158] = 8'b0;
    XRAM[51159] = 8'b0;
    XRAM[51160] = 8'b0;
    XRAM[51161] = 8'b0;
    XRAM[51162] = 8'b0;
    XRAM[51163] = 8'b0;
    XRAM[51164] = 8'b0;
    XRAM[51165] = 8'b0;
    XRAM[51166] = 8'b0;
    XRAM[51167] = 8'b0;
    XRAM[51168] = 8'b0;
    XRAM[51169] = 8'b0;
    XRAM[51170] = 8'b0;
    XRAM[51171] = 8'b0;
    XRAM[51172] = 8'b0;
    XRAM[51173] = 8'b0;
    XRAM[51174] = 8'b0;
    XRAM[51175] = 8'b0;
    XRAM[51176] = 8'b0;
    XRAM[51177] = 8'b0;
    XRAM[51178] = 8'b0;
    XRAM[51179] = 8'b0;
    XRAM[51180] = 8'b0;
    XRAM[51181] = 8'b0;
    XRAM[51182] = 8'b0;
    XRAM[51183] = 8'b0;
    XRAM[51184] = 8'b0;
    XRAM[51185] = 8'b0;
    XRAM[51186] = 8'b0;
    XRAM[51187] = 8'b0;
    XRAM[51188] = 8'b0;
    XRAM[51189] = 8'b0;
    XRAM[51190] = 8'b0;
    XRAM[51191] = 8'b0;
    XRAM[51192] = 8'b0;
    XRAM[51193] = 8'b0;
    XRAM[51194] = 8'b0;
    XRAM[51195] = 8'b0;
    XRAM[51196] = 8'b0;
    XRAM[51197] = 8'b0;
    XRAM[51198] = 8'b0;
    XRAM[51199] = 8'b0;
    XRAM[51200] = 8'b0;
    XRAM[51201] = 8'b0;
    XRAM[51202] = 8'b0;
    XRAM[51203] = 8'b0;
    XRAM[51204] = 8'b0;
    XRAM[51205] = 8'b0;
    XRAM[51206] = 8'b0;
    XRAM[51207] = 8'b0;
    XRAM[51208] = 8'b0;
    XRAM[51209] = 8'b0;
    XRAM[51210] = 8'b0;
    XRAM[51211] = 8'b0;
    XRAM[51212] = 8'b0;
    XRAM[51213] = 8'b0;
    XRAM[51214] = 8'b0;
    XRAM[51215] = 8'b0;
    XRAM[51216] = 8'b0;
    XRAM[51217] = 8'b0;
    XRAM[51218] = 8'b0;
    XRAM[51219] = 8'b0;
    XRAM[51220] = 8'b0;
    XRAM[51221] = 8'b0;
    XRAM[51222] = 8'b0;
    XRAM[51223] = 8'b0;
    XRAM[51224] = 8'b0;
    XRAM[51225] = 8'b0;
    XRAM[51226] = 8'b0;
    XRAM[51227] = 8'b0;
    XRAM[51228] = 8'b0;
    XRAM[51229] = 8'b0;
    XRAM[51230] = 8'b0;
    XRAM[51231] = 8'b0;
    XRAM[51232] = 8'b0;
    XRAM[51233] = 8'b0;
    XRAM[51234] = 8'b0;
    XRAM[51235] = 8'b0;
    XRAM[51236] = 8'b0;
    XRAM[51237] = 8'b0;
    XRAM[51238] = 8'b0;
    XRAM[51239] = 8'b0;
    XRAM[51240] = 8'b0;
    XRAM[51241] = 8'b0;
    XRAM[51242] = 8'b0;
    XRAM[51243] = 8'b0;
    XRAM[51244] = 8'b0;
    XRAM[51245] = 8'b0;
    XRAM[51246] = 8'b0;
    XRAM[51247] = 8'b0;
    XRAM[51248] = 8'b0;
    XRAM[51249] = 8'b0;
    XRAM[51250] = 8'b0;
    XRAM[51251] = 8'b0;
    XRAM[51252] = 8'b0;
    XRAM[51253] = 8'b0;
    XRAM[51254] = 8'b0;
    XRAM[51255] = 8'b0;
    XRAM[51256] = 8'b0;
    XRAM[51257] = 8'b0;
    XRAM[51258] = 8'b0;
    XRAM[51259] = 8'b0;
    XRAM[51260] = 8'b0;
    XRAM[51261] = 8'b0;
    XRAM[51262] = 8'b0;
    XRAM[51263] = 8'b0;
    XRAM[51264] = 8'b0;
    XRAM[51265] = 8'b0;
    XRAM[51266] = 8'b0;
    XRAM[51267] = 8'b0;
    XRAM[51268] = 8'b0;
    XRAM[51269] = 8'b0;
    XRAM[51270] = 8'b0;
    XRAM[51271] = 8'b0;
    XRAM[51272] = 8'b0;
    XRAM[51273] = 8'b0;
    XRAM[51274] = 8'b0;
    XRAM[51275] = 8'b0;
    XRAM[51276] = 8'b0;
    XRAM[51277] = 8'b0;
    XRAM[51278] = 8'b0;
    XRAM[51279] = 8'b0;
    XRAM[51280] = 8'b0;
    XRAM[51281] = 8'b0;
    XRAM[51282] = 8'b0;
    XRAM[51283] = 8'b0;
    XRAM[51284] = 8'b0;
    XRAM[51285] = 8'b0;
    XRAM[51286] = 8'b0;
    XRAM[51287] = 8'b0;
    XRAM[51288] = 8'b0;
    XRAM[51289] = 8'b0;
    XRAM[51290] = 8'b0;
    XRAM[51291] = 8'b0;
    XRAM[51292] = 8'b0;
    XRAM[51293] = 8'b0;
    XRAM[51294] = 8'b0;
    XRAM[51295] = 8'b0;
    XRAM[51296] = 8'b0;
    XRAM[51297] = 8'b0;
    XRAM[51298] = 8'b0;
    XRAM[51299] = 8'b0;
    XRAM[51300] = 8'b0;
    XRAM[51301] = 8'b0;
    XRAM[51302] = 8'b0;
    XRAM[51303] = 8'b0;
    XRAM[51304] = 8'b0;
    XRAM[51305] = 8'b0;
    XRAM[51306] = 8'b0;
    XRAM[51307] = 8'b0;
    XRAM[51308] = 8'b0;
    XRAM[51309] = 8'b0;
    XRAM[51310] = 8'b0;
    XRAM[51311] = 8'b0;
    XRAM[51312] = 8'b0;
    XRAM[51313] = 8'b0;
    XRAM[51314] = 8'b0;
    XRAM[51315] = 8'b0;
    XRAM[51316] = 8'b0;
    XRAM[51317] = 8'b0;
    XRAM[51318] = 8'b0;
    XRAM[51319] = 8'b0;
    XRAM[51320] = 8'b0;
    XRAM[51321] = 8'b0;
    XRAM[51322] = 8'b0;
    XRAM[51323] = 8'b0;
    XRAM[51324] = 8'b0;
    XRAM[51325] = 8'b0;
    XRAM[51326] = 8'b0;
    XRAM[51327] = 8'b0;
    XRAM[51328] = 8'b0;
    XRAM[51329] = 8'b0;
    XRAM[51330] = 8'b0;
    XRAM[51331] = 8'b0;
    XRAM[51332] = 8'b0;
    XRAM[51333] = 8'b0;
    XRAM[51334] = 8'b0;
    XRAM[51335] = 8'b0;
    XRAM[51336] = 8'b0;
    XRAM[51337] = 8'b0;
    XRAM[51338] = 8'b0;
    XRAM[51339] = 8'b0;
    XRAM[51340] = 8'b0;
    XRAM[51341] = 8'b0;
    XRAM[51342] = 8'b0;
    XRAM[51343] = 8'b0;
    XRAM[51344] = 8'b0;
    XRAM[51345] = 8'b0;
    XRAM[51346] = 8'b0;
    XRAM[51347] = 8'b0;
    XRAM[51348] = 8'b0;
    XRAM[51349] = 8'b0;
    XRAM[51350] = 8'b0;
    XRAM[51351] = 8'b0;
    XRAM[51352] = 8'b0;
    XRAM[51353] = 8'b0;
    XRAM[51354] = 8'b0;
    XRAM[51355] = 8'b0;
    XRAM[51356] = 8'b0;
    XRAM[51357] = 8'b0;
    XRAM[51358] = 8'b0;
    XRAM[51359] = 8'b0;
    XRAM[51360] = 8'b0;
    XRAM[51361] = 8'b0;
    XRAM[51362] = 8'b0;
    XRAM[51363] = 8'b0;
    XRAM[51364] = 8'b0;
    XRAM[51365] = 8'b0;
    XRAM[51366] = 8'b0;
    XRAM[51367] = 8'b0;
    XRAM[51368] = 8'b0;
    XRAM[51369] = 8'b0;
    XRAM[51370] = 8'b0;
    XRAM[51371] = 8'b0;
    XRAM[51372] = 8'b0;
    XRAM[51373] = 8'b0;
    XRAM[51374] = 8'b0;
    XRAM[51375] = 8'b0;
    XRAM[51376] = 8'b0;
    XRAM[51377] = 8'b0;
    XRAM[51378] = 8'b0;
    XRAM[51379] = 8'b0;
    XRAM[51380] = 8'b0;
    XRAM[51381] = 8'b0;
    XRAM[51382] = 8'b0;
    XRAM[51383] = 8'b0;
    XRAM[51384] = 8'b0;
    XRAM[51385] = 8'b0;
    XRAM[51386] = 8'b0;
    XRAM[51387] = 8'b0;
    XRAM[51388] = 8'b0;
    XRAM[51389] = 8'b0;
    XRAM[51390] = 8'b0;
    XRAM[51391] = 8'b0;
    XRAM[51392] = 8'b0;
    XRAM[51393] = 8'b0;
    XRAM[51394] = 8'b0;
    XRAM[51395] = 8'b0;
    XRAM[51396] = 8'b0;
    XRAM[51397] = 8'b0;
    XRAM[51398] = 8'b0;
    XRAM[51399] = 8'b0;
    XRAM[51400] = 8'b0;
    XRAM[51401] = 8'b0;
    XRAM[51402] = 8'b0;
    XRAM[51403] = 8'b0;
    XRAM[51404] = 8'b0;
    XRAM[51405] = 8'b0;
    XRAM[51406] = 8'b0;
    XRAM[51407] = 8'b0;
    XRAM[51408] = 8'b0;
    XRAM[51409] = 8'b0;
    XRAM[51410] = 8'b0;
    XRAM[51411] = 8'b0;
    XRAM[51412] = 8'b0;
    XRAM[51413] = 8'b0;
    XRAM[51414] = 8'b0;
    XRAM[51415] = 8'b0;
    XRAM[51416] = 8'b0;
    XRAM[51417] = 8'b0;
    XRAM[51418] = 8'b0;
    XRAM[51419] = 8'b0;
    XRAM[51420] = 8'b0;
    XRAM[51421] = 8'b0;
    XRAM[51422] = 8'b0;
    XRAM[51423] = 8'b0;
    XRAM[51424] = 8'b0;
    XRAM[51425] = 8'b0;
    XRAM[51426] = 8'b0;
    XRAM[51427] = 8'b0;
    XRAM[51428] = 8'b0;
    XRAM[51429] = 8'b0;
    XRAM[51430] = 8'b0;
    XRAM[51431] = 8'b0;
    XRAM[51432] = 8'b0;
    XRAM[51433] = 8'b0;
    XRAM[51434] = 8'b0;
    XRAM[51435] = 8'b0;
    XRAM[51436] = 8'b0;
    XRAM[51437] = 8'b0;
    XRAM[51438] = 8'b0;
    XRAM[51439] = 8'b0;
    XRAM[51440] = 8'b0;
    XRAM[51441] = 8'b0;
    XRAM[51442] = 8'b0;
    XRAM[51443] = 8'b0;
    XRAM[51444] = 8'b0;
    XRAM[51445] = 8'b0;
    XRAM[51446] = 8'b0;
    XRAM[51447] = 8'b0;
    XRAM[51448] = 8'b0;
    XRAM[51449] = 8'b0;
    XRAM[51450] = 8'b0;
    XRAM[51451] = 8'b0;
    XRAM[51452] = 8'b0;
    XRAM[51453] = 8'b0;
    XRAM[51454] = 8'b0;
    XRAM[51455] = 8'b0;
    XRAM[51456] = 8'b0;
    XRAM[51457] = 8'b0;
    XRAM[51458] = 8'b0;
    XRAM[51459] = 8'b0;
    XRAM[51460] = 8'b0;
    XRAM[51461] = 8'b0;
    XRAM[51462] = 8'b0;
    XRAM[51463] = 8'b0;
    XRAM[51464] = 8'b0;
    XRAM[51465] = 8'b0;
    XRAM[51466] = 8'b0;
    XRAM[51467] = 8'b0;
    XRAM[51468] = 8'b0;
    XRAM[51469] = 8'b0;
    XRAM[51470] = 8'b0;
    XRAM[51471] = 8'b0;
    XRAM[51472] = 8'b0;
    XRAM[51473] = 8'b0;
    XRAM[51474] = 8'b0;
    XRAM[51475] = 8'b0;
    XRAM[51476] = 8'b0;
    XRAM[51477] = 8'b0;
    XRAM[51478] = 8'b0;
    XRAM[51479] = 8'b0;
    XRAM[51480] = 8'b0;
    XRAM[51481] = 8'b0;
    XRAM[51482] = 8'b0;
    XRAM[51483] = 8'b0;
    XRAM[51484] = 8'b0;
    XRAM[51485] = 8'b0;
    XRAM[51486] = 8'b0;
    XRAM[51487] = 8'b0;
    XRAM[51488] = 8'b0;
    XRAM[51489] = 8'b0;
    XRAM[51490] = 8'b0;
    XRAM[51491] = 8'b0;
    XRAM[51492] = 8'b0;
    XRAM[51493] = 8'b0;
    XRAM[51494] = 8'b0;
    XRAM[51495] = 8'b0;
    XRAM[51496] = 8'b0;
    XRAM[51497] = 8'b0;
    XRAM[51498] = 8'b0;
    XRAM[51499] = 8'b0;
    XRAM[51500] = 8'b0;
    XRAM[51501] = 8'b0;
    XRAM[51502] = 8'b0;
    XRAM[51503] = 8'b0;
    XRAM[51504] = 8'b0;
    XRAM[51505] = 8'b0;
    XRAM[51506] = 8'b0;
    XRAM[51507] = 8'b0;
    XRAM[51508] = 8'b0;
    XRAM[51509] = 8'b0;
    XRAM[51510] = 8'b0;
    XRAM[51511] = 8'b0;
    XRAM[51512] = 8'b0;
    XRAM[51513] = 8'b0;
    XRAM[51514] = 8'b0;
    XRAM[51515] = 8'b0;
    XRAM[51516] = 8'b0;
    XRAM[51517] = 8'b0;
    XRAM[51518] = 8'b0;
    XRAM[51519] = 8'b0;
    XRAM[51520] = 8'b0;
    XRAM[51521] = 8'b0;
    XRAM[51522] = 8'b0;
    XRAM[51523] = 8'b0;
    XRAM[51524] = 8'b0;
    XRAM[51525] = 8'b0;
    XRAM[51526] = 8'b0;
    XRAM[51527] = 8'b0;
    XRAM[51528] = 8'b0;
    XRAM[51529] = 8'b0;
    XRAM[51530] = 8'b0;
    XRAM[51531] = 8'b0;
    XRAM[51532] = 8'b0;
    XRAM[51533] = 8'b0;
    XRAM[51534] = 8'b0;
    XRAM[51535] = 8'b0;
    XRAM[51536] = 8'b0;
    XRAM[51537] = 8'b0;
    XRAM[51538] = 8'b0;
    XRAM[51539] = 8'b0;
    XRAM[51540] = 8'b0;
    XRAM[51541] = 8'b0;
    XRAM[51542] = 8'b0;
    XRAM[51543] = 8'b0;
    XRAM[51544] = 8'b0;
    XRAM[51545] = 8'b0;
    XRAM[51546] = 8'b0;
    XRAM[51547] = 8'b0;
    XRAM[51548] = 8'b0;
    XRAM[51549] = 8'b0;
    XRAM[51550] = 8'b0;
    XRAM[51551] = 8'b0;
    XRAM[51552] = 8'b0;
    XRAM[51553] = 8'b0;
    XRAM[51554] = 8'b0;
    XRAM[51555] = 8'b0;
    XRAM[51556] = 8'b0;
    XRAM[51557] = 8'b0;
    XRAM[51558] = 8'b0;
    XRAM[51559] = 8'b0;
    XRAM[51560] = 8'b0;
    XRAM[51561] = 8'b0;
    XRAM[51562] = 8'b0;
    XRAM[51563] = 8'b0;
    XRAM[51564] = 8'b0;
    XRAM[51565] = 8'b0;
    XRAM[51566] = 8'b0;
    XRAM[51567] = 8'b0;
    XRAM[51568] = 8'b0;
    XRAM[51569] = 8'b0;
    XRAM[51570] = 8'b0;
    XRAM[51571] = 8'b0;
    XRAM[51572] = 8'b0;
    XRAM[51573] = 8'b0;
    XRAM[51574] = 8'b0;
    XRAM[51575] = 8'b0;
    XRAM[51576] = 8'b0;
    XRAM[51577] = 8'b0;
    XRAM[51578] = 8'b0;
    XRAM[51579] = 8'b0;
    XRAM[51580] = 8'b0;
    XRAM[51581] = 8'b0;
    XRAM[51582] = 8'b0;
    XRAM[51583] = 8'b0;
    XRAM[51584] = 8'b0;
    XRAM[51585] = 8'b0;
    XRAM[51586] = 8'b0;
    XRAM[51587] = 8'b0;
    XRAM[51588] = 8'b0;
    XRAM[51589] = 8'b0;
    XRAM[51590] = 8'b0;
    XRAM[51591] = 8'b0;
    XRAM[51592] = 8'b0;
    XRAM[51593] = 8'b0;
    XRAM[51594] = 8'b0;
    XRAM[51595] = 8'b0;
    XRAM[51596] = 8'b0;
    XRAM[51597] = 8'b0;
    XRAM[51598] = 8'b0;
    XRAM[51599] = 8'b0;
    XRAM[51600] = 8'b0;
    XRAM[51601] = 8'b0;
    XRAM[51602] = 8'b0;
    XRAM[51603] = 8'b0;
    XRAM[51604] = 8'b0;
    XRAM[51605] = 8'b0;
    XRAM[51606] = 8'b0;
    XRAM[51607] = 8'b0;
    XRAM[51608] = 8'b0;
    XRAM[51609] = 8'b0;
    XRAM[51610] = 8'b0;
    XRAM[51611] = 8'b0;
    XRAM[51612] = 8'b0;
    XRAM[51613] = 8'b0;
    XRAM[51614] = 8'b0;
    XRAM[51615] = 8'b0;
    XRAM[51616] = 8'b0;
    XRAM[51617] = 8'b0;
    XRAM[51618] = 8'b0;
    XRAM[51619] = 8'b0;
    XRAM[51620] = 8'b0;
    XRAM[51621] = 8'b0;
    XRAM[51622] = 8'b0;
    XRAM[51623] = 8'b0;
    XRAM[51624] = 8'b0;
    XRAM[51625] = 8'b0;
    XRAM[51626] = 8'b0;
    XRAM[51627] = 8'b0;
    XRAM[51628] = 8'b0;
    XRAM[51629] = 8'b0;
    XRAM[51630] = 8'b0;
    XRAM[51631] = 8'b0;
    XRAM[51632] = 8'b0;
    XRAM[51633] = 8'b0;
    XRAM[51634] = 8'b0;
    XRAM[51635] = 8'b0;
    XRAM[51636] = 8'b0;
    XRAM[51637] = 8'b0;
    XRAM[51638] = 8'b0;
    XRAM[51639] = 8'b0;
    XRAM[51640] = 8'b0;
    XRAM[51641] = 8'b0;
    XRAM[51642] = 8'b0;
    XRAM[51643] = 8'b0;
    XRAM[51644] = 8'b0;
    XRAM[51645] = 8'b0;
    XRAM[51646] = 8'b0;
    XRAM[51647] = 8'b0;
    XRAM[51648] = 8'b0;
    XRAM[51649] = 8'b0;
    XRAM[51650] = 8'b0;
    XRAM[51651] = 8'b0;
    XRAM[51652] = 8'b0;
    XRAM[51653] = 8'b0;
    XRAM[51654] = 8'b0;
    XRAM[51655] = 8'b0;
    XRAM[51656] = 8'b0;
    XRAM[51657] = 8'b0;
    XRAM[51658] = 8'b0;
    XRAM[51659] = 8'b0;
    XRAM[51660] = 8'b0;
    XRAM[51661] = 8'b0;
    XRAM[51662] = 8'b0;
    XRAM[51663] = 8'b0;
    XRAM[51664] = 8'b0;
    XRAM[51665] = 8'b0;
    XRAM[51666] = 8'b0;
    XRAM[51667] = 8'b0;
    XRAM[51668] = 8'b0;
    XRAM[51669] = 8'b0;
    XRAM[51670] = 8'b0;
    XRAM[51671] = 8'b0;
    XRAM[51672] = 8'b0;
    XRAM[51673] = 8'b0;
    XRAM[51674] = 8'b0;
    XRAM[51675] = 8'b0;
    XRAM[51676] = 8'b0;
    XRAM[51677] = 8'b0;
    XRAM[51678] = 8'b0;
    XRAM[51679] = 8'b0;
    XRAM[51680] = 8'b0;
    XRAM[51681] = 8'b0;
    XRAM[51682] = 8'b0;
    XRAM[51683] = 8'b0;
    XRAM[51684] = 8'b0;
    XRAM[51685] = 8'b0;
    XRAM[51686] = 8'b0;
    XRAM[51687] = 8'b0;
    XRAM[51688] = 8'b0;
    XRAM[51689] = 8'b0;
    XRAM[51690] = 8'b0;
    XRAM[51691] = 8'b0;
    XRAM[51692] = 8'b0;
    XRAM[51693] = 8'b0;
    XRAM[51694] = 8'b0;
    XRAM[51695] = 8'b0;
    XRAM[51696] = 8'b0;
    XRAM[51697] = 8'b0;
    XRAM[51698] = 8'b0;
    XRAM[51699] = 8'b0;
    XRAM[51700] = 8'b0;
    XRAM[51701] = 8'b0;
    XRAM[51702] = 8'b0;
    XRAM[51703] = 8'b0;
    XRAM[51704] = 8'b0;
    XRAM[51705] = 8'b0;
    XRAM[51706] = 8'b0;
    XRAM[51707] = 8'b0;
    XRAM[51708] = 8'b0;
    XRAM[51709] = 8'b0;
    XRAM[51710] = 8'b0;
    XRAM[51711] = 8'b0;
    XRAM[51712] = 8'b0;
    XRAM[51713] = 8'b0;
    XRAM[51714] = 8'b0;
    XRAM[51715] = 8'b0;
    XRAM[51716] = 8'b0;
    XRAM[51717] = 8'b0;
    XRAM[51718] = 8'b0;
    XRAM[51719] = 8'b0;
    XRAM[51720] = 8'b0;
    XRAM[51721] = 8'b0;
    XRAM[51722] = 8'b0;
    XRAM[51723] = 8'b0;
    XRAM[51724] = 8'b0;
    XRAM[51725] = 8'b0;
    XRAM[51726] = 8'b0;
    XRAM[51727] = 8'b0;
    XRAM[51728] = 8'b0;
    XRAM[51729] = 8'b0;
    XRAM[51730] = 8'b0;
    XRAM[51731] = 8'b0;
    XRAM[51732] = 8'b0;
    XRAM[51733] = 8'b0;
    XRAM[51734] = 8'b0;
    XRAM[51735] = 8'b0;
    XRAM[51736] = 8'b0;
    XRAM[51737] = 8'b0;
    XRAM[51738] = 8'b0;
    XRAM[51739] = 8'b0;
    XRAM[51740] = 8'b0;
    XRAM[51741] = 8'b0;
    XRAM[51742] = 8'b0;
    XRAM[51743] = 8'b0;
    XRAM[51744] = 8'b0;
    XRAM[51745] = 8'b0;
    XRAM[51746] = 8'b0;
    XRAM[51747] = 8'b0;
    XRAM[51748] = 8'b0;
    XRAM[51749] = 8'b0;
    XRAM[51750] = 8'b0;
    XRAM[51751] = 8'b0;
    XRAM[51752] = 8'b0;
    XRAM[51753] = 8'b0;
    XRAM[51754] = 8'b0;
    XRAM[51755] = 8'b0;
    XRAM[51756] = 8'b0;
    XRAM[51757] = 8'b0;
    XRAM[51758] = 8'b0;
    XRAM[51759] = 8'b0;
    XRAM[51760] = 8'b0;
    XRAM[51761] = 8'b0;
    XRAM[51762] = 8'b0;
    XRAM[51763] = 8'b0;
    XRAM[51764] = 8'b0;
    XRAM[51765] = 8'b0;
    XRAM[51766] = 8'b0;
    XRAM[51767] = 8'b0;
    XRAM[51768] = 8'b0;
    XRAM[51769] = 8'b0;
    XRAM[51770] = 8'b0;
    XRAM[51771] = 8'b0;
    XRAM[51772] = 8'b0;
    XRAM[51773] = 8'b0;
    XRAM[51774] = 8'b0;
    XRAM[51775] = 8'b0;
    XRAM[51776] = 8'b0;
    XRAM[51777] = 8'b0;
    XRAM[51778] = 8'b0;
    XRAM[51779] = 8'b0;
    XRAM[51780] = 8'b0;
    XRAM[51781] = 8'b0;
    XRAM[51782] = 8'b0;
    XRAM[51783] = 8'b0;
    XRAM[51784] = 8'b0;
    XRAM[51785] = 8'b0;
    XRAM[51786] = 8'b0;
    XRAM[51787] = 8'b0;
    XRAM[51788] = 8'b0;
    XRAM[51789] = 8'b0;
    XRAM[51790] = 8'b0;
    XRAM[51791] = 8'b0;
    XRAM[51792] = 8'b0;
    XRAM[51793] = 8'b0;
    XRAM[51794] = 8'b0;
    XRAM[51795] = 8'b0;
    XRAM[51796] = 8'b0;
    XRAM[51797] = 8'b0;
    XRAM[51798] = 8'b0;
    XRAM[51799] = 8'b0;
    XRAM[51800] = 8'b0;
    XRAM[51801] = 8'b0;
    XRAM[51802] = 8'b0;
    XRAM[51803] = 8'b0;
    XRAM[51804] = 8'b0;
    XRAM[51805] = 8'b0;
    XRAM[51806] = 8'b0;
    XRAM[51807] = 8'b0;
    XRAM[51808] = 8'b0;
    XRAM[51809] = 8'b0;
    XRAM[51810] = 8'b0;
    XRAM[51811] = 8'b0;
    XRAM[51812] = 8'b0;
    XRAM[51813] = 8'b0;
    XRAM[51814] = 8'b0;
    XRAM[51815] = 8'b0;
    XRAM[51816] = 8'b0;
    XRAM[51817] = 8'b0;
    XRAM[51818] = 8'b0;
    XRAM[51819] = 8'b0;
    XRAM[51820] = 8'b0;
    XRAM[51821] = 8'b0;
    XRAM[51822] = 8'b0;
    XRAM[51823] = 8'b0;
    XRAM[51824] = 8'b0;
    XRAM[51825] = 8'b0;
    XRAM[51826] = 8'b0;
    XRAM[51827] = 8'b0;
    XRAM[51828] = 8'b0;
    XRAM[51829] = 8'b0;
    XRAM[51830] = 8'b0;
    XRAM[51831] = 8'b0;
    XRAM[51832] = 8'b0;
    XRAM[51833] = 8'b0;
    XRAM[51834] = 8'b0;
    XRAM[51835] = 8'b0;
    XRAM[51836] = 8'b0;
    XRAM[51837] = 8'b0;
    XRAM[51838] = 8'b0;
    XRAM[51839] = 8'b0;
    XRAM[51840] = 8'b0;
    XRAM[51841] = 8'b0;
    XRAM[51842] = 8'b0;
    XRAM[51843] = 8'b0;
    XRAM[51844] = 8'b0;
    XRAM[51845] = 8'b0;
    XRAM[51846] = 8'b0;
    XRAM[51847] = 8'b0;
    XRAM[51848] = 8'b0;
    XRAM[51849] = 8'b0;
    XRAM[51850] = 8'b0;
    XRAM[51851] = 8'b0;
    XRAM[51852] = 8'b0;
    XRAM[51853] = 8'b0;
    XRAM[51854] = 8'b0;
    XRAM[51855] = 8'b0;
    XRAM[51856] = 8'b0;
    XRAM[51857] = 8'b0;
    XRAM[51858] = 8'b0;
    XRAM[51859] = 8'b0;
    XRAM[51860] = 8'b0;
    XRAM[51861] = 8'b0;
    XRAM[51862] = 8'b0;
    XRAM[51863] = 8'b0;
    XRAM[51864] = 8'b0;
    XRAM[51865] = 8'b0;
    XRAM[51866] = 8'b0;
    XRAM[51867] = 8'b0;
    XRAM[51868] = 8'b0;
    XRAM[51869] = 8'b0;
    XRAM[51870] = 8'b0;
    XRAM[51871] = 8'b0;
    XRAM[51872] = 8'b0;
    XRAM[51873] = 8'b0;
    XRAM[51874] = 8'b0;
    XRAM[51875] = 8'b0;
    XRAM[51876] = 8'b0;
    XRAM[51877] = 8'b0;
    XRAM[51878] = 8'b0;
    XRAM[51879] = 8'b0;
    XRAM[51880] = 8'b0;
    XRAM[51881] = 8'b0;
    XRAM[51882] = 8'b0;
    XRAM[51883] = 8'b0;
    XRAM[51884] = 8'b0;
    XRAM[51885] = 8'b0;
    XRAM[51886] = 8'b0;
    XRAM[51887] = 8'b0;
    XRAM[51888] = 8'b0;
    XRAM[51889] = 8'b0;
    XRAM[51890] = 8'b0;
    XRAM[51891] = 8'b0;
    XRAM[51892] = 8'b0;
    XRAM[51893] = 8'b0;
    XRAM[51894] = 8'b0;
    XRAM[51895] = 8'b0;
    XRAM[51896] = 8'b0;
    XRAM[51897] = 8'b0;
    XRAM[51898] = 8'b0;
    XRAM[51899] = 8'b0;
    XRAM[51900] = 8'b0;
    XRAM[51901] = 8'b0;
    XRAM[51902] = 8'b0;
    XRAM[51903] = 8'b0;
    XRAM[51904] = 8'b0;
    XRAM[51905] = 8'b0;
    XRAM[51906] = 8'b0;
    XRAM[51907] = 8'b0;
    XRAM[51908] = 8'b0;
    XRAM[51909] = 8'b0;
    XRAM[51910] = 8'b0;
    XRAM[51911] = 8'b0;
    XRAM[51912] = 8'b0;
    XRAM[51913] = 8'b0;
    XRAM[51914] = 8'b0;
    XRAM[51915] = 8'b0;
    XRAM[51916] = 8'b0;
    XRAM[51917] = 8'b0;
    XRAM[51918] = 8'b0;
    XRAM[51919] = 8'b0;
    XRAM[51920] = 8'b0;
    XRAM[51921] = 8'b0;
    XRAM[51922] = 8'b0;
    XRAM[51923] = 8'b0;
    XRAM[51924] = 8'b0;
    XRAM[51925] = 8'b0;
    XRAM[51926] = 8'b0;
    XRAM[51927] = 8'b0;
    XRAM[51928] = 8'b0;
    XRAM[51929] = 8'b0;
    XRAM[51930] = 8'b0;
    XRAM[51931] = 8'b0;
    XRAM[51932] = 8'b0;
    XRAM[51933] = 8'b0;
    XRAM[51934] = 8'b0;
    XRAM[51935] = 8'b0;
    XRAM[51936] = 8'b0;
    XRAM[51937] = 8'b0;
    XRAM[51938] = 8'b0;
    XRAM[51939] = 8'b0;
    XRAM[51940] = 8'b0;
    XRAM[51941] = 8'b0;
    XRAM[51942] = 8'b0;
    XRAM[51943] = 8'b0;
    XRAM[51944] = 8'b0;
    XRAM[51945] = 8'b0;
    XRAM[51946] = 8'b0;
    XRAM[51947] = 8'b0;
    XRAM[51948] = 8'b0;
    XRAM[51949] = 8'b0;
    XRAM[51950] = 8'b0;
    XRAM[51951] = 8'b0;
    XRAM[51952] = 8'b0;
    XRAM[51953] = 8'b0;
    XRAM[51954] = 8'b0;
    XRAM[51955] = 8'b0;
    XRAM[51956] = 8'b0;
    XRAM[51957] = 8'b0;
    XRAM[51958] = 8'b0;
    XRAM[51959] = 8'b0;
    XRAM[51960] = 8'b0;
    XRAM[51961] = 8'b0;
    XRAM[51962] = 8'b0;
    XRAM[51963] = 8'b0;
    XRAM[51964] = 8'b0;
    XRAM[51965] = 8'b0;
    XRAM[51966] = 8'b0;
    XRAM[51967] = 8'b0;
    XRAM[51968] = 8'b0;
    XRAM[51969] = 8'b0;
    XRAM[51970] = 8'b0;
    XRAM[51971] = 8'b0;
    XRAM[51972] = 8'b0;
    XRAM[51973] = 8'b0;
    XRAM[51974] = 8'b0;
    XRAM[51975] = 8'b0;
    XRAM[51976] = 8'b0;
    XRAM[51977] = 8'b0;
    XRAM[51978] = 8'b0;
    XRAM[51979] = 8'b0;
    XRAM[51980] = 8'b0;
    XRAM[51981] = 8'b0;
    XRAM[51982] = 8'b0;
    XRAM[51983] = 8'b0;
    XRAM[51984] = 8'b0;
    XRAM[51985] = 8'b0;
    XRAM[51986] = 8'b0;
    XRAM[51987] = 8'b0;
    XRAM[51988] = 8'b0;
    XRAM[51989] = 8'b0;
    XRAM[51990] = 8'b0;
    XRAM[51991] = 8'b0;
    XRAM[51992] = 8'b0;
    XRAM[51993] = 8'b0;
    XRAM[51994] = 8'b0;
    XRAM[51995] = 8'b0;
    XRAM[51996] = 8'b0;
    XRAM[51997] = 8'b0;
    XRAM[51998] = 8'b0;
    XRAM[51999] = 8'b0;
    XRAM[52000] = 8'b0;
    XRAM[52001] = 8'b0;
    XRAM[52002] = 8'b0;
    XRAM[52003] = 8'b0;
    XRAM[52004] = 8'b0;
    XRAM[52005] = 8'b0;
    XRAM[52006] = 8'b0;
    XRAM[52007] = 8'b0;
    XRAM[52008] = 8'b0;
    XRAM[52009] = 8'b0;
    XRAM[52010] = 8'b0;
    XRAM[52011] = 8'b0;
    XRAM[52012] = 8'b0;
    XRAM[52013] = 8'b0;
    XRAM[52014] = 8'b0;
    XRAM[52015] = 8'b0;
    XRAM[52016] = 8'b0;
    XRAM[52017] = 8'b0;
    XRAM[52018] = 8'b0;
    XRAM[52019] = 8'b0;
    XRAM[52020] = 8'b0;
    XRAM[52021] = 8'b0;
    XRAM[52022] = 8'b0;
    XRAM[52023] = 8'b0;
    XRAM[52024] = 8'b0;
    XRAM[52025] = 8'b0;
    XRAM[52026] = 8'b0;
    XRAM[52027] = 8'b0;
    XRAM[52028] = 8'b0;
    XRAM[52029] = 8'b0;
    XRAM[52030] = 8'b0;
    XRAM[52031] = 8'b0;
    XRAM[52032] = 8'b0;
    XRAM[52033] = 8'b0;
    XRAM[52034] = 8'b0;
    XRAM[52035] = 8'b0;
    XRAM[52036] = 8'b0;
    XRAM[52037] = 8'b0;
    XRAM[52038] = 8'b0;
    XRAM[52039] = 8'b0;
    XRAM[52040] = 8'b0;
    XRAM[52041] = 8'b0;
    XRAM[52042] = 8'b0;
    XRAM[52043] = 8'b0;
    XRAM[52044] = 8'b0;
    XRAM[52045] = 8'b0;
    XRAM[52046] = 8'b0;
    XRAM[52047] = 8'b0;
    XRAM[52048] = 8'b0;
    XRAM[52049] = 8'b0;
    XRAM[52050] = 8'b0;
    XRAM[52051] = 8'b0;
    XRAM[52052] = 8'b0;
    XRAM[52053] = 8'b0;
    XRAM[52054] = 8'b0;
    XRAM[52055] = 8'b0;
    XRAM[52056] = 8'b0;
    XRAM[52057] = 8'b0;
    XRAM[52058] = 8'b0;
    XRAM[52059] = 8'b0;
    XRAM[52060] = 8'b0;
    XRAM[52061] = 8'b0;
    XRAM[52062] = 8'b0;
    XRAM[52063] = 8'b0;
    XRAM[52064] = 8'b0;
    XRAM[52065] = 8'b0;
    XRAM[52066] = 8'b0;
    XRAM[52067] = 8'b0;
    XRAM[52068] = 8'b0;
    XRAM[52069] = 8'b0;
    XRAM[52070] = 8'b0;
    XRAM[52071] = 8'b0;
    XRAM[52072] = 8'b0;
    XRAM[52073] = 8'b0;
    XRAM[52074] = 8'b0;
    XRAM[52075] = 8'b0;
    XRAM[52076] = 8'b0;
    XRAM[52077] = 8'b0;
    XRAM[52078] = 8'b0;
    XRAM[52079] = 8'b0;
    XRAM[52080] = 8'b0;
    XRAM[52081] = 8'b0;
    XRAM[52082] = 8'b0;
    XRAM[52083] = 8'b0;
    XRAM[52084] = 8'b0;
    XRAM[52085] = 8'b0;
    XRAM[52086] = 8'b0;
    XRAM[52087] = 8'b0;
    XRAM[52088] = 8'b0;
    XRAM[52089] = 8'b0;
    XRAM[52090] = 8'b0;
    XRAM[52091] = 8'b0;
    XRAM[52092] = 8'b0;
    XRAM[52093] = 8'b0;
    XRAM[52094] = 8'b0;
    XRAM[52095] = 8'b0;
    XRAM[52096] = 8'b0;
    XRAM[52097] = 8'b0;
    XRAM[52098] = 8'b0;
    XRAM[52099] = 8'b0;
    XRAM[52100] = 8'b0;
    XRAM[52101] = 8'b0;
    XRAM[52102] = 8'b0;
    XRAM[52103] = 8'b0;
    XRAM[52104] = 8'b0;
    XRAM[52105] = 8'b0;
    XRAM[52106] = 8'b0;
    XRAM[52107] = 8'b0;
    XRAM[52108] = 8'b0;
    XRAM[52109] = 8'b0;
    XRAM[52110] = 8'b0;
    XRAM[52111] = 8'b0;
    XRAM[52112] = 8'b0;
    XRAM[52113] = 8'b0;
    XRAM[52114] = 8'b0;
    XRAM[52115] = 8'b0;
    XRAM[52116] = 8'b0;
    XRAM[52117] = 8'b0;
    XRAM[52118] = 8'b0;
    XRAM[52119] = 8'b0;
    XRAM[52120] = 8'b0;
    XRAM[52121] = 8'b0;
    XRAM[52122] = 8'b0;
    XRAM[52123] = 8'b0;
    XRAM[52124] = 8'b0;
    XRAM[52125] = 8'b0;
    XRAM[52126] = 8'b0;
    XRAM[52127] = 8'b0;
    XRAM[52128] = 8'b0;
    XRAM[52129] = 8'b0;
    XRAM[52130] = 8'b0;
    XRAM[52131] = 8'b0;
    XRAM[52132] = 8'b0;
    XRAM[52133] = 8'b0;
    XRAM[52134] = 8'b0;
    XRAM[52135] = 8'b0;
    XRAM[52136] = 8'b0;
    XRAM[52137] = 8'b0;
    XRAM[52138] = 8'b0;
    XRAM[52139] = 8'b0;
    XRAM[52140] = 8'b0;
    XRAM[52141] = 8'b0;
    XRAM[52142] = 8'b0;
    XRAM[52143] = 8'b0;
    XRAM[52144] = 8'b0;
    XRAM[52145] = 8'b0;
    XRAM[52146] = 8'b0;
    XRAM[52147] = 8'b0;
    XRAM[52148] = 8'b0;
    XRAM[52149] = 8'b0;
    XRAM[52150] = 8'b0;
    XRAM[52151] = 8'b0;
    XRAM[52152] = 8'b0;
    XRAM[52153] = 8'b0;
    XRAM[52154] = 8'b0;
    XRAM[52155] = 8'b0;
    XRAM[52156] = 8'b0;
    XRAM[52157] = 8'b0;
    XRAM[52158] = 8'b0;
    XRAM[52159] = 8'b0;
    XRAM[52160] = 8'b0;
    XRAM[52161] = 8'b0;
    XRAM[52162] = 8'b0;
    XRAM[52163] = 8'b0;
    XRAM[52164] = 8'b0;
    XRAM[52165] = 8'b0;
    XRAM[52166] = 8'b0;
    XRAM[52167] = 8'b0;
    XRAM[52168] = 8'b0;
    XRAM[52169] = 8'b0;
    XRAM[52170] = 8'b0;
    XRAM[52171] = 8'b0;
    XRAM[52172] = 8'b0;
    XRAM[52173] = 8'b0;
    XRAM[52174] = 8'b0;
    XRAM[52175] = 8'b0;
    XRAM[52176] = 8'b0;
    XRAM[52177] = 8'b0;
    XRAM[52178] = 8'b0;
    XRAM[52179] = 8'b0;
    XRAM[52180] = 8'b0;
    XRAM[52181] = 8'b0;
    XRAM[52182] = 8'b0;
    XRAM[52183] = 8'b0;
    XRAM[52184] = 8'b0;
    XRAM[52185] = 8'b0;
    XRAM[52186] = 8'b0;
    XRAM[52187] = 8'b0;
    XRAM[52188] = 8'b0;
    XRAM[52189] = 8'b0;
    XRAM[52190] = 8'b0;
    XRAM[52191] = 8'b0;
    XRAM[52192] = 8'b0;
    XRAM[52193] = 8'b0;
    XRAM[52194] = 8'b0;
    XRAM[52195] = 8'b0;
    XRAM[52196] = 8'b0;
    XRAM[52197] = 8'b0;
    XRAM[52198] = 8'b0;
    XRAM[52199] = 8'b0;
    XRAM[52200] = 8'b0;
    XRAM[52201] = 8'b0;
    XRAM[52202] = 8'b0;
    XRAM[52203] = 8'b0;
    XRAM[52204] = 8'b0;
    XRAM[52205] = 8'b0;
    XRAM[52206] = 8'b0;
    XRAM[52207] = 8'b0;
    XRAM[52208] = 8'b0;
    XRAM[52209] = 8'b0;
    XRAM[52210] = 8'b0;
    XRAM[52211] = 8'b0;
    XRAM[52212] = 8'b0;
    XRAM[52213] = 8'b0;
    XRAM[52214] = 8'b0;
    XRAM[52215] = 8'b0;
    XRAM[52216] = 8'b0;
    XRAM[52217] = 8'b0;
    XRAM[52218] = 8'b0;
    XRAM[52219] = 8'b0;
    XRAM[52220] = 8'b0;
    XRAM[52221] = 8'b0;
    XRAM[52222] = 8'b0;
    XRAM[52223] = 8'b0;
    XRAM[52224] = 8'b0;
    XRAM[52225] = 8'b0;
    XRAM[52226] = 8'b0;
    XRAM[52227] = 8'b0;
    XRAM[52228] = 8'b0;
    XRAM[52229] = 8'b0;
    XRAM[52230] = 8'b0;
    XRAM[52231] = 8'b0;
    XRAM[52232] = 8'b0;
    XRAM[52233] = 8'b0;
    XRAM[52234] = 8'b0;
    XRAM[52235] = 8'b0;
    XRAM[52236] = 8'b0;
    XRAM[52237] = 8'b0;
    XRAM[52238] = 8'b0;
    XRAM[52239] = 8'b0;
    XRAM[52240] = 8'b0;
    XRAM[52241] = 8'b0;
    XRAM[52242] = 8'b0;
    XRAM[52243] = 8'b0;
    XRAM[52244] = 8'b0;
    XRAM[52245] = 8'b0;
    XRAM[52246] = 8'b0;
    XRAM[52247] = 8'b0;
    XRAM[52248] = 8'b0;
    XRAM[52249] = 8'b0;
    XRAM[52250] = 8'b0;
    XRAM[52251] = 8'b0;
    XRAM[52252] = 8'b0;
    XRAM[52253] = 8'b0;
    XRAM[52254] = 8'b0;
    XRAM[52255] = 8'b0;
    XRAM[52256] = 8'b0;
    XRAM[52257] = 8'b0;
    XRAM[52258] = 8'b0;
    XRAM[52259] = 8'b0;
    XRAM[52260] = 8'b0;
    XRAM[52261] = 8'b0;
    XRAM[52262] = 8'b0;
    XRAM[52263] = 8'b0;
    XRAM[52264] = 8'b0;
    XRAM[52265] = 8'b0;
    XRAM[52266] = 8'b0;
    XRAM[52267] = 8'b0;
    XRAM[52268] = 8'b0;
    XRAM[52269] = 8'b0;
    XRAM[52270] = 8'b0;
    XRAM[52271] = 8'b0;
    XRAM[52272] = 8'b0;
    XRAM[52273] = 8'b0;
    XRAM[52274] = 8'b0;
    XRAM[52275] = 8'b0;
    XRAM[52276] = 8'b0;
    XRAM[52277] = 8'b0;
    XRAM[52278] = 8'b0;
    XRAM[52279] = 8'b0;
    XRAM[52280] = 8'b0;
    XRAM[52281] = 8'b0;
    XRAM[52282] = 8'b0;
    XRAM[52283] = 8'b0;
    XRAM[52284] = 8'b0;
    XRAM[52285] = 8'b0;
    XRAM[52286] = 8'b0;
    XRAM[52287] = 8'b0;
    XRAM[52288] = 8'b0;
    XRAM[52289] = 8'b0;
    XRAM[52290] = 8'b0;
    XRAM[52291] = 8'b0;
    XRAM[52292] = 8'b0;
    XRAM[52293] = 8'b0;
    XRAM[52294] = 8'b0;
    XRAM[52295] = 8'b0;
    XRAM[52296] = 8'b0;
    XRAM[52297] = 8'b0;
    XRAM[52298] = 8'b0;
    XRAM[52299] = 8'b0;
    XRAM[52300] = 8'b0;
    XRAM[52301] = 8'b0;
    XRAM[52302] = 8'b0;
    XRAM[52303] = 8'b0;
    XRAM[52304] = 8'b0;
    XRAM[52305] = 8'b0;
    XRAM[52306] = 8'b0;
    XRAM[52307] = 8'b0;
    XRAM[52308] = 8'b0;
    XRAM[52309] = 8'b0;
    XRAM[52310] = 8'b0;
    XRAM[52311] = 8'b0;
    XRAM[52312] = 8'b0;
    XRAM[52313] = 8'b0;
    XRAM[52314] = 8'b0;
    XRAM[52315] = 8'b0;
    XRAM[52316] = 8'b0;
    XRAM[52317] = 8'b0;
    XRAM[52318] = 8'b0;
    XRAM[52319] = 8'b0;
    XRAM[52320] = 8'b0;
    XRAM[52321] = 8'b0;
    XRAM[52322] = 8'b0;
    XRAM[52323] = 8'b0;
    XRAM[52324] = 8'b0;
    XRAM[52325] = 8'b0;
    XRAM[52326] = 8'b0;
    XRAM[52327] = 8'b0;
    XRAM[52328] = 8'b0;
    XRAM[52329] = 8'b0;
    XRAM[52330] = 8'b0;
    XRAM[52331] = 8'b0;
    XRAM[52332] = 8'b0;
    XRAM[52333] = 8'b0;
    XRAM[52334] = 8'b0;
    XRAM[52335] = 8'b0;
    XRAM[52336] = 8'b0;
    XRAM[52337] = 8'b0;
    XRAM[52338] = 8'b0;
    XRAM[52339] = 8'b0;
    XRAM[52340] = 8'b0;
    XRAM[52341] = 8'b0;
    XRAM[52342] = 8'b0;
    XRAM[52343] = 8'b0;
    XRAM[52344] = 8'b0;
    XRAM[52345] = 8'b0;
    XRAM[52346] = 8'b0;
    XRAM[52347] = 8'b0;
    XRAM[52348] = 8'b0;
    XRAM[52349] = 8'b0;
    XRAM[52350] = 8'b0;
    XRAM[52351] = 8'b0;
    XRAM[52352] = 8'b0;
    XRAM[52353] = 8'b0;
    XRAM[52354] = 8'b0;
    XRAM[52355] = 8'b0;
    XRAM[52356] = 8'b0;
    XRAM[52357] = 8'b0;
    XRAM[52358] = 8'b0;
    XRAM[52359] = 8'b0;
    XRAM[52360] = 8'b0;
    XRAM[52361] = 8'b0;
    XRAM[52362] = 8'b0;
    XRAM[52363] = 8'b0;
    XRAM[52364] = 8'b0;
    XRAM[52365] = 8'b0;
    XRAM[52366] = 8'b0;
    XRAM[52367] = 8'b0;
    XRAM[52368] = 8'b0;
    XRAM[52369] = 8'b0;
    XRAM[52370] = 8'b0;
    XRAM[52371] = 8'b0;
    XRAM[52372] = 8'b0;
    XRAM[52373] = 8'b0;
    XRAM[52374] = 8'b0;
    XRAM[52375] = 8'b0;
    XRAM[52376] = 8'b0;
    XRAM[52377] = 8'b0;
    XRAM[52378] = 8'b0;
    XRAM[52379] = 8'b0;
    XRAM[52380] = 8'b0;
    XRAM[52381] = 8'b0;
    XRAM[52382] = 8'b0;
    XRAM[52383] = 8'b0;
    XRAM[52384] = 8'b0;
    XRAM[52385] = 8'b0;
    XRAM[52386] = 8'b0;
    XRAM[52387] = 8'b0;
    XRAM[52388] = 8'b0;
    XRAM[52389] = 8'b0;
    XRAM[52390] = 8'b0;
    XRAM[52391] = 8'b0;
    XRAM[52392] = 8'b0;
    XRAM[52393] = 8'b0;
    XRAM[52394] = 8'b0;
    XRAM[52395] = 8'b0;
    XRAM[52396] = 8'b0;
    XRAM[52397] = 8'b0;
    XRAM[52398] = 8'b0;
    XRAM[52399] = 8'b0;
    XRAM[52400] = 8'b0;
    XRAM[52401] = 8'b0;
    XRAM[52402] = 8'b0;
    XRAM[52403] = 8'b0;
    XRAM[52404] = 8'b0;
    XRAM[52405] = 8'b0;
    XRAM[52406] = 8'b0;
    XRAM[52407] = 8'b0;
    XRAM[52408] = 8'b0;
    XRAM[52409] = 8'b0;
    XRAM[52410] = 8'b0;
    XRAM[52411] = 8'b0;
    XRAM[52412] = 8'b0;
    XRAM[52413] = 8'b0;
    XRAM[52414] = 8'b0;
    XRAM[52415] = 8'b0;
    XRAM[52416] = 8'b0;
    XRAM[52417] = 8'b0;
    XRAM[52418] = 8'b0;
    XRAM[52419] = 8'b0;
    XRAM[52420] = 8'b0;
    XRAM[52421] = 8'b0;
    XRAM[52422] = 8'b0;
    XRAM[52423] = 8'b0;
    XRAM[52424] = 8'b0;
    XRAM[52425] = 8'b0;
    XRAM[52426] = 8'b0;
    XRAM[52427] = 8'b0;
    XRAM[52428] = 8'b0;
    XRAM[52429] = 8'b0;
    XRAM[52430] = 8'b0;
    XRAM[52431] = 8'b0;
    XRAM[52432] = 8'b0;
    XRAM[52433] = 8'b0;
    XRAM[52434] = 8'b0;
    XRAM[52435] = 8'b0;
    XRAM[52436] = 8'b0;
    XRAM[52437] = 8'b0;
    XRAM[52438] = 8'b0;
    XRAM[52439] = 8'b0;
    XRAM[52440] = 8'b0;
    XRAM[52441] = 8'b0;
    XRAM[52442] = 8'b0;
    XRAM[52443] = 8'b0;
    XRAM[52444] = 8'b0;
    XRAM[52445] = 8'b0;
    XRAM[52446] = 8'b0;
    XRAM[52447] = 8'b0;
    XRAM[52448] = 8'b0;
    XRAM[52449] = 8'b0;
    XRAM[52450] = 8'b0;
    XRAM[52451] = 8'b0;
    XRAM[52452] = 8'b0;
    XRAM[52453] = 8'b0;
    XRAM[52454] = 8'b0;
    XRAM[52455] = 8'b0;
    XRAM[52456] = 8'b0;
    XRAM[52457] = 8'b0;
    XRAM[52458] = 8'b0;
    XRAM[52459] = 8'b0;
    XRAM[52460] = 8'b0;
    XRAM[52461] = 8'b0;
    XRAM[52462] = 8'b0;
    XRAM[52463] = 8'b0;
    XRAM[52464] = 8'b0;
    XRAM[52465] = 8'b0;
    XRAM[52466] = 8'b0;
    XRAM[52467] = 8'b0;
    XRAM[52468] = 8'b0;
    XRAM[52469] = 8'b0;
    XRAM[52470] = 8'b0;
    XRAM[52471] = 8'b0;
    XRAM[52472] = 8'b0;
    XRAM[52473] = 8'b0;
    XRAM[52474] = 8'b0;
    XRAM[52475] = 8'b0;
    XRAM[52476] = 8'b0;
    XRAM[52477] = 8'b0;
    XRAM[52478] = 8'b0;
    XRAM[52479] = 8'b0;
    XRAM[52480] = 8'b0;
    XRAM[52481] = 8'b0;
    XRAM[52482] = 8'b0;
    XRAM[52483] = 8'b0;
    XRAM[52484] = 8'b0;
    XRAM[52485] = 8'b0;
    XRAM[52486] = 8'b0;
    XRAM[52487] = 8'b0;
    XRAM[52488] = 8'b0;
    XRAM[52489] = 8'b0;
    XRAM[52490] = 8'b0;
    XRAM[52491] = 8'b0;
    XRAM[52492] = 8'b0;
    XRAM[52493] = 8'b0;
    XRAM[52494] = 8'b0;
    XRAM[52495] = 8'b0;
    XRAM[52496] = 8'b0;
    XRAM[52497] = 8'b0;
    XRAM[52498] = 8'b0;
    XRAM[52499] = 8'b0;
    XRAM[52500] = 8'b0;
    XRAM[52501] = 8'b0;
    XRAM[52502] = 8'b0;
    XRAM[52503] = 8'b0;
    XRAM[52504] = 8'b0;
    XRAM[52505] = 8'b0;
    XRAM[52506] = 8'b0;
    XRAM[52507] = 8'b0;
    XRAM[52508] = 8'b0;
    XRAM[52509] = 8'b0;
    XRAM[52510] = 8'b0;
    XRAM[52511] = 8'b0;
    XRAM[52512] = 8'b0;
    XRAM[52513] = 8'b0;
    XRAM[52514] = 8'b0;
    XRAM[52515] = 8'b0;
    XRAM[52516] = 8'b0;
    XRAM[52517] = 8'b0;
    XRAM[52518] = 8'b0;
    XRAM[52519] = 8'b0;
    XRAM[52520] = 8'b0;
    XRAM[52521] = 8'b0;
    XRAM[52522] = 8'b0;
    XRAM[52523] = 8'b0;
    XRAM[52524] = 8'b0;
    XRAM[52525] = 8'b0;
    XRAM[52526] = 8'b0;
    XRAM[52527] = 8'b0;
    XRAM[52528] = 8'b0;
    XRAM[52529] = 8'b0;
    XRAM[52530] = 8'b0;
    XRAM[52531] = 8'b0;
    XRAM[52532] = 8'b0;
    XRAM[52533] = 8'b0;
    XRAM[52534] = 8'b0;
    XRAM[52535] = 8'b0;
    XRAM[52536] = 8'b0;
    XRAM[52537] = 8'b0;
    XRAM[52538] = 8'b0;
    XRAM[52539] = 8'b0;
    XRAM[52540] = 8'b0;
    XRAM[52541] = 8'b0;
    XRAM[52542] = 8'b0;
    XRAM[52543] = 8'b0;
    XRAM[52544] = 8'b0;
    XRAM[52545] = 8'b0;
    XRAM[52546] = 8'b0;
    XRAM[52547] = 8'b0;
    XRAM[52548] = 8'b0;
    XRAM[52549] = 8'b0;
    XRAM[52550] = 8'b0;
    XRAM[52551] = 8'b0;
    XRAM[52552] = 8'b0;
    XRAM[52553] = 8'b0;
    XRAM[52554] = 8'b0;
    XRAM[52555] = 8'b0;
    XRAM[52556] = 8'b0;
    XRAM[52557] = 8'b0;
    XRAM[52558] = 8'b0;
    XRAM[52559] = 8'b0;
    XRAM[52560] = 8'b0;
    XRAM[52561] = 8'b0;
    XRAM[52562] = 8'b0;
    XRAM[52563] = 8'b0;
    XRAM[52564] = 8'b0;
    XRAM[52565] = 8'b0;
    XRAM[52566] = 8'b0;
    XRAM[52567] = 8'b0;
    XRAM[52568] = 8'b0;
    XRAM[52569] = 8'b0;
    XRAM[52570] = 8'b0;
    XRAM[52571] = 8'b0;
    XRAM[52572] = 8'b0;
    XRAM[52573] = 8'b0;
    XRAM[52574] = 8'b0;
    XRAM[52575] = 8'b0;
    XRAM[52576] = 8'b0;
    XRAM[52577] = 8'b0;
    XRAM[52578] = 8'b0;
    XRAM[52579] = 8'b0;
    XRAM[52580] = 8'b0;
    XRAM[52581] = 8'b0;
    XRAM[52582] = 8'b0;
    XRAM[52583] = 8'b0;
    XRAM[52584] = 8'b0;
    XRAM[52585] = 8'b0;
    XRAM[52586] = 8'b0;
    XRAM[52587] = 8'b0;
    XRAM[52588] = 8'b0;
    XRAM[52589] = 8'b0;
    XRAM[52590] = 8'b0;
    XRAM[52591] = 8'b0;
    XRAM[52592] = 8'b0;
    XRAM[52593] = 8'b0;
    XRAM[52594] = 8'b0;
    XRAM[52595] = 8'b0;
    XRAM[52596] = 8'b0;
    XRAM[52597] = 8'b0;
    XRAM[52598] = 8'b0;
    XRAM[52599] = 8'b0;
    XRAM[52600] = 8'b0;
    XRAM[52601] = 8'b0;
    XRAM[52602] = 8'b0;
    XRAM[52603] = 8'b0;
    XRAM[52604] = 8'b0;
    XRAM[52605] = 8'b0;
    XRAM[52606] = 8'b0;
    XRAM[52607] = 8'b0;
    XRAM[52608] = 8'b0;
    XRAM[52609] = 8'b0;
    XRAM[52610] = 8'b0;
    XRAM[52611] = 8'b0;
    XRAM[52612] = 8'b0;
    XRAM[52613] = 8'b0;
    XRAM[52614] = 8'b0;
    XRAM[52615] = 8'b0;
    XRAM[52616] = 8'b0;
    XRAM[52617] = 8'b0;
    XRAM[52618] = 8'b0;
    XRAM[52619] = 8'b0;
    XRAM[52620] = 8'b0;
    XRAM[52621] = 8'b0;
    XRAM[52622] = 8'b0;
    XRAM[52623] = 8'b0;
    XRAM[52624] = 8'b0;
    XRAM[52625] = 8'b0;
    XRAM[52626] = 8'b0;
    XRAM[52627] = 8'b0;
    XRAM[52628] = 8'b0;
    XRAM[52629] = 8'b0;
    XRAM[52630] = 8'b0;
    XRAM[52631] = 8'b0;
    XRAM[52632] = 8'b0;
    XRAM[52633] = 8'b0;
    XRAM[52634] = 8'b0;
    XRAM[52635] = 8'b0;
    XRAM[52636] = 8'b0;
    XRAM[52637] = 8'b0;
    XRAM[52638] = 8'b0;
    XRAM[52639] = 8'b0;
    XRAM[52640] = 8'b0;
    XRAM[52641] = 8'b0;
    XRAM[52642] = 8'b0;
    XRAM[52643] = 8'b0;
    XRAM[52644] = 8'b0;
    XRAM[52645] = 8'b0;
    XRAM[52646] = 8'b0;
    XRAM[52647] = 8'b0;
    XRAM[52648] = 8'b0;
    XRAM[52649] = 8'b0;
    XRAM[52650] = 8'b0;
    XRAM[52651] = 8'b0;
    XRAM[52652] = 8'b0;
    XRAM[52653] = 8'b0;
    XRAM[52654] = 8'b0;
    XRAM[52655] = 8'b0;
    XRAM[52656] = 8'b0;
    XRAM[52657] = 8'b0;
    XRAM[52658] = 8'b0;
    XRAM[52659] = 8'b0;
    XRAM[52660] = 8'b0;
    XRAM[52661] = 8'b0;
    XRAM[52662] = 8'b0;
    XRAM[52663] = 8'b0;
    XRAM[52664] = 8'b0;
    XRAM[52665] = 8'b0;
    XRAM[52666] = 8'b0;
    XRAM[52667] = 8'b0;
    XRAM[52668] = 8'b0;
    XRAM[52669] = 8'b0;
    XRAM[52670] = 8'b0;
    XRAM[52671] = 8'b0;
    XRAM[52672] = 8'b0;
    XRAM[52673] = 8'b0;
    XRAM[52674] = 8'b0;
    XRAM[52675] = 8'b0;
    XRAM[52676] = 8'b0;
    XRAM[52677] = 8'b0;
    XRAM[52678] = 8'b0;
    XRAM[52679] = 8'b0;
    XRAM[52680] = 8'b0;
    XRAM[52681] = 8'b0;
    XRAM[52682] = 8'b0;
    XRAM[52683] = 8'b0;
    XRAM[52684] = 8'b0;
    XRAM[52685] = 8'b0;
    XRAM[52686] = 8'b0;
    XRAM[52687] = 8'b0;
    XRAM[52688] = 8'b0;
    XRAM[52689] = 8'b0;
    XRAM[52690] = 8'b0;
    XRAM[52691] = 8'b0;
    XRAM[52692] = 8'b0;
    XRAM[52693] = 8'b0;
    XRAM[52694] = 8'b0;
    XRAM[52695] = 8'b0;
    XRAM[52696] = 8'b0;
    XRAM[52697] = 8'b0;
    XRAM[52698] = 8'b0;
    XRAM[52699] = 8'b0;
    XRAM[52700] = 8'b0;
    XRAM[52701] = 8'b0;
    XRAM[52702] = 8'b0;
    XRAM[52703] = 8'b0;
    XRAM[52704] = 8'b0;
    XRAM[52705] = 8'b0;
    XRAM[52706] = 8'b0;
    XRAM[52707] = 8'b0;
    XRAM[52708] = 8'b0;
    XRAM[52709] = 8'b0;
    XRAM[52710] = 8'b0;
    XRAM[52711] = 8'b0;
    XRAM[52712] = 8'b0;
    XRAM[52713] = 8'b0;
    XRAM[52714] = 8'b0;
    XRAM[52715] = 8'b0;
    XRAM[52716] = 8'b0;
    XRAM[52717] = 8'b0;
    XRAM[52718] = 8'b0;
    XRAM[52719] = 8'b0;
    XRAM[52720] = 8'b0;
    XRAM[52721] = 8'b0;
    XRAM[52722] = 8'b0;
    XRAM[52723] = 8'b0;
    XRAM[52724] = 8'b0;
    XRAM[52725] = 8'b0;
    XRAM[52726] = 8'b0;
    XRAM[52727] = 8'b0;
    XRAM[52728] = 8'b0;
    XRAM[52729] = 8'b0;
    XRAM[52730] = 8'b0;
    XRAM[52731] = 8'b0;
    XRAM[52732] = 8'b0;
    XRAM[52733] = 8'b0;
    XRAM[52734] = 8'b0;
    XRAM[52735] = 8'b0;
    XRAM[52736] = 8'b0;
    XRAM[52737] = 8'b0;
    XRAM[52738] = 8'b0;
    XRAM[52739] = 8'b0;
    XRAM[52740] = 8'b0;
    XRAM[52741] = 8'b0;
    XRAM[52742] = 8'b0;
    XRAM[52743] = 8'b0;
    XRAM[52744] = 8'b0;
    XRAM[52745] = 8'b0;
    XRAM[52746] = 8'b0;
    XRAM[52747] = 8'b0;
    XRAM[52748] = 8'b0;
    XRAM[52749] = 8'b0;
    XRAM[52750] = 8'b0;
    XRAM[52751] = 8'b0;
    XRAM[52752] = 8'b0;
    XRAM[52753] = 8'b0;
    XRAM[52754] = 8'b0;
    XRAM[52755] = 8'b0;
    XRAM[52756] = 8'b0;
    XRAM[52757] = 8'b0;
    XRAM[52758] = 8'b0;
    XRAM[52759] = 8'b0;
    XRAM[52760] = 8'b0;
    XRAM[52761] = 8'b0;
    XRAM[52762] = 8'b0;
    XRAM[52763] = 8'b0;
    XRAM[52764] = 8'b0;
    XRAM[52765] = 8'b0;
    XRAM[52766] = 8'b0;
    XRAM[52767] = 8'b0;
    XRAM[52768] = 8'b0;
    XRAM[52769] = 8'b0;
    XRAM[52770] = 8'b0;
    XRAM[52771] = 8'b0;
    XRAM[52772] = 8'b0;
    XRAM[52773] = 8'b0;
    XRAM[52774] = 8'b0;
    XRAM[52775] = 8'b0;
    XRAM[52776] = 8'b0;
    XRAM[52777] = 8'b0;
    XRAM[52778] = 8'b0;
    XRAM[52779] = 8'b0;
    XRAM[52780] = 8'b0;
    XRAM[52781] = 8'b0;
    XRAM[52782] = 8'b0;
    XRAM[52783] = 8'b0;
    XRAM[52784] = 8'b0;
    XRAM[52785] = 8'b0;
    XRAM[52786] = 8'b0;
    XRAM[52787] = 8'b0;
    XRAM[52788] = 8'b0;
    XRAM[52789] = 8'b0;
    XRAM[52790] = 8'b0;
    XRAM[52791] = 8'b0;
    XRAM[52792] = 8'b0;
    XRAM[52793] = 8'b0;
    XRAM[52794] = 8'b0;
    XRAM[52795] = 8'b0;
    XRAM[52796] = 8'b0;
    XRAM[52797] = 8'b0;
    XRAM[52798] = 8'b0;
    XRAM[52799] = 8'b0;
    XRAM[52800] = 8'b0;
    XRAM[52801] = 8'b0;
    XRAM[52802] = 8'b0;
    XRAM[52803] = 8'b0;
    XRAM[52804] = 8'b0;
    XRAM[52805] = 8'b0;
    XRAM[52806] = 8'b0;
    XRAM[52807] = 8'b0;
    XRAM[52808] = 8'b0;
    XRAM[52809] = 8'b0;
    XRAM[52810] = 8'b0;
    XRAM[52811] = 8'b0;
    XRAM[52812] = 8'b0;
    XRAM[52813] = 8'b0;
    XRAM[52814] = 8'b0;
    XRAM[52815] = 8'b0;
    XRAM[52816] = 8'b0;
    XRAM[52817] = 8'b0;
    XRAM[52818] = 8'b0;
    XRAM[52819] = 8'b0;
    XRAM[52820] = 8'b0;
    XRAM[52821] = 8'b0;
    XRAM[52822] = 8'b0;
    XRAM[52823] = 8'b0;
    XRAM[52824] = 8'b0;
    XRAM[52825] = 8'b0;
    XRAM[52826] = 8'b0;
    XRAM[52827] = 8'b0;
    XRAM[52828] = 8'b0;
    XRAM[52829] = 8'b0;
    XRAM[52830] = 8'b0;
    XRAM[52831] = 8'b0;
    XRAM[52832] = 8'b0;
    XRAM[52833] = 8'b0;
    XRAM[52834] = 8'b0;
    XRAM[52835] = 8'b0;
    XRAM[52836] = 8'b0;
    XRAM[52837] = 8'b0;
    XRAM[52838] = 8'b0;
    XRAM[52839] = 8'b0;
    XRAM[52840] = 8'b0;
    XRAM[52841] = 8'b0;
    XRAM[52842] = 8'b0;
    XRAM[52843] = 8'b0;
    XRAM[52844] = 8'b0;
    XRAM[52845] = 8'b0;
    XRAM[52846] = 8'b0;
    XRAM[52847] = 8'b0;
    XRAM[52848] = 8'b0;
    XRAM[52849] = 8'b0;
    XRAM[52850] = 8'b0;
    XRAM[52851] = 8'b0;
    XRAM[52852] = 8'b0;
    XRAM[52853] = 8'b0;
    XRAM[52854] = 8'b0;
    XRAM[52855] = 8'b0;
    XRAM[52856] = 8'b0;
    XRAM[52857] = 8'b0;
    XRAM[52858] = 8'b0;
    XRAM[52859] = 8'b0;
    XRAM[52860] = 8'b0;
    XRAM[52861] = 8'b0;
    XRAM[52862] = 8'b0;
    XRAM[52863] = 8'b0;
    XRAM[52864] = 8'b0;
    XRAM[52865] = 8'b0;
    XRAM[52866] = 8'b0;
    XRAM[52867] = 8'b0;
    XRAM[52868] = 8'b0;
    XRAM[52869] = 8'b0;
    XRAM[52870] = 8'b0;
    XRAM[52871] = 8'b0;
    XRAM[52872] = 8'b0;
    XRAM[52873] = 8'b0;
    XRAM[52874] = 8'b0;
    XRAM[52875] = 8'b0;
    XRAM[52876] = 8'b0;
    XRAM[52877] = 8'b0;
    XRAM[52878] = 8'b0;
    XRAM[52879] = 8'b0;
    XRAM[52880] = 8'b0;
    XRAM[52881] = 8'b0;
    XRAM[52882] = 8'b0;
    XRAM[52883] = 8'b0;
    XRAM[52884] = 8'b0;
    XRAM[52885] = 8'b0;
    XRAM[52886] = 8'b0;
    XRAM[52887] = 8'b0;
    XRAM[52888] = 8'b0;
    XRAM[52889] = 8'b0;
    XRAM[52890] = 8'b0;
    XRAM[52891] = 8'b0;
    XRAM[52892] = 8'b0;
    XRAM[52893] = 8'b0;
    XRAM[52894] = 8'b0;
    XRAM[52895] = 8'b0;
    XRAM[52896] = 8'b0;
    XRAM[52897] = 8'b0;
    XRAM[52898] = 8'b0;
    XRAM[52899] = 8'b0;
    XRAM[52900] = 8'b0;
    XRAM[52901] = 8'b0;
    XRAM[52902] = 8'b0;
    XRAM[52903] = 8'b0;
    XRAM[52904] = 8'b0;
    XRAM[52905] = 8'b0;
    XRAM[52906] = 8'b0;
    XRAM[52907] = 8'b0;
    XRAM[52908] = 8'b0;
    XRAM[52909] = 8'b0;
    XRAM[52910] = 8'b0;
    XRAM[52911] = 8'b0;
    XRAM[52912] = 8'b0;
    XRAM[52913] = 8'b0;
    XRAM[52914] = 8'b0;
    XRAM[52915] = 8'b0;
    XRAM[52916] = 8'b0;
    XRAM[52917] = 8'b0;
    XRAM[52918] = 8'b0;
    XRAM[52919] = 8'b0;
    XRAM[52920] = 8'b0;
    XRAM[52921] = 8'b0;
    XRAM[52922] = 8'b0;
    XRAM[52923] = 8'b0;
    XRAM[52924] = 8'b0;
    XRAM[52925] = 8'b0;
    XRAM[52926] = 8'b0;
    XRAM[52927] = 8'b0;
    XRAM[52928] = 8'b0;
    XRAM[52929] = 8'b0;
    XRAM[52930] = 8'b0;
    XRAM[52931] = 8'b0;
    XRAM[52932] = 8'b0;
    XRAM[52933] = 8'b0;
    XRAM[52934] = 8'b0;
    XRAM[52935] = 8'b0;
    XRAM[52936] = 8'b0;
    XRAM[52937] = 8'b0;
    XRAM[52938] = 8'b0;
    XRAM[52939] = 8'b0;
    XRAM[52940] = 8'b0;
    XRAM[52941] = 8'b0;
    XRAM[52942] = 8'b0;
    XRAM[52943] = 8'b0;
    XRAM[52944] = 8'b0;
    XRAM[52945] = 8'b0;
    XRAM[52946] = 8'b0;
    XRAM[52947] = 8'b0;
    XRAM[52948] = 8'b0;
    XRAM[52949] = 8'b0;
    XRAM[52950] = 8'b0;
    XRAM[52951] = 8'b0;
    XRAM[52952] = 8'b0;
    XRAM[52953] = 8'b0;
    XRAM[52954] = 8'b0;
    XRAM[52955] = 8'b0;
    XRAM[52956] = 8'b0;
    XRAM[52957] = 8'b0;
    XRAM[52958] = 8'b0;
    XRAM[52959] = 8'b0;
    XRAM[52960] = 8'b0;
    XRAM[52961] = 8'b0;
    XRAM[52962] = 8'b0;
    XRAM[52963] = 8'b0;
    XRAM[52964] = 8'b0;
    XRAM[52965] = 8'b0;
    XRAM[52966] = 8'b0;
    XRAM[52967] = 8'b0;
    XRAM[52968] = 8'b0;
    XRAM[52969] = 8'b0;
    XRAM[52970] = 8'b0;
    XRAM[52971] = 8'b0;
    XRAM[52972] = 8'b0;
    XRAM[52973] = 8'b0;
    XRAM[52974] = 8'b0;
    XRAM[52975] = 8'b0;
    XRAM[52976] = 8'b0;
    XRAM[52977] = 8'b0;
    XRAM[52978] = 8'b0;
    XRAM[52979] = 8'b0;
    XRAM[52980] = 8'b0;
    XRAM[52981] = 8'b0;
    XRAM[52982] = 8'b0;
    XRAM[52983] = 8'b0;
    XRAM[52984] = 8'b0;
    XRAM[52985] = 8'b0;
    XRAM[52986] = 8'b0;
    XRAM[52987] = 8'b0;
    XRAM[52988] = 8'b0;
    XRAM[52989] = 8'b0;
    XRAM[52990] = 8'b0;
    XRAM[52991] = 8'b0;
    XRAM[52992] = 8'b0;
    XRAM[52993] = 8'b0;
    XRAM[52994] = 8'b0;
    XRAM[52995] = 8'b0;
    XRAM[52996] = 8'b0;
    XRAM[52997] = 8'b0;
    XRAM[52998] = 8'b0;
    XRAM[52999] = 8'b0;
    XRAM[53000] = 8'b0;
    XRAM[53001] = 8'b0;
    XRAM[53002] = 8'b0;
    XRAM[53003] = 8'b0;
    XRAM[53004] = 8'b0;
    XRAM[53005] = 8'b0;
    XRAM[53006] = 8'b0;
    XRAM[53007] = 8'b0;
    XRAM[53008] = 8'b0;
    XRAM[53009] = 8'b0;
    XRAM[53010] = 8'b0;
    XRAM[53011] = 8'b0;
    XRAM[53012] = 8'b0;
    XRAM[53013] = 8'b0;
    XRAM[53014] = 8'b0;
    XRAM[53015] = 8'b0;
    XRAM[53016] = 8'b0;
    XRAM[53017] = 8'b0;
    XRAM[53018] = 8'b0;
    XRAM[53019] = 8'b0;
    XRAM[53020] = 8'b0;
    XRAM[53021] = 8'b0;
    XRAM[53022] = 8'b0;
    XRAM[53023] = 8'b0;
    XRAM[53024] = 8'b0;
    XRAM[53025] = 8'b0;
    XRAM[53026] = 8'b0;
    XRAM[53027] = 8'b0;
    XRAM[53028] = 8'b0;
    XRAM[53029] = 8'b0;
    XRAM[53030] = 8'b0;
    XRAM[53031] = 8'b0;
    XRAM[53032] = 8'b0;
    XRAM[53033] = 8'b0;
    XRAM[53034] = 8'b0;
    XRAM[53035] = 8'b0;
    XRAM[53036] = 8'b0;
    XRAM[53037] = 8'b0;
    XRAM[53038] = 8'b0;
    XRAM[53039] = 8'b0;
    XRAM[53040] = 8'b0;
    XRAM[53041] = 8'b0;
    XRAM[53042] = 8'b0;
    XRAM[53043] = 8'b0;
    XRAM[53044] = 8'b0;
    XRAM[53045] = 8'b0;
    XRAM[53046] = 8'b0;
    XRAM[53047] = 8'b0;
    XRAM[53048] = 8'b0;
    XRAM[53049] = 8'b0;
    XRAM[53050] = 8'b0;
    XRAM[53051] = 8'b0;
    XRAM[53052] = 8'b0;
    XRAM[53053] = 8'b0;
    XRAM[53054] = 8'b0;
    XRAM[53055] = 8'b0;
    XRAM[53056] = 8'b0;
    XRAM[53057] = 8'b0;
    XRAM[53058] = 8'b0;
    XRAM[53059] = 8'b0;
    XRAM[53060] = 8'b0;
    XRAM[53061] = 8'b0;
    XRAM[53062] = 8'b0;
    XRAM[53063] = 8'b0;
    XRAM[53064] = 8'b0;
    XRAM[53065] = 8'b0;
    XRAM[53066] = 8'b0;
    XRAM[53067] = 8'b0;
    XRAM[53068] = 8'b0;
    XRAM[53069] = 8'b0;
    XRAM[53070] = 8'b0;
    XRAM[53071] = 8'b0;
    XRAM[53072] = 8'b0;
    XRAM[53073] = 8'b0;
    XRAM[53074] = 8'b0;
    XRAM[53075] = 8'b0;
    XRAM[53076] = 8'b0;
    XRAM[53077] = 8'b0;
    XRAM[53078] = 8'b0;
    XRAM[53079] = 8'b0;
    XRAM[53080] = 8'b0;
    XRAM[53081] = 8'b0;
    XRAM[53082] = 8'b0;
    XRAM[53083] = 8'b0;
    XRAM[53084] = 8'b0;
    XRAM[53085] = 8'b0;
    XRAM[53086] = 8'b0;
    XRAM[53087] = 8'b0;
    XRAM[53088] = 8'b0;
    XRAM[53089] = 8'b0;
    XRAM[53090] = 8'b0;
    XRAM[53091] = 8'b0;
    XRAM[53092] = 8'b0;
    XRAM[53093] = 8'b0;
    XRAM[53094] = 8'b0;
    XRAM[53095] = 8'b0;
    XRAM[53096] = 8'b0;
    XRAM[53097] = 8'b0;
    XRAM[53098] = 8'b0;
    XRAM[53099] = 8'b0;
    XRAM[53100] = 8'b0;
    XRAM[53101] = 8'b0;
    XRAM[53102] = 8'b0;
    XRAM[53103] = 8'b0;
    XRAM[53104] = 8'b0;
    XRAM[53105] = 8'b0;
    XRAM[53106] = 8'b0;
    XRAM[53107] = 8'b0;
    XRAM[53108] = 8'b0;
    XRAM[53109] = 8'b0;
    XRAM[53110] = 8'b0;
    XRAM[53111] = 8'b0;
    XRAM[53112] = 8'b0;
    XRAM[53113] = 8'b0;
    XRAM[53114] = 8'b0;
    XRAM[53115] = 8'b0;
    XRAM[53116] = 8'b0;
    XRAM[53117] = 8'b0;
    XRAM[53118] = 8'b0;
    XRAM[53119] = 8'b0;
    XRAM[53120] = 8'b0;
    XRAM[53121] = 8'b0;
    XRAM[53122] = 8'b0;
    XRAM[53123] = 8'b0;
    XRAM[53124] = 8'b0;
    XRAM[53125] = 8'b0;
    XRAM[53126] = 8'b0;
    XRAM[53127] = 8'b0;
    XRAM[53128] = 8'b0;
    XRAM[53129] = 8'b0;
    XRAM[53130] = 8'b0;
    XRAM[53131] = 8'b0;
    XRAM[53132] = 8'b0;
    XRAM[53133] = 8'b0;
    XRAM[53134] = 8'b0;
    XRAM[53135] = 8'b0;
    XRAM[53136] = 8'b0;
    XRAM[53137] = 8'b0;
    XRAM[53138] = 8'b0;
    XRAM[53139] = 8'b0;
    XRAM[53140] = 8'b0;
    XRAM[53141] = 8'b0;
    XRAM[53142] = 8'b0;
    XRAM[53143] = 8'b0;
    XRAM[53144] = 8'b0;
    XRAM[53145] = 8'b0;
    XRAM[53146] = 8'b0;
    XRAM[53147] = 8'b0;
    XRAM[53148] = 8'b0;
    XRAM[53149] = 8'b0;
    XRAM[53150] = 8'b0;
    XRAM[53151] = 8'b0;
    XRAM[53152] = 8'b0;
    XRAM[53153] = 8'b0;
    XRAM[53154] = 8'b0;
    XRAM[53155] = 8'b0;
    XRAM[53156] = 8'b0;
    XRAM[53157] = 8'b0;
    XRAM[53158] = 8'b0;
    XRAM[53159] = 8'b0;
    XRAM[53160] = 8'b0;
    XRAM[53161] = 8'b0;
    XRAM[53162] = 8'b0;
    XRAM[53163] = 8'b0;
    XRAM[53164] = 8'b0;
    XRAM[53165] = 8'b0;
    XRAM[53166] = 8'b0;
    XRAM[53167] = 8'b0;
    XRAM[53168] = 8'b0;
    XRAM[53169] = 8'b0;
    XRAM[53170] = 8'b0;
    XRAM[53171] = 8'b0;
    XRAM[53172] = 8'b0;
    XRAM[53173] = 8'b0;
    XRAM[53174] = 8'b0;
    XRAM[53175] = 8'b0;
    XRAM[53176] = 8'b0;
    XRAM[53177] = 8'b0;
    XRAM[53178] = 8'b0;
    XRAM[53179] = 8'b0;
    XRAM[53180] = 8'b0;
    XRAM[53181] = 8'b0;
    XRAM[53182] = 8'b0;
    XRAM[53183] = 8'b0;
    XRAM[53184] = 8'b0;
    XRAM[53185] = 8'b0;
    XRAM[53186] = 8'b0;
    XRAM[53187] = 8'b0;
    XRAM[53188] = 8'b0;
    XRAM[53189] = 8'b0;
    XRAM[53190] = 8'b0;
    XRAM[53191] = 8'b0;
    XRAM[53192] = 8'b0;
    XRAM[53193] = 8'b0;
    XRAM[53194] = 8'b0;
    XRAM[53195] = 8'b0;
    XRAM[53196] = 8'b0;
    XRAM[53197] = 8'b0;
    XRAM[53198] = 8'b0;
    XRAM[53199] = 8'b0;
    XRAM[53200] = 8'b0;
    XRAM[53201] = 8'b0;
    XRAM[53202] = 8'b0;
    XRAM[53203] = 8'b0;
    XRAM[53204] = 8'b0;
    XRAM[53205] = 8'b0;
    XRAM[53206] = 8'b0;
    XRAM[53207] = 8'b0;
    XRAM[53208] = 8'b0;
    XRAM[53209] = 8'b0;
    XRAM[53210] = 8'b0;
    XRAM[53211] = 8'b0;
    XRAM[53212] = 8'b0;
    XRAM[53213] = 8'b0;
    XRAM[53214] = 8'b0;
    XRAM[53215] = 8'b0;
    XRAM[53216] = 8'b0;
    XRAM[53217] = 8'b0;
    XRAM[53218] = 8'b0;
    XRAM[53219] = 8'b0;
    XRAM[53220] = 8'b0;
    XRAM[53221] = 8'b0;
    XRAM[53222] = 8'b0;
    XRAM[53223] = 8'b0;
    XRAM[53224] = 8'b0;
    XRAM[53225] = 8'b0;
    XRAM[53226] = 8'b0;
    XRAM[53227] = 8'b0;
    XRAM[53228] = 8'b0;
    XRAM[53229] = 8'b0;
    XRAM[53230] = 8'b0;
    XRAM[53231] = 8'b0;
    XRAM[53232] = 8'b0;
    XRAM[53233] = 8'b0;
    XRAM[53234] = 8'b0;
    XRAM[53235] = 8'b0;
    XRAM[53236] = 8'b0;
    XRAM[53237] = 8'b0;
    XRAM[53238] = 8'b0;
    XRAM[53239] = 8'b0;
    XRAM[53240] = 8'b0;
    XRAM[53241] = 8'b0;
    XRAM[53242] = 8'b0;
    XRAM[53243] = 8'b0;
    XRAM[53244] = 8'b0;
    XRAM[53245] = 8'b0;
    XRAM[53246] = 8'b0;
    XRAM[53247] = 8'b0;
    XRAM[53248] = 8'b0;
    XRAM[53249] = 8'b0;
    XRAM[53250] = 8'b0;
    XRAM[53251] = 8'b0;
    XRAM[53252] = 8'b0;
    XRAM[53253] = 8'b0;
    XRAM[53254] = 8'b0;
    XRAM[53255] = 8'b0;
    XRAM[53256] = 8'b0;
    XRAM[53257] = 8'b0;
    XRAM[53258] = 8'b0;
    XRAM[53259] = 8'b0;
    XRAM[53260] = 8'b0;
    XRAM[53261] = 8'b0;
    XRAM[53262] = 8'b0;
    XRAM[53263] = 8'b0;
    XRAM[53264] = 8'b0;
    XRAM[53265] = 8'b0;
    XRAM[53266] = 8'b0;
    XRAM[53267] = 8'b0;
    XRAM[53268] = 8'b0;
    XRAM[53269] = 8'b0;
    XRAM[53270] = 8'b0;
    XRAM[53271] = 8'b0;
    XRAM[53272] = 8'b0;
    XRAM[53273] = 8'b0;
    XRAM[53274] = 8'b0;
    XRAM[53275] = 8'b0;
    XRAM[53276] = 8'b0;
    XRAM[53277] = 8'b0;
    XRAM[53278] = 8'b0;
    XRAM[53279] = 8'b0;
    XRAM[53280] = 8'b0;
    XRAM[53281] = 8'b0;
    XRAM[53282] = 8'b0;
    XRAM[53283] = 8'b0;
    XRAM[53284] = 8'b0;
    XRAM[53285] = 8'b0;
    XRAM[53286] = 8'b0;
    XRAM[53287] = 8'b0;
    XRAM[53288] = 8'b0;
    XRAM[53289] = 8'b0;
    XRAM[53290] = 8'b0;
    XRAM[53291] = 8'b0;
    XRAM[53292] = 8'b0;
    XRAM[53293] = 8'b0;
    XRAM[53294] = 8'b0;
    XRAM[53295] = 8'b0;
    XRAM[53296] = 8'b0;
    XRAM[53297] = 8'b0;
    XRAM[53298] = 8'b0;
    XRAM[53299] = 8'b0;
    XRAM[53300] = 8'b0;
    XRAM[53301] = 8'b0;
    XRAM[53302] = 8'b0;
    XRAM[53303] = 8'b0;
    XRAM[53304] = 8'b0;
    XRAM[53305] = 8'b0;
    XRAM[53306] = 8'b0;
    XRAM[53307] = 8'b0;
    XRAM[53308] = 8'b0;
    XRAM[53309] = 8'b0;
    XRAM[53310] = 8'b0;
    XRAM[53311] = 8'b0;
    XRAM[53312] = 8'b0;
    XRAM[53313] = 8'b0;
    XRAM[53314] = 8'b0;
    XRAM[53315] = 8'b0;
    XRAM[53316] = 8'b0;
    XRAM[53317] = 8'b0;
    XRAM[53318] = 8'b0;
    XRAM[53319] = 8'b0;
    XRAM[53320] = 8'b0;
    XRAM[53321] = 8'b0;
    XRAM[53322] = 8'b0;
    XRAM[53323] = 8'b0;
    XRAM[53324] = 8'b0;
    XRAM[53325] = 8'b0;
    XRAM[53326] = 8'b0;
    XRAM[53327] = 8'b0;
    XRAM[53328] = 8'b0;
    XRAM[53329] = 8'b0;
    XRAM[53330] = 8'b0;
    XRAM[53331] = 8'b0;
    XRAM[53332] = 8'b0;
    XRAM[53333] = 8'b0;
    XRAM[53334] = 8'b0;
    XRAM[53335] = 8'b0;
    XRAM[53336] = 8'b0;
    XRAM[53337] = 8'b0;
    XRAM[53338] = 8'b0;
    XRAM[53339] = 8'b0;
    XRAM[53340] = 8'b0;
    XRAM[53341] = 8'b0;
    XRAM[53342] = 8'b0;
    XRAM[53343] = 8'b0;
    XRAM[53344] = 8'b0;
    XRAM[53345] = 8'b0;
    XRAM[53346] = 8'b0;
    XRAM[53347] = 8'b0;
    XRAM[53348] = 8'b0;
    XRAM[53349] = 8'b0;
    XRAM[53350] = 8'b0;
    XRAM[53351] = 8'b0;
    XRAM[53352] = 8'b0;
    XRAM[53353] = 8'b0;
    XRAM[53354] = 8'b0;
    XRAM[53355] = 8'b0;
    XRAM[53356] = 8'b0;
    XRAM[53357] = 8'b0;
    XRAM[53358] = 8'b0;
    XRAM[53359] = 8'b0;
    XRAM[53360] = 8'b0;
    XRAM[53361] = 8'b0;
    XRAM[53362] = 8'b0;
    XRAM[53363] = 8'b0;
    XRAM[53364] = 8'b0;
    XRAM[53365] = 8'b0;
    XRAM[53366] = 8'b0;
    XRAM[53367] = 8'b0;
    XRAM[53368] = 8'b0;
    XRAM[53369] = 8'b0;
    XRAM[53370] = 8'b0;
    XRAM[53371] = 8'b0;
    XRAM[53372] = 8'b0;
    XRAM[53373] = 8'b0;
    XRAM[53374] = 8'b0;
    XRAM[53375] = 8'b0;
    XRAM[53376] = 8'b0;
    XRAM[53377] = 8'b0;
    XRAM[53378] = 8'b0;
    XRAM[53379] = 8'b0;
    XRAM[53380] = 8'b0;
    XRAM[53381] = 8'b0;
    XRAM[53382] = 8'b0;
    XRAM[53383] = 8'b0;
    XRAM[53384] = 8'b0;
    XRAM[53385] = 8'b0;
    XRAM[53386] = 8'b0;
    XRAM[53387] = 8'b0;
    XRAM[53388] = 8'b0;
    XRAM[53389] = 8'b0;
    XRAM[53390] = 8'b0;
    XRAM[53391] = 8'b0;
    XRAM[53392] = 8'b0;
    XRAM[53393] = 8'b0;
    XRAM[53394] = 8'b0;
    XRAM[53395] = 8'b0;
    XRAM[53396] = 8'b0;
    XRAM[53397] = 8'b0;
    XRAM[53398] = 8'b0;
    XRAM[53399] = 8'b0;
    XRAM[53400] = 8'b0;
    XRAM[53401] = 8'b0;
    XRAM[53402] = 8'b0;
    XRAM[53403] = 8'b0;
    XRAM[53404] = 8'b0;
    XRAM[53405] = 8'b0;
    XRAM[53406] = 8'b0;
    XRAM[53407] = 8'b0;
    XRAM[53408] = 8'b0;
    XRAM[53409] = 8'b0;
    XRAM[53410] = 8'b0;
    XRAM[53411] = 8'b0;
    XRAM[53412] = 8'b0;
    XRAM[53413] = 8'b0;
    XRAM[53414] = 8'b0;
    XRAM[53415] = 8'b0;
    XRAM[53416] = 8'b0;
    XRAM[53417] = 8'b0;
    XRAM[53418] = 8'b0;
    XRAM[53419] = 8'b0;
    XRAM[53420] = 8'b0;
    XRAM[53421] = 8'b0;
    XRAM[53422] = 8'b0;
    XRAM[53423] = 8'b0;
    XRAM[53424] = 8'b0;
    XRAM[53425] = 8'b0;
    XRAM[53426] = 8'b0;
    XRAM[53427] = 8'b0;
    XRAM[53428] = 8'b0;
    XRAM[53429] = 8'b0;
    XRAM[53430] = 8'b0;
    XRAM[53431] = 8'b0;
    XRAM[53432] = 8'b0;
    XRAM[53433] = 8'b0;
    XRAM[53434] = 8'b0;
    XRAM[53435] = 8'b0;
    XRAM[53436] = 8'b0;
    XRAM[53437] = 8'b0;
    XRAM[53438] = 8'b0;
    XRAM[53439] = 8'b0;
    XRAM[53440] = 8'b0;
    XRAM[53441] = 8'b0;
    XRAM[53442] = 8'b0;
    XRAM[53443] = 8'b0;
    XRAM[53444] = 8'b0;
    XRAM[53445] = 8'b0;
    XRAM[53446] = 8'b0;
    XRAM[53447] = 8'b0;
    XRAM[53448] = 8'b0;
    XRAM[53449] = 8'b0;
    XRAM[53450] = 8'b0;
    XRAM[53451] = 8'b0;
    XRAM[53452] = 8'b0;
    XRAM[53453] = 8'b0;
    XRAM[53454] = 8'b0;
    XRAM[53455] = 8'b0;
    XRAM[53456] = 8'b0;
    XRAM[53457] = 8'b0;
    XRAM[53458] = 8'b0;
    XRAM[53459] = 8'b0;
    XRAM[53460] = 8'b0;
    XRAM[53461] = 8'b0;
    XRAM[53462] = 8'b0;
    XRAM[53463] = 8'b0;
    XRAM[53464] = 8'b0;
    XRAM[53465] = 8'b0;
    XRAM[53466] = 8'b0;
    XRAM[53467] = 8'b0;
    XRAM[53468] = 8'b0;
    XRAM[53469] = 8'b0;
    XRAM[53470] = 8'b0;
    XRAM[53471] = 8'b0;
    XRAM[53472] = 8'b0;
    XRAM[53473] = 8'b0;
    XRAM[53474] = 8'b0;
    XRAM[53475] = 8'b0;
    XRAM[53476] = 8'b0;
    XRAM[53477] = 8'b0;
    XRAM[53478] = 8'b0;
    XRAM[53479] = 8'b0;
    XRAM[53480] = 8'b0;
    XRAM[53481] = 8'b0;
    XRAM[53482] = 8'b0;
    XRAM[53483] = 8'b0;
    XRAM[53484] = 8'b0;
    XRAM[53485] = 8'b0;
    XRAM[53486] = 8'b0;
    XRAM[53487] = 8'b0;
    XRAM[53488] = 8'b0;
    XRAM[53489] = 8'b0;
    XRAM[53490] = 8'b0;
    XRAM[53491] = 8'b0;
    XRAM[53492] = 8'b0;
    XRAM[53493] = 8'b0;
    XRAM[53494] = 8'b0;
    XRAM[53495] = 8'b0;
    XRAM[53496] = 8'b0;
    XRAM[53497] = 8'b0;
    XRAM[53498] = 8'b0;
    XRAM[53499] = 8'b0;
    XRAM[53500] = 8'b0;
    XRAM[53501] = 8'b0;
    XRAM[53502] = 8'b0;
    XRAM[53503] = 8'b0;
    XRAM[53504] = 8'b0;
    XRAM[53505] = 8'b0;
    XRAM[53506] = 8'b0;
    XRAM[53507] = 8'b0;
    XRAM[53508] = 8'b0;
    XRAM[53509] = 8'b0;
    XRAM[53510] = 8'b0;
    XRAM[53511] = 8'b0;
    XRAM[53512] = 8'b0;
    XRAM[53513] = 8'b0;
    XRAM[53514] = 8'b0;
    XRAM[53515] = 8'b0;
    XRAM[53516] = 8'b0;
    XRAM[53517] = 8'b0;
    XRAM[53518] = 8'b0;
    XRAM[53519] = 8'b0;
    XRAM[53520] = 8'b0;
    XRAM[53521] = 8'b0;
    XRAM[53522] = 8'b0;
    XRAM[53523] = 8'b0;
    XRAM[53524] = 8'b0;
    XRAM[53525] = 8'b0;
    XRAM[53526] = 8'b0;
    XRAM[53527] = 8'b0;
    XRAM[53528] = 8'b0;
    XRAM[53529] = 8'b0;
    XRAM[53530] = 8'b0;
    XRAM[53531] = 8'b0;
    XRAM[53532] = 8'b0;
    XRAM[53533] = 8'b0;
    XRAM[53534] = 8'b0;
    XRAM[53535] = 8'b0;
    XRAM[53536] = 8'b0;
    XRAM[53537] = 8'b0;
    XRAM[53538] = 8'b0;
    XRAM[53539] = 8'b0;
    XRAM[53540] = 8'b0;
    XRAM[53541] = 8'b0;
    XRAM[53542] = 8'b0;
    XRAM[53543] = 8'b0;
    XRAM[53544] = 8'b0;
    XRAM[53545] = 8'b0;
    XRAM[53546] = 8'b0;
    XRAM[53547] = 8'b0;
    XRAM[53548] = 8'b0;
    XRAM[53549] = 8'b0;
    XRAM[53550] = 8'b0;
    XRAM[53551] = 8'b0;
    XRAM[53552] = 8'b0;
    XRAM[53553] = 8'b0;
    XRAM[53554] = 8'b0;
    XRAM[53555] = 8'b0;
    XRAM[53556] = 8'b0;
    XRAM[53557] = 8'b0;
    XRAM[53558] = 8'b0;
    XRAM[53559] = 8'b0;
    XRAM[53560] = 8'b0;
    XRAM[53561] = 8'b0;
    XRAM[53562] = 8'b0;
    XRAM[53563] = 8'b0;
    XRAM[53564] = 8'b0;
    XRAM[53565] = 8'b0;
    XRAM[53566] = 8'b0;
    XRAM[53567] = 8'b0;
    XRAM[53568] = 8'b0;
    XRAM[53569] = 8'b0;
    XRAM[53570] = 8'b0;
    XRAM[53571] = 8'b0;
    XRAM[53572] = 8'b0;
    XRAM[53573] = 8'b0;
    XRAM[53574] = 8'b0;
    XRAM[53575] = 8'b0;
    XRAM[53576] = 8'b0;
    XRAM[53577] = 8'b0;
    XRAM[53578] = 8'b0;
    XRAM[53579] = 8'b0;
    XRAM[53580] = 8'b0;
    XRAM[53581] = 8'b0;
    XRAM[53582] = 8'b0;
    XRAM[53583] = 8'b0;
    XRAM[53584] = 8'b0;
    XRAM[53585] = 8'b0;
    XRAM[53586] = 8'b0;
    XRAM[53587] = 8'b0;
    XRAM[53588] = 8'b0;
    XRAM[53589] = 8'b0;
    XRAM[53590] = 8'b0;
    XRAM[53591] = 8'b0;
    XRAM[53592] = 8'b0;
    XRAM[53593] = 8'b0;
    XRAM[53594] = 8'b0;
    XRAM[53595] = 8'b0;
    XRAM[53596] = 8'b0;
    XRAM[53597] = 8'b0;
    XRAM[53598] = 8'b0;
    XRAM[53599] = 8'b0;
    XRAM[53600] = 8'b0;
    XRAM[53601] = 8'b0;
    XRAM[53602] = 8'b0;
    XRAM[53603] = 8'b0;
    XRAM[53604] = 8'b0;
    XRAM[53605] = 8'b0;
    XRAM[53606] = 8'b0;
    XRAM[53607] = 8'b0;
    XRAM[53608] = 8'b0;
    XRAM[53609] = 8'b0;
    XRAM[53610] = 8'b0;
    XRAM[53611] = 8'b0;
    XRAM[53612] = 8'b0;
    XRAM[53613] = 8'b0;
    XRAM[53614] = 8'b0;
    XRAM[53615] = 8'b0;
    XRAM[53616] = 8'b0;
    XRAM[53617] = 8'b0;
    XRAM[53618] = 8'b0;
    XRAM[53619] = 8'b0;
    XRAM[53620] = 8'b0;
    XRAM[53621] = 8'b0;
    XRAM[53622] = 8'b0;
    XRAM[53623] = 8'b0;
    XRAM[53624] = 8'b0;
    XRAM[53625] = 8'b0;
    XRAM[53626] = 8'b0;
    XRAM[53627] = 8'b0;
    XRAM[53628] = 8'b0;
    XRAM[53629] = 8'b0;
    XRAM[53630] = 8'b0;
    XRAM[53631] = 8'b0;
    XRAM[53632] = 8'b0;
    XRAM[53633] = 8'b0;
    XRAM[53634] = 8'b0;
    XRAM[53635] = 8'b0;
    XRAM[53636] = 8'b0;
    XRAM[53637] = 8'b0;
    XRAM[53638] = 8'b0;
    XRAM[53639] = 8'b0;
    XRAM[53640] = 8'b0;
    XRAM[53641] = 8'b0;
    XRAM[53642] = 8'b0;
    XRAM[53643] = 8'b0;
    XRAM[53644] = 8'b0;
    XRAM[53645] = 8'b0;
    XRAM[53646] = 8'b0;
    XRAM[53647] = 8'b0;
    XRAM[53648] = 8'b0;
    XRAM[53649] = 8'b0;
    XRAM[53650] = 8'b0;
    XRAM[53651] = 8'b0;
    XRAM[53652] = 8'b0;
    XRAM[53653] = 8'b0;
    XRAM[53654] = 8'b0;
    XRAM[53655] = 8'b0;
    XRAM[53656] = 8'b0;
    XRAM[53657] = 8'b0;
    XRAM[53658] = 8'b0;
    XRAM[53659] = 8'b0;
    XRAM[53660] = 8'b0;
    XRAM[53661] = 8'b0;
    XRAM[53662] = 8'b0;
    XRAM[53663] = 8'b0;
    XRAM[53664] = 8'b0;
    XRAM[53665] = 8'b0;
    XRAM[53666] = 8'b0;
    XRAM[53667] = 8'b0;
    XRAM[53668] = 8'b0;
    XRAM[53669] = 8'b0;
    XRAM[53670] = 8'b0;
    XRAM[53671] = 8'b0;
    XRAM[53672] = 8'b0;
    XRAM[53673] = 8'b0;
    XRAM[53674] = 8'b0;
    XRAM[53675] = 8'b0;
    XRAM[53676] = 8'b0;
    XRAM[53677] = 8'b0;
    XRAM[53678] = 8'b0;
    XRAM[53679] = 8'b0;
    XRAM[53680] = 8'b0;
    XRAM[53681] = 8'b0;
    XRAM[53682] = 8'b0;
    XRAM[53683] = 8'b0;
    XRAM[53684] = 8'b0;
    XRAM[53685] = 8'b0;
    XRAM[53686] = 8'b0;
    XRAM[53687] = 8'b0;
    XRAM[53688] = 8'b0;
    XRAM[53689] = 8'b0;
    XRAM[53690] = 8'b0;
    XRAM[53691] = 8'b0;
    XRAM[53692] = 8'b0;
    XRAM[53693] = 8'b0;
    XRAM[53694] = 8'b0;
    XRAM[53695] = 8'b0;
    XRAM[53696] = 8'b0;
    XRAM[53697] = 8'b0;
    XRAM[53698] = 8'b0;
    XRAM[53699] = 8'b0;
    XRAM[53700] = 8'b0;
    XRAM[53701] = 8'b0;
    XRAM[53702] = 8'b0;
    XRAM[53703] = 8'b0;
    XRAM[53704] = 8'b0;
    XRAM[53705] = 8'b0;
    XRAM[53706] = 8'b0;
    XRAM[53707] = 8'b0;
    XRAM[53708] = 8'b0;
    XRAM[53709] = 8'b0;
    XRAM[53710] = 8'b0;
    XRAM[53711] = 8'b0;
    XRAM[53712] = 8'b0;
    XRAM[53713] = 8'b0;
    XRAM[53714] = 8'b0;
    XRAM[53715] = 8'b0;
    XRAM[53716] = 8'b0;
    XRAM[53717] = 8'b0;
    XRAM[53718] = 8'b0;
    XRAM[53719] = 8'b0;
    XRAM[53720] = 8'b0;
    XRAM[53721] = 8'b0;
    XRAM[53722] = 8'b0;
    XRAM[53723] = 8'b0;
    XRAM[53724] = 8'b0;
    XRAM[53725] = 8'b0;
    XRAM[53726] = 8'b0;
    XRAM[53727] = 8'b0;
    XRAM[53728] = 8'b0;
    XRAM[53729] = 8'b0;
    XRAM[53730] = 8'b0;
    XRAM[53731] = 8'b0;
    XRAM[53732] = 8'b0;
    XRAM[53733] = 8'b0;
    XRAM[53734] = 8'b0;
    XRAM[53735] = 8'b0;
    XRAM[53736] = 8'b0;
    XRAM[53737] = 8'b0;
    XRAM[53738] = 8'b0;
    XRAM[53739] = 8'b0;
    XRAM[53740] = 8'b0;
    XRAM[53741] = 8'b0;
    XRAM[53742] = 8'b0;
    XRAM[53743] = 8'b0;
    XRAM[53744] = 8'b0;
    XRAM[53745] = 8'b0;
    XRAM[53746] = 8'b0;
    XRAM[53747] = 8'b0;
    XRAM[53748] = 8'b0;
    XRAM[53749] = 8'b0;
    XRAM[53750] = 8'b0;
    XRAM[53751] = 8'b0;
    XRAM[53752] = 8'b0;
    XRAM[53753] = 8'b0;
    XRAM[53754] = 8'b0;
    XRAM[53755] = 8'b0;
    XRAM[53756] = 8'b0;
    XRAM[53757] = 8'b0;
    XRAM[53758] = 8'b0;
    XRAM[53759] = 8'b0;
    XRAM[53760] = 8'b0;
    XRAM[53761] = 8'b0;
    XRAM[53762] = 8'b0;
    XRAM[53763] = 8'b0;
    XRAM[53764] = 8'b0;
    XRAM[53765] = 8'b0;
    XRAM[53766] = 8'b0;
    XRAM[53767] = 8'b0;
    XRAM[53768] = 8'b0;
    XRAM[53769] = 8'b0;
    XRAM[53770] = 8'b0;
    XRAM[53771] = 8'b0;
    XRAM[53772] = 8'b0;
    XRAM[53773] = 8'b0;
    XRAM[53774] = 8'b0;
    XRAM[53775] = 8'b0;
    XRAM[53776] = 8'b0;
    XRAM[53777] = 8'b0;
    XRAM[53778] = 8'b0;
    XRAM[53779] = 8'b0;
    XRAM[53780] = 8'b0;
    XRAM[53781] = 8'b0;
    XRAM[53782] = 8'b0;
    XRAM[53783] = 8'b0;
    XRAM[53784] = 8'b0;
    XRAM[53785] = 8'b0;
    XRAM[53786] = 8'b0;
    XRAM[53787] = 8'b0;
    XRAM[53788] = 8'b0;
    XRAM[53789] = 8'b0;
    XRAM[53790] = 8'b0;
    XRAM[53791] = 8'b0;
    XRAM[53792] = 8'b0;
    XRAM[53793] = 8'b0;
    XRAM[53794] = 8'b0;
    XRAM[53795] = 8'b0;
    XRAM[53796] = 8'b0;
    XRAM[53797] = 8'b0;
    XRAM[53798] = 8'b0;
    XRAM[53799] = 8'b0;
    XRAM[53800] = 8'b0;
    XRAM[53801] = 8'b0;
    XRAM[53802] = 8'b0;
    XRAM[53803] = 8'b0;
    XRAM[53804] = 8'b0;
    XRAM[53805] = 8'b0;
    XRAM[53806] = 8'b0;
    XRAM[53807] = 8'b0;
    XRAM[53808] = 8'b0;
    XRAM[53809] = 8'b0;
    XRAM[53810] = 8'b0;
    XRAM[53811] = 8'b0;
    XRAM[53812] = 8'b0;
    XRAM[53813] = 8'b0;
    XRAM[53814] = 8'b0;
    XRAM[53815] = 8'b0;
    XRAM[53816] = 8'b0;
    XRAM[53817] = 8'b0;
    XRAM[53818] = 8'b0;
    XRAM[53819] = 8'b0;
    XRAM[53820] = 8'b0;
    XRAM[53821] = 8'b0;
    XRAM[53822] = 8'b0;
    XRAM[53823] = 8'b0;
    XRAM[53824] = 8'b0;
    XRAM[53825] = 8'b0;
    XRAM[53826] = 8'b0;
    XRAM[53827] = 8'b0;
    XRAM[53828] = 8'b0;
    XRAM[53829] = 8'b0;
    XRAM[53830] = 8'b0;
    XRAM[53831] = 8'b0;
    XRAM[53832] = 8'b0;
    XRAM[53833] = 8'b0;
    XRAM[53834] = 8'b0;
    XRAM[53835] = 8'b0;
    XRAM[53836] = 8'b0;
    XRAM[53837] = 8'b0;
    XRAM[53838] = 8'b0;
    XRAM[53839] = 8'b0;
    XRAM[53840] = 8'b0;
    XRAM[53841] = 8'b0;
    XRAM[53842] = 8'b0;
    XRAM[53843] = 8'b0;
    XRAM[53844] = 8'b0;
    XRAM[53845] = 8'b0;
    XRAM[53846] = 8'b0;
    XRAM[53847] = 8'b0;
    XRAM[53848] = 8'b0;
    XRAM[53849] = 8'b0;
    XRAM[53850] = 8'b0;
    XRAM[53851] = 8'b0;
    XRAM[53852] = 8'b0;
    XRAM[53853] = 8'b0;
    XRAM[53854] = 8'b0;
    XRAM[53855] = 8'b0;
    XRAM[53856] = 8'b0;
    XRAM[53857] = 8'b0;
    XRAM[53858] = 8'b0;
    XRAM[53859] = 8'b0;
    XRAM[53860] = 8'b0;
    XRAM[53861] = 8'b0;
    XRAM[53862] = 8'b0;
    XRAM[53863] = 8'b0;
    XRAM[53864] = 8'b0;
    XRAM[53865] = 8'b0;
    XRAM[53866] = 8'b0;
    XRAM[53867] = 8'b0;
    XRAM[53868] = 8'b0;
    XRAM[53869] = 8'b0;
    XRAM[53870] = 8'b0;
    XRAM[53871] = 8'b0;
    XRAM[53872] = 8'b0;
    XRAM[53873] = 8'b0;
    XRAM[53874] = 8'b0;
    XRAM[53875] = 8'b0;
    XRAM[53876] = 8'b0;
    XRAM[53877] = 8'b0;
    XRAM[53878] = 8'b0;
    XRAM[53879] = 8'b0;
    XRAM[53880] = 8'b0;
    XRAM[53881] = 8'b0;
    XRAM[53882] = 8'b0;
    XRAM[53883] = 8'b0;
    XRAM[53884] = 8'b0;
    XRAM[53885] = 8'b0;
    XRAM[53886] = 8'b0;
    XRAM[53887] = 8'b0;
    XRAM[53888] = 8'b0;
    XRAM[53889] = 8'b0;
    XRAM[53890] = 8'b0;
    XRAM[53891] = 8'b0;
    XRAM[53892] = 8'b0;
    XRAM[53893] = 8'b0;
    XRAM[53894] = 8'b0;
    XRAM[53895] = 8'b0;
    XRAM[53896] = 8'b0;
    XRAM[53897] = 8'b0;
    XRAM[53898] = 8'b0;
    XRAM[53899] = 8'b0;
    XRAM[53900] = 8'b0;
    XRAM[53901] = 8'b0;
    XRAM[53902] = 8'b0;
    XRAM[53903] = 8'b0;
    XRAM[53904] = 8'b0;
    XRAM[53905] = 8'b0;
    XRAM[53906] = 8'b0;
    XRAM[53907] = 8'b0;
    XRAM[53908] = 8'b0;
    XRAM[53909] = 8'b0;
    XRAM[53910] = 8'b0;
    XRAM[53911] = 8'b0;
    XRAM[53912] = 8'b0;
    XRAM[53913] = 8'b0;
    XRAM[53914] = 8'b0;
    XRAM[53915] = 8'b0;
    XRAM[53916] = 8'b0;
    XRAM[53917] = 8'b0;
    XRAM[53918] = 8'b0;
    XRAM[53919] = 8'b0;
    XRAM[53920] = 8'b0;
    XRAM[53921] = 8'b0;
    XRAM[53922] = 8'b0;
    XRAM[53923] = 8'b0;
    XRAM[53924] = 8'b0;
    XRAM[53925] = 8'b0;
    XRAM[53926] = 8'b0;
    XRAM[53927] = 8'b0;
    XRAM[53928] = 8'b0;
    XRAM[53929] = 8'b0;
    XRAM[53930] = 8'b0;
    XRAM[53931] = 8'b0;
    XRAM[53932] = 8'b0;
    XRAM[53933] = 8'b0;
    XRAM[53934] = 8'b0;
    XRAM[53935] = 8'b0;
    XRAM[53936] = 8'b0;
    XRAM[53937] = 8'b0;
    XRAM[53938] = 8'b0;
    XRAM[53939] = 8'b0;
    XRAM[53940] = 8'b0;
    XRAM[53941] = 8'b0;
    XRAM[53942] = 8'b0;
    XRAM[53943] = 8'b0;
    XRAM[53944] = 8'b0;
    XRAM[53945] = 8'b0;
    XRAM[53946] = 8'b0;
    XRAM[53947] = 8'b0;
    XRAM[53948] = 8'b0;
    XRAM[53949] = 8'b0;
    XRAM[53950] = 8'b0;
    XRAM[53951] = 8'b0;
    XRAM[53952] = 8'b0;
    XRAM[53953] = 8'b0;
    XRAM[53954] = 8'b0;
    XRAM[53955] = 8'b0;
    XRAM[53956] = 8'b0;
    XRAM[53957] = 8'b0;
    XRAM[53958] = 8'b0;
    XRAM[53959] = 8'b0;
    XRAM[53960] = 8'b0;
    XRAM[53961] = 8'b0;
    XRAM[53962] = 8'b0;
    XRAM[53963] = 8'b0;
    XRAM[53964] = 8'b0;
    XRAM[53965] = 8'b0;
    XRAM[53966] = 8'b0;
    XRAM[53967] = 8'b0;
    XRAM[53968] = 8'b0;
    XRAM[53969] = 8'b0;
    XRAM[53970] = 8'b0;
    XRAM[53971] = 8'b0;
    XRAM[53972] = 8'b0;
    XRAM[53973] = 8'b0;
    XRAM[53974] = 8'b0;
    XRAM[53975] = 8'b0;
    XRAM[53976] = 8'b0;
    XRAM[53977] = 8'b0;
    XRAM[53978] = 8'b0;
    XRAM[53979] = 8'b0;
    XRAM[53980] = 8'b0;
    XRAM[53981] = 8'b0;
    XRAM[53982] = 8'b0;
    XRAM[53983] = 8'b0;
    XRAM[53984] = 8'b0;
    XRAM[53985] = 8'b0;
    XRAM[53986] = 8'b0;
    XRAM[53987] = 8'b0;
    XRAM[53988] = 8'b0;
    XRAM[53989] = 8'b0;
    XRAM[53990] = 8'b0;
    XRAM[53991] = 8'b0;
    XRAM[53992] = 8'b0;
    XRAM[53993] = 8'b0;
    XRAM[53994] = 8'b0;
    XRAM[53995] = 8'b0;
    XRAM[53996] = 8'b0;
    XRAM[53997] = 8'b0;
    XRAM[53998] = 8'b0;
    XRAM[53999] = 8'b0;
    XRAM[54000] = 8'b0;
    XRAM[54001] = 8'b0;
    XRAM[54002] = 8'b0;
    XRAM[54003] = 8'b0;
    XRAM[54004] = 8'b0;
    XRAM[54005] = 8'b0;
    XRAM[54006] = 8'b0;
    XRAM[54007] = 8'b0;
    XRAM[54008] = 8'b0;
    XRAM[54009] = 8'b0;
    XRAM[54010] = 8'b0;
    XRAM[54011] = 8'b0;
    XRAM[54012] = 8'b0;
    XRAM[54013] = 8'b0;
    XRAM[54014] = 8'b0;
    XRAM[54015] = 8'b0;
    XRAM[54016] = 8'b0;
    XRAM[54017] = 8'b0;
    XRAM[54018] = 8'b0;
    XRAM[54019] = 8'b0;
    XRAM[54020] = 8'b0;
    XRAM[54021] = 8'b0;
    XRAM[54022] = 8'b0;
    XRAM[54023] = 8'b0;
    XRAM[54024] = 8'b0;
    XRAM[54025] = 8'b0;
    XRAM[54026] = 8'b0;
    XRAM[54027] = 8'b0;
    XRAM[54028] = 8'b0;
    XRAM[54029] = 8'b0;
    XRAM[54030] = 8'b0;
    XRAM[54031] = 8'b0;
    XRAM[54032] = 8'b0;
    XRAM[54033] = 8'b0;
    XRAM[54034] = 8'b0;
    XRAM[54035] = 8'b0;
    XRAM[54036] = 8'b0;
    XRAM[54037] = 8'b0;
    XRAM[54038] = 8'b0;
    XRAM[54039] = 8'b0;
    XRAM[54040] = 8'b0;
    XRAM[54041] = 8'b0;
    XRAM[54042] = 8'b0;
    XRAM[54043] = 8'b0;
    XRAM[54044] = 8'b0;
    XRAM[54045] = 8'b0;
    XRAM[54046] = 8'b0;
    XRAM[54047] = 8'b0;
    XRAM[54048] = 8'b0;
    XRAM[54049] = 8'b0;
    XRAM[54050] = 8'b0;
    XRAM[54051] = 8'b0;
    XRAM[54052] = 8'b0;
    XRAM[54053] = 8'b0;
    XRAM[54054] = 8'b0;
    XRAM[54055] = 8'b0;
    XRAM[54056] = 8'b0;
    XRAM[54057] = 8'b0;
    XRAM[54058] = 8'b0;
    XRAM[54059] = 8'b0;
    XRAM[54060] = 8'b0;
    XRAM[54061] = 8'b0;
    XRAM[54062] = 8'b0;
    XRAM[54063] = 8'b0;
    XRAM[54064] = 8'b0;
    XRAM[54065] = 8'b0;
    XRAM[54066] = 8'b0;
    XRAM[54067] = 8'b0;
    XRAM[54068] = 8'b0;
    XRAM[54069] = 8'b0;
    XRAM[54070] = 8'b0;
    XRAM[54071] = 8'b0;
    XRAM[54072] = 8'b0;
    XRAM[54073] = 8'b0;
    XRAM[54074] = 8'b0;
    XRAM[54075] = 8'b0;
    XRAM[54076] = 8'b0;
    XRAM[54077] = 8'b0;
    XRAM[54078] = 8'b0;
    XRAM[54079] = 8'b0;
    XRAM[54080] = 8'b0;
    XRAM[54081] = 8'b0;
    XRAM[54082] = 8'b0;
    XRAM[54083] = 8'b0;
    XRAM[54084] = 8'b0;
    XRAM[54085] = 8'b0;
    XRAM[54086] = 8'b0;
    XRAM[54087] = 8'b0;
    XRAM[54088] = 8'b0;
    XRAM[54089] = 8'b0;
    XRAM[54090] = 8'b0;
    XRAM[54091] = 8'b0;
    XRAM[54092] = 8'b0;
    XRAM[54093] = 8'b0;
    XRAM[54094] = 8'b0;
    XRAM[54095] = 8'b0;
    XRAM[54096] = 8'b0;
    XRAM[54097] = 8'b0;
    XRAM[54098] = 8'b0;
    XRAM[54099] = 8'b0;
    XRAM[54100] = 8'b0;
    XRAM[54101] = 8'b0;
    XRAM[54102] = 8'b0;
    XRAM[54103] = 8'b0;
    XRAM[54104] = 8'b0;
    XRAM[54105] = 8'b0;
    XRAM[54106] = 8'b0;
    XRAM[54107] = 8'b0;
    XRAM[54108] = 8'b0;
    XRAM[54109] = 8'b0;
    XRAM[54110] = 8'b0;
    XRAM[54111] = 8'b0;
    XRAM[54112] = 8'b0;
    XRAM[54113] = 8'b0;
    XRAM[54114] = 8'b0;
    XRAM[54115] = 8'b0;
    XRAM[54116] = 8'b0;
    XRAM[54117] = 8'b0;
    XRAM[54118] = 8'b0;
    XRAM[54119] = 8'b0;
    XRAM[54120] = 8'b0;
    XRAM[54121] = 8'b0;
    XRAM[54122] = 8'b0;
    XRAM[54123] = 8'b0;
    XRAM[54124] = 8'b0;
    XRAM[54125] = 8'b0;
    XRAM[54126] = 8'b0;
    XRAM[54127] = 8'b0;
    XRAM[54128] = 8'b0;
    XRAM[54129] = 8'b0;
    XRAM[54130] = 8'b0;
    XRAM[54131] = 8'b0;
    XRAM[54132] = 8'b0;
    XRAM[54133] = 8'b0;
    XRAM[54134] = 8'b0;
    XRAM[54135] = 8'b0;
    XRAM[54136] = 8'b0;
    XRAM[54137] = 8'b0;
    XRAM[54138] = 8'b0;
    XRAM[54139] = 8'b0;
    XRAM[54140] = 8'b0;
    XRAM[54141] = 8'b0;
    XRAM[54142] = 8'b0;
    XRAM[54143] = 8'b0;
    XRAM[54144] = 8'b0;
    XRAM[54145] = 8'b0;
    XRAM[54146] = 8'b0;
    XRAM[54147] = 8'b0;
    XRAM[54148] = 8'b0;
    XRAM[54149] = 8'b0;
    XRAM[54150] = 8'b0;
    XRAM[54151] = 8'b0;
    XRAM[54152] = 8'b0;
    XRAM[54153] = 8'b0;
    XRAM[54154] = 8'b0;
    XRAM[54155] = 8'b0;
    XRAM[54156] = 8'b0;
    XRAM[54157] = 8'b0;
    XRAM[54158] = 8'b0;
    XRAM[54159] = 8'b0;
    XRAM[54160] = 8'b0;
    XRAM[54161] = 8'b0;
    XRAM[54162] = 8'b0;
    XRAM[54163] = 8'b0;
    XRAM[54164] = 8'b0;
    XRAM[54165] = 8'b0;
    XRAM[54166] = 8'b0;
    XRAM[54167] = 8'b0;
    XRAM[54168] = 8'b0;
    XRAM[54169] = 8'b0;
    XRAM[54170] = 8'b0;
    XRAM[54171] = 8'b0;
    XRAM[54172] = 8'b0;
    XRAM[54173] = 8'b0;
    XRAM[54174] = 8'b0;
    XRAM[54175] = 8'b0;
    XRAM[54176] = 8'b0;
    XRAM[54177] = 8'b0;
    XRAM[54178] = 8'b0;
    XRAM[54179] = 8'b0;
    XRAM[54180] = 8'b0;
    XRAM[54181] = 8'b0;
    XRAM[54182] = 8'b0;
    XRAM[54183] = 8'b0;
    XRAM[54184] = 8'b0;
    XRAM[54185] = 8'b0;
    XRAM[54186] = 8'b0;
    XRAM[54187] = 8'b0;
    XRAM[54188] = 8'b0;
    XRAM[54189] = 8'b0;
    XRAM[54190] = 8'b0;
    XRAM[54191] = 8'b0;
    XRAM[54192] = 8'b0;
    XRAM[54193] = 8'b0;
    XRAM[54194] = 8'b0;
    XRAM[54195] = 8'b0;
    XRAM[54196] = 8'b0;
    XRAM[54197] = 8'b0;
    XRAM[54198] = 8'b0;
    XRAM[54199] = 8'b0;
    XRAM[54200] = 8'b0;
    XRAM[54201] = 8'b0;
    XRAM[54202] = 8'b0;
    XRAM[54203] = 8'b0;
    XRAM[54204] = 8'b0;
    XRAM[54205] = 8'b0;
    XRAM[54206] = 8'b0;
    XRAM[54207] = 8'b0;
    XRAM[54208] = 8'b0;
    XRAM[54209] = 8'b0;
    XRAM[54210] = 8'b0;
    XRAM[54211] = 8'b0;
    XRAM[54212] = 8'b0;
    XRAM[54213] = 8'b0;
    XRAM[54214] = 8'b0;
    XRAM[54215] = 8'b0;
    XRAM[54216] = 8'b0;
    XRAM[54217] = 8'b0;
    XRAM[54218] = 8'b0;
    XRAM[54219] = 8'b0;
    XRAM[54220] = 8'b0;
    XRAM[54221] = 8'b0;
    XRAM[54222] = 8'b0;
    XRAM[54223] = 8'b0;
    XRAM[54224] = 8'b0;
    XRAM[54225] = 8'b0;
    XRAM[54226] = 8'b0;
    XRAM[54227] = 8'b0;
    XRAM[54228] = 8'b0;
    XRAM[54229] = 8'b0;
    XRAM[54230] = 8'b0;
    XRAM[54231] = 8'b0;
    XRAM[54232] = 8'b0;
    XRAM[54233] = 8'b0;
    XRAM[54234] = 8'b0;
    XRAM[54235] = 8'b0;
    XRAM[54236] = 8'b0;
    XRAM[54237] = 8'b0;
    XRAM[54238] = 8'b0;
    XRAM[54239] = 8'b0;
    XRAM[54240] = 8'b0;
    XRAM[54241] = 8'b0;
    XRAM[54242] = 8'b0;
    XRAM[54243] = 8'b0;
    XRAM[54244] = 8'b0;
    XRAM[54245] = 8'b0;
    XRAM[54246] = 8'b0;
    XRAM[54247] = 8'b0;
    XRAM[54248] = 8'b0;
    XRAM[54249] = 8'b0;
    XRAM[54250] = 8'b0;
    XRAM[54251] = 8'b0;
    XRAM[54252] = 8'b0;
    XRAM[54253] = 8'b0;
    XRAM[54254] = 8'b0;
    XRAM[54255] = 8'b0;
    XRAM[54256] = 8'b0;
    XRAM[54257] = 8'b0;
    XRAM[54258] = 8'b0;
    XRAM[54259] = 8'b0;
    XRAM[54260] = 8'b0;
    XRAM[54261] = 8'b0;
    XRAM[54262] = 8'b0;
    XRAM[54263] = 8'b0;
    XRAM[54264] = 8'b0;
    XRAM[54265] = 8'b0;
    XRAM[54266] = 8'b0;
    XRAM[54267] = 8'b0;
    XRAM[54268] = 8'b0;
    XRAM[54269] = 8'b0;
    XRAM[54270] = 8'b0;
    XRAM[54271] = 8'b0;
    XRAM[54272] = 8'b0;
    XRAM[54273] = 8'b0;
    XRAM[54274] = 8'b0;
    XRAM[54275] = 8'b0;
    XRAM[54276] = 8'b0;
    XRAM[54277] = 8'b0;
    XRAM[54278] = 8'b0;
    XRAM[54279] = 8'b0;
    XRAM[54280] = 8'b0;
    XRAM[54281] = 8'b0;
    XRAM[54282] = 8'b0;
    XRAM[54283] = 8'b0;
    XRAM[54284] = 8'b0;
    XRAM[54285] = 8'b0;
    XRAM[54286] = 8'b0;
    XRAM[54287] = 8'b0;
    XRAM[54288] = 8'b0;
    XRAM[54289] = 8'b0;
    XRAM[54290] = 8'b0;
    XRAM[54291] = 8'b0;
    XRAM[54292] = 8'b0;
    XRAM[54293] = 8'b0;
    XRAM[54294] = 8'b0;
    XRAM[54295] = 8'b0;
    XRAM[54296] = 8'b0;
    XRAM[54297] = 8'b0;
    XRAM[54298] = 8'b0;
    XRAM[54299] = 8'b0;
    XRAM[54300] = 8'b0;
    XRAM[54301] = 8'b0;
    XRAM[54302] = 8'b0;
    XRAM[54303] = 8'b0;
    XRAM[54304] = 8'b0;
    XRAM[54305] = 8'b0;
    XRAM[54306] = 8'b0;
    XRAM[54307] = 8'b0;
    XRAM[54308] = 8'b0;
    XRAM[54309] = 8'b0;
    XRAM[54310] = 8'b0;
    XRAM[54311] = 8'b0;
    XRAM[54312] = 8'b0;
    XRAM[54313] = 8'b0;
    XRAM[54314] = 8'b0;
    XRAM[54315] = 8'b0;
    XRAM[54316] = 8'b0;
    XRAM[54317] = 8'b0;
    XRAM[54318] = 8'b0;
    XRAM[54319] = 8'b0;
    XRAM[54320] = 8'b0;
    XRAM[54321] = 8'b0;
    XRAM[54322] = 8'b0;
    XRAM[54323] = 8'b0;
    XRAM[54324] = 8'b0;
    XRAM[54325] = 8'b0;
    XRAM[54326] = 8'b0;
    XRAM[54327] = 8'b0;
    XRAM[54328] = 8'b0;
    XRAM[54329] = 8'b0;
    XRAM[54330] = 8'b0;
    XRAM[54331] = 8'b0;
    XRAM[54332] = 8'b0;
    XRAM[54333] = 8'b0;
    XRAM[54334] = 8'b0;
    XRAM[54335] = 8'b0;
    XRAM[54336] = 8'b0;
    XRAM[54337] = 8'b0;
    XRAM[54338] = 8'b0;
    XRAM[54339] = 8'b0;
    XRAM[54340] = 8'b0;
    XRAM[54341] = 8'b0;
    XRAM[54342] = 8'b0;
    XRAM[54343] = 8'b0;
    XRAM[54344] = 8'b0;
    XRAM[54345] = 8'b0;
    XRAM[54346] = 8'b0;
    XRAM[54347] = 8'b0;
    XRAM[54348] = 8'b0;
    XRAM[54349] = 8'b0;
    XRAM[54350] = 8'b0;
    XRAM[54351] = 8'b0;
    XRAM[54352] = 8'b0;
    XRAM[54353] = 8'b0;
    XRAM[54354] = 8'b0;
    XRAM[54355] = 8'b0;
    XRAM[54356] = 8'b0;
    XRAM[54357] = 8'b0;
    XRAM[54358] = 8'b0;
    XRAM[54359] = 8'b0;
    XRAM[54360] = 8'b0;
    XRAM[54361] = 8'b0;
    XRAM[54362] = 8'b0;
    XRAM[54363] = 8'b0;
    XRAM[54364] = 8'b0;
    XRAM[54365] = 8'b0;
    XRAM[54366] = 8'b0;
    XRAM[54367] = 8'b0;
    XRAM[54368] = 8'b0;
    XRAM[54369] = 8'b0;
    XRAM[54370] = 8'b0;
    XRAM[54371] = 8'b0;
    XRAM[54372] = 8'b0;
    XRAM[54373] = 8'b0;
    XRAM[54374] = 8'b0;
    XRAM[54375] = 8'b0;
    XRAM[54376] = 8'b0;
    XRAM[54377] = 8'b0;
    XRAM[54378] = 8'b0;
    XRAM[54379] = 8'b0;
    XRAM[54380] = 8'b0;
    XRAM[54381] = 8'b0;
    XRAM[54382] = 8'b0;
    XRAM[54383] = 8'b0;
    XRAM[54384] = 8'b0;
    XRAM[54385] = 8'b0;
    XRAM[54386] = 8'b0;
    XRAM[54387] = 8'b0;
    XRAM[54388] = 8'b0;
    XRAM[54389] = 8'b0;
    XRAM[54390] = 8'b0;
    XRAM[54391] = 8'b0;
    XRAM[54392] = 8'b0;
    XRAM[54393] = 8'b0;
    XRAM[54394] = 8'b0;
    XRAM[54395] = 8'b0;
    XRAM[54396] = 8'b0;
    XRAM[54397] = 8'b0;
    XRAM[54398] = 8'b0;
    XRAM[54399] = 8'b0;
    XRAM[54400] = 8'b0;
    XRAM[54401] = 8'b0;
    XRAM[54402] = 8'b0;
    XRAM[54403] = 8'b0;
    XRAM[54404] = 8'b0;
    XRAM[54405] = 8'b0;
    XRAM[54406] = 8'b0;
    XRAM[54407] = 8'b0;
    XRAM[54408] = 8'b0;
    XRAM[54409] = 8'b0;
    XRAM[54410] = 8'b0;
    XRAM[54411] = 8'b0;
    XRAM[54412] = 8'b0;
    XRAM[54413] = 8'b0;
    XRAM[54414] = 8'b0;
    XRAM[54415] = 8'b0;
    XRAM[54416] = 8'b0;
    XRAM[54417] = 8'b0;
    XRAM[54418] = 8'b0;
    XRAM[54419] = 8'b0;
    XRAM[54420] = 8'b0;
    XRAM[54421] = 8'b0;
    XRAM[54422] = 8'b0;
    XRAM[54423] = 8'b0;
    XRAM[54424] = 8'b0;
    XRAM[54425] = 8'b0;
    XRAM[54426] = 8'b0;
    XRAM[54427] = 8'b0;
    XRAM[54428] = 8'b0;
    XRAM[54429] = 8'b0;
    XRAM[54430] = 8'b0;
    XRAM[54431] = 8'b0;
    XRAM[54432] = 8'b0;
    XRAM[54433] = 8'b0;
    XRAM[54434] = 8'b0;
    XRAM[54435] = 8'b0;
    XRAM[54436] = 8'b0;
    XRAM[54437] = 8'b0;
    XRAM[54438] = 8'b0;
    XRAM[54439] = 8'b0;
    XRAM[54440] = 8'b0;
    XRAM[54441] = 8'b0;
    XRAM[54442] = 8'b0;
    XRAM[54443] = 8'b0;
    XRAM[54444] = 8'b0;
    XRAM[54445] = 8'b0;
    XRAM[54446] = 8'b0;
    XRAM[54447] = 8'b0;
    XRAM[54448] = 8'b0;
    XRAM[54449] = 8'b0;
    XRAM[54450] = 8'b0;
    XRAM[54451] = 8'b0;
    XRAM[54452] = 8'b0;
    XRAM[54453] = 8'b0;
    XRAM[54454] = 8'b0;
    XRAM[54455] = 8'b0;
    XRAM[54456] = 8'b0;
    XRAM[54457] = 8'b0;
    XRAM[54458] = 8'b0;
    XRAM[54459] = 8'b0;
    XRAM[54460] = 8'b0;
    XRAM[54461] = 8'b0;
    XRAM[54462] = 8'b0;
    XRAM[54463] = 8'b0;
    XRAM[54464] = 8'b0;
    XRAM[54465] = 8'b0;
    XRAM[54466] = 8'b0;
    XRAM[54467] = 8'b0;
    XRAM[54468] = 8'b0;
    XRAM[54469] = 8'b0;
    XRAM[54470] = 8'b0;
    XRAM[54471] = 8'b0;
    XRAM[54472] = 8'b0;
    XRAM[54473] = 8'b0;
    XRAM[54474] = 8'b0;
    XRAM[54475] = 8'b0;
    XRAM[54476] = 8'b0;
    XRAM[54477] = 8'b0;
    XRAM[54478] = 8'b0;
    XRAM[54479] = 8'b0;
    XRAM[54480] = 8'b0;
    XRAM[54481] = 8'b0;
    XRAM[54482] = 8'b0;
    XRAM[54483] = 8'b0;
    XRAM[54484] = 8'b0;
    XRAM[54485] = 8'b0;
    XRAM[54486] = 8'b0;
    XRAM[54487] = 8'b0;
    XRAM[54488] = 8'b0;
    XRAM[54489] = 8'b0;
    XRAM[54490] = 8'b0;
    XRAM[54491] = 8'b0;
    XRAM[54492] = 8'b0;
    XRAM[54493] = 8'b0;
    XRAM[54494] = 8'b0;
    XRAM[54495] = 8'b0;
    XRAM[54496] = 8'b0;
    XRAM[54497] = 8'b0;
    XRAM[54498] = 8'b0;
    XRAM[54499] = 8'b0;
    XRAM[54500] = 8'b0;
    XRAM[54501] = 8'b0;
    XRAM[54502] = 8'b0;
    XRAM[54503] = 8'b0;
    XRAM[54504] = 8'b0;
    XRAM[54505] = 8'b0;
    XRAM[54506] = 8'b0;
    XRAM[54507] = 8'b0;
    XRAM[54508] = 8'b0;
    XRAM[54509] = 8'b0;
    XRAM[54510] = 8'b0;
    XRAM[54511] = 8'b0;
    XRAM[54512] = 8'b0;
    XRAM[54513] = 8'b0;
    XRAM[54514] = 8'b0;
    XRAM[54515] = 8'b0;
    XRAM[54516] = 8'b0;
    XRAM[54517] = 8'b0;
    XRAM[54518] = 8'b0;
    XRAM[54519] = 8'b0;
    XRAM[54520] = 8'b0;
    XRAM[54521] = 8'b0;
    XRAM[54522] = 8'b0;
    XRAM[54523] = 8'b0;
    XRAM[54524] = 8'b0;
    XRAM[54525] = 8'b0;
    XRAM[54526] = 8'b0;
    XRAM[54527] = 8'b0;
    XRAM[54528] = 8'b0;
    XRAM[54529] = 8'b0;
    XRAM[54530] = 8'b0;
    XRAM[54531] = 8'b0;
    XRAM[54532] = 8'b0;
    XRAM[54533] = 8'b0;
    XRAM[54534] = 8'b0;
    XRAM[54535] = 8'b0;
    XRAM[54536] = 8'b0;
    XRAM[54537] = 8'b0;
    XRAM[54538] = 8'b0;
    XRAM[54539] = 8'b0;
    XRAM[54540] = 8'b0;
    XRAM[54541] = 8'b0;
    XRAM[54542] = 8'b0;
    XRAM[54543] = 8'b0;
    XRAM[54544] = 8'b0;
    XRAM[54545] = 8'b0;
    XRAM[54546] = 8'b0;
    XRAM[54547] = 8'b0;
    XRAM[54548] = 8'b0;
    XRAM[54549] = 8'b0;
    XRAM[54550] = 8'b0;
    XRAM[54551] = 8'b0;
    XRAM[54552] = 8'b0;
    XRAM[54553] = 8'b0;
    XRAM[54554] = 8'b0;
    XRAM[54555] = 8'b0;
    XRAM[54556] = 8'b0;
    XRAM[54557] = 8'b0;
    XRAM[54558] = 8'b0;
    XRAM[54559] = 8'b0;
    XRAM[54560] = 8'b0;
    XRAM[54561] = 8'b0;
    XRAM[54562] = 8'b0;
    XRAM[54563] = 8'b0;
    XRAM[54564] = 8'b0;
    XRAM[54565] = 8'b0;
    XRAM[54566] = 8'b0;
    XRAM[54567] = 8'b0;
    XRAM[54568] = 8'b0;
    XRAM[54569] = 8'b0;
    XRAM[54570] = 8'b0;
    XRAM[54571] = 8'b0;
    XRAM[54572] = 8'b0;
    XRAM[54573] = 8'b0;
    XRAM[54574] = 8'b0;
    XRAM[54575] = 8'b0;
    XRAM[54576] = 8'b0;
    XRAM[54577] = 8'b0;
    XRAM[54578] = 8'b0;
    XRAM[54579] = 8'b0;
    XRAM[54580] = 8'b0;
    XRAM[54581] = 8'b0;
    XRAM[54582] = 8'b0;
    XRAM[54583] = 8'b0;
    XRAM[54584] = 8'b0;
    XRAM[54585] = 8'b0;
    XRAM[54586] = 8'b0;
    XRAM[54587] = 8'b0;
    XRAM[54588] = 8'b0;
    XRAM[54589] = 8'b0;
    XRAM[54590] = 8'b0;
    XRAM[54591] = 8'b0;
    XRAM[54592] = 8'b0;
    XRAM[54593] = 8'b0;
    XRAM[54594] = 8'b0;
    XRAM[54595] = 8'b0;
    XRAM[54596] = 8'b0;
    XRAM[54597] = 8'b0;
    XRAM[54598] = 8'b0;
    XRAM[54599] = 8'b0;
    XRAM[54600] = 8'b0;
    XRAM[54601] = 8'b0;
    XRAM[54602] = 8'b0;
    XRAM[54603] = 8'b0;
    XRAM[54604] = 8'b0;
    XRAM[54605] = 8'b0;
    XRAM[54606] = 8'b0;
    XRAM[54607] = 8'b0;
    XRAM[54608] = 8'b0;
    XRAM[54609] = 8'b0;
    XRAM[54610] = 8'b0;
    XRAM[54611] = 8'b0;
    XRAM[54612] = 8'b0;
    XRAM[54613] = 8'b0;
    XRAM[54614] = 8'b0;
    XRAM[54615] = 8'b0;
    XRAM[54616] = 8'b0;
    XRAM[54617] = 8'b0;
    XRAM[54618] = 8'b0;
    XRAM[54619] = 8'b0;
    XRAM[54620] = 8'b0;
    XRAM[54621] = 8'b0;
    XRAM[54622] = 8'b0;
    XRAM[54623] = 8'b0;
    XRAM[54624] = 8'b0;
    XRAM[54625] = 8'b0;
    XRAM[54626] = 8'b0;
    XRAM[54627] = 8'b0;
    XRAM[54628] = 8'b0;
    XRAM[54629] = 8'b0;
    XRAM[54630] = 8'b0;
    XRAM[54631] = 8'b0;
    XRAM[54632] = 8'b0;
    XRAM[54633] = 8'b0;
    XRAM[54634] = 8'b0;
    XRAM[54635] = 8'b0;
    XRAM[54636] = 8'b0;
    XRAM[54637] = 8'b0;
    XRAM[54638] = 8'b0;
    XRAM[54639] = 8'b0;
    XRAM[54640] = 8'b0;
    XRAM[54641] = 8'b0;
    XRAM[54642] = 8'b0;
    XRAM[54643] = 8'b0;
    XRAM[54644] = 8'b0;
    XRAM[54645] = 8'b0;
    XRAM[54646] = 8'b0;
    XRAM[54647] = 8'b0;
    XRAM[54648] = 8'b0;
    XRAM[54649] = 8'b0;
    XRAM[54650] = 8'b0;
    XRAM[54651] = 8'b0;
    XRAM[54652] = 8'b0;
    XRAM[54653] = 8'b0;
    XRAM[54654] = 8'b0;
    XRAM[54655] = 8'b0;
    XRAM[54656] = 8'b0;
    XRAM[54657] = 8'b0;
    XRAM[54658] = 8'b0;
    XRAM[54659] = 8'b0;
    XRAM[54660] = 8'b0;
    XRAM[54661] = 8'b0;
    XRAM[54662] = 8'b0;
    XRAM[54663] = 8'b0;
    XRAM[54664] = 8'b0;
    XRAM[54665] = 8'b0;
    XRAM[54666] = 8'b0;
    XRAM[54667] = 8'b0;
    XRAM[54668] = 8'b0;
    XRAM[54669] = 8'b0;
    XRAM[54670] = 8'b0;
    XRAM[54671] = 8'b0;
    XRAM[54672] = 8'b0;
    XRAM[54673] = 8'b0;
    XRAM[54674] = 8'b0;
    XRAM[54675] = 8'b0;
    XRAM[54676] = 8'b0;
    XRAM[54677] = 8'b0;
    XRAM[54678] = 8'b0;
    XRAM[54679] = 8'b0;
    XRAM[54680] = 8'b0;
    XRAM[54681] = 8'b0;
    XRAM[54682] = 8'b0;
    XRAM[54683] = 8'b0;
    XRAM[54684] = 8'b0;
    XRAM[54685] = 8'b0;
    XRAM[54686] = 8'b0;
    XRAM[54687] = 8'b0;
    XRAM[54688] = 8'b0;
    XRAM[54689] = 8'b0;
    XRAM[54690] = 8'b0;
    XRAM[54691] = 8'b0;
    XRAM[54692] = 8'b0;
    XRAM[54693] = 8'b0;
    XRAM[54694] = 8'b0;
    XRAM[54695] = 8'b0;
    XRAM[54696] = 8'b0;
    XRAM[54697] = 8'b0;
    XRAM[54698] = 8'b0;
    XRAM[54699] = 8'b0;
    XRAM[54700] = 8'b0;
    XRAM[54701] = 8'b0;
    XRAM[54702] = 8'b0;
    XRAM[54703] = 8'b0;
    XRAM[54704] = 8'b0;
    XRAM[54705] = 8'b0;
    XRAM[54706] = 8'b0;
    XRAM[54707] = 8'b0;
    XRAM[54708] = 8'b0;
    XRAM[54709] = 8'b0;
    XRAM[54710] = 8'b0;
    XRAM[54711] = 8'b0;
    XRAM[54712] = 8'b0;
    XRAM[54713] = 8'b0;
    XRAM[54714] = 8'b0;
    XRAM[54715] = 8'b0;
    XRAM[54716] = 8'b0;
    XRAM[54717] = 8'b0;
    XRAM[54718] = 8'b0;
    XRAM[54719] = 8'b0;
    XRAM[54720] = 8'b0;
    XRAM[54721] = 8'b0;
    XRAM[54722] = 8'b0;
    XRAM[54723] = 8'b0;
    XRAM[54724] = 8'b0;
    XRAM[54725] = 8'b0;
    XRAM[54726] = 8'b0;
    XRAM[54727] = 8'b0;
    XRAM[54728] = 8'b0;
    XRAM[54729] = 8'b0;
    XRAM[54730] = 8'b0;
    XRAM[54731] = 8'b0;
    XRAM[54732] = 8'b0;
    XRAM[54733] = 8'b0;
    XRAM[54734] = 8'b0;
    XRAM[54735] = 8'b0;
    XRAM[54736] = 8'b0;
    XRAM[54737] = 8'b0;
    XRAM[54738] = 8'b0;
    XRAM[54739] = 8'b0;
    XRAM[54740] = 8'b0;
    XRAM[54741] = 8'b0;
    XRAM[54742] = 8'b0;
    XRAM[54743] = 8'b0;
    XRAM[54744] = 8'b0;
    XRAM[54745] = 8'b0;
    XRAM[54746] = 8'b0;
    XRAM[54747] = 8'b0;
    XRAM[54748] = 8'b0;
    XRAM[54749] = 8'b0;
    XRAM[54750] = 8'b0;
    XRAM[54751] = 8'b0;
    XRAM[54752] = 8'b0;
    XRAM[54753] = 8'b0;
    XRAM[54754] = 8'b0;
    XRAM[54755] = 8'b0;
    XRAM[54756] = 8'b0;
    XRAM[54757] = 8'b0;
    XRAM[54758] = 8'b0;
    XRAM[54759] = 8'b0;
    XRAM[54760] = 8'b0;
    XRAM[54761] = 8'b0;
    XRAM[54762] = 8'b0;
    XRAM[54763] = 8'b0;
    XRAM[54764] = 8'b0;
    XRAM[54765] = 8'b0;
    XRAM[54766] = 8'b0;
    XRAM[54767] = 8'b0;
    XRAM[54768] = 8'b0;
    XRAM[54769] = 8'b0;
    XRAM[54770] = 8'b0;
    XRAM[54771] = 8'b0;
    XRAM[54772] = 8'b0;
    XRAM[54773] = 8'b0;
    XRAM[54774] = 8'b0;
    XRAM[54775] = 8'b0;
    XRAM[54776] = 8'b0;
    XRAM[54777] = 8'b0;
    XRAM[54778] = 8'b0;
    XRAM[54779] = 8'b0;
    XRAM[54780] = 8'b0;
    XRAM[54781] = 8'b0;
    XRAM[54782] = 8'b0;
    XRAM[54783] = 8'b0;
    XRAM[54784] = 8'b0;
    XRAM[54785] = 8'b0;
    XRAM[54786] = 8'b0;
    XRAM[54787] = 8'b0;
    XRAM[54788] = 8'b0;
    XRAM[54789] = 8'b0;
    XRAM[54790] = 8'b0;
    XRAM[54791] = 8'b0;
    XRAM[54792] = 8'b0;
    XRAM[54793] = 8'b0;
    XRAM[54794] = 8'b0;
    XRAM[54795] = 8'b0;
    XRAM[54796] = 8'b0;
    XRAM[54797] = 8'b0;
    XRAM[54798] = 8'b0;
    XRAM[54799] = 8'b0;
    XRAM[54800] = 8'b0;
    XRAM[54801] = 8'b0;
    XRAM[54802] = 8'b0;
    XRAM[54803] = 8'b0;
    XRAM[54804] = 8'b0;
    XRAM[54805] = 8'b0;
    XRAM[54806] = 8'b0;
    XRAM[54807] = 8'b0;
    XRAM[54808] = 8'b0;
    XRAM[54809] = 8'b0;
    XRAM[54810] = 8'b0;
    XRAM[54811] = 8'b0;
    XRAM[54812] = 8'b0;
    XRAM[54813] = 8'b0;
    XRAM[54814] = 8'b0;
    XRAM[54815] = 8'b0;
    XRAM[54816] = 8'b0;
    XRAM[54817] = 8'b0;
    XRAM[54818] = 8'b0;
    XRAM[54819] = 8'b0;
    XRAM[54820] = 8'b0;
    XRAM[54821] = 8'b0;
    XRAM[54822] = 8'b0;
    XRAM[54823] = 8'b0;
    XRAM[54824] = 8'b0;
    XRAM[54825] = 8'b0;
    XRAM[54826] = 8'b0;
    XRAM[54827] = 8'b0;
    XRAM[54828] = 8'b0;
    XRAM[54829] = 8'b0;
    XRAM[54830] = 8'b0;
    XRAM[54831] = 8'b0;
    XRAM[54832] = 8'b0;
    XRAM[54833] = 8'b0;
    XRAM[54834] = 8'b0;
    XRAM[54835] = 8'b0;
    XRAM[54836] = 8'b0;
    XRAM[54837] = 8'b0;
    XRAM[54838] = 8'b0;
    XRAM[54839] = 8'b0;
    XRAM[54840] = 8'b0;
    XRAM[54841] = 8'b0;
    XRAM[54842] = 8'b0;
    XRAM[54843] = 8'b0;
    XRAM[54844] = 8'b0;
    XRAM[54845] = 8'b0;
    XRAM[54846] = 8'b0;
    XRAM[54847] = 8'b0;
    XRAM[54848] = 8'b0;
    XRAM[54849] = 8'b0;
    XRAM[54850] = 8'b0;
    XRAM[54851] = 8'b0;
    XRAM[54852] = 8'b0;
    XRAM[54853] = 8'b0;
    XRAM[54854] = 8'b0;
    XRAM[54855] = 8'b0;
    XRAM[54856] = 8'b0;
    XRAM[54857] = 8'b0;
    XRAM[54858] = 8'b0;
    XRAM[54859] = 8'b0;
    XRAM[54860] = 8'b0;
    XRAM[54861] = 8'b0;
    XRAM[54862] = 8'b0;
    XRAM[54863] = 8'b0;
    XRAM[54864] = 8'b0;
    XRAM[54865] = 8'b0;
    XRAM[54866] = 8'b0;
    XRAM[54867] = 8'b0;
    XRAM[54868] = 8'b0;
    XRAM[54869] = 8'b0;
    XRAM[54870] = 8'b0;
    XRAM[54871] = 8'b0;
    XRAM[54872] = 8'b0;
    XRAM[54873] = 8'b0;
    XRAM[54874] = 8'b0;
    XRAM[54875] = 8'b0;
    XRAM[54876] = 8'b0;
    XRAM[54877] = 8'b0;
    XRAM[54878] = 8'b0;
    XRAM[54879] = 8'b0;
    XRAM[54880] = 8'b0;
    XRAM[54881] = 8'b0;
    XRAM[54882] = 8'b0;
    XRAM[54883] = 8'b0;
    XRAM[54884] = 8'b0;
    XRAM[54885] = 8'b0;
    XRAM[54886] = 8'b0;
    XRAM[54887] = 8'b0;
    XRAM[54888] = 8'b0;
    XRAM[54889] = 8'b0;
    XRAM[54890] = 8'b0;
    XRAM[54891] = 8'b0;
    XRAM[54892] = 8'b0;
    XRAM[54893] = 8'b0;
    XRAM[54894] = 8'b0;
    XRAM[54895] = 8'b0;
    XRAM[54896] = 8'b0;
    XRAM[54897] = 8'b0;
    XRAM[54898] = 8'b0;
    XRAM[54899] = 8'b0;
    XRAM[54900] = 8'b0;
    XRAM[54901] = 8'b0;
    XRAM[54902] = 8'b0;
    XRAM[54903] = 8'b0;
    XRAM[54904] = 8'b0;
    XRAM[54905] = 8'b0;
    XRAM[54906] = 8'b0;
    XRAM[54907] = 8'b0;
    XRAM[54908] = 8'b0;
    XRAM[54909] = 8'b0;
    XRAM[54910] = 8'b0;
    XRAM[54911] = 8'b0;
    XRAM[54912] = 8'b0;
    XRAM[54913] = 8'b0;
    XRAM[54914] = 8'b0;
    XRAM[54915] = 8'b0;
    XRAM[54916] = 8'b0;
    XRAM[54917] = 8'b0;
    XRAM[54918] = 8'b0;
    XRAM[54919] = 8'b0;
    XRAM[54920] = 8'b0;
    XRAM[54921] = 8'b0;
    XRAM[54922] = 8'b0;
    XRAM[54923] = 8'b0;
    XRAM[54924] = 8'b0;
    XRAM[54925] = 8'b0;
    XRAM[54926] = 8'b0;
    XRAM[54927] = 8'b0;
    XRAM[54928] = 8'b0;
    XRAM[54929] = 8'b0;
    XRAM[54930] = 8'b0;
    XRAM[54931] = 8'b0;
    XRAM[54932] = 8'b0;
    XRAM[54933] = 8'b0;
    XRAM[54934] = 8'b0;
    XRAM[54935] = 8'b0;
    XRAM[54936] = 8'b0;
    XRAM[54937] = 8'b0;
    XRAM[54938] = 8'b0;
    XRAM[54939] = 8'b0;
    XRAM[54940] = 8'b0;
    XRAM[54941] = 8'b0;
    XRAM[54942] = 8'b0;
    XRAM[54943] = 8'b0;
    XRAM[54944] = 8'b0;
    XRAM[54945] = 8'b0;
    XRAM[54946] = 8'b0;
    XRAM[54947] = 8'b0;
    XRAM[54948] = 8'b0;
    XRAM[54949] = 8'b0;
    XRAM[54950] = 8'b0;
    XRAM[54951] = 8'b0;
    XRAM[54952] = 8'b0;
    XRAM[54953] = 8'b0;
    XRAM[54954] = 8'b0;
    XRAM[54955] = 8'b0;
    XRAM[54956] = 8'b0;
    XRAM[54957] = 8'b0;
    XRAM[54958] = 8'b0;
    XRAM[54959] = 8'b0;
    XRAM[54960] = 8'b0;
    XRAM[54961] = 8'b0;
    XRAM[54962] = 8'b0;
    XRAM[54963] = 8'b0;
    XRAM[54964] = 8'b0;
    XRAM[54965] = 8'b0;
    XRAM[54966] = 8'b0;
    XRAM[54967] = 8'b0;
    XRAM[54968] = 8'b0;
    XRAM[54969] = 8'b0;
    XRAM[54970] = 8'b0;
    XRAM[54971] = 8'b0;
    XRAM[54972] = 8'b0;
    XRAM[54973] = 8'b0;
    XRAM[54974] = 8'b0;
    XRAM[54975] = 8'b0;
    XRAM[54976] = 8'b0;
    XRAM[54977] = 8'b0;
    XRAM[54978] = 8'b0;
    XRAM[54979] = 8'b0;
    XRAM[54980] = 8'b0;
    XRAM[54981] = 8'b0;
    XRAM[54982] = 8'b0;
    XRAM[54983] = 8'b0;
    XRAM[54984] = 8'b0;
    XRAM[54985] = 8'b0;
    XRAM[54986] = 8'b0;
    XRAM[54987] = 8'b0;
    XRAM[54988] = 8'b0;
    XRAM[54989] = 8'b0;
    XRAM[54990] = 8'b0;
    XRAM[54991] = 8'b0;
    XRAM[54992] = 8'b0;
    XRAM[54993] = 8'b0;
    XRAM[54994] = 8'b0;
    XRAM[54995] = 8'b0;
    XRAM[54996] = 8'b0;
    XRAM[54997] = 8'b0;
    XRAM[54998] = 8'b0;
    XRAM[54999] = 8'b0;
    XRAM[55000] = 8'b0;
    XRAM[55001] = 8'b0;
    XRAM[55002] = 8'b0;
    XRAM[55003] = 8'b0;
    XRAM[55004] = 8'b0;
    XRAM[55005] = 8'b0;
    XRAM[55006] = 8'b0;
    XRAM[55007] = 8'b0;
    XRAM[55008] = 8'b0;
    XRAM[55009] = 8'b0;
    XRAM[55010] = 8'b0;
    XRAM[55011] = 8'b0;
    XRAM[55012] = 8'b0;
    XRAM[55013] = 8'b0;
    XRAM[55014] = 8'b0;
    XRAM[55015] = 8'b0;
    XRAM[55016] = 8'b0;
    XRAM[55017] = 8'b0;
    XRAM[55018] = 8'b0;
    XRAM[55019] = 8'b0;
    XRAM[55020] = 8'b0;
    XRAM[55021] = 8'b0;
    XRAM[55022] = 8'b0;
    XRAM[55023] = 8'b0;
    XRAM[55024] = 8'b0;
    XRAM[55025] = 8'b0;
    XRAM[55026] = 8'b0;
    XRAM[55027] = 8'b0;
    XRAM[55028] = 8'b0;
    XRAM[55029] = 8'b0;
    XRAM[55030] = 8'b0;
    XRAM[55031] = 8'b0;
    XRAM[55032] = 8'b0;
    XRAM[55033] = 8'b0;
    XRAM[55034] = 8'b0;
    XRAM[55035] = 8'b0;
    XRAM[55036] = 8'b0;
    XRAM[55037] = 8'b0;
    XRAM[55038] = 8'b0;
    XRAM[55039] = 8'b0;
    XRAM[55040] = 8'b0;
    XRAM[55041] = 8'b0;
    XRAM[55042] = 8'b0;
    XRAM[55043] = 8'b0;
    XRAM[55044] = 8'b0;
    XRAM[55045] = 8'b0;
    XRAM[55046] = 8'b0;
    XRAM[55047] = 8'b0;
    XRAM[55048] = 8'b0;
    XRAM[55049] = 8'b0;
    XRAM[55050] = 8'b0;
    XRAM[55051] = 8'b0;
    XRAM[55052] = 8'b0;
    XRAM[55053] = 8'b0;
    XRAM[55054] = 8'b0;
    XRAM[55055] = 8'b0;
    XRAM[55056] = 8'b0;
    XRAM[55057] = 8'b0;
    XRAM[55058] = 8'b0;
    XRAM[55059] = 8'b0;
    XRAM[55060] = 8'b0;
    XRAM[55061] = 8'b0;
    XRAM[55062] = 8'b0;
    XRAM[55063] = 8'b0;
    XRAM[55064] = 8'b0;
    XRAM[55065] = 8'b0;
    XRAM[55066] = 8'b0;
    XRAM[55067] = 8'b0;
    XRAM[55068] = 8'b0;
    XRAM[55069] = 8'b0;
    XRAM[55070] = 8'b0;
    XRAM[55071] = 8'b0;
    XRAM[55072] = 8'b0;
    XRAM[55073] = 8'b0;
    XRAM[55074] = 8'b0;
    XRAM[55075] = 8'b0;
    XRAM[55076] = 8'b0;
    XRAM[55077] = 8'b0;
    XRAM[55078] = 8'b0;
    XRAM[55079] = 8'b0;
    XRAM[55080] = 8'b0;
    XRAM[55081] = 8'b0;
    XRAM[55082] = 8'b0;
    XRAM[55083] = 8'b0;
    XRAM[55084] = 8'b0;
    XRAM[55085] = 8'b0;
    XRAM[55086] = 8'b0;
    XRAM[55087] = 8'b0;
    XRAM[55088] = 8'b0;
    XRAM[55089] = 8'b0;
    XRAM[55090] = 8'b0;
    XRAM[55091] = 8'b0;
    XRAM[55092] = 8'b0;
    XRAM[55093] = 8'b0;
    XRAM[55094] = 8'b0;
    XRAM[55095] = 8'b0;
    XRAM[55096] = 8'b0;
    XRAM[55097] = 8'b0;
    XRAM[55098] = 8'b0;
    XRAM[55099] = 8'b0;
    XRAM[55100] = 8'b0;
    XRAM[55101] = 8'b0;
    XRAM[55102] = 8'b0;
    XRAM[55103] = 8'b0;
    XRAM[55104] = 8'b0;
    XRAM[55105] = 8'b0;
    XRAM[55106] = 8'b0;
    XRAM[55107] = 8'b0;
    XRAM[55108] = 8'b0;
    XRAM[55109] = 8'b0;
    XRAM[55110] = 8'b0;
    XRAM[55111] = 8'b0;
    XRAM[55112] = 8'b0;
    XRAM[55113] = 8'b0;
    XRAM[55114] = 8'b0;
    XRAM[55115] = 8'b0;
    XRAM[55116] = 8'b0;
    XRAM[55117] = 8'b0;
    XRAM[55118] = 8'b0;
    XRAM[55119] = 8'b0;
    XRAM[55120] = 8'b0;
    XRAM[55121] = 8'b0;
    XRAM[55122] = 8'b0;
    XRAM[55123] = 8'b0;
    XRAM[55124] = 8'b0;
    XRAM[55125] = 8'b0;
    XRAM[55126] = 8'b0;
    XRAM[55127] = 8'b0;
    XRAM[55128] = 8'b0;
    XRAM[55129] = 8'b0;
    XRAM[55130] = 8'b0;
    XRAM[55131] = 8'b0;
    XRAM[55132] = 8'b0;
    XRAM[55133] = 8'b0;
    XRAM[55134] = 8'b0;
    XRAM[55135] = 8'b0;
    XRAM[55136] = 8'b0;
    XRAM[55137] = 8'b0;
    XRAM[55138] = 8'b0;
    XRAM[55139] = 8'b0;
    XRAM[55140] = 8'b0;
    XRAM[55141] = 8'b0;
    XRAM[55142] = 8'b0;
    XRAM[55143] = 8'b0;
    XRAM[55144] = 8'b0;
    XRAM[55145] = 8'b0;
    XRAM[55146] = 8'b0;
    XRAM[55147] = 8'b0;
    XRAM[55148] = 8'b0;
    XRAM[55149] = 8'b0;
    XRAM[55150] = 8'b0;
    XRAM[55151] = 8'b0;
    XRAM[55152] = 8'b0;
    XRAM[55153] = 8'b0;
    XRAM[55154] = 8'b0;
    XRAM[55155] = 8'b0;
    XRAM[55156] = 8'b0;
    XRAM[55157] = 8'b0;
    XRAM[55158] = 8'b0;
    XRAM[55159] = 8'b0;
    XRAM[55160] = 8'b0;
    XRAM[55161] = 8'b0;
    XRAM[55162] = 8'b0;
    XRAM[55163] = 8'b0;
    XRAM[55164] = 8'b0;
    XRAM[55165] = 8'b0;
    XRAM[55166] = 8'b0;
    XRAM[55167] = 8'b0;
    XRAM[55168] = 8'b0;
    XRAM[55169] = 8'b0;
    XRAM[55170] = 8'b0;
    XRAM[55171] = 8'b0;
    XRAM[55172] = 8'b0;
    XRAM[55173] = 8'b0;
    XRAM[55174] = 8'b0;
    XRAM[55175] = 8'b0;
    XRAM[55176] = 8'b0;
    XRAM[55177] = 8'b0;
    XRAM[55178] = 8'b0;
    XRAM[55179] = 8'b0;
    XRAM[55180] = 8'b0;
    XRAM[55181] = 8'b0;
    XRAM[55182] = 8'b0;
    XRAM[55183] = 8'b0;
    XRAM[55184] = 8'b0;
    XRAM[55185] = 8'b0;
    XRAM[55186] = 8'b0;
    XRAM[55187] = 8'b0;
    XRAM[55188] = 8'b0;
    XRAM[55189] = 8'b0;
    XRAM[55190] = 8'b0;
    XRAM[55191] = 8'b0;
    XRAM[55192] = 8'b0;
    XRAM[55193] = 8'b0;
    XRAM[55194] = 8'b0;
    XRAM[55195] = 8'b0;
    XRAM[55196] = 8'b0;
    XRAM[55197] = 8'b0;
    XRAM[55198] = 8'b0;
    XRAM[55199] = 8'b0;
    XRAM[55200] = 8'b0;
    XRAM[55201] = 8'b0;
    XRAM[55202] = 8'b0;
    XRAM[55203] = 8'b0;
    XRAM[55204] = 8'b0;
    XRAM[55205] = 8'b0;
    XRAM[55206] = 8'b0;
    XRAM[55207] = 8'b0;
    XRAM[55208] = 8'b0;
    XRAM[55209] = 8'b0;
    XRAM[55210] = 8'b0;
    XRAM[55211] = 8'b0;
    XRAM[55212] = 8'b0;
    XRAM[55213] = 8'b0;
    XRAM[55214] = 8'b0;
    XRAM[55215] = 8'b0;
    XRAM[55216] = 8'b0;
    XRAM[55217] = 8'b0;
    XRAM[55218] = 8'b0;
    XRAM[55219] = 8'b0;
    XRAM[55220] = 8'b0;
    XRAM[55221] = 8'b0;
    XRAM[55222] = 8'b0;
    XRAM[55223] = 8'b0;
    XRAM[55224] = 8'b0;
    XRAM[55225] = 8'b0;
    XRAM[55226] = 8'b0;
    XRAM[55227] = 8'b0;
    XRAM[55228] = 8'b0;
    XRAM[55229] = 8'b0;
    XRAM[55230] = 8'b0;
    XRAM[55231] = 8'b0;
    XRAM[55232] = 8'b0;
    XRAM[55233] = 8'b0;
    XRAM[55234] = 8'b0;
    XRAM[55235] = 8'b0;
    XRAM[55236] = 8'b0;
    XRAM[55237] = 8'b0;
    XRAM[55238] = 8'b0;
    XRAM[55239] = 8'b0;
    XRAM[55240] = 8'b0;
    XRAM[55241] = 8'b0;
    XRAM[55242] = 8'b0;
    XRAM[55243] = 8'b0;
    XRAM[55244] = 8'b0;
    XRAM[55245] = 8'b0;
    XRAM[55246] = 8'b0;
    XRAM[55247] = 8'b0;
    XRAM[55248] = 8'b0;
    XRAM[55249] = 8'b0;
    XRAM[55250] = 8'b0;
    XRAM[55251] = 8'b0;
    XRAM[55252] = 8'b0;
    XRAM[55253] = 8'b0;
    XRAM[55254] = 8'b0;
    XRAM[55255] = 8'b0;
    XRAM[55256] = 8'b0;
    XRAM[55257] = 8'b0;
    XRAM[55258] = 8'b0;
    XRAM[55259] = 8'b0;
    XRAM[55260] = 8'b0;
    XRAM[55261] = 8'b0;
    XRAM[55262] = 8'b0;
    XRAM[55263] = 8'b0;
    XRAM[55264] = 8'b0;
    XRAM[55265] = 8'b0;
    XRAM[55266] = 8'b0;
    XRAM[55267] = 8'b0;
    XRAM[55268] = 8'b0;
    XRAM[55269] = 8'b0;
    XRAM[55270] = 8'b0;
    XRAM[55271] = 8'b0;
    XRAM[55272] = 8'b0;
    XRAM[55273] = 8'b0;
    XRAM[55274] = 8'b0;
    XRAM[55275] = 8'b0;
    XRAM[55276] = 8'b0;
    XRAM[55277] = 8'b0;
    XRAM[55278] = 8'b0;
    XRAM[55279] = 8'b0;
    XRAM[55280] = 8'b0;
    XRAM[55281] = 8'b0;
    XRAM[55282] = 8'b0;
    XRAM[55283] = 8'b0;
    XRAM[55284] = 8'b0;
    XRAM[55285] = 8'b0;
    XRAM[55286] = 8'b0;
    XRAM[55287] = 8'b0;
    XRAM[55288] = 8'b0;
    XRAM[55289] = 8'b0;
    XRAM[55290] = 8'b0;
    XRAM[55291] = 8'b0;
    XRAM[55292] = 8'b0;
    XRAM[55293] = 8'b0;
    XRAM[55294] = 8'b0;
    XRAM[55295] = 8'b0;
    XRAM[55296] = 8'b0;
    XRAM[55297] = 8'b0;
    XRAM[55298] = 8'b0;
    XRAM[55299] = 8'b0;
    XRAM[55300] = 8'b0;
    XRAM[55301] = 8'b0;
    XRAM[55302] = 8'b0;
    XRAM[55303] = 8'b0;
    XRAM[55304] = 8'b0;
    XRAM[55305] = 8'b0;
    XRAM[55306] = 8'b0;
    XRAM[55307] = 8'b0;
    XRAM[55308] = 8'b0;
    XRAM[55309] = 8'b0;
    XRAM[55310] = 8'b0;
    XRAM[55311] = 8'b0;
    XRAM[55312] = 8'b0;
    XRAM[55313] = 8'b0;
    XRAM[55314] = 8'b0;
    XRAM[55315] = 8'b0;
    XRAM[55316] = 8'b0;
    XRAM[55317] = 8'b0;
    XRAM[55318] = 8'b0;
    XRAM[55319] = 8'b0;
    XRAM[55320] = 8'b0;
    XRAM[55321] = 8'b0;
    XRAM[55322] = 8'b0;
    XRAM[55323] = 8'b0;
    XRAM[55324] = 8'b0;
    XRAM[55325] = 8'b0;
    XRAM[55326] = 8'b0;
    XRAM[55327] = 8'b0;
    XRAM[55328] = 8'b0;
    XRAM[55329] = 8'b0;
    XRAM[55330] = 8'b0;
    XRAM[55331] = 8'b0;
    XRAM[55332] = 8'b0;
    XRAM[55333] = 8'b0;
    XRAM[55334] = 8'b0;
    XRAM[55335] = 8'b0;
    XRAM[55336] = 8'b0;
    XRAM[55337] = 8'b0;
    XRAM[55338] = 8'b0;
    XRAM[55339] = 8'b0;
    XRAM[55340] = 8'b0;
    XRAM[55341] = 8'b0;
    XRAM[55342] = 8'b0;
    XRAM[55343] = 8'b0;
    XRAM[55344] = 8'b0;
    XRAM[55345] = 8'b0;
    XRAM[55346] = 8'b0;
    XRAM[55347] = 8'b0;
    XRAM[55348] = 8'b0;
    XRAM[55349] = 8'b0;
    XRAM[55350] = 8'b0;
    XRAM[55351] = 8'b0;
    XRAM[55352] = 8'b0;
    XRAM[55353] = 8'b0;
    XRAM[55354] = 8'b0;
    XRAM[55355] = 8'b0;
    XRAM[55356] = 8'b0;
    XRAM[55357] = 8'b0;
    XRAM[55358] = 8'b0;
    XRAM[55359] = 8'b0;
    XRAM[55360] = 8'b0;
    XRAM[55361] = 8'b0;
    XRAM[55362] = 8'b0;
    XRAM[55363] = 8'b0;
    XRAM[55364] = 8'b0;
    XRAM[55365] = 8'b0;
    XRAM[55366] = 8'b0;
    XRAM[55367] = 8'b0;
    XRAM[55368] = 8'b0;
    XRAM[55369] = 8'b0;
    XRAM[55370] = 8'b0;
    XRAM[55371] = 8'b0;
    XRAM[55372] = 8'b0;
    XRAM[55373] = 8'b0;
    XRAM[55374] = 8'b0;
    XRAM[55375] = 8'b0;
    XRAM[55376] = 8'b0;
    XRAM[55377] = 8'b0;
    XRAM[55378] = 8'b0;
    XRAM[55379] = 8'b0;
    XRAM[55380] = 8'b0;
    XRAM[55381] = 8'b0;
    XRAM[55382] = 8'b0;
    XRAM[55383] = 8'b0;
    XRAM[55384] = 8'b0;
    XRAM[55385] = 8'b0;
    XRAM[55386] = 8'b0;
    XRAM[55387] = 8'b0;
    XRAM[55388] = 8'b0;
    XRAM[55389] = 8'b0;
    XRAM[55390] = 8'b0;
    XRAM[55391] = 8'b0;
    XRAM[55392] = 8'b0;
    XRAM[55393] = 8'b0;
    XRAM[55394] = 8'b0;
    XRAM[55395] = 8'b0;
    XRAM[55396] = 8'b0;
    XRAM[55397] = 8'b0;
    XRAM[55398] = 8'b0;
    XRAM[55399] = 8'b0;
    XRAM[55400] = 8'b0;
    XRAM[55401] = 8'b0;
    XRAM[55402] = 8'b0;
    XRAM[55403] = 8'b0;
    XRAM[55404] = 8'b0;
    XRAM[55405] = 8'b0;
    XRAM[55406] = 8'b0;
    XRAM[55407] = 8'b0;
    XRAM[55408] = 8'b0;
    XRAM[55409] = 8'b0;
    XRAM[55410] = 8'b0;
    XRAM[55411] = 8'b0;
    XRAM[55412] = 8'b0;
    XRAM[55413] = 8'b0;
    XRAM[55414] = 8'b0;
    XRAM[55415] = 8'b0;
    XRAM[55416] = 8'b0;
    XRAM[55417] = 8'b0;
    XRAM[55418] = 8'b0;
    XRAM[55419] = 8'b0;
    XRAM[55420] = 8'b0;
    XRAM[55421] = 8'b0;
    XRAM[55422] = 8'b0;
    XRAM[55423] = 8'b0;
    XRAM[55424] = 8'b0;
    XRAM[55425] = 8'b0;
    XRAM[55426] = 8'b0;
    XRAM[55427] = 8'b0;
    XRAM[55428] = 8'b0;
    XRAM[55429] = 8'b0;
    XRAM[55430] = 8'b0;
    XRAM[55431] = 8'b0;
    XRAM[55432] = 8'b0;
    XRAM[55433] = 8'b0;
    XRAM[55434] = 8'b0;
    XRAM[55435] = 8'b0;
    XRAM[55436] = 8'b0;
    XRAM[55437] = 8'b0;
    XRAM[55438] = 8'b0;
    XRAM[55439] = 8'b0;
    XRAM[55440] = 8'b0;
    XRAM[55441] = 8'b0;
    XRAM[55442] = 8'b0;
    XRAM[55443] = 8'b0;
    XRAM[55444] = 8'b0;
    XRAM[55445] = 8'b0;
    XRAM[55446] = 8'b0;
    XRAM[55447] = 8'b0;
    XRAM[55448] = 8'b0;
    XRAM[55449] = 8'b0;
    XRAM[55450] = 8'b0;
    XRAM[55451] = 8'b0;
    XRAM[55452] = 8'b0;
    XRAM[55453] = 8'b0;
    XRAM[55454] = 8'b0;
    XRAM[55455] = 8'b0;
    XRAM[55456] = 8'b0;
    XRAM[55457] = 8'b0;
    XRAM[55458] = 8'b0;
    XRAM[55459] = 8'b0;
    XRAM[55460] = 8'b0;
    XRAM[55461] = 8'b0;
    XRAM[55462] = 8'b0;
    XRAM[55463] = 8'b0;
    XRAM[55464] = 8'b0;
    XRAM[55465] = 8'b0;
    XRAM[55466] = 8'b0;
    XRAM[55467] = 8'b0;
    XRAM[55468] = 8'b0;
    XRAM[55469] = 8'b0;
    XRAM[55470] = 8'b0;
    XRAM[55471] = 8'b0;
    XRAM[55472] = 8'b0;
    XRAM[55473] = 8'b0;
    XRAM[55474] = 8'b0;
    XRAM[55475] = 8'b0;
    XRAM[55476] = 8'b0;
    XRAM[55477] = 8'b0;
    XRAM[55478] = 8'b0;
    XRAM[55479] = 8'b0;
    XRAM[55480] = 8'b0;
    XRAM[55481] = 8'b0;
    XRAM[55482] = 8'b0;
    XRAM[55483] = 8'b0;
    XRAM[55484] = 8'b0;
    XRAM[55485] = 8'b0;
    XRAM[55486] = 8'b0;
    XRAM[55487] = 8'b0;
    XRAM[55488] = 8'b0;
    XRAM[55489] = 8'b0;
    XRAM[55490] = 8'b0;
    XRAM[55491] = 8'b0;
    XRAM[55492] = 8'b0;
    XRAM[55493] = 8'b0;
    XRAM[55494] = 8'b0;
    XRAM[55495] = 8'b0;
    XRAM[55496] = 8'b0;
    XRAM[55497] = 8'b0;
    XRAM[55498] = 8'b0;
    XRAM[55499] = 8'b0;
    XRAM[55500] = 8'b0;
    XRAM[55501] = 8'b0;
    XRAM[55502] = 8'b0;
    XRAM[55503] = 8'b0;
    XRAM[55504] = 8'b0;
    XRAM[55505] = 8'b0;
    XRAM[55506] = 8'b0;
    XRAM[55507] = 8'b0;
    XRAM[55508] = 8'b0;
    XRAM[55509] = 8'b0;
    XRAM[55510] = 8'b0;
    XRAM[55511] = 8'b0;
    XRAM[55512] = 8'b0;
    XRAM[55513] = 8'b0;
    XRAM[55514] = 8'b0;
    XRAM[55515] = 8'b0;
    XRAM[55516] = 8'b0;
    XRAM[55517] = 8'b0;
    XRAM[55518] = 8'b0;
    XRAM[55519] = 8'b0;
    XRAM[55520] = 8'b0;
    XRAM[55521] = 8'b0;
    XRAM[55522] = 8'b0;
    XRAM[55523] = 8'b0;
    XRAM[55524] = 8'b0;
    XRAM[55525] = 8'b0;
    XRAM[55526] = 8'b0;
    XRAM[55527] = 8'b0;
    XRAM[55528] = 8'b0;
    XRAM[55529] = 8'b0;
    XRAM[55530] = 8'b0;
    XRAM[55531] = 8'b0;
    XRAM[55532] = 8'b0;
    XRAM[55533] = 8'b0;
    XRAM[55534] = 8'b0;
    XRAM[55535] = 8'b0;
    XRAM[55536] = 8'b0;
    XRAM[55537] = 8'b0;
    XRAM[55538] = 8'b0;
    XRAM[55539] = 8'b0;
    XRAM[55540] = 8'b0;
    XRAM[55541] = 8'b0;
    XRAM[55542] = 8'b0;
    XRAM[55543] = 8'b0;
    XRAM[55544] = 8'b0;
    XRAM[55545] = 8'b0;
    XRAM[55546] = 8'b0;
    XRAM[55547] = 8'b0;
    XRAM[55548] = 8'b0;
    XRAM[55549] = 8'b0;
    XRAM[55550] = 8'b0;
    XRAM[55551] = 8'b0;
    XRAM[55552] = 8'b0;
    XRAM[55553] = 8'b0;
    XRAM[55554] = 8'b0;
    XRAM[55555] = 8'b0;
    XRAM[55556] = 8'b0;
    XRAM[55557] = 8'b0;
    XRAM[55558] = 8'b0;
    XRAM[55559] = 8'b0;
    XRAM[55560] = 8'b0;
    XRAM[55561] = 8'b0;
    XRAM[55562] = 8'b0;
    XRAM[55563] = 8'b0;
    XRAM[55564] = 8'b0;
    XRAM[55565] = 8'b0;
    XRAM[55566] = 8'b0;
    XRAM[55567] = 8'b0;
    XRAM[55568] = 8'b0;
    XRAM[55569] = 8'b0;
    XRAM[55570] = 8'b0;
    XRAM[55571] = 8'b0;
    XRAM[55572] = 8'b0;
    XRAM[55573] = 8'b0;
    XRAM[55574] = 8'b0;
    XRAM[55575] = 8'b0;
    XRAM[55576] = 8'b0;
    XRAM[55577] = 8'b0;
    XRAM[55578] = 8'b0;
    XRAM[55579] = 8'b0;
    XRAM[55580] = 8'b0;
    XRAM[55581] = 8'b0;
    XRAM[55582] = 8'b0;
    XRAM[55583] = 8'b0;
    XRAM[55584] = 8'b0;
    XRAM[55585] = 8'b0;
    XRAM[55586] = 8'b0;
    XRAM[55587] = 8'b0;
    XRAM[55588] = 8'b0;
    XRAM[55589] = 8'b0;
    XRAM[55590] = 8'b0;
    XRAM[55591] = 8'b0;
    XRAM[55592] = 8'b0;
    XRAM[55593] = 8'b0;
    XRAM[55594] = 8'b0;
    XRAM[55595] = 8'b0;
    XRAM[55596] = 8'b0;
    XRAM[55597] = 8'b0;
    XRAM[55598] = 8'b0;
    XRAM[55599] = 8'b0;
    XRAM[55600] = 8'b0;
    XRAM[55601] = 8'b0;
    XRAM[55602] = 8'b0;
    XRAM[55603] = 8'b0;
    XRAM[55604] = 8'b0;
    XRAM[55605] = 8'b0;
    XRAM[55606] = 8'b0;
    XRAM[55607] = 8'b0;
    XRAM[55608] = 8'b0;
    XRAM[55609] = 8'b0;
    XRAM[55610] = 8'b0;
    XRAM[55611] = 8'b0;
    XRAM[55612] = 8'b0;
    XRAM[55613] = 8'b0;
    XRAM[55614] = 8'b0;
    XRAM[55615] = 8'b0;
    XRAM[55616] = 8'b0;
    XRAM[55617] = 8'b0;
    XRAM[55618] = 8'b0;
    XRAM[55619] = 8'b0;
    XRAM[55620] = 8'b0;
    XRAM[55621] = 8'b0;
    XRAM[55622] = 8'b0;
    XRAM[55623] = 8'b0;
    XRAM[55624] = 8'b0;
    XRAM[55625] = 8'b0;
    XRAM[55626] = 8'b0;
    XRAM[55627] = 8'b0;
    XRAM[55628] = 8'b0;
    XRAM[55629] = 8'b0;
    XRAM[55630] = 8'b0;
    XRAM[55631] = 8'b0;
    XRAM[55632] = 8'b0;
    XRAM[55633] = 8'b0;
    XRAM[55634] = 8'b0;
    XRAM[55635] = 8'b0;
    XRAM[55636] = 8'b0;
    XRAM[55637] = 8'b0;
    XRAM[55638] = 8'b0;
    XRAM[55639] = 8'b0;
    XRAM[55640] = 8'b0;
    XRAM[55641] = 8'b0;
    XRAM[55642] = 8'b0;
    XRAM[55643] = 8'b0;
    XRAM[55644] = 8'b0;
    XRAM[55645] = 8'b0;
    XRAM[55646] = 8'b0;
    XRAM[55647] = 8'b0;
    XRAM[55648] = 8'b0;
    XRAM[55649] = 8'b0;
    XRAM[55650] = 8'b0;
    XRAM[55651] = 8'b0;
    XRAM[55652] = 8'b0;
    XRAM[55653] = 8'b0;
    XRAM[55654] = 8'b0;
    XRAM[55655] = 8'b0;
    XRAM[55656] = 8'b0;
    XRAM[55657] = 8'b0;
    XRAM[55658] = 8'b0;
    XRAM[55659] = 8'b0;
    XRAM[55660] = 8'b0;
    XRAM[55661] = 8'b0;
    XRAM[55662] = 8'b0;
    XRAM[55663] = 8'b0;
    XRAM[55664] = 8'b0;
    XRAM[55665] = 8'b0;
    XRAM[55666] = 8'b0;
    XRAM[55667] = 8'b0;
    XRAM[55668] = 8'b0;
    XRAM[55669] = 8'b0;
    XRAM[55670] = 8'b0;
    XRAM[55671] = 8'b0;
    XRAM[55672] = 8'b0;
    XRAM[55673] = 8'b0;
    XRAM[55674] = 8'b0;
    XRAM[55675] = 8'b0;
    XRAM[55676] = 8'b0;
    XRAM[55677] = 8'b0;
    XRAM[55678] = 8'b0;
    XRAM[55679] = 8'b0;
    XRAM[55680] = 8'b0;
    XRAM[55681] = 8'b0;
    XRAM[55682] = 8'b0;
    XRAM[55683] = 8'b0;
    XRAM[55684] = 8'b0;
    XRAM[55685] = 8'b0;
    XRAM[55686] = 8'b0;
    XRAM[55687] = 8'b0;
    XRAM[55688] = 8'b0;
    XRAM[55689] = 8'b0;
    XRAM[55690] = 8'b0;
    XRAM[55691] = 8'b0;
    XRAM[55692] = 8'b0;
    XRAM[55693] = 8'b0;
    XRAM[55694] = 8'b0;
    XRAM[55695] = 8'b0;
    XRAM[55696] = 8'b0;
    XRAM[55697] = 8'b0;
    XRAM[55698] = 8'b0;
    XRAM[55699] = 8'b0;
    XRAM[55700] = 8'b0;
    XRAM[55701] = 8'b0;
    XRAM[55702] = 8'b0;
    XRAM[55703] = 8'b0;
    XRAM[55704] = 8'b0;
    XRAM[55705] = 8'b0;
    XRAM[55706] = 8'b0;
    XRAM[55707] = 8'b0;
    XRAM[55708] = 8'b0;
    XRAM[55709] = 8'b0;
    XRAM[55710] = 8'b0;
    XRAM[55711] = 8'b0;
    XRAM[55712] = 8'b0;
    XRAM[55713] = 8'b0;
    XRAM[55714] = 8'b0;
    XRAM[55715] = 8'b0;
    XRAM[55716] = 8'b0;
    XRAM[55717] = 8'b0;
    XRAM[55718] = 8'b0;
    XRAM[55719] = 8'b0;
    XRAM[55720] = 8'b0;
    XRAM[55721] = 8'b0;
    XRAM[55722] = 8'b0;
    XRAM[55723] = 8'b0;
    XRAM[55724] = 8'b0;
    XRAM[55725] = 8'b0;
    XRAM[55726] = 8'b0;
    XRAM[55727] = 8'b0;
    XRAM[55728] = 8'b0;
    XRAM[55729] = 8'b0;
    XRAM[55730] = 8'b0;
    XRAM[55731] = 8'b0;
    XRAM[55732] = 8'b0;
    XRAM[55733] = 8'b0;
    XRAM[55734] = 8'b0;
    XRAM[55735] = 8'b0;
    XRAM[55736] = 8'b0;
    XRAM[55737] = 8'b0;
    XRAM[55738] = 8'b0;
    XRAM[55739] = 8'b0;
    XRAM[55740] = 8'b0;
    XRAM[55741] = 8'b0;
    XRAM[55742] = 8'b0;
    XRAM[55743] = 8'b0;
    XRAM[55744] = 8'b0;
    XRAM[55745] = 8'b0;
    XRAM[55746] = 8'b0;
    XRAM[55747] = 8'b0;
    XRAM[55748] = 8'b0;
    XRAM[55749] = 8'b0;
    XRAM[55750] = 8'b0;
    XRAM[55751] = 8'b0;
    XRAM[55752] = 8'b0;
    XRAM[55753] = 8'b0;
    XRAM[55754] = 8'b0;
    XRAM[55755] = 8'b0;
    XRAM[55756] = 8'b0;
    XRAM[55757] = 8'b0;
    XRAM[55758] = 8'b0;
    XRAM[55759] = 8'b0;
    XRAM[55760] = 8'b0;
    XRAM[55761] = 8'b0;
    XRAM[55762] = 8'b0;
    XRAM[55763] = 8'b0;
    XRAM[55764] = 8'b0;
    XRAM[55765] = 8'b0;
    XRAM[55766] = 8'b0;
    XRAM[55767] = 8'b0;
    XRAM[55768] = 8'b0;
    XRAM[55769] = 8'b0;
    XRAM[55770] = 8'b0;
    XRAM[55771] = 8'b0;
    XRAM[55772] = 8'b0;
    XRAM[55773] = 8'b0;
    XRAM[55774] = 8'b0;
    XRAM[55775] = 8'b0;
    XRAM[55776] = 8'b0;
    XRAM[55777] = 8'b0;
    XRAM[55778] = 8'b0;
    XRAM[55779] = 8'b0;
    XRAM[55780] = 8'b0;
    XRAM[55781] = 8'b0;
    XRAM[55782] = 8'b0;
    XRAM[55783] = 8'b0;
    XRAM[55784] = 8'b0;
    XRAM[55785] = 8'b0;
    XRAM[55786] = 8'b0;
    XRAM[55787] = 8'b0;
    XRAM[55788] = 8'b0;
    XRAM[55789] = 8'b0;
    XRAM[55790] = 8'b0;
    XRAM[55791] = 8'b0;
    XRAM[55792] = 8'b0;
    XRAM[55793] = 8'b0;
    XRAM[55794] = 8'b0;
    XRAM[55795] = 8'b0;
    XRAM[55796] = 8'b0;
    XRAM[55797] = 8'b0;
    XRAM[55798] = 8'b0;
    XRAM[55799] = 8'b0;
    XRAM[55800] = 8'b0;
    XRAM[55801] = 8'b0;
    XRAM[55802] = 8'b0;
    XRAM[55803] = 8'b0;
    XRAM[55804] = 8'b0;
    XRAM[55805] = 8'b0;
    XRAM[55806] = 8'b0;
    XRAM[55807] = 8'b0;
    XRAM[55808] = 8'b0;
    XRAM[55809] = 8'b0;
    XRAM[55810] = 8'b0;
    XRAM[55811] = 8'b0;
    XRAM[55812] = 8'b0;
    XRAM[55813] = 8'b0;
    XRAM[55814] = 8'b0;
    XRAM[55815] = 8'b0;
    XRAM[55816] = 8'b0;
    XRAM[55817] = 8'b0;
    XRAM[55818] = 8'b0;
    XRAM[55819] = 8'b0;
    XRAM[55820] = 8'b0;
    XRAM[55821] = 8'b0;
    XRAM[55822] = 8'b0;
    XRAM[55823] = 8'b0;
    XRAM[55824] = 8'b0;
    XRAM[55825] = 8'b0;
    XRAM[55826] = 8'b0;
    XRAM[55827] = 8'b0;
    XRAM[55828] = 8'b0;
    XRAM[55829] = 8'b0;
    XRAM[55830] = 8'b0;
    XRAM[55831] = 8'b0;
    XRAM[55832] = 8'b0;
    XRAM[55833] = 8'b0;
    XRAM[55834] = 8'b0;
    XRAM[55835] = 8'b0;
    XRAM[55836] = 8'b0;
    XRAM[55837] = 8'b0;
    XRAM[55838] = 8'b0;
    XRAM[55839] = 8'b0;
    XRAM[55840] = 8'b0;
    XRAM[55841] = 8'b0;
    XRAM[55842] = 8'b0;
    XRAM[55843] = 8'b0;
    XRAM[55844] = 8'b0;
    XRAM[55845] = 8'b0;
    XRAM[55846] = 8'b0;
    XRAM[55847] = 8'b0;
    XRAM[55848] = 8'b0;
    XRAM[55849] = 8'b0;
    XRAM[55850] = 8'b0;
    XRAM[55851] = 8'b0;
    XRAM[55852] = 8'b0;
    XRAM[55853] = 8'b0;
    XRAM[55854] = 8'b0;
    XRAM[55855] = 8'b0;
    XRAM[55856] = 8'b0;
    XRAM[55857] = 8'b0;
    XRAM[55858] = 8'b0;
    XRAM[55859] = 8'b0;
    XRAM[55860] = 8'b0;
    XRAM[55861] = 8'b0;
    XRAM[55862] = 8'b0;
    XRAM[55863] = 8'b0;
    XRAM[55864] = 8'b0;
    XRAM[55865] = 8'b0;
    XRAM[55866] = 8'b0;
    XRAM[55867] = 8'b0;
    XRAM[55868] = 8'b0;
    XRAM[55869] = 8'b0;
    XRAM[55870] = 8'b0;
    XRAM[55871] = 8'b0;
    XRAM[55872] = 8'b0;
    XRAM[55873] = 8'b0;
    XRAM[55874] = 8'b0;
    XRAM[55875] = 8'b0;
    XRAM[55876] = 8'b0;
    XRAM[55877] = 8'b0;
    XRAM[55878] = 8'b0;
    XRAM[55879] = 8'b0;
    XRAM[55880] = 8'b0;
    XRAM[55881] = 8'b0;
    XRAM[55882] = 8'b0;
    XRAM[55883] = 8'b0;
    XRAM[55884] = 8'b0;
    XRAM[55885] = 8'b0;
    XRAM[55886] = 8'b0;
    XRAM[55887] = 8'b0;
    XRAM[55888] = 8'b0;
    XRAM[55889] = 8'b0;
    XRAM[55890] = 8'b0;
    XRAM[55891] = 8'b0;
    XRAM[55892] = 8'b0;
    XRAM[55893] = 8'b0;
    XRAM[55894] = 8'b0;
    XRAM[55895] = 8'b0;
    XRAM[55896] = 8'b0;
    XRAM[55897] = 8'b0;
    XRAM[55898] = 8'b0;
    XRAM[55899] = 8'b0;
    XRAM[55900] = 8'b0;
    XRAM[55901] = 8'b0;
    XRAM[55902] = 8'b0;
    XRAM[55903] = 8'b0;
    XRAM[55904] = 8'b0;
    XRAM[55905] = 8'b0;
    XRAM[55906] = 8'b0;
    XRAM[55907] = 8'b0;
    XRAM[55908] = 8'b0;
    XRAM[55909] = 8'b0;
    XRAM[55910] = 8'b0;
    XRAM[55911] = 8'b0;
    XRAM[55912] = 8'b0;
    XRAM[55913] = 8'b0;
    XRAM[55914] = 8'b0;
    XRAM[55915] = 8'b0;
    XRAM[55916] = 8'b0;
    XRAM[55917] = 8'b0;
    XRAM[55918] = 8'b0;
    XRAM[55919] = 8'b0;
    XRAM[55920] = 8'b0;
    XRAM[55921] = 8'b0;
    XRAM[55922] = 8'b0;
    XRAM[55923] = 8'b0;
    XRAM[55924] = 8'b0;
    XRAM[55925] = 8'b0;
    XRAM[55926] = 8'b0;
    XRAM[55927] = 8'b0;
    XRAM[55928] = 8'b0;
    XRAM[55929] = 8'b0;
    XRAM[55930] = 8'b0;
    XRAM[55931] = 8'b0;
    XRAM[55932] = 8'b0;
    XRAM[55933] = 8'b0;
    XRAM[55934] = 8'b0;
    XRAM[55935] = 8'b0;
    XRAM[55936] = 8'b0;
    XRAM[55937] = 8'b0;
    XRAM[55938] = 8'b0;
    XRAM[55939] = 8'b0;
    XRAM[55940] = 8'b0;
    XRAM[55941] = 8'b0;
    XRAM[55942] = 8'b0;
    XRAM[55943] = 8'b0;
    XRAM[55944] = 8'b0;
    XRAM[55945] = 8'b0;
    XRAM[55946] = 8'b0;
    XRAM[55947] = 8'b0;
    XRAM[55948] = 8'b0;
    XRAM[55949] = 8'b0;
    XRAM[55950] = 8'b0;
    XRAM[55951] = 8'b0;
    XRAM[55952] = 8'b0;
    XRAM[55953] = 8'b0;
    XRAM[55954] = 8'b0;
    XRAM[55955] = 8'b0;
    XRAM[55956] = 8'b0;
    XRAM[55957] = 8'b0;
    XRAM[55958] = 8'b0;
    XRAM[55959] = 8'b0;
    XRAM[55960] = 8'b0;
    XRAM[55961] = 8'b0;
    XRAM[55962] = 8'b0;
    XRAM[55963] = 8'b0;
    XRAM[55964] = 8'b0;
    XRAM[55965] = 8'b0;
    XRAM[55966] = 8'b0;
    XRAM[55967] = 8'b0;
    XRAM[55968] = 8'b0;
    XRAM[55969] = 8'b0;
    XRAM[55970] = 8'b0;
    XRAM[55971] = 8'b0;
    XRAM[55972] = 8'b0;
    XRAM[55973] = 8'b0;
    XRAM[55974] = 8'b0;
    XRAM[55975] = 8'b0;
    XRAM[55976] = 8'b0;
    XRAM[55977] = 8'b0;
    XRAM[55978] = 8'b0;
    XRAM[55979] = 8'b0;
    XRAM[55980] = 8'b0;
    XRAM[55981] = 8'b0;
    XRAM[55982] = 8'b0;
    XRAM[55983] = 8'b0;
    XRAM[55984] = 8'b0;
    XRAM[55985] = 8'b0;
    XRAM[55986] = 8'b0;
    XRAM[55987] = 8'b0;
    XRAM[55988] = 8'b0;
    XRAM[55989] = 8'b0;
    XRAM[55990] = 8'b0;
    XRAM[55991] = 8'b0;
    XRAM[55992] = 8'b0;
    XRAM[55993] = 8'b0;
    XRAM[55994] = 8'b0;
    XRAM[55995] = 8'b0;
    XRAM[55996] = 8'b0;
    XRAM[55997] = 8'b0;
    XRAM[55998] = 8'b0;
    XRAM[55999] = 8'b0;
    XRAM[56000] = 8'b0;
    XRAM[56001] = 8'b0;
    XRAM[56002] = 8'b0;
    XRAM[56003] = 8'b0;
    XRAM[56004] = 8'b0;
    XRAM[56005] = 8'b0;
    XRAM[56006] = 8'b0;
    XRAM[56007] = 8'b0;
    XRAM[56008] = 8'b0;
    XRAM[56009] = 8'b0;
    XRAM[56010] = 8'b0;
    XRAM[56011] = 8'b0;
    XRAM[56012] = 8'b0;
    XRAM[56013] = 8'b0;
    XRAM[56014] = 8'b0;
    XRAM[56015] = 8'b0;
    XRAM[56016] = 8'b0;
    XRAM[56017] = 8'b0;
    XRAM[56018] = 8'b0;
    XRAM[56019] = 8'b0;
    XRAM[56020] = 8'b0;
    XRAM[56021] = 8'b0;
    XRAM[56022] = 8'b0;
    XRAM[56023] = 8'b0;
    XRAM[56024] = 8'b0;
    XRAM[56025] = 8'b0;
    XRAM[56026] = 8'b0;
    XRAM[56027] = 8'b0;
    XRAM[56028] = 8'b0;
    XRAM[56029] = 8'b0;
    XRAM[56030] = 8'b0;
    XRAM[56031] = 8'b0;
    XRAM[56032] = 8'b0;
    XRAM[56033] = 8'b0;
    XRAM[56034] = 8'b0;
    XRAM[56035] = 8'b0;
    XRAM[56036] = 8'b0;
    XRAM[56037] = 8'b0;
    XRAM[56038] = 8'b0;
    XRAM[56039] = 8'b0;
    XRAM[56040] = 8'b0;
    XRAM[56041] = 8'b0;
    XRAM[56042] = 8'b0;
    XRAM[56043] = 8'b0;
    XRAM[56044] = 8'b0;
    XRAM[56045] = 8'b0;
    XRAM[56046] = 8'b0;
    XRAM[56047] = 8'b0;
    XRAM[56048] = 8'b0;
    XRAM[56049] = 8'b0;
    XRAM[56050] = 8'b0;
    XRAM[56051] = 8'b0;
    XRAM[56052] = 8'b0;
    XRAM[56053] = 8'b0;
    XRAM[56054] = 8'b0;
    XRAM[56055] = 8'b0;
    XRAM[56056] = 8'b0;
    XRAM[56057] = 8'b0;
    XRAM[56058] = 8'b0;
    XRAM[56059] = 8'b0;
    XRAM[56060] = 8'b0;
    XRAM[56061] = 8'b0;
    XRAM[56062] = 8'b0;
    XRAM[56063] = 8'b0;
    XRAM[56064] = 8'b0;
    XRAM[56065] = 8'b0;
    XRAM[56066] = 8'b0;
    XRAM[56067] = 8'b0;
    XRAM[56068] = 8'b0;
    XRAM[56069] = 8'b0;
    XRAM[56070] = 8'b0;
    XRAM[56071] = 8'b0;
    XRAM[56072] = 8'b0;
    XRAM[56073] = 8'b0;
    XRAM[56074] = 8'b0;
    XRAM[56075] = 8'b0;
    XRAM[56076] = 8'b0;
    XRAM[56077] = 8'b0;
    XRAM[56078] = 8'b0;
    XRAM[56079] = 8'b0;
    XRAM[56080] = 8'b0;
    XRAM[56081] = 8'b0;
    XRAM[56082] = 8'b0;
    XRAM[56083] = 8'b0;
    XRAM[56084] = 8'b0;
    XRAM[56085] = 8'b0;
    XRAM[56086] = 8'b0;
    XRAM[56087] = 8'b0;
    XRAM[56088] = 8'b0;
    XRAM[56089] = 8'b0;
    XRAM[56090] = 8'b0;
    XRAM[56091] = 8'b0;
    XRAM[56092] = 8'b0;
    XRAM[56093] = 8'b0;
    XRAM[56094] = 8'b0;
    XRAM[56095] = 8'b0;
    XRAM[56096] = 8'b0;
    XRAM[56097] = 8'b0;
    XRAM[56098] = 8'b0;
    XRAM[56099] = 8'b0;
    XRAM[56100] = 8'b0;
    XRAM[56101] = 8'b0;
    XRAM[56102] = 8'b0;
    XRAM[56103] = 8'b0;
    XRAM[56104] = 8'b0;
    XRAM[56105] = 8'b0;
    XRAM[56106] = 8'b0;
    XRAM[56107] = 8'b0;
    XRAM[56108] = 8'b0;
    XRAM[56109] = 8'b0;
    XRAM[56110] = 8'b0;
    XRAM[56111] = 8'b0;
    XRAM[56112] = 8'b0;
    XRAM[56113] = 8'b0;
    XRAM[56114] = 8'b0;
    XRAM[56115] = 8'b0;
    XRAM[56116] = 8'b0;
    XRAM[56117] = 8'b0;
    XRAM[56118] = 8'b0;
    XRAM[56119] = 8'b0;
    XRAM[56120] = 8'b0;
    XRAM[56121] = 8'b0;
    XRAM[56122] = 8'b0;
    XRAM[56123] = 8'b0;
    XRAM[56124] = 8'b0;
    XRAM[56125] = 8'b0;
    XRAM[56126] = 8'b0;
    XRAM[56127] = 8'b0;
    XRAM[56128] = 8'b0;
    XRAM[56129] = 8'b0;
    XRAM[56130] = 8'b0;
    XRAM[56131] = 8'b0;
    XRAM[56132] = 8'b0;
    XRAM[56133] = 8'b0;
    XRAM[56134] = 8'b0;
    XRAM[56135] = 8'b0;
    XRAM[56136] = 8'b0;
    XRAM[56137] = 8'b0;
    XRAM[56138] = 8'b0;
    XRAM[56139] = 8'b0;
    XRAM[56140] = 8'b0;
    XRAM[56141] = 8'b0;
    XRAM[56142] = 8'b0;
    XRAM[56143] = 8'b0;
    XRAM[56144] = 8'b0;
    XRAM[56145] = 8'b0;
    XRAM[56146] = 8'b0;
    XRAM[56147] = 8'b0;
    XRAM[56148] = 8'b0;
    XRAM[56149] = 8'b0;
    XRAM[56150] = 8'b0;
    XRAM[56151] = 8'b0;
    XRAM[56152] = 8'b0;
    XRAM[56153] = 8'b0;
    XRAM[56154] = 8'b0;
    XRAM[56155] = 8'b0;
    XRAM[56156] = 8'b0;
    XRAM[56157] = 8'b0;
    XRAM[56158] = 8'b0;
    XRAM[56159] = 8'b0;
    XRAM[56160] = 8'b0;
    XRAM[56161] = 8'b0;
    XRAM[56162] = 8'b0;
    XRAM[56163] = 8'b0;
    XRAM[56164] = 8'b0;
    XRAM[56165] = 8'b0;
    XRAM[56166] = 8'b0;
    XRAM[56167] = 8'b0;
    XRAM[56168] = 8'b0;
    XRAM[56169] = 8'b0;
    XRAM[56170] = 8'b0;
    XRAM[56171] = 8'b0;
    XRAM[56172] = 8'b0;
    XRAM[56173] = 8'b0;
    XRAM[56174] = 8'b0;
    XRAM[56175] = 8'b0;
    XRAM[56176] = 8'b0;
    XRAM[56177] = 8'b0;
    XRAM[56178] = 8'b0;
    XRAM[56179] = 8'b0;
    XRAM[56180] = 8'b0;
    XRAM[56181] = 8'b0;
    XRAM[56182] = 8'b0;
    XRAM[56183] = 8'b0;
    XRAM[56184] = 8'b0;
    XRAM[56185] = 8'b0;
    XRAM[56186] = 8'b0;
    XRAM[56187] = 8'b0;
    XRAM[56188] = 8'b0;
    XRAM[56189] = 8'b0;
    XRAM[56190] = 8'b0;
    XRAM[56191] = 8'b0;
    XRAM[56192] = 8'b0;
    XRAM[56193] = 8'b0;
    XRAM[56194] = 8'b0;
    XRAM[56195] = 8'b0;
    XRAM[56196] = 8'b0;
    XRAM[56197] = 8'b0;
    XRAM[56198] = 8'b0;
    XRAM[56199] = 8'b0;
    XRAM[56200] = 8'b0;
    XRAM[56201] = 8'b0;
    XRAM[56202] = 8'b0;
    XRAM[56203] = 8'b0;
    XRAM[56204] = 8'b0;
    XRAM[56205] = 8'b0;
    XRAM[56206] = 8'b0;
    XRAM[56207] = 8'b0;
    XRAM[56208] = 8'b0;
    XRAM[56209] = 8'b0;
    XRAM[56210] = 8'b0;
    XRAM[56211] = 8'b0;
    XRAM[56212] = 8'b0;
    XRAM[56213] = 8'b0;
    XRAM[56214] = 8'b0;
    XRAM[56215] = 8'b0;
    XRAM[56216] = 8'b0;
    XRAM[56217] = 8'b0;
    XRAM[56218] = 8'b0;
    XRAM[56219] = 8'b0;
    XRAM[56220] = 8'b0;
    XRAM[56221] = 8'b0;
    XRAM[56222] = 8'b0;
    XRAM[56223] = 8'b0;
    XRAM[56224] = 8'b0;
    XRAM[56225] = 8'b0;
    XRAM[56226] = 8'b0;
    XRAM[56227] = 8'b0;
    XRAM[56228] = 8'b0;
    XRAM[56229] = 8'b0;
    XRAM[56230] = 8'b0;
    XRAM[56231] = 8'b0;
    XRAM[56232] = 8'b0;
    XRAM[56233] = 8'b0;
    XRAM[56234] = 8'b0;
    XRAM[56235] = 8'b0;
    XRAM[56236] = 8'b0;
    XRAM[56237] = 8'b0;
    XRAM[56238] = 8'b0;
    XRAM[56239] = 8'b0;
    XRAM[56240] = 8'b0;
    XRAM[56241] = 8'b0;
    XRAM[56242] = 8'b0;
    XRAM[56243] = 8'b0;
    XRAM[56244] = 8'b0;
    XRAM[56245] = 8'b0;
    XRAM[56246] = 8'b0;
    XRAM[56247] = 8'b0;
    XRAM[56248] = 8'b0;
    XRAM[56249] = 8'b0;
    XRAM[56250] = 8'b0;
    XRAM[56251] = 8'b0;
    XRAM[56252] = 8'b0;
    XRAM[56253] = 8'b0;
    XRAM[56254] = 8'b0;
    XRAM[56255] = 8'b0;
    XRAM[56256] = 8'b0;
    XRAM[56257] = 8'b0;
    XRAM[56258] = 8'b0;
    XRAM[56259] = 8'b0;
    XRAM[56260] = 8'b0;
    XRAM[56261] = 8'b0;
    XRAM[56262] = 8'b0;
    XRAM[56263] = 8'b0;
    XRAM[56264] = 8'b0;
    XRAM[56265] = 8'b0;
    XRAM[56266] = 8'b0;
    XRAM[56267] = 8'b0;
    XRAM[56268] = 8'b0;
    XRAM[56269] = 8'b0;
    XRAM[56270] = 8'b0;
    XRAM[56271] = 8'b0;
    XRAM[56272] = 8'b0;
    XRAM[56273] = 8'b0;
    XRAM[56274] = 8'b0;
    XRAM[56275] = 8'b0;
    XRAM[56276] = 8'b0;
    XRAM[56277] = 8'b0;
    XRAM[56278] = 8'b0;
    XRAM[56279] = 8'b0;
    XRAM[56280] = 8'b0;
    XRAM[56281] = 8'b0;
    XRAM[56282] = 8'b0;
    XRAM[56283] = 8'b0;
    XRAM[56284] = 8'b0;
    XRAM[56285] = 8'b0;
    XRAM[56286] = 8'b0;
    XRAM[56287] = 8'b0;
    XRAM[56288] = 8'b0;
    XRAM[56289] = 8'b0;
    XRAM[56290] = 8'b0;
    XRAM[56291] = 8'b0;
    XRAM[56292] = 8'b0;
    XRAM[56293] = 8'b0;
    XRAM[56294] = 8'b0;
    XRAM[56295] = 8'b0;
    XRAM[56296] = 8'b0;
    XRAM[56297] = 8'b0;
    XRAM[56298] = 8'b0;
    XRAM[56299] = 8'b0;
    XRAM[56300] = 8'b0;
    XRAM[56301] = 8'b0;
    XRAM[56302] = 8'b0;
    XRAM[56303] = 8'b0;
    XRAM[56304] = 8'b0;
    XRAM[56305] = 8'b0;
    XRAM[56306] = 8'b0;
    XRAM[56307] = 8'b0;
    XRAM[56308] = 8'b0;
    XRAM[56309] = 8'b0;
    XRAM[56310] = 8'b0;
    XRAM[56311] = 8'b0;
    XRAM[56312] = 8'b0;
    XRAM[56313] = 8'b0;
    XRAM[56314] = 8'b0;
    XRAM[56315] = 8'b0;
    XRAM[56316] = 8'b0;
    XRAM[56317] = 8'b0;
    XRAM[56318] = 8'b0;
    XRAM[56319] = 8'b0;
    XRAM[56320] = 8'b0;
    XRAM[56321] = 8'b0;
    XRAM[56322] = 8'b0;
    XRAM[56323] = 8'b0;
    XRAM[56324] = 8'b0;
    XRAM[56325] = 8'b0;
    XRAM[56326] = 8'b0;
    XRAM[56327] = 8'b0;
    XRAM[56328] = 8'b0;
    XRAM[56329] = 8'b0;
    XRAM[56330] = 8'b0;
    XRAM[56331] = 8'b0;
    XRAM[56332] = 8'b0;
    XRAM[56333] = 8'b0;
    XRAM[56334] = 8'b0;
    XRAM[56335] = 8'b0;
    XRAM[56336] = 8'b0;
    XRAM[56337] = 8'b0;
    XRAM[56338] = 8'b0;
    XRAM[56339] = 8'b0;
    XRAM[56340] = 8'b0;
    XRAM[56341] = 8'b0;
    XRAM[56342] = 8'b0;
    XRAM[56343] = 8'b0;
    XRAM[56344] = 8'b0;
    XRAM[56345] = 8'b0;
    XRAM[56346] = 8'b0;
    XRAM[56347] = 8'b0;
    XRAM[56348] = 8'b0;
    XRAM[56349] = 8'b0;
    XRAM[56350] = 8'b0;
    XRAM[56351] = 8'b0;
    XRAM[56352] = 8'b0;
    XRAM[56353] = 8'b0;
    XRAM[56354] = 8'b0;
    XRAM[56355] = 8'b0;
    XRAM[56356] = 8'b0;
    XRAM[56357] = 8'b0;
    XRAM[56358] = 8'b0;
    XRAM[56359] = 8'b0;
    XRAM[56360] = 8'b0;
    XRAM[56361] = 8'b0;
    XRAM[56362] = 8'b0;
    XRAM[56363] = 8'b0;
    XRAM[56364] = 8'b0;
    XRAM[56365] = 8'b0;
    XRAM[56366] = 8'b0;
    XRAM[56367] = 8'b0;
    XRAM[56368] = 8'b0;
    XRAM[56369] = 8'b0;
    XRAM[56370] = 8'b0;
    XRAM[56371] = 8'b0;
    XRAM[56372] = 8'b0;
    XRAM[56373] = 8'b0;
    XRAM[56374] = 8'b0;
    XRAM[56375] = 8'b0;
    XRAM[56376] = 8'b0;
    XRAM[56377] = 8'b0;
    XRAM[56378] = 8'b0;
    XRAM[56379] = 8'b0;
    XRAM[56380] = 8'b0;
    XRAM[56381] = 8'b0;
    XRAM[56382] = 8'b0;
    XRAM[56383] = 8'b0;
    XRAM[56384] = 8'b0;
    XRAM[56385] = 8'b0;
    XRAM[56386] = 8'b0;
    XRAM[56387] = 8'b0;
    XRAM[56388] = 8'b0;
    XRAM[56389] = 8'b0;
    XRAM[56390] = 8'b0;
    XRAM[56391] = 8'b0;
    XRAM[56392] = 8'b0;
    XRAM[56393] = 8'b0;
    XRAM[56394] = 8'b0;
    XRAM[56395] = 8'b0;
    XRAM[56396] = 8'b0;
    XRAM[56397] = 8'b0;
    XRAM[56398] = 8'b0;
    XRAM[56399] = 8'b0;
    XRAM[56400] = 8'b0;
    XRAM[56401] = 8'b0;
    XRAM[56402] = 8'b0;
    XRAM[56403] = 8'b0;
    XRAM[56404] = 8'b0;
    XRAM[56405] = 8'b0;
    XRAM[56406] = 8'b0;
    XRAM[56407] = 8'b0;
    XRAM[56408] = 8'b0;
    XRAM[56409] = 8'b0;
    XRAM[56410] = 8'b0;
    XRAM[56411] = 8'b0;
    XRAM[56412] = 8'b0;
    XRAM[56413] = 8'b0;
    XRAM[56414] = 8'b0;
    XRAM[56415] = 8'b0;
    XRAM[56416] = 8'b0;
    XRAM[56417] = 8'b0;
    XRAM[56418] = 8'b0;
    XRAM[56419] = 8'b0;
    XRAM[56420] = 8'b0;
    XRAM[56421] = 8'b0;
    XRAM[56422] = 8'b0;
    XRAM[56423] = 8'b0;
    XRAM[56424] = 8'b0;
    XRAM[56425] = 8'b0;
    XRAM[56426] = 8'b0;
    XRAM[56427] = 8'b0;
    XRAM[56428] = 8'b0;
    XRAM[56429] = 8'b0;
    XRAM[56430] = 8'b0;
    XRAM[56431] = 8'b0;
    XRAM[56432] = 8'b0;
    XRAM[56433] = 8'b0;
    XRAM[56434] = 8'b0;
    XRAM[56435] = 8'b0;
    XRAM[56436] = 8'b0;
    XRAM[56437] = 8'b0;
    XRAM[56438] = 8'b0;
    XRAM[56439] = 8'b0;
    XRAM[56440] = 8'b0;
    XRAM[56441] = 8'b0;
    XRAM[56442] = 8'b0;
    XRAM[56443] = 8'b0;
    XRAM[56444] = 8'b0;
    XRAM[56445] = 8'b0;
    XRAM[56446] = 8'b0;
    XRAM[56447] = 8'b0;
    XRAM[56448] = 8'b0;
    XRAM[56449] = 8'b0;
    XRAM[56450] = 8'b0;
    XRAM[56451] = 8'b0;
    XRAM[56452] = 8'b0;
    XRAM[56453] = 8'b0;
    XRAM[56454] = 8'b0;
    XRAM[56455] = 8'b0;
    XRAM[56456] = 8'b0;
    XRAM[56457] = 8'b0;
    XRAM[56458] = 8'b0;
    XRAM[56459] = 8'b0;
    XRAM[56460] = 8'b0;
    XRAM[56461] = 8'b0;
    XRAM[56462] = 8'b0;
    XRAM[56463] = 8'b0;
    XRAM[56464] = 8'b0;
    XRAM[56465] = 8'b0;
    XRAM[56466] = 8'b0;
    XRAM[56467] = 8'b0;
    XRAM[56468] = 8'b0;
    XRAM[56469] = 8'b0;
    XRAM[56470] = 8'b0;
    XRAM[56471] = 8'b0;
    XRAM[56472] = 8'b0;
    XRAM[56473] = 8'b0;
    XRAM[56474] = 8'b0;
    XRAM[56475] = 8'b0;
    XRAM[56476] = 8'b0;
    XRAM[56477] = 8'b0;
    XRAM[56478] = 8'b0;
    XRAM[56479] = 8'b0;
    XRAM[56480] = 8'b0;
    XRAM[56481] = 8'b0;
    XRAM[56482] = 8'b0;
    XRAM[56483] = 8'b0;
    XRAM[56484] = 8'b0;
    XRAM[56485] = 8'b0;
    XRAM[56486] = 8'b0;
    XRAM[56487] = 8'b0;
    XRAM[56488] = 8'b0;
    XRAM[56489] = 8'b0;
    XRAM[56490] = 8'b0;
    XRAM[56491] = 8'b0;
    XRAM[56492] = 8'b0;
    XRAM[56493] = 8'b0;
    XRAM[56494] = 8'b0;
    XRAM[56495] = 8'b0;
    XRAM[56496] = 8'b0;
    XRAM[56497] = 8'b0;
    XRAM[56498] = 8'b0;
    XRAM[56499] = 8'b0;
    XRAM[56500] = 8'b0;
    XRAM[56501] = 8'b0;
    XRAM[56502] = 8'b0;
    XRAM[56503] = 8'b0;
    XRAM[56504] = 8'b0;
    XRAM[56505] = 8'b0;
    XRAM[56506] = 8'b0;
    XRAM[56507] = 8'b0;
    XRAM[56508] = 8'b0;
    XRAM[56509] = 8'b0;
    XRAM[56510] = 8'b0;
    XRAM[56511] = 8'b0;
    XRAM[56512] = 8'b0;
    XRAM[56513] = 8'b0;
    XRAM[56514] = 8'b0;
    XRAM[56515] = 8'b0;
    XRAM[56516] = 8'b0;
    XRAM[56517] = 8'b0;
    XRAM[56518] = 8'b0;
    XRAM[56519] = 8'b0;
    XRAM[56520] = 8'b0;
    XRAM[56521] = 8'b0;
    XRAM[56522] = 8'b0;
    XRAM[56523] = 8'b0;
    XRAM[56524] = 8'b0;
    XRAM[56525] = 8'b0;
    XRAM[56526] = 8'b0;
    XRAM[56527] = 8'b0;
    XRAM[56528] = 8'b0;
    XRAM[56529] = 8'b0;
    XRAM[56530] = 8'b0;
    XRAM[56531] = 8'b0;
    XRAM[56532] = 8'b0;
    XRAM[56533] = 8'b0;
    XRAM[56534] = 8'b0;
    XRAM[56535] = 8'b0;
    XRAM[56536] = 8'b0;
    XRAM[56537] = 8'b0;
    XRAM[56538] = 8'b0;
    XRAM[56539] = 8'b0;
    XRAM[56540] = 8'b0;
    XRAM[56541] = 8'b0;
    XRAM[56542] = 8'b0;
    XRAM[56543] = 8'b0;
    XRAM[56544] = 8'b0;
    XRAM[56545] = 8'b0;
    XRAM[56546] = 8'b0;
    XRAM[56547] = 8'b0;
    XRAM[56548] = 8'b0;
    XRAM[56549] = 8'b0;
    XRAM[56550] = 8'b0;
    XRAM[56551] = 8'b0;
    XRAM[56552] = 8'b0;
    XRAM[56553] = 8'b0;
    XRAM[56554] = 8'b0;
    XRAM[56555] = 8'b0;
    XRAM[56556] = 8'b0;
    XRAM[56557] = 8'b0;
    XRAM[56558] = 8'b0;
    XRAM[56559] = 8'b0;
    XRAM[56560] = 8'b0;
    XRAM[56561] = 8'b0;
    XRAM[56562] = 8'b0;
    XRAM[56563] = 8'b0;
    XRAM[56564] = 8'b0;
    XRAM[56565] = 8'b0;
    XRAM[56566] = 8'b0;
    XRAM[56567] = 8'b0;
    XRAM[56568] = 8'b0;
    XRAM[56569] = 8'b0;
    XRAM[56570] = 8'b0;
    XRAM[56571] = 8'b0;
    XRAM[56572] = 8'b0;
    XRAM[56573] = 8'b0;
    XRAM[56574] = 8'b0;
    XRAM[56575] = 8'b0;
    XRAM[56576] = 8'b0;
    XRAM[56577] = 8'b0;
    XRAM[56578] = 8'b0;
    XRAM[56579] = 8'b0;
    XRAM[56580] = 8'b0;
    XRAM[56581] = 8'b0;
    XRAM[56582] = 8'b0;
    XRAM[56583] = 8'b0;
    XRAM[56584] = 8'b0;
    XRAM[56585] = 8'b0;
    XRAM[56586] = 8'b0;
    XRAM[56587] = 8'b0;
    XRAM[56588] = 8'b0;
    XRAM[56589] = 8'b0;
    XRAM[56590] = 8'b0;
    XRAM[56591] = 8'b0;
    XRAM[56592] = 8'b0;
    XRAM[56593] = 8'b0;
    XRAM[56594] = 8'b0;
    XRAM[56595] = 8'b0;
    XRAM[56596] = 8'b0;
    XRAM[56597] = 8'b0;
    XRAM[56598] = 8'b0;
    XRAM[56599] = 8'b0;
    XRAM[56600] = 8'b0;
    XRAM[56601] = 8'b0;
    XRAM[56602] = 8'b0;
    XRAM[56603] = 8'b0;
    XRAM[56604] = 8'b0;
    XRAM[56605] = 8'b0;
    XRAM[56606] = 8'b0;
    XRAM[56607] = 8'b0;
    XRAM[56608] = 8'b0;
    XRAM[56609] = 8'b0;
    XRAM[56610] = 8'b0;
    XRAM[56611] = 8'b0;
    XRAM[56612] = 8'b0;
    XRAM[56613] = 8'b0;
    XRAM[56614] = 8'b0;
    XRAM[56615] = 8'b0;
    XRAM[56616] = 8'b0;
    XRAM[56617] = 8'b0;
    XRAM[56618] = 8'b0;
    XRAM[56619] = 8'b0;
    XRAM[56620] = 8'b0;
    XRAM[56621] = 8'b0;
    XRAM[56622] = 8'b0;
    XRAM[56623] = 8'b0;
    XRAM[56624] = 8'b0;
    XRAM[56625] = 8'b0;
    XRAM[56626] = 8'b0;
    XRAM[56627] = 8'b0;
    XRAM[56628] = 8'b0;
    XRAM[56629] = 8'b0;
    XRAM[56630] = 8'b0;
    XRAM[56631] = 8'b0;
    XRAM[56632] = 8'b0;
    XRAM[56633] = 8'b0;
    XRAM[56634] = 8'b0;
    XRAM[56635] = 8'b0;
    XRAM[56636] = 8'b0;
    XRAM[56637] = 8'b0;
    XRAM[56638] = 8'b0;
    XRAM[56639] = 8'b0;
    XRAM[56640] = 8'b0;
    XRAM[56641] = 8'b0;
    XRAM[56642] = 8'b0;
    XRAM[56643] = 8'b0;
    XRAM[56644] = 8'b0;
    XRAM[56645] = 8'b0;
    XRAM[56646] = 8'b0;
    XRAM[56647] = 8'b0;
    XRAM[56648] = 8'b0;
    XRAM[56649] = 8'b0;
    XRAM[56650] = 8'b0;
    XRAM[56651] = 8'b0;
    XRAM[56652] = 8'b0;
    XRAM[56653] = 8'b0;
    XRAM[56654] = 8'b0;
    XRAM[56655] = 8'b0;
    XRAM[56656] = 8'b0;
    XRAM[56657] = 8'b0;
    XRAM[56658] = 8'b0;
    XRAM[56659] = 8'b0;
    XRAM[56660] = 8'b0;
    XRAM[56661] = 8'b0;
    XRAM[56662] = 8'b0;
    XRAM[56663] = 8'b0;
    XRAM[56664] = 8'b0;
    XRAM[56665] = 8'b0;
    XRAM[56666] = 8'b0;
    XRAM[56667] = 8'b0;
    XRAM[56668] = 8'b0;
    XRAM[56669] = 8'b0;
    XRAM[56670] = 8'b0;
    XRAM[56671] = 8'b0;
    XRAM[56672] = 8'b0;
    XRAM[56673] = 8'b0;
    XRAM[56674] = 8'b0;
    XRAM[56675] = 8'b0;
    XRAM[56676] = 8'b0;
    XRAM[56677] = 8'b0;
    XRAM[56678] = 8'b0;
    XRAM[56679] = 8'b0;
    XRAM[56680] = 8'b0;
    XRAM[56681] = 8'b0;
    XRAM[56682] = 8'b0;
    XRAM[56683] = 8'b0;
    XRAM[56684] = 8'b0;
    XRAM[56685] = 8'b0;
    XRAM[56686] = 8'b0;
    XRAM[56687] = 8'b0;
    XRAM[56688] = 8'b0;
    XRAM[56689] = 8'b0;
    XRAM[56690] = 8'b0;
    XRAM[56691] = 8'b0;
    XRAM[56692] = 8'b0;
    XRAM[56693] = 8'b0;
    XRAM[56694] = 8'b0;
    XRAM[56695] = 8'b0;
    XRAM[56696] = 8'b0;
    XRAM[56697] = 8'b0;
    XRAM[56698] = 8'b0;
    XRAM[56699] = 8'b0;
    XRAM[56700] = 8'b0;
    XRAM[56701] = 8'b0;
    XRAM[56702] = 8'b0;
    XRAM[56703] = 8'b0;
    XRAM[56704] = 8'b0;
    XRAM[56705] = 8'b0;
    XRAM[56706] = 8'b0;
    XRAM[56707] = 8'b0;
    XRAM[56708] = 8'b0;
    XRAM[56709] = 8'b0;
    XRAM[56710] = 8'b0;
    XRAM[56711] = 8'b0;
    XRAM[56712] = 8'b0;
    XRAM[56713] = 8'b0;
    XRAM[56714] = 8'b0;
    XRAM[56715] = 8'b0;
    XRAM[56716] = 8'b0;
    XRAM[56717] = 8'b0;
    XRAM[56718] = 8'b0;
    XRAM[56719] = 8'b0;
    XRAM[56720] = 8'b0;
    XRAM[56721] = 8'b0;
    XRAM[56722] = 8'b0;
    XRAM[56723] = 8'b0;
    XRAM[56724] = 8'b0;
    XRAM[56725] = 8'b0;
    XRAM[56726] = 8'b0;
    XRAM[56727] = 8'b0;
    XRAM[56728] = 8'b0;
    XRAM[56729] = 8'b0;
    XRAM[56730] = 8'b0;
    XRAM[56731] = 8'b0;
    XRAM[56732] = 8'b0;
    XRAM[56733] = 8'b0;
    XRAM[56734] = 8'b0;
    XRAM[56735] = 8'b0;
    XRAM[56736] = 8'b0;
    XRAM[56737] = 8'b0;
    XRAM[56738] = 8'b0;
    XRAM[56739] = 8'b0;
    XRAM[56740] = 8'b0;
    XRAM[56741] = 8'b0;
    XRAM[56742] = 8'b0;
    XRAM[56743] = 8'b0;
    XRAM[56744] = 8'b0;
    XRAM[56745] = 8'b0;
    XRAM[56746] = 8'b0;
    XRAM[56747] = 8'b0;
    XRAM[56748] = 8'b0;
    XRAM[56749] = 8'b0;
    XRAM[56750] = 8'b0;
    XRAM[56751] = 8'b0;
    XRAM[56752] = 8'b0;
    XRAM[56753] = 8'b0;
    XRAM[56754] = 8'b0;
    XRAM[56755] = 8'b0;
    XRAM[56756] = 8'b0;
    XRAM[56757] = 8'b0;
    XRAM[56758] = 8'b0;
    XRAM[56759] = 8'b0;
    XRAM[56760] = 8'b0;
    XRAM[56761] = 8'b0;
    XRAM[56762] = 8'b0;
    XRAM[56763] = 8'b0;
    XRAM[56764] = 8'b0;
    XRAM[56765] = 8'b0;
    XRAM[56766] = 8'b0;
    XRAM[56767] = 8'b0;
    XRAM[56768] = 8'b0;
    XRAM[56769] = 8'b0;
    XRAM[56770] = 8'b0;
    XRAM[56771] = 8'b0;
    XRAM[56772] = 8'b0;
    XRAM[56773] = 8'b0;
    XRAM[56774] = 8'b0;
    XRAM[56775] = 8'b0;
    XRAM[56776] = 8'b0;
    XRAM[56777] = 8'b0;
    XRAM[56778] = 8'b0;
    XRAM[56779] = 8'b0;
    XRAM[56780] = 8'b0;
    XRAM[56781] = 8'b0;
    XRAM[56782] = 8'b0;
    XRAM[56783] = 8'b0;
    XRAM[56784] = 8'b0;
    XRAM[56785] = 8'b0;
    XRAM[56786] = 8'b0;
    XRAM[56787] = 8'b0;
    XRAM[56788] = 8'b0;
    XRAM[56789] = 8'b0;
    XRAM[56790] = 8'b0;
    XRAM[56791] = 8'b0;
    XRAM[56792] = 8'b0;
    XRAM[56793] = 8'b0;
    XRAM[56794] = 8'b0;
    XRAM[56795] = 8'b0;
    XRAM[56796] = 8'b0;
    XRAM[56797] = 8'b0;
    XRAM[56798] = 8'b0;
    XRAM[56799] = 8'b0;
    XRAM[56800] = 8'b0;
    XRAM[56801] = 8'b0;
    XRAM[56802] = 8'b0;
    XRAM[56803] = 8'b0;
    XRAM[56804] = 8'b0;
    XRAM[56805] = 8'b0;
    XRAM[56806] = 8'b0;
    XRAM[56807] = 8'b0;
    XRAM[56808] = 8'b0;
    XRAM[56809] = 8'b0;
    XRAM[56810] = 8'b0;
    XRAM[56811] = 8'b0;
    XRAM[56812] = 8'b0;
    XRAM[56813] = 8'b0;
    XRAM[56814] = 8'b0;
    XRAM[56815] = 8'b0;
    XRAM[56816] = 8'b0;
    XRAM[56817] = 8'b0;
    XRAM[56818] = 8'b0;
    XRAM[56819] = 8'b0;
    XRAM[56820] = 8'b0;
    XRAM[56821] = 8'b0;
    XRAM[56822] = 8'b0;
    XRAM[56823] = 8'b0;
    XRAM[56824] = 8'b0;
    XRAM[56825] = 8'b0;
    XRAM[56826] = 8'b0;
    XRAM[56827] = 8'b0;
    XRAM[56828] = 8'b0;
    XRAM[56829] = 8'b0;
    XRAM[56830] = 8'b0;
    XRAM[56831] = 8'b0;
    XRAM[56832] = 8'b0;
    XRAM[56833] = 8'b0;
    XRAM[56834] = 8'b0;
    XRAM[56835] = 8'b0;
    XRAM[56836] = 8'b0;
    XRAM[56837] = 8'b0;
    XRAM[56838] = 8'b0;
    XRAM[56839] = 8'b0;
    XRAM[56840] = 8'b0;
    XRAM[56841] = 8'b0;
    XRAM[56842] = 8'b0;
    XRAM[56843] = 8'b0;
    XRAM[56844] = 8'b0;
    XRAM[56845] = 8'b0;
    XRAM[56846] = 8'b0;
    XRAM[56847] = 8'b0;
    XRAM[56848] = 8'b0;
    XRAM[56849] = 8'b0;
    XRAM[56850] = 8'b0;
    XRAM[56851] = 8'b0;
    XRAM[56852] = 8'b0;
    XRAM[56853] = 8'b0;
    XRAM[56854] = 8'b0;
    XRAM[56855] = 8'b0;
    XRAM[56856] = 8'b0;
    XRAM[56857] = 8'b0;
    XRAM[56858] = 8'b0;
    XRAM[56859] = 8'b0;
    XRAM[56860] = 8'b0;
    XRAM[56861] = 8'b0;
    XRAM[56862] = 8'b0;
    XRAM[56863] = 8'b0;
    XRAM[56864] = 8'b0;
    XRAM[56865] = 8'b0;
    XRAM[56866] = 8'b0;
    XRAM[56867] = 8'b0;
    XRAM[56868] = 8'b0;
    XRAM[56869] = 8'b0;
    XRAM[56870] = 8'b0;
    XRAM[56871] = 8'b0;
    XRAM[56872] = 8'b0;
    XRAM[56873] = 8'b0;
    XRAM[56874] = 8'b0;
    XRAM[56875] = 8'b0;
    XRAM[56876] = 8'b0;
    XRAM[56877] = 8'b0;
    XRAM[56878] = 8'b0;
    XRAM[56879] = 8'b0;
    XRAM[56880] = 8'b0;
    XRAM[56881] = 8'b0;
    XRAM[56882] = 8'b0;
    XRAM[56883] = 8'b0;
    XRAM[56884] = 8'b0;
    XRAM[56885] = 8'b0;
    XRAM[56886] = 8'b0;
    XRAM[56887] = 8'b0;
    XRAM[56888] = 8'b0;
    XRAM[56889] = 8'b0;
    XRAM[56890] = 8'b0;
    XRAM[56891] = 8'b0;
    XRAM[56892] = 8'b0;
    XRAM[56893] = 8'b0;
    XRAM[56894] = 8'b0;
    XRAM[56895] = 8'b0;
    XRAM[56896] = 8'b0;
    XRAM[56897] = 8'b0;
    XRAM[56898] = 8'b0;
    XRAM[56899] = 8'b0;
    XRAM[56900] = 8'b0;
    XRAM[56901] = 8'b0;
    XRAM[56902] = 8'b0;
    XRAM[56903] = 8'b0;
    XRAM[56904] = 8'b0;
    XRAM[56905] = 8'b0;
    XRAM[56906] = 8'b0;
    XRAM[56907] = 8'b0;
    XRAM[56908] = 8'b0;
    XRAM[56909] = 8'b0;
    XRAM[56910] = 8'b0;
    XRAM[56911] = 8'b0;
    XRAM[56912] = 8'b0;
    XRAM[56913] = 8'b0;
    XRAM[56914] = 8'b0;
    XRAM[56915] = 8'b0;
    XRAM[56916] = 8'b0;
    XRAM[56917] = 8'b0;
    XRAM[56918] = 8'b0;
    XRAM[56919] = 8'b0;
    XRAM[56920] = 8'b0;
    XRAM[56921] = 8'b0;
    XRAM[56922] = 8'b0;
    XRAM[56923] = 8'b0;
    XRAM[56924] = 8'b0;
    XRAM[56925] = 8'b0;
    XRAM[56926] = 8'b0;
    XRAM[56927] = 8'b0;
    XRAM[56928] = 8'b0;
    XRAM[56929] = 8'b0;
    XRAM[56930] = 8'b0;
    XRAM[56931] = 8'b0;
    XRAM[56932] = 8'b0;
    XRAM[56933] = 8'b0;
    XRAM[56934] = 8'b0;
    XRAM[56935] = 8'b0;
    XRAM[56936] = 8'b0;
    XRAM[56937] = 8'b0;
    XRAM[56938] = 8'b0;
    XRAM[56939] = 8'b0;
    XRAM[56940] = 8'b0;
    XRAM[56941] = 8'b0;
    XRAM[56942] = 8'b0;
    XRAM[56943] = 8'b0;
    XRAM[56944] = 8'b0;
    XRAM[56945] = 8'b0;
    XRAM[56946] = 8'b0;
    XRAM[56947] = 8'b0;
    XRAM[56948] = 8'b0;
    XRAM[56949] = 8'b0;
    XRAM[56950] = 8'b0;
    XRAM[56951] = 8'b0;
    XRAM[56952] = 8'b0;
    XRAM[56953] = 8'b0;
    XRAM[56954] = 8'b0;
    XRAM[56955] = 8'b0;
    XRAM[56956] = 8'b0;
    XRAM[56957] = 8'b0;
    XRAM[56958] = 8'b0;
    XRAM[56959] = 8'b0;
    XRAM[56960] = 8'b0;
    XRAM[56961] = 8'b0;
    XRAM[56962] = 8'b0;
    XRAM[56963] = 8'b0;
    XRAM[56964] = 8'b0;
    XRAM[56965] = 8'b0;
    XRAM[56966] = 8'b0;
    XRAM[56967] = 8'b0;
    XRAM[56968] = 8'b0;
    XRAM[56969] = 8'b0;
    XRAM[56970] = 8'b0;
    XRAM[56971] = 8'b0;
    XRAM[56972] = 8'b0;
    XRAM[56973] = 8'b0;
    XRAM[56974] = 8'b0;
    XRAM[56975] = 8'b0;
    XRAM[56976] = 8'b0;
    XRAM[56977] = 8'b0;
    XRAM[56978] = 8'b0;
    XRAM[56979] = 8'b0;
    XRAM[56980] = 8'b0;
    XRAM[56981] = 8'b0;
    XRAM[56982] = 8'b0;
    XRAM[56983] = 8'b0;
    XRAM[56984] = 8'b0;
    XRAM[56985] = 8'b0;
    XRAM[56986] = 8'b0;
    XRAM[56987] = 8'b0;
    XRAM[56988] = 8'b0;
    XRAM[56989] = 8'b0;
    XRAM[56990] = 8'b0;
    XRAM[56991] = 8'b0;
    XRAM[56992] = 8'b0;
    XRAM[56993] = 8'b0;
    XRAM[56994] = 8'b0;
    XRAM[56995] = 8'b0;
    XRAM[56996] = 8'b0;
    XRAM[56997] = 8'b0;
    XRAM[56998] = 8'b0;
    XRAM[56999] = 8'b0;
    XRAM[57000] = 8'b0;
    XRAM[57001] = 8'b0;
    XRAM[57002] = 8'b0;
    XRAM[57003] = 8'b0;
    XRAM[57004] = 8'b0;
    XRAM[57005] = 8'b0;
    XRAM[57006] = 8'b0;
    XRAM[57007] = 8'b0;
    XRAM[57008] = 8'b0;
    XRAM[57009] = 8'b0;
    XRAM[57010] = 8'b0;
    XRAM[57011] = 8'b0;
    XRAM[57012] = 8'b0;
    XRAM[57013] = 8'b0;
    XRAM[57014] = 8'b0;
    XRAM[57015] = 8'b0;
    XRAM[57016] = 8'b0;
    XRAM[57017] = 8'b0;
    XRAM[57018] = 8'b0;
    XRAM[57019] = 8'b0;
    XRAM[57020] = 8'b0;
    XRAM[57021] = 8'b0;
    XRAM[57022] = 8'b0;
    XRAM[57023] = 8'b0;
    XRAM[57024] = 8'b0;
    XRAM[57025] = 8'b0;
    XRAM[57026] = 8'b0;
    XRAM[57027] = 8'b0;
    XRAM[57028] = 8'b0;
    XRAM[57029] = 8'b0;
    XRAM[57030] = 8'b0;
    XRAM[57031] = 8'b0;
    XRAM[57032] = 8'b0;
    XRAM[57033] = 8'b0;
    XRAM[57034] = 8'b0;
    XRAM[57035] = 8'b0;
    XRAM[57036] = 8'b0;
    XRAM[57037] = 8'b0;
    XRAM[57038] = 8'b0;
    XRAM[57039] = 8'b0;
    XRAM[57040] = 8'b0;
    XRAM[57041] = 8'b0;
    XRAM[57042] = 8'b0;
    XRAM[57043] = 8'b0;
    XRAM[57044] = 8'b0;
    XRAM[57045] = 8'b0;
    XRAM[57046] = 8'b0;
    XRAM[57047] = 8'b0;
    XRAM[57048] = 8'b0;
    XRAM[57049] = 8'b0;
    XRAM[57050] = 8'b0;
    XRAM[57051] = 8'b0;
    XRAM[57052] = 8'b0;
    XRAM[57053] = 8'b0;
    XRAM[57054] = 8'b0;
    XRAM[57055] = 8'b0;
    XRAM[57056] = 8'b0;
    XRAM[57057] = 8'b0;
    XRAM[57058] = 8'b0;
    XRAM[57059] = 8'b0;
    XRAM[57060] = 8'b0;
    XRAM[57061] = 8'b0;
    XRAM[57062] = 8'b0;
    XRAM[57063] = 8'b0;
    XRAM[57064] = 8'b0;
    XRAM[57065] = 8'b0;
    XRAM[57066] = 8'b0;
    XRAM[57067] = 8'b0;
    XRAM[57068] = 8'b0;
    XRAM[57069] = 8'b0;
    XRAM[57070] = 8'b0;
    XRAM[57071] = 8'b0;
    XRAM[57072] = 8'b0;
    XRAM[57073] = 8'b0;
    XRAM[57074] = 8'b0;
    XRAM[57075] = 8'b0;
    XRAM[57076] = 8'b0;
    XRAM[57077] = 8'b0;
    XRAM[57078] = 8'b0;
    XRAM[57079] = 8'b0;
    XRAM[57080] = 8'b0;
    XRAM[57081] = 8'b0;
    XRAM[57082] = 8'b0;
    XRAM[57083] = 8'b0;
    XRAM[57084] = 8'b0;
    XRAM[57085] = 8'b0;
    XRAM[57086] = 8'b0;
    XRAM[57087] = 8'b0;
    XRAM[57088] = 8'b0;
    XRAM[57089] = 8'b0;
    XRAM[57090] = 8'b0;
    XRAM[57091] = 8'b0;
    XRAM[57092] = 8'b0;
    XRAM[57093] = 8'b0;
    XRAM[57094] = 8'b0;
    XRAM[57095] = 8'b0;
    XRAM[57096] = 8'b0;
    XRAM[57097] = 8'b0;
    XRAM[57098] = 8'b0;
    XRAM[57099] = 8'b0;
    XRAM[57100] = 8'b0;
    XRAM[57101] = 8'b0;
    XRAM[57102] = 8'b0;
    XRAM[57103] = 8'b0;
    XRAM[57104] = 8'b0;
    XRAM[57105] = 8'b0;
    XRAM[57106] = 8'b0;
    XRAM[57107] = 8'b0;
    XRAM[57108] = 8'b0;
    XRAM[57109] = 8'b0;
    XRAM[57110] = 8'b0;
    XRAM[57111] = 8'b0;
    XRAM[57112] = 8'b0;
    XRAM[57113] = 8'b0;
    XRAM[57114] = 8'b0;
    XRAM[57115] = 8'b0;
    XRAM[57116] = 8'b0;
    XRAM[57117] = 8'b0;
    XRAM[57118] = 8'b0;
    XRAM[57119] = 8'b0;
    XRAM[57120] = 8'b0;
    XRAM[57121] = 8'b0;
    XRAM[57122] = 8'b0;
    XRAM[57123] = 8'b0;
    XRAM[57124] = 8'b0;
    XRAM[57125] = 8'b0;
    XRAM[57126] = 8'b0;
    XRAM[57127] = 8'b0;
    XRAM[57128] = 8'b0;
    XRAM[57129] = 8'b0;
    XRAM[57130] = 8'b0;
    XRAM[57131] = 8'b0;
    XRAM[57132] = 8'b0;
    XRAM[57133] = 8'b0;
    XRAM[57134] = 8'b0;
    XRAM[57135] = 8'b0;
    XRAM[57136] = 8'b0;
    XRAM[57137] = 8'b0;
    XRAM[57138] = 8'b0;
    XRAM[57139] = 8'b0;
    XRAM[57140] = 8'b0;
    XRAM[57141] = 8'b0;
    XRAM[57142] = 8'b0;
    XRAM[57143] = 8'b0;
    XRAM[57144] = 8'b0;
    XRAM[57145] = 8'b0;
    XRAM[57146] = 8'b0;
    XRAM[57147] = 8'b0;
    XRAM[57148] = 8'b0;
    XRAM[57149] = 8'b0;
    XRAM[57150] = 8'b0;
    XRAM[57151] = 8'b0;
    XRAM[57152] = 8'b0;
    XRAM[57153] = 8'b0;
    XRAM[57154] = 8'b0;
    XRAM[57155] = 8'b0;
    XRAM[57156] = 8'b0;
    XRAM[57157] = 8'b0;
    XRAM[57158] = 8'b0;
    XRAM[57159] = 8'b0;
    XRAM[57160] = 8'b0;
    XRAM[57161] = 8'b0;
    XRAM[57162] = 8'b0;
    XRAM[57163] = 8'b0;
    XRAM[57164] = 8'b0;
    XRAM[57165] = 8'b0;
    XRAM[57166] = 8'b0;
    XRAM[57167] = 8'b0;
    XRAM[57168] = 8'b0;
    XRAM[57169] = 8'b0;
    XRAM[57170] = 8'b0;
    XRAM[57171] = 8'b0;
    XRAM[57172] = 8'b0;
    XRAM[57173] = 8'b0;
    XRAM[57174] = 8'b0;
    XRAM[57175] = 8'b0;
    XRAM[57176] = 8'b0;
    XRAM[57177] = 8'b0;
    XRAM[57178] = 8'b0;
    XRAM[57179] = 8'b0;
    XRAM[57180] = 8'b0;
    XRAM[57181] = 8'b0;
    XRAM[57182] = 8'b0;
    XRAM[57183] = 8'b0;
    XRAM[57184] = 8'b0;
    XRAM[57185] = 8'b0;
    XRAM[57186] = 8'b0;
    XRAM[57187] = 8'b0;
    XRAM[57188] = 8'b0;
    XRAM[57189] = 8'b0;
    XRAM[57190] = 8'b0;
    XRAM[57191] = 8'b0;
    XRAM[57192] = 8'b0;
    XRAM[57193] = 8'b0;
    XRAM[57194] = 8'b0;
    XRAM[57195] = 8'b0;
    XRAM[57196] = 8'b0;
    XRAM[57197] = 8'b0;
    XRAM[57198] = 8'b0;
    XRAM[57199] = 8'b0;
    XRAM[57200] = 8'b0;
    XRAM[57201] = 8'b0;
    XRAM[57202] = 8'b0;
    XRAM[57203] = 8'b0;
    XRAM[57204] = 8'b0;
    XRAM[57205] = 8'b0;
    XRAM[57206] = 8'b0;
    XRAM[57207] = 8'b0;
    XRAM[57208] = 8'b0;
    XRAM[57209] = 8'b0;
    XRAM[57210] = 8'b0;
    XRAM[57211] = 8'b0;
    XRAM[57212] = 8'b0;
    XRAM[57213] = 8'b0;
    XRAM[57214] = 8'b0;
    XRAM[57215] = 8'b0;
    XRAM[57216] = 8'b0;
    XRAM[57217] = 8'b0;
    XRAM[57218] = 8'b0;
    XRAM[57219] = 8'b0;
    XRAM[57220] = 8'b0;
    XRAM[57221] = 8'b0;
    XRAM[57222] = 8'b0;
    XRAM[57223] = 8'b0;
    XRAM[57224] = 8'b0;
    XRAM[57225] = 8'b0;
    XRAM[57226] = 8'b0;
    XRAM[57227] = 8'b0;
    XRAM[57228] = 8'b0;
    XRAM[57229] = 8'b0;
    XRAM[57230] = 8'b0;
    XRAM[57231] = 8'b0;
    XRAM[57232] = 8'b0;
    XRAM[57233] = 8'b0;
    XRAM[57234] = 8'b0;
    XRAM[57235] = 8'b0;
    XRAM[57236] = 8'b0;
    XRAM[57237] = 8'b0;
    XRAM[57238] = 8'b0;
    XRAM[57239] = 8'b0;
    XRAM[57240] = 8'b0;
    XRAM[57241] = 8'b0;
    XRAM[57242] = 8'b0;
    XRAM[57243] = 8'b0;
    XRAM[57244] = 8'b0;
    XRAM[57245] = 8'b0;
    XRAM[57246] = 8'b0;
    XRAM[57247] = 8'b0;
    XRAM[57248] = 8'b0;
    XRAM[57249] = 8'b0;
    XRAM[57250] = 8'b0;
    XRAM[57251] = 8'b0;
    XRAM[57252] = 8'b0;
    XRAM[57253] = 8'b0;
    XRAM[57254] = 8'b0;
    XRAM[57255] = 8'b0;
    XRAM[57256] = 8'b0;
    XRAM[57257] = 8'b0;
    XRAM[57258] = 8'b0;
    XRAM[57259] = 8'b0;
    XRAM[57260] = 8'b0;
    XRAM[57261] = 8'b0;
    XRAM[57262] = 8'b0;
    XRAM[57263] = 8'b0;
    XRAM[57264] = 8'b0;
    XRAM[57265] = 8'b0;
    XRAM[57266] = 8'b0;
    XRAM[57267] = 8'b0;
    XRAM[57268] = 8'b0;
    XRAM[57269] = 8'b0;
    XRAM[57270] = 8'b0;
    XRAM[57271] = 8'b0;
    XRAM[57272] = 8'b0;
    XRAM[57273] = 8'b0;
    XRAM[57274] = 8'b0;
    XRAM[57275] = 8'b0;
    XRAM[57276] = 8'b0;
    XRAM[57277] = 8'b0;
    XRAM[57278] = 8'b0;
    XRAM[57279] = 8'b0;
    XRAM[57280] = 8'b0;
    XRAM[57281] = 8'b0;
    XRAM[57282] = 8'b0;
    XRAM[57283] = 8'b0;
    XRAM[57284] = 8'b0;
    XRAM[57285] = 8'b0;
    XRAM[57286] = 8'b0;
    XRAM[57287] = 8'b0;
    XRAM[57288] = 8'b0;
    XRAM[57289] = 8'b0;
    XRAM[57290] = 8'b0;
    XRAM[57291] = 8'b0;
    XRAM[57292] = 8'b0;
    XRAM[57293] = 8'b0;
    XRAM[57294] = 8'b0;
    XRAM[57295] = 8'b0;
    XRAM[57296] = 8'b0;
    XRAM[57297] = 8'b0;
    XRAM[57298] = 8'b0;
    XRAM[57299] = 8'b0;
    XRAM[57300] = 8'b0;
    XRAM[57301] = 8'b0;
    XRAM[57302] = 8'b0;
    XRAM[57303] = 8'b0;
    XRAM[57304] = 8'b0;
    XRAM[57305] = 8'b0;
    XRAM[57306] = 8'b0;
    XRAM[57307] = 8'b0;
    XRAM[57308] = 8'b0;
    XRAM[57309] = 8'b0;
    XRAM[57310] = 8'b0;
    XRAM[57311] = 8'b0;
    XRAM[57312] = 8'b0;
    XRAM[57313] = 8'b0;
    XRAM[57314] = 8'b0;
    XRAM[57315] = 8'b0;
    XRAM[57316] = 8'b0;
    XRAM[57317] = 8'b0;
    XRAM[57318] = 8'b0;
    XRAM[57319] = 8'b0;
    XRAM[57320] = 8'b0;
    XRAM[57321] = 8'b0;
    XRAM[57322] = 8'b0;
    XRAM[57323] = 8'b0;
    XRAM[57324] = 8'b0;
    XRAM[57325] = 8'b0;
    XRAM[57326] = 8'b0;
    XRAM[57327] = 8'b0;
    XRAM[57328] = 8'b0;
    XRAM[57329] = 8'b0;
    XRAM[57330] = 8'b0;
    XRAM[57331] = 8'b0;
    XRAM[57332] = 8'b0;
    XRAM[57333] = 8'b0;
    XRAM[57334] = 8'b0;
    XRAM[57335] = 8'b0;
    XRAM[57336] = 8'b0;
    XRAM[57337] = 8'b0;
    XRAM[57338] = 8'b0;
    XRAM[57339] = 8'b0;
    XRAM[57340] = 8'b0;
    XRAM[57341] = 8'b0;
    XRAM[57342] = 8'b0;
    XRAM[57343] = 8'b0;
    XRAM[57344] = 8'b0;
    XRAM[57345] = 8'b0;
    XRAM[57346] = 8'b0;
    XRAM[57347] = 8'b0;
    XRAM[57348] = 8'b0;
    XRAM[57349] = 8'b0;
    XRAM[57350] = 8'b0;
    XRAM[57351] = 8'b0;
    XRAM[57352] = 8'b0;
    XRAM[57353] = 8'b0;
    XRAM[57354] = 8'b0;
    XRAM[57355] = 8'b0;
    XRAM[57356] = 8'b0;
    XRAM[57357] = 8'b0;
    XRAM[57358] = 8'b0;
    XRAM[57359] = 8'b0;
    XRAM[57360] = 8'b0;
    XRAM[57361] = 8'b0;
    XRAM[57362] = 8'b0;
    XRAM[57363] = 8'b0;
    XRAM[57364] = 8'b0;
    XRAM[57365] = 8'b0;
    XRAM[57366] = 8'b0;
    XRAM[57367] = 8'b0;
    XRAM[57368] = 8'b0;
    XRAM[57369] = 8'b0;
    XRAM[57370] = 8'b0;
    XRAM[57371] = 8'b0;
    XRAM[57372] = 8'b0;
    XRAM[57373] = 8'b0;
    XRAM[57374] = 8'b0;
    XRAM[57375] = 8'b0;
    XRAM[57376] = 8'b0;
    XRAM[57377] = 8'b0;
    XRAM[57378] = 8'b0;
    XRAM[57379] = 8'b0;
    XRAM[57380] = 8'b0;
    XRAM[57381] = 8'b0;
    XRAM[57382] = 8'b0;
    XRAM[57383] = 8'b0;
    XRAM[57384] = 8'b0;
    XRAM[57385] = 8'b0;
    XRAM[57386] = 8'b0;
    XRAM[57387] = 8'b0;
    XRAM[57388] = 8'b0;
    XRAM[57389] = 8'b0;
    XRAM[57390] = 8'b0;
    XRAM[57391] = 8'b0;
    XRAM[57392] = 8'b0;
    XRAM[57393] = 8'b0;
    XRAM[57394] = 8'b0;
    XRAM[57395] = 8'b0;
    XRAM[57396] = 8'b0;
    XRAM[57397] = 8'b0;
    XRAM[57398] = 8'b0;
    XRAM[57399] = 8'b0;
    XRAM[57400] = 8'b0;
    XRAM[57401] = 8'b0;
    XRAM[57402] = 8'b0;
    XRAM[57403] = 8'b0;
    XRAM[57404] = 8'b0;
    XRAM[57405] = 8'b0;
    XRAM[57406] = 8'b0;
    XRAM[57407] = 8'b0;
    XRAM[57408] = 8'b0;
    XRAM[57409] = 8'b0;
    XRAM[57410] = 8'b0;
    XRAM[57411] = 8'b0;
    XRAM[57412] = 8'b0;
    XRAM[57413] = 8'b0;
    XRAM[57414] = 8'b0;
    XRAM[57415] = 8'b0;
    XRAM[57416] = 8'b0;
    XRAM[57417] = 8'b0;
    XRAM[57418] = 8'b0;
    XRAM[57419] = 8'b0;
    XRAM[57420] = 8'b0;
    XRAM[57421] = 8'b0;
    XRAM[57422] = 8'b0;
    XRAM[57423] = 8'b0;
    XRAM[57424] = 8'b0;
    XRAM[57425] = 8'b0;
    XRAM[57426] = 8'b0;
    XRAM[57427] = 8'b0;
    XRAM[57428] = 8'b0;
    XRAM[57429] = 8'b0;
    XRAM[57430] = 8'b0;
    XRAM[57431] = 8'b0;
    XRAM[57432] = 8'b0;
    XRAM[57433] = 8'b0;
    XRAM[57434] = 8'b0;
    XRAM[57435] = 8'b0;
    XRAM[57436] = 8'b0;
    XRAM[57437] = 8'b0;
    XRAM[57438] = 8'b0;
    XRAM[57439] = 8'b0;
    XRAM[57440] = 8'b0;
    XRAM[57441] = 8'b0;
    XRAM[57442] = 8'b0;
    XRAM[57443] = 8'b0;
    XRAM[57444] = 8'b0;
    XRAM[57445] = 8'b0;
    XRAM[57446] = 8'b0;
    XRAM[57447] = 8'b0;
    XRAM[57448] = 8'b0;
    XRAM[57449] = 8'b0;
    XRAM[57450] = 8'b0;
    XRAM[57451] = 8'b0;
    XRAM[57452] = 8'b0;
    XRAM[57453] = 8'b0;
    XRAM[57454] = 8'b0;
    XRAM[57455] = 8'b0;
    XRAM[57456] = 8'b0;
    XRAM[57457] = 8'b0;
    XRAM[57458] = 8'b0;
    XRAM[57459] = 8'b0;
    XRAM[57460] = 8'b0;
    XRAM[57461] = 8'b0;
    XRAM[57462] = 8'b0;
    XRAM[57463] = 8'b0;
    XRAM[57464] = 8'b0;
    XRAM[57465] = 8'b0;
    XRAM[57466] = 8'b0;
    XRAM[57467] = 8'b0;
    XRAM[57468] = 8'b0;
    XRAM[57469] = 8'b0;
    XRAM[57470] = 8'b0;
    XRAM[57471] = 8'b0;
    XRAM[57472] = 8'b0;
    XRAM[57473] = 8'b0;
    XRAM[57474] = 8'b0;
    XRAM[57475] = 8'b0;
    XRAM[57476] = 8'b0;
    XRAM[57477] = 8'b0;
    XRAM[57478] = 8'b0;
    XRAM[57479] = 8'b0;
    XRAM[57480] = 8'b0;
    XRAM[57481] = 8'b0;
    XRAM[57482] = 8'b0;
    XRAM[57483] = 8'b0;
    XRAM[57484] = 8'b0;
    XRAM[57485] = 8'b0;
    XRAM[57486] = 8'b0;
    XRAM[57487] = 8'b0;
    XRAM[57488] = 8'b0;
    XRAM[57489] = 8'b0;
    XRAM[57490] = 8'b0;
    XRAM[57491] = 8'b0;
    XRAM[57492] = 8'b0;
    XRAM[57493] = 8'b0;
    XRAM[57494] = 8'b0;
    XRAM[57495] = 8'b0;
    XRAM[57496] = 8'b0;
    XRAM[57497] = 8'b0;
    XRAM[57498] = 8'b0;
    XRAM[57499] = 8'b0;
    XRAM[57500] = 8'b0;
    XRAM[57501] = 8'b0;
    XRAM[57502] = 8'b0;
    XRAM[57503] = 8'b0;
    XRAM[57504] = 8'b0;
    XRAM[57505] = 8'b0;
    XRAM[57506] = 8'b0;
    XRAM[57507] = 8'b0;
    XRAM[57508] = 8'b0;
    XRAM[57509] = 8'b0;
    XRAM[57510] = 8'b0;
    XRAM[57511] = 8'b0;
    XRAM[57512] = 8'b0;
    XRAM[57513] = 8'b0;
    XRAM[57514] = 8'b0;
    XRAM[57515] = 8'b0;
    XRAM[57516] = 8'b0;
    XRAM[57517] = 8'b0;
    XRAM[57518] = 8'b0;
    XRAM[57519] = 8'b0;
    XRAM[57520] = 8'b0;
    XRAM[57521] = 8'b0;
    XRAM[57522] = 8'b0;
    XRAM[57523] = 8'b0;
    XRAM[57524] = 8'b0;
    XRAM[57525] = 8'b0;
    XRAM[57526] = 8'b0;
    XRAM[57527] = 8'b0;
    XRAM[57528] = 8'b0;
    XRAM[57529] = 8'b0;
    XRAM[57530] = 8'b0;
    XRAM[57531] = 8'b0;
    XRAM[57532] = 8'b0;
    XRAM[57533] = 8'b0;
    XRAM[57534] = 8'b0;
    XRAM[57535] = 8'b0;
    XRAM[57536] = 8'b0;
    XRAM[57537] = 8'b0;
    XRAM[57538] = 8'b0;
    XRAM[57539] = 8'b0;
    XRAM[57540] = 8'b0;
    XRAM[57541] = 8'b0;
    XRAM[57542] = 8'b0;
    XRAM[57543] = 8'b0;
    XRAM[57544] = 8'b0;
    XRAM[57545] = 8'b0;
    XRAM[57546] = 8'b0;
    XRAM[57547] = 8'b0;
    XRAM[57548] = 8'b0;
    XRAM[57549] = 8'b0;
    XRAM[57550] = 8'b0;
    XRAM[57551] = 8'b0;
    XRAM[57552] = 8'b0;
    XRAM[57553] = 8'b0;
    XRAM[57554] = 8'b0;
    XRAM[57555] = 8'b0;
    XRAM[57556] = 8'b0;
    XRAM[57557] = 8'b0;
    XRAM[57558] = 8'b0;
    XRAM[57559] = 8'b0;
    XRAM[57560] = 8'b0;
    XRAM[57561] = 8'b0;
    XRAM[57562] = 8'b0;
    XRAM[57563] = 8'b0;
    XRAM[57564] = 8'b0;
    XRAM[57565] = 8'b0;
    XRAM[57566] = 8'b0;
    XRAM[57567] = 8'b0;
    XRAM[57568] = 8'b0;
    XRAM[57569] = 8'b0;
    XRAM[57570] = 8'b0;
    XRAM[57571] = 8'b0;
    XRAM[57572] = 8'b0;
    XRAM[57573] = 8'b0;
    XRAM[57574] = 8'b0;
    XRAM[57575] = 8'b0;
    XRAM[57576] = 8'b0;
    XRAM[57577] = 8'b0;
    XRAM[57578] = 8'b0;
    XRAM[57579] = 8'b0;
    XRAM[57580] = 8'b0;
    XRAM[57581] = 8'b0;
    XRAM[57582] = 8'b0;
    XRAM[57583] = 8'b0;
    XRAM[57584] = 8'b0;
    XRAM[57585] = 8'b0;
    XRAM[57586] = 8'b0;
    XRAM[57587] = 8'b0;
    XRAM[57588] = 8'b0;
    XRAM[57589] = 8'b0;
    XRAM[57590] = 8'b0;
    XRAM[57591] = 8'b0;
    XRAM[57592] = 8'b0;
    XRAM[57593] = 8'b0;
    XRAM[57594] = 8'b0;
    XRAM[57595] = 8'b0;
    XRAM[57596] = 8'b0;
    XRAM[57597] = 8'b0;
    XRAM[57598] = 8'b0;
    XRAM[57599] = 8'b0;
    XRAM[57600] = 8'b0;
    XRAM[57601] = 8'b0;
    XRAM[57602] = 8'b0;
    XRAM[57603] = 8'b0;
    XRAM[57604] = 8'b0;
    XRAM[57605] = 8'b0;
    XRAM[57606] = 8'b0;
    XRAM[57607] = 8'b0;
    XRAM[57608] = 8'b0;
    XRAM[57609] = 8'b0;
    XRAM[57610] = 8'b0;
    XRAM[57611] = 8'b0;
    XRAM[57612] = 8'b0;
    XRAM[57613] = 8'b0;
    XRAM[57614] = 8'b0;
    XRAM[57615] = 8'b0;
    XRAM[57616] = 8'b0;
    XRAM[57617] = 8'b0;
    XRAM[57618] = 8'b0;
    XRAM[57619] = 8'b0;
    XRAM[57620] = 8'b0;
    XRAM[57621] = 8'b0;
    XRAM[57622] = 8'b0;
    XRAM[57623] = 8'b0;
    XRAM[57624] = 8'b0;
    XRAM[57625] = 8'b0;
    XRAM[57626] = 8'b0;
    XRAM[57627] = 8'b0;
    XRAM[57628] = 8'b0;
    XRAM[57629] = 8'b0;
    XRAM[57630] = 8'b0;
    XRAM[57631] = 8'b0;
    XRAM[57632] = 8'b0;
    XRAM[57633] = 8'b0;
    XRAM[57634] = 8'b0;
    XRAM[57635] = 8'b0;
    XRAM[57636] = 8'b0;
    XRAM[57637] = 8'b0;
    XRAM[57638] = 8'b0;
    XRAM[57639] = 8'b0;
    XRAM[57640] = 8'b0;
    XRAM[57641] = 8'b0;
    XRAM[57642] = 8'b0;
    XRAM[57643] = 8'b0;
    XRAM[57644] = 8'b0;
    XRAM[57645] = 8'b0;
    XRAM[57646] = 8'b0;
    XRAM[57647] = 8'b0;
    XRAM[57648] = 8'b0;
    XRAM[57649] = 8'b0;
    XRAM[57650] = 8'b0;
    XRAM[57651] = 8'b0;
    XRAM[57652] = 8'b0;
    XRAM[57653] = 8'b0;
    XRAM[57654] = 8'b0;
    XRAM[57655] = 8'b0;
    XRAM[57656] = 8'b0;
    XRAM[57657] = 8'b0;
    XRAM[57658] = 8'b0;
    XRAM[57659] = 8'b0;
    XRAM[57660] = 8'b0;
    XRAM[57661] = 8'b0;
    XRAM[57662] = 8'b0;
    XRAM[57663] = 8'b0;
    XRAM[57664] = 8'b0;
    XRAM[57665] = 8'b0;
    XRAM[57666] = 8'b0;
    XRAM[57667] = 8'b0;
    XRAM[57668] = 8'b0;
    XRAM[57669] = 8'b0;
    XRAM[57670] = 8'b0;
    XRAM[57671] = 8'b0;
    XRAM[57672] = 8'b0;
    XRAM[57673] = 8'b0;
    XRAM[57674] = 8'b0;
    XRAM[57675] = 8'b0;
    XRAM[57676] = 8'b0;
    XRAM[57677] = 8'b0;
    XRAM[57678] = 8'b0;
    XRAM[57679] = 8'b0;
    XRAM[57680] = 8'b0;
    XRAM[57681] = 8'b0;
    XRAM[57682] = 8'b0;
    XRAM[57683] = 8'b0;
    XRAM[57684] = 8'b0;
    XRAM[57685] = 8'b0;
    XRAM[57686] = 8'b0;
    XRAM[57687] = 8'b0;
    XRAM[57688] = 8'b0;
    XRAM[57689] = 8'b0;
    XRAM[57690] = 8'b0;
    XRAM[57691] = 8'b0;
    XRAM[57692] = 8'b0;
    XRAM[57693] = 8'b0;
    XRAM[57694] = 8'b0;
    XRAM[57695] = 8'b0;
    XRAM[57696] = 8'b0;
    XRAM[57697] = 8'b0;
    XRAM[57698] = 8'b0;
    XRAM[57699] = 8'b0;
    XRAM[57700] = 8'b0;
    XRAM[57701] = 8'b0;
    XRAM[57702] = 8'b0;
    XRAM[57703] = 8'b0;
    XRAM[57704] = 8'b0;
    XRAM[57705] = 8'b0;
    XRAM[57706] = 8'b0;
    XRAM[57707] = 8'b0;
    XRAM[57708] = 8'b0;
    XRAM[57709] = 8'b0;
    XRAM[57710] = 8'b0;
    XRAM[57711] = 8'b0;
    XRAM[57712] = 8'b0;
    XRAM[57713] = 8'b0;
    XRAM[57714] = 8'b0;
    XRAM[57715] = 8'b0;
    XRAM[57716] = 8'b0;
    XRAM[57717] = 8'b0;
    XRAM[57718] = 8'b0;
    XRAM[57719] = 8'b0;
    XRAM[57720] = 8'b0;
    XRAM[57721] = 8'b0;
    XRAM[57722] = 8'b0;
    XRAM[57723] = 8'b0;
    XRAM[57724] = 8'b0;
    XRAM[57725] = 8'b0;
    XRAM[57726] = 8'b0;
    XRAM[57727] = 8'b0;
    XRAM[57728] = 8'b0;
    XRAM[57729] = 8'b0;
    XRAM[57730] = 8'b0;
    XRAM[57731] = 8'b0;
    XRAM[57732] = 8'b0;
    XRAM[57733] = 8'b0;
    XRAM[57734] = 8'b0;
    XRAM[57735] = 8'b0;
    XRAM[57736] = 8'b0;
    XRAM[57737] = 8'b0;
    XRAM[57738] = 8'b0;
    XRAM[57739] = 8'b0;
    XRAM[57740] = 8'b0;
    XRAM[57741] = 8'b0;
    XRAM[57742] = 8'b0;
    XRAM[57743] = 8'b0;
    XRAM[57744] = 8'b0;
    XRAM[57745] = 8'b0;
    XRAM[57746] = 8'b0;
    XRAM[57747] = 8'b0;
    XRAM[57748] = 8'b0;
    XRAM[57749] = 8'b0;
    XRAM[57750] = 8'b0;
    XRAM[57751] = 8'b0;
    XRAM[57752] = 8'b0;
    XRAM[57753] = 8'b0;
    XRAM[57754] = 8'b0;
    XRAM[57755] = 8'b0;
    XRAM[57756] = 8'b0;
    XRAM[57757] = 8'b0;
    XRAM[57758] = 8'b0;
    XRAM[57759] = 8'b0;
    XRAM[57760] = 8'b0;
    XRAM[57761] = 8'b0;
    XRAM[57762] = 8'b0;
    XRAM[57763] = 8'b0;
    XRAM[57764] = 8'b0;
    XRAM[57765] = 8'b0;
    XRAM[57766] = 8'b0;
    XRAM[57767] = 8'b0;
    XRAM[57768] = 8'b0;
    XRAM[57769] = 8'b0;
    XRAM[57770] = 8'b0;
    XRAM[57771] = 8'b0;
    XRAM[57772] = 8'b0;
    XRAM[57773] = 8'b0;
    XRAM[57774] = 8'b0;
    XRAM[57775] = 8'b0;
    XRAM[57776] = 8'b0;
    XRAM[57777] = 8'b0;
    XRAM[57778] = 8'b0;
    XRAM[57779] = 8'b0;
    XRAM[57780] = 8'b0;
    XRAM[57781] = 8'b0;
    XRAM[57782] = 8'b0;
    XRAM[57783] = 8'b0;
    XRAM[57784] = 8'b0;
    XRAM[57785] = 8'b0;
    XRAM[57786] = 8'b0;
    XRAM[57787] = 8'b0;
    XRAM[57788] = 8'b0;
    XRAM[57789] = 8'b0;
    XRAM[57790] = 8'b0;
    XRAM[57791] = 8'b0;
    XRAM[57792] = 8'b0;
    XRAM[57793] = 8'b0;
    XRAM[57794] = 8'b0;
    XRAM[57795] = 8'b0;
    XRAM[57796] = 8'b0;
    XRAM[57797] = 8'b0;
    XRAM[57798] = 8'b0;
    XRAM[57799] = 8'b0;
    XRAM[57800] = 8'b0;
    XRAM[57801] = 8'b0;
    XRAM[57802] = 8'b0;
    XRAM[57803] = 8'b0;
    XRAM[57804] = 8'b0;
    XRAM[57805] = 8'b0;
    XRAM[57806] = 8'b0;
    XRAM[57807] = 8'b0;
    XRAM[57808] = 8'b0;
    XRAM[57809] = 8'b0;
    XRAM[57810] = 8'b0;
    XRAM[57811] = 8'b0;
    XRAM[57812] = 8'b0;
    XRAM[57813] = 8'b0;
    XRAM[57814] = 8'b0;
    XRAM[57815] = 8'b0;
    XRAM[57816] = 8'b0;
    XRAM[57817] = 8'b0;
    XRAM[57818] = 8'b0;
    XRAM[57819] = 8'b0;
    XRAM[57820] = 8'b0;
    XRAM[57821] = 8'b0;
    XRAM[57822] = 8'b0;
    XRAM[57823] = 8'b0;
    XRAM[57824] = 8'b0;
    XRAM[57825] = 8'b0;
    XRAM[57826] = 8'b0;
    XRAM[57827] = 8'b0;
    XRAM[57828] = 8'b0;
    XRAM[57829] = 8'b0;
    XRAM[57830] = 8'b0;
    XRAM[57831] = 8'b0;
    XRAM[57832] = 8'b0;
    XRAM[57833] = 8'b0;
    XRAM[57834] = 8'b0;
    XRAM[57835] = 8'b0;
    XRAM[57836] = 8'b0;
    XRAM[57837] = 8'b0;
    XRAM[57838] = 8'b0;
    XRAM[57839] = 8'b0;
    XRAM[57840] = 8'b0;
    XRAM[57841] = 8'b0;
    XRAM[57842] = 8'b0;
    XRAM[57843] = 8'b0;
    XRAM[57844] = 8'b0;
    XRAM[57845] = 8'b0;
    XRAM[57846] = 8'b0;
    XRAM[57847] = 8'b0;
    XRAM[57848] = 8'b0;
    XRAM[57849] = 8'b0;
    XRAM[57850] = 8'b0;
    XRAM[57851] = 8'b0;
    XRAM[57852] = 8'b0;
    XRAM[57853] = 8'b0;
    XRAM[57854] = 8'b0;
    XRAM[57855] = 8'b0;
    XRAM[57856] = 8'b0;
    XRAM[57857] = 8'b0;
    XRAM[57858] = 8'b0;
    XRAM[57859] = 8'b0;
    XRAM[57860] = 8'b0;
    XRAM[57861] = 8'b0;
    XRAM[57862] = 8'b0;
    XRAM[57863] = 8'b0;
    XRAM[57864] = 8'b0;
    XRAM[57865] = 8'b0;
    XRAM[57866] = 8'b0;
    XRAM[57867] = 8'b0;
    XRAM[57868] = 8'b0;
    XRAM[57869] = 8'b0;
    XRAM[57870] = 8'b0;
    XRAM[57871] = 8'b0;
    XRAM[57872] = 8'b0;
    XRAM[57873] = 8'b0;
    XRAM[57874] = 8'b0;
    XRAM[57875] = 8'b0;
    XRAM[57876] = 8'b0;
    XRAM[57877] = 8'b0;
    XRAM[57878] = 8'b0;
    XRAM[57879] = 8'b0;
    XRAM[57880] = 8'b0;
    XRAM[57881] = 8'b0;
    XRAM[57882] = 8'b0;
    XRAM[57883] = 8'b0;
    XRAM[57884] = 8'b0;
    XRAM[57885] = 8'b0;
    XRAM[57886] = 8'b0;
    XRAM[57887] = 8'b0;
    XRAM[57888] = 8'b0;
    XRAM[57889] = 8'b0;
    XRAM[57890] = 8'b0;
    XRAM[57891] = 8'b0;
    XRAM[57892] = 8'b0;
    XRAM[57893] = 8'b0;
    XRAM[57894] = 8'b0;
    XRAM[57895] = 8'b0;
    XRAM[57896] = 8'b0;
    XRAM[57897] = 8'b0;
    XRAM[57898] = 8'b0;
    XRAM[57899] = 8'b0;
    XRAM[57900] = 8'b0;
    XRAM[57901] = 8'b0;
    XRAM[57902] = 8'b0;
    XRAM[57903] = 8'b0;
    XRAM[57904] = 8'b0;
    XRAM[57905] = 8'b0;
    XRAM[57906] = 8'b0;
    XRAM[57907] = 8'b0;
    XRAM[57908] = 8'b0;
    XRAM[57909] = 8'b0;
    XRAM[57910] = 8'b0;
    XRAM[57911] = 8'b0;
    XRAM[57912] = 8'b0;
    XRAM[57913] = 8'b0;
    XRAM[57914] = 8'b0;
    XRAM[57915] = 8'b0;
    XRAM[57916] = 8'b0;
    XRAM[57917] = 8'b0;
    XRAM[57918] = 8'b0;
    XRAM[57919] = 8'b0;
    XRAM[57920] = 8'b0;
    XRAM[57921] = 8'b0;
    XRAM[57922] = 8'b0;
    XRAM[57923] = 8'b0;
    XRAM[57924] = 8'b0;
    XRAM[57925] = 8'b0;
    XRAM[57926] = 8'b0;
    XRAM[57927] = 8'b0;
    XRAM[57928] = 8'b0;
    XRAM[57929] = 8'b0;
    XRAM[57930] = 8'b0;
    XRAM[57931] = 8'b0;
    XRAM[57932] = 8'b0;
    XRAM[57933] = 8'b0;
    XRAM[57934] = 8'b0;
    XRAM[57935] = 8'b0;
    XRAM[57936] = 8'b0;
    XRAM[57937] = 8'b0;
    XRAM[57938] = 8'b0;
    XRAM[57939] = 8'b0;
    XRAM[57940] = 8'b0;
    XRAM[57941] = 8'b0;
    XRAM[57942] = 8'b0;
    XRAM[57943] = 8'b0;
    XRAM[57944] = 8'b0;
    XRAM[57945] = 8'b0;
    XRAM[57946] = 8'b0;
    XRAM[57947] = 8'b0;
    XRAM[57948] = 8'b0;
    XRAM[57949] = 8'b0;
    XRAM[57950] = 8'b0;
    XRAM[57951] = 8'b0;
    XRAM[57952] = 8'b0;
    XRAM[57953] = 8'b0;
    XRAM[57954] = 8'b0;
    XRAM[57955] = 8'b0;
    XRAM[57956] = 8'b0;
    XRAM[57957] = 8'b0;
    XRAM[57958] = 8'b0;
    XRAM[57959] = 8'b0;
    XRAM[57960] = 8'b0;
    XRAM[57961] = 8'b0;
    XRAM[57962] = 8'b0;
    XRAM[57963] = 8'b0;
    XRAM[57964] = 8'b0;
    XRAM[57965] = 8'b0;
    XRAM[57966] = 8'b0;
    XRAM[57967] = 8'b0;
    XRAM[57968] = 8'b0;
    XRAM[57969] = 8'b0;
    XRAM[57970] = 8'b0;
    XRAM[57971] = 8'b0;
    XRAM[57972] = 8'b0;
    XRAM[57973] = 8'b0;
    XRAM[57974] = 8'b0;
    XRAM[57975] = 8'b0;
    XRAM[57976] = 8'b0;
    XRAM[57977] = 8'b0;
    XRAM[57978] = 8'b0;
    XRAM[57979] = 8'b0;
    XRAM[57980] = 8'b0;
    XRAM[57981] = 8'b0;
    XRAM[57982] = 8'b0;
    XRAM[57983] = 8'b0;
    XRAM[57984] = 8'b0;
    XRAM[57985] = 8'b0;
    XRAM[57986] = 8'b0;
    XRAM[57987] = 8'b0;
    XRAM[57988] = 8'b0;
    XRAM[57989] = 8'b0;
    XRAM[57990] = 8'b0;
    XRAM[57991] = 8'b0;
    XRAM[57992] = 8'b0;
    XRAM[57993] = 8'b0;
    XRAM[57994] = 8'b0;
    XRAM[57995] = 8'b0;
    XRAM[57996] = 8'b0;
    XRAM[57997] = 8'b0;
    XRAM[57998] = 8'b0;
    XRAM[57999] = 8'b0;
    XRAM[58000] = 8'b0;
    XRAM[58001] = 8'b0;
    XRAM[58002] = 8'b0;
    XRAM[58003] = 8'b0;
    XRAM[58004] = 8'b0;
    XRAM[58005] = 8'b0;
    XRAM[58006] = 8'b0;
    XRAM[58007] = 8'b0;
    XRAM[58008] = 8'b0;
    XRAM[58009] = 8'b0;
    XRAM[58010] = 8'b0;
    XRAM[58011] = 8'b0;
    XRAM[58012] = 8'b0;
    XRAM[58013] = 8'b0;
    XRAM[58014] = 8'b0;
    XRAM[58015] = 8'b0;
    XRAM[58016] = 8'b0;
    XRAM[58017] = 8'b0;
    XRAM[58018] = 8'b0;
    XRAM[58019] = 8'b0;
    XRAM[58020] = 8'b0;
    XRAM[58021] = 8'b0;
    XRAM[58022] = 8'b0;
    XRAM[58023] = 8'b0;
    XRAM[58024] = 8'b0;
    XRAM[58025] = 8'b0;
    XRAM[58026] = 8'b0;
    XRAM[58027] = 8'b0;
    XRAM[58028] = 8'b0;
    XRAM[58029] = 8'b0;
    XRAM[58030] = 8'b0;
    XRAM[58031] = 8'b0;
    XRAM[58032] = 8'b0;
    XRAM[58033] = 8'b0;
    XRAM[58034] = 8'b0;
    XRAM[58035] = 8'b0;
    XRAM[58036] = 8'b0;
    XRAM[58037] = 8'b0;
    XRAM[58038] = 8'b0;
    XRAM[58039] = 8'b0;
    XRAM[58040] = 8'b0;
    XRAM[58041] = 8'b0;
    XRAM[58042] = 8'b0;
    XRAM[58043] = 8'b0;
    XRAM[58044] = 8'b0;
    XRAM[58045] = 8'b0;
    XRAM[58046] = 8'b0;
    XRAM[58047] = 8'b0;
    XRAM[58048] = 8'b0;
    XRAM[58049] = 8'b0;
    XRAM[58050] = 8'b0;
    XRAM[58051] = 8'b0;
    XRAM[58052] = 8'b0;
    XRAM[58053] = 8'b0;
    XRAM[58054] = 8'b0;
    XRAM[58055] = 8'b0;
    XRAM[58056] = 8'b0;
    XRAM[58057] = 8'b0;
    XRAM[58058] = 8'b0;
    XRAM[58059] = 8'b0;
    XRAM[58060] = 8'b0;
    XRAM[58061] = 8'b0;
    XRAM[58062] = 8'b0;
    XRAM[58063] = 8'b0;
    XRAM[58064] = 8'b0;
    XRAM[58065] = 8'b0;
    XRAM[58066] = 8'b0;
    XRAM[58067] = 8'b0;
    XRAM[58068] = 8'b0;
    XRAM[58069] = 8'b0;
    XRAM[58070] = 8'b0;
    XRAM[58071] = 8'b0;
    XRAM[58072] = 8'b0;
    XRAM[58073] = 8'b0;
    XRAM[58074] = 8'b0;
    XRAM[58075] = 8'b0;
    XRAM[58076] = 8'b0;
    XRAM[58077] = 8'b0;
    XRAM[58078] = 8'b0;
    XRAM[58079] = 8'b0;
    XRAM[58080] = 8'b0;
    XRAM[58081] = 8'b0;
    XRAM[58082] = 8'b0;
    XRAM[58083] = 8'b0;
    XRAM[58084] = 8'b0;
    XRAM[58085] = 8'b0;
    XRAM[58086] = 8'b0;
    XRAM[58087] = 8'b0;
    XRAM[58088] = 8'b0;
    XRAM[58089] = 8'b0;
    XRAM[58090] = 8'b0;
    XRAM[58091] = 8'b0;
    XRAM[58092] = 8'b0;
    XRAM[58093] = 8'b0;
    XRAM[58094] = 8'b0;
    XRAM[58095] = 8'b0;
    XRAM[58096] = 8'b0;
    XRAM[58097] = 8'b0;
    XRAM[58098] = 8'b0;
    XRAM[58099] = 8'b0;
    XRAM[58100] = 8'b0;
    XRAM[58101] = 8'b0;
    XRAM[58102] = 8'b0;
    XRAM[58103] = 8'b0;
    XRAM[58104] = 8'b0;
    XRAM[58105] = 8'b0;
    XRAM[58106] = 8'b0;
    XRAM[58107] = 8'b0;
    XRAM[58108] = 8'b0;
    XRAM[58109] = 8'b0;
    XRAM[58110] = 8'b0;
    XRAM[58111] = 8'b0;
    XRAM[58112] = 8'b0;
    XRAM[58113] = 8'b0;
    XRAM[58114] = 8'b0;
    XRAM[58115] = 8'b0;
    XRAM[58116] = 8'b0;
    XRAM[58117] = 8'b0;
    XRAM[58118] = 8'b0;
    XRAM[58119] = 8'b0;
    XRAM[58120] = 8'b0;
    XRAM[58121] = 8'b0;
    XRAM[58122] = 8'b0;
    XRAM[58123] = 8'b0;
    XRAM[58124] = 8'b0;
    XRAM[58125] = 8'b0;
    XRAM[58126] = 8'b0;
    XRAM[58127] = 8'b0;
    XRAM[58128] = 8'b0;
    XRAM[58129] = 8'b0;
    XRAM[58130] = 8'b0;
    XRAM[58131] = 8'b0;
    XRAM[58132] = 8'b0;
    XRAM[58133] = 8'b0;
    XRAM[58134] = 8'b0;
    XRAM[58135] = 8'b0;
    XRAM[58136] = 8'b0;
    XRAM[58137] = 8'b0;
    XRAM[58138] = 8'b0;
    XRAM[58139] = 8'b0;
    XRAM[58140] = 8'b0;
    XRAM[58141] = 8'b0;
    XRAM[58142] = 8'b0;
    XRAM[58143] = 8'b0;
    XRAM[58144] = 8'b0;
    XRAM[58145] = 8'b0;
    XRAM[58146] = 8'b0;
    XRAM[58147] = 8'b0;
    XRAM[58148] = 8'b0;
    XRAM[58149] = 8'b0;
    XRAM[58150] = 8'b0;
    XRAM[58151] = 8'b0;
    XRAM[58152] = 8'b0;
    XRAM[58153] = 8'b0;
    XRAM[58154] = 8'b0;
    XRAM[58155] = 8'b0;
    XRAM[58156] = 8'b0;
    XRAM[58157] = 8'b0;
    XRAM[58158] = 8'b0;
    XRAM[58159] = 8'b0;
    XRAM[58160] = 8'b0;
    XRAM[58161] = 8'b0;
    XRAM[58162] = 8'b0;
    XRAM[58163] = 8'b0;
    XRAM[58164] = 8'b0;
    XRAM[58165] = 8'b0;
    XRAM[58166] = 8'b0;
    XRAM[58167] = 8'b0;
    XRAM[58168] = 8'b0;
    XRAM[58169] = 8'b0;
    XRAM[58170] = 8'b0;
    XRAM[58171] = 8'b0;
    XRAM[58172] = 8'b0;
    XRAM[58173] = 8'b0;
    XRAM[58174] = 8'b0;
    XRAM[58175] = 8'b0;
    XRAM[58176] = 8'b0;
    XRAM[58177] = 8'b0;
    XRAM[58178] = 8'b0;
    XRAM[58179] = 8'b0;
    XRAM[58180] = 8'b0;
    XRAM[58181] = 8'b0;
    XRAM[58182] = 8'b0;
    XRAM[58183] = 8'b0;
    XRAM[58184] = 8'b0;
    XRAM[58185] = 8'b0;
    XRAM[58186] = 8'b0;
    XRAM[58187] = 8'b0;
    XRAM[58188] = 8'b0;
    XRAM[58189] = 8'b0;
    XRAM[58190] = 8'b0;
    XRAM[58191] = 8'b0;
    XRAM[58192] = 8'b0;
    XRAM[58193] = 8'b0;
    XRAM[58194] = 8'b0;
    XRAM[58195] = 8'b0;
    XRAM[58196] = 8'b0;
    XRAM[58197] = 8'b0;
    XRAM[58198] = 8'b0;
    XRAM[58199] = 8'b0;
    XRAM[58200] = 8'b0;
    XRAM[58201] = 8'b0;
    XRAM[58202] = 8'b0;
    XRAM[58203] = 8'b0;
    XRAM[58204] = 8'b0;
    XRAM[58205] = 8'b0;
    XRAM[58206] = 8'b0;
    XRAM[58207] = 8'b0;
    XRAM[58208] = 8'b0;
    XRAM[58209] = 8'b0;
    XRAM[58210] = 8'b0;
    XRAM[58211] = 8'b0;
    XRAM[58212] = 8'b0;
    XRAM[58213] = 8'b0;
    XRAM[58214] = 8'b0;
    XRAM[58215] = 8'b0;
    XRAM[58216] = 8'b0;
    XRAM[58217] = 8'b0;
    XRAM[58218] = 8'b0;
    XRAM[58219] = 8'b0;
    XRAM[58220] = 8'b0;
    XRAM[58221] = 8'b0;
    XRAM[58222] = 8'b0;
    XRAM[58223] = 8'b0;
    XRAM[58224] = 8'b0;
    XRAM[58225] = 8'b0;
    XRAM[58226] = 8'b0;
    XRAM[58227] = 8'b0;
    XRAM[58228] = 8'b0;
    XRAM[58229] = 8'b0;
    XRAM[58230] = 8'b0;
    XRAM[58231] = 8'b0;
    XRAM[58232] = 8'b0;
    XRAM[58233] = 8'b0;
    XRAM[58234] = 8'b0;
    XRAM[58235] = 8'b0;
    XRAM[58236] = 8'b0;
    XRAM[58237] = 8'b0;
    XRAM[58238] = 8'b0;
    XRAM[58239] = 8'b0;
    XRAM[58240] = 8'b0;
    XRAM[58241] = 8'b0;
    XRAM[58242] = 8'b0;
    XRAM[58243] = 8'b0;
    XRAM[58244] = 8'b0;
    XRAM[58245] = 8'b0;
    XRAM[58246] = 8'b0;
    XRAM[58247] = 8'b0;
    XRAM[58248] = 8'b0;
    XRAM[58249] = 8'b0;
    XRAM[58250] = 8'b0;
    XRAM[58251] = 8'b0;
    XRAM[58252] = 8'b0;
    XRAM[58253] = 8'b0;
    XRAM[58254] = 8'b0;
    XRAM[58255] = 8'b0;
    XRAM[58256] = 8'b0;
    XRAM[58257] = 8'b0;
    XRAM[58258] = 8'b0;
    XRAM[58259] = 8'b0;
    XRAM[58260] = 8'b0;
    XRAM[58261] = 8'b0;
    XRAM[58262] = 8'b0;
    XRAM[58263] = 8'b0;
    XRAM[58264] = 8'b0;
    XRAM[58265] = 8'b0;
    XRAM[58266] = 8'b0;
    XRAM[58267] = 8'b0;
    XRAM[58268] = 8'b0;
    XRAM[58269] = 8'b0;
    XRAM[58270] = 8'b0;
    XRAM[58271] = 8'b0;
    XRAM[58272] = 8'b0;
    XRAM[58273] = 8'b0;
    XRAM[58274] = 8'b0;
    XRAM[58275] = 8'b0;
    XRAM[58276] = 8'b0;
    XRAM[58277] = 8'b0;
    XRAM[58278] = 8'b0;
    XRAM[58279] = 8'b0;
    XRAM[58280] = 8'b0;
    XRAM[58281] = 8'b0;
    XRAM[58282] = 8'b0;
    XRAM[58283] = 8'b0;
    XRAM[58284] = 8'b0;
    XRAM[58285] = 8'b0;
    XRAM[58286] = 8'b0;
    XRAM[58287] = 8'b0;
    XRAM[58288] = 8'b0;
    XRAM[58289] = 8'b0;
    XRAM[58290] = 8'b0;
    XRAM[58291] = 8'b0;
    XRAM[58292] = 8'b0;
    XRAM[58293] = 8'b0;
    XRAM[58294] = 8'b0;
    XRAM[58295] = 8'b0;
    XRAM[58296] = 8'b0;
    XRAM[58297] = 8'b0;
    XRAM[58298] = 8'b0;
    XRAM[58299] = 8'b0;
    XRAM[58300] = 8'b0;
    XRAM[58301] = 8'b0;
    XRAM[58302] = 8'b0;
    XRAM[58303] = 8'b0;
    XRAM[58304] = 8'b0;
    XRAM[58305] = 8'b0;
    XRAM[58306] = 8'b0;
    XRAM[58307] = 8'b0;
    XRAM[58308] = 8'b0;
    XRAM[58309] = 8'b0;
    XRAM[58310] = 8'b0;
    XRAM[58311] = 8'b0;
    XRAM[58312] = 8'b0;
    XRAM[58313] = 8'b0;
    XRAM[58314] = 8'b0;
    XRAM[58315] = 8'b0;
    XRAM[58316] = 8'b0;
    XRAM[58317] = 8'b0;
    XRAM[58318] = 8'b0;
    XRAM[58319] = 8'b0;
    XRAM[58320] = 8'b0;
    XRAM[58321] = 8'b0;
    XRAM[58322] = 8'b0;
    XRAM[58323] = 8'b0;
    XRAM[58324] = 8'b0;
    XRAM[58325] = 8'b0;
    XRAM[58326] = 8'b0;
    XRAM[58327] = 8'b0;
    XRAM[58328] = 8'b0;
    XRAM[58329] = 8'b0;
    XRAM[58330] = 8'b0;
    XRAM[58331] = 8'b0;
    XRAM[58332] = 8'b0;
    XRAM[58333] = 8'b0;
    XRAM[58334] = 8'b0;
    XRAM[58335] = 8'b0;
    XRAM[58336] = 8'b0;
    XRAM[58337] = 8'b0;
    XRAM[58338] = 8'b0;
    XRAM[58339] = 8'b0;
    XRAM[58340] = 8'b0;
    XRAM[58341] = 8'b0;
    XRAM[58342] = 8'b0;
    XRAM[58343] = 8'b0;
    XRAM[58344] = 8'b0;
    XRAM[58345] = 8'b0;
    XRAM[58346] = 8'b0;
    XRAM[58347] = 8'b0;
    XRAM[58348] = 8'b0;
    XRAM[58349] = 8'b0;
    XRAM[58350] = 8'b0;
    XRAM[58351] = 8'b0;
    XRAM[58352] = 8'b0;
    XRAM[58353] = 8'b0;
    XRAM[58354] = 8'b0;
    XRAM[58355] = 8'b0;
    XRAM[58356] = 8'b0;
    XRAM[58357] = 8'b0;
    XRAM[58358] = 8'b0;
    XRAM[58359] = 8'b0;
    XRAM[58360] = 8'b0;
    XRAM[58361] = 8'b0;
    XRAM[58362] = 8'b0;
    XRAM[58363] = 8'b0;
    XRAM[58364] = 8'b0;
    XRAM[58365] = 8'b0;
    XRAM[58366] = 8'b0;
    XRAM[58367] = 8'b0;
    XRAM[58368] = 8'b0;
    XRAM[58369] = 8'b0;
    XRAM[58370] = 8'b0;
    XRAM[58371] = 8'b0;
    XRAM[58372] = 8'b0;
    XRAM[58373] = 8'b0;
    XRAM[58374] = 8'b0;
    XRAM[58375] = 8'b0;
    XRAM[58376] = 8'b0;
    XRAM[58377] = 8'b0;
    XRAM[58378] = 8'b0;
    XRAM[58379] = 8'b0;
    XRAM[58380] = 8'b0;
    XRAM[58381] = 8'b0;
    XRAM[58382] = 8'b0;
    XRAM[58383] = 8'b0;
    XRAM[58384] = 8'b0;
    XRAM[58385] = 8'b0;
    XRAM[58386] = 8'b0;
    XRAM[58387] = 8'b0;
    XRAM[58388] = 8'b0;
    XRAM[58389] = 8'b0;
    XRAM[58390] = 8'b0;
    XRAM[58391] = 8'b0;
    XRAM[58392] = 8'b0;
    XRAM[58393] = 8'b0;
    XRAM[58394] = 8'b0;
    XRAM[58395] = 8'b0;
    XRAM[58396] = 8'b0;
    XRAM[58397] = 8'b0;
    XRAM[58398] = 8'b0;
    XRAM[58399] = 8'b0;
    XRAM[58400] = 8'b0;
    XRAM[58401] = 8'b0;
    XRAM[58402] = 8'b0;
    XRAM[58403] = 8'b0;
    XRAM[58404] = 8'b0;
    XRAM[58405] = 8'b0;
    XRAM[58406] = 8'b0;
    XRAM[58407] = 8'b0;
    XRAM[58408] = 8'b0;
    XRAM[58409] = 8'b0;
    XRAM[58410] = 8'b0;
    XRAM[58411] = 8'b0;
    XRAM[58412] = 8'b0;
    XRAM[58413] = 8'b0;
    XRAM[58414] = 8'b0;
    XRAM[58415] = 8'b0;
    XRAM[58416] = 8'b0;
    XRAM[58417] = 8'b0;
    XRAM[58418] = 8'b0;
    XRAM[58419] = 8'b0;
    XRAM[58420] = 8'b0;
    XRAM[58421] = 8'b0;
    XRAM[58422] = 8'b0;
    XRAM[58423] = 8'b0;
    XRAM[58424] = 8'b0;
    XRAM[58425] = 8'b0;
    XRAM[58426] = 8'b0;
    XRAM[58427] = 8'b0;
    XRAM[58428] = 8'b0;
    XRAM[58429] = 8'b0;
    XRAM[58430] = 8'b0;
    XRAM[58431] = 8'b0;
    XRAM[58432] = 8'b0;
    XRAM[58433] = 8'b0;
    XRAM[58434] = 8'b0;
    XRAM[58435] = 8'b0;
    XRAM[58436] = 8'b0;
    XRAM[58437] = 8'b0;
    XRAM[58438] = 8'b0;
    XRAM[58439] = 8'b0;
    XRAM[58440] = 8'b0;
    XRAM[58441] = 8'b0;
    XRAM[58442] = 8'b0;
    XRAM[58443] = 8'b0;
    XRAM[58444] = 8'b0;
    XRAM[58445] = 8'b0;
    XRAM[58446] = 8'b0;
    XRAM[58447] = 8'b0;
    XRAM[58448] = 8'b0;
    XRAM[58449] = 8'b0;
    XRAM[58450] = 8'b0;
    XRAM[58451] = 8'b0;
    XRAM[58452] = 8'b0;
    XRAM[58453] = 8'b0;
    XRAM[58454] = 8'b0;
    XRAM[58455] = 8'b0;
    XRAM[58456] = 8'b0;
    XRAM[58457] = 8'b0;
    XRAM[58458] = 8'b0;
    XRAM[58459] = 8'b0;
    XRAM[58460] = 8'b0;
    XRAM[58461] = 8'b0;
    XRAM[58462] = 8'b0;
    XRAM[58463] = 8'b0;
    XRAM[58464] = 8'b0;
    XRAM[58465] = 8'b0;
    XRAM[58466] = 8'b0;
    XRAM[58467] = 8'b0;
    XRAM[58468] = 8'b0;
    XRAM[58469] = 8'b0;
    XRAM[58470] = 8'b0;
    XRAM[58471] = 8'b0;
    XRAM[58472] = 8'b0;
    XRAM[58473] = 8'b0;
    XRAM[58474] = 8'b0;
    XRAM[58475] = 8'b0;
    XRAM[58476] = 8'b0;
    XRAM[58477] = 8'b0;
    XRAM[58478] = 8'b0;
    XRAM[58479] = 8'b0;
    XRAM[58480] = 8'b0;
    XRAM[58481] = 8'b0;
    XRAM[58482] = 8'b0;
    XRAM[58483] = 8'b0;
    XRAM[58484] = 8'b0;
    XRAM[58485] = 8'b0;
    XRAM[58486] = 8'b0;
    XRAM[58487] = 8'b0;
    XRAM[58488] = 8'b0;
    XRAM[58489] = 8'b0;
    XRAM[58490] = 8'b0;
    XRAM[58491] = 8'b0;
    XRAM[58492] = 8'b0;
    XRAM[58493] = 8'b0;
    XRAM[58494] = 8'b0;
    XRAM[58495] = 8'b0;
    XRAM[58496] = 8'b0;
    XRAM[58497] = 8'b0;
    XRAM[58498] = 8'b0;
    XRAM[58499] = 8'b0;
    XRAM[58500] = 8'b0;
    XRAM[58501] = 8'b0;
    XRAM[58502] = 8'b0;
    XRAM[58503] = 8'b0;
    XRAM[58504] = 8'b0;
    XRAM[58505] = 8'b0;
    XRAM[58506] = 8'b0;
    XRAM[58507] = 8'b0;
    XRAM[58508] = 8'b0;
    XRAM[58509] = 8'b0;
    XRAM[58510] = 8'b0;
    XRAM[58511] = 8'b0;
    XRAM[58512] = 8'b0;
    XRAM[58513] = 8'b0;
    XRAM[58514] = 8'b0;
    XRAM[58515] = 8'b0;
    XRAM[58516] = 8'b0;
    XRAM[58517] = 8'b0;
    XRAM[58518] = 8'b0;
    XRAM[58519] = 8'b0;
    XRAM[58520] = 8'b0;
    XRAM[58521] = 8'b0;
    XRAM[58522] = 8'b0;
    XRAM[58523] = 8'b0;
    XRAM[58524] = 8'b0;
    XRAM[58525] = 8'b0;
    XRAM[58526] = 8'b0;
    XRAM[58527] = 8'b0;
    XRAM[58528] = 8'b0;
    XRAM[58529] = 8'b0;
    XRAM[58530] = 8'b0;
    XRAM[58531] = 8'b0;
    XRAM[58532] = 8'b0;
    XRAM[58533] = 8'b0;
    XRAM[58534] = 8'b0;
    XRAM[58535] = 8'b0;
    XRAM[58536] = 8'b0;
    XRAM[58537] = 8'b0;
    XRAM[58538] = 8'b0;
    XRAM[58539] = 8'b0;
    XRAM[58540] = 8'b0;
    XRAM[58541] = 8'b0;
    XRAM[58542] = 8'b0;
    XRAM[58543] = 8'b0;
    XRAM[58544] = 8'b0;
    XRAM[58545] = 8'b0;
    XRAM[58546] = 8'b0;
    XRAM[58547] = 8'b0;
    XRAM[58548] = 8'b0;
    XRAM[58549] = 8'b0;
    XRAM[58550] = 8'b0;
    XRAM[58551] = 8'b0;
    XRAM[58552] = 8'b0;
    XRAM[58553] = 8'b0;
    XRAM[58554] = 8'b0;
    XRAM[58555] = 8'b0;
    XRAM[58556] = 8'b0;
    XRAM[58557] = 8'b0;
    XRAM[58558] = 8'b0;
    XRAM[58559] = 8'b0;
    XRAM[58560] = 8'b0;
    XRAM[58561] = 8'b0;
    XRAM[58562] = 8'b0;
    XRAM[58563] = 8'b0;
    XRAM[58564] = 8'b0;
    XRAM[58565] = 8'b0;
    XRAM[58566] = 8'b0;
    XRAM[58567] = 8'b0;
    XRAM[58568] = 8'b0;
    XRAM[58569] = 8'b0;
    XRAM[58570] = 8'b0;
    XRAM[58571] = 8'b0;
    XRAM[58572] = 8'b0;
    XRAM[58573] = 8'b0;
    XRAM[58574] = 8'b0;
    XRAM[58575] = 8'b0;
    XRAM[58576] = 8'b0;
    XRAM[58577] = 8'b0;
    XRAM[58578] = 8'b0;
    XRAM[58579] = 8'b0;
    XRAM[58580] = 8'b0;
    XRAM[58581] = 8'b0;
    XRAM[58582] = 8'b0;
    XRAM[58583] = 8'b0;
    XRAM[58584] = 8'b0;
    XRAM[58585] = 8'b0;
    XRAM[58586] = 8'b0;
    XRAM[58587] = 8'b0;
    XRAM[58588] = 8'b0;
    XRAM[58589] = 8'b0;
    XRAM[58590] = 8'b0;
    XRAM[58591] = 8'b0;
    XRAM[58592] = 8'b0;
    XRAM[58593] = 8'b0;
    XRAM[58594] = 8'b0;
    XRAM[58595] = 8'b0;
    XRAM[58596] = 8'b0;
    XRAM[58597] = 8'b0;
    XRAM[58598] = 8'b0;
    XRAM[58599] = 8'b0;
    XRAM[58600] = 8'b0;
    XRAM[58601] = 8'b0;
    XRAM[58602] = 8'b0;
    XRAM[58603] = 8'b0;
    XRAM[58604] = 8'b0;
    XRAM[58605] = 8'b0;
    XRAM[58606] = 8'b0;
    XRAM[58607] = 8'b0;
    XRAM[58608] = 8'b0;
    XRAM[58609] = 8'b0;
    XRAM[58610] = 8'b0;
    XRAM[58611] = 8'b0;
    XRAM[58612] = 8'b0;
    XRAM[58613] = 8'b0;
    XRAM[58614] = 8'b0;
    XRAM[58615] = 8'b0;
    XRAM[58616] = 8'b0;
    XRAM[58617] = 8'b0;
    XRAM[58618] = 8'b0;
    XRAM[58619] = 8'b0;
    XRAM[58620] = 8'b0;
    XRAM[58621] = 8'b0;
    XRAM[58622] = 8'b0;
    XRAM[58623] = 8'b0;
    XRAM[58624] = 8'b0;
    XRAM[58625] = 8'b0;
    XRAM[58626] = 8'b0;
    XRAM[58627] = 8'b0;
    XRAM[58628] = 8'b0;
    XRAM[58629] = 8'b0;
    XRAM[58630] = 8'b0;
    XRAM[58631] = 8'b0;
    XRAM[58632] = 8'b0;
    XRAM[58633] = 8'b0;
    XRAM[58634] = 8'b0;
    XRAM[58635] = 8'b0;
    XRAM[58636] = 8'b0;
    XRAM[58637] = 8'b0;
    XRAM[58638] = 8'b0;
    XRAM[58639] = 8'b0;
    XRAM[58640] = 8'b0;
    XRAM[58641] = 8'b0;
    XRAM[58642] = 8'b0;
    XRAM[58643] = 8'b0;
    XRAM[58644] = 8'b0;
    XRAM[58645] = 8'b0;
    XRAM[58646] = 8'b0;
    XRAM[58647] = 8'b0;
    XRAM[58648] = 8'b0;
    XRAM[58649] = 8'b0;
    XRAM[58650] = 8'b0;
    XRAM[58651] = 8'b0;
    XRAM[58652] = 8'b0;
    XRAM[58653] = 8'b0;
    XRAM[58654] = 8'b0;
    XRAM[58655] = 8'b0;
    XRAM[58656] = 8'b0;
    XRAM[58657] = 8'b0;
    XRAM[58658] = 8'b0;
    XRAM[58659] = 8'b0;
    XRAM[58660] = 8'b0;
    XRAM[58661] = 8'b0;
    XRAM[58662] = 8'b0;
    XRAM[58663] = 8'b0;
    XRAM[58664] = 8'b0;
    XRAM[58665] = 8'b0;
    XRAM[58666] = 8'b0;
    XRAM[58667] = 8'b0;
    XRAM[58668] = 8'b0;
    XRAM[58669] = 8'b0;
    XRAM[58670] = 8'b0;
    XRAM[58671] = 8'b0;
    XRAM[58672] = 8'b0;
    XRAM[58673] = 8'b0;
    XRAM[58674] = 8'b0;
    XRAM[58675] = 8'b0;
    XRAM[58676] = 8'b0;
    XRAM[58677] = 8'b0;
    XRAM[58678] = 8'b0;
    XRAM[58679] = 8'b0;
    XRAM[58680] = 8'b0;
    XRAM[58681] = 8'b0;
    XRAM[58682] = 8'b0;
    XRAM[58683] = 8'b0;
    XRAM[58684] = 8'b0;
    XRAM[58685] = 8'b0;
    XRAM[58686] = 8'b0;
    XRAM[58687] = 8'b0;
    XRAM[58688] = 8'b0;
    XRAM[58689] = 8'b0;
    XRAM[58690] = 8'b0;
    XRAM[58691] = 8'b0;
    XRAM[58692] = 8'b0;
    XRAM[58693] = 8'b0;
    XRAM[58694] = 8'b0;
    XRAM[58695] = 8'b0;
    XRAM[58696] = 8'b0;
    XRAM[58697] = 8'b0;
    XRAM[58698] = 8'b0;
    XRAM[58699] = 8'b0;
    XRAM[58700] = 8'b0;
    XRAM[58701] = 8'b0;
    XRAM[58702] = 8'b0;
    XRAM[58703] = 8'b0;
    XRAM[58704] = 8'b0;
    XRAM[58705] = 8'b0;
    XRAM[58706] = 8'b0;
    XRAM[58707] = 8'b0;
    XRAM[58708] = 8'b0;
    XRAM[58709] = 8'b0;
    XRAM[58710] = 8'b0;
    XRAM[58711] = 8'b0;
    XRAM[58712] = 8'b0;
    XRAM[58713] = 8'b0;
    XRAM[58714] = 8'b0;
    XRAM[58715] = 8'b0;
    XRAM[58716] = 8'b0;
    XRAM[58717] = 8'b0;
    XRAM[58718] = 8'b0;
    XRAM[58719] = 8'b0;
    XRAM[58720] = 8'b0;
    XRAM[58721] = 8'b0;
    XRAM[58722] = 8'b0;
    XRAM[58723] = 8'b0;
    XRAM[58724] = 8'b0;
    XRAM[58725] = 8'b0;
    XRAM[58726] = 8'b0;
    XRAM[58727] = 8'b0;
    XRAM[58728] = 8'b0;
    XRAM[58729] = 8'b0;
    XRAM[58730] = 8'b0;
    XRAM[58731] = 8'b0;
    XRAM[58732] = 8'b0;
    XRAM[58733] = 8'b0;
    XRAM[58734] = 8'b0;
    XRAM[58735] = 8'b0;
    XRAM[58736] = 8'b0;
    XRAM[58737] = 8'b0;
    XRAM[58738] = 8'b0;
    XRAM[58739] = 8'b0;
    XRAM[58740] = 8'b0;
    XRAM[58741] = 8'b0;
    XRAM[58742] = 8'b0;
    XRAM[58743] = 8'b0;
    XRAM[58744] = 8'b0;
    XRAM[58745] = 8'b0;
    XRAM[58746] = 8'b0;
    XRAM[58747] = 8'b0;
    XRAM[58748] = 8'b0;
    XRAM[58749] = 8'b0;
    XRAM[58750] = 8'b0;
    XRAM[58751] = 8'b0;
    XRAM[58752] = 8'b0;
    XRAM[58753] = 8'b0;
    XRAM[58754] = 8'b0;
    XRAM[58755] = 8'b0;
    XRAM[58756] = 8'b0;
    XRAM[58757] = 8'b0;
    XRAM[58758] = 8'b0;
    XRAM[58759] = 8'b0;
    XRAM[58760] = 8'b0;
    XRAM[58761] = 8'b0;
    XRAM[58762] = 8'b0;
    XRAM[58763] = 8'b0;
    XRAM[58764] = 8'b0;
    XRAM[58765] = 8'b0;
    XRAM[58766] = 8'b0;
    XRAM[58767] = 8'b0;
    XRAM[58768] = 8'b0;
    XRAM[58769] = 8'b0;
    XRAM[58770] = 8'b0;
    XRAM[58771] = 8'b0;
    XRAM[58772] = 8'b0;
    XRAM[58773] = 8'b0;
    XRAM[58774] = 8'b0;
    XRAM[58775] = 8'b0;
    XRAM[58776] = 8'b0;
    XRAM[58777] = 8'b0;
    XRAM[58778] = 8'b0;
    XRAM[58779] = 8'b0;
    XRAM[58780] = 8'b0;
    XRAM[58781] = 8'b0;
    XRAM[58782] = 8'b0;
    XRAM[58783] = 8'b0;
    XRAM[58784] = 8'b0;
    XRAM[58785] = 8'b0;
    XRAM[58786] = 8'b0;
    XRAM[58787] = 8'b0;
    XRAM[58788] = 8'b0;
    XRAM[58789] = 8'b0;
    XRAM[58790] = 8'b0;
    XRAM[58791] = 8'b0;
    XRAM[58792] = 8'b0;
    XRAM[58793] = 8'b0;
    XRAM[58794] = 8'b0;
    XRAM[58795] = 8'b0;
    XRAM[58796] = 8'b0;
    XRAM[58797] = 8'b0;
    XRAM[58798] = 8'b0;
    XRAM[58799] = 8'b0;
    XRAM[58800] = 8'b0;
    XRAM[58801] = 8'b0;
    XRAM[58802] = 8'b0;
    XRAM[58803] = 8'b0;
    XRAM[58804] = 8'b0;
    XRAM[58805] = 8'b0;
    XRAM[58806] = 8'b0;
    XRAM[58807] = 8'b0;
    XRAM[58808] = 8'b0;
    XRAM[58809] = 8'b0;
    XRAM[58810] = 8'b0;
    XRAM[58811] = 8'b0;
    XRAM[58812] = 8'b0;
    XRAM[58813] = 8'b0;
    XRAM[58814] = 8'b0;
    XRAM[58815] = 8'b0;
    XRAM[58816] = 8'b0;
    XRAM[58817] = 8'b0;
    XRAM[58818] = 8'b0;
    XRAM[58819] = 8'b0;
    XRAM[58820] = 8'b0;
    XRAM[58821] = 8'b0;
    XRAM[58822] = 8'b0;
    XRAM[58823] = 8'b0;
    XRAM[58824] = 8'b0;
    XRAM[58825] = 8'b0;
    XRAM[58826] = 8'b0;
    XRAM[58827] = 8'b0;
    XRAM[58828] = 8'b0;
    XRAM[58829] = 8'b0;
    XRAM[58830] = 8'b0;
    XRAM[58831] = 8'b0;
    XRAM[58832] = 8'b0;
    XRAM[58833] = 8'b0;
    XRAM[58834] = 8'b0;
    XRAM[58835] = 8'b0;
    XRAM[58836] = 8'b0;
    XRAM[58837] = 8'b0;
    XRAM[58838] = 8'b0;
    XRAM[58839] = 8'b0;
    XRAM[58840] = 8'b0;
    XRAM[58841] = 8'b0;
    XRAM[58842] = 8'b0;
    XRAM[58843] = 8'b0;
    XRAM[58844] = 8'b0;
    XRAM[58845] = 8'b0;
    XRAM[58846] = 8'b0;
    XRAM[58847] = 8'b0;
    XRAM[58848] = 8'b0;
    XRAM[58849] = 8'b0;
    XRAM[58850] = 8'b0;
    XRAM[58851] = 8'b0;
    XRAM[58852] = 8'b0;
    XRAM[58853] = 8'b0;
    XRAM[58854] = 8'b0;
    XRAM[58855] = 8'b0;
    XRAM[58856] = 8'b0;
    XRAM[58857] = 8'b0;
    XRAM[58858] = 8'b0;
    XRAM[58859] = 8'b0;
    XRAM[58860] = 8'b0;
    XRAM[58861] = 8'b0;
    XRAM[58862] = 8'b0;
    XRAM[58863] = 8'b0;
    XRAM[58864] = 8'b0;
    XRAM[58865] = 8'b0;
    XRAM[58866] = 8'b0;
    XRAM[58867] = 8'b0;
    XRAM[58868] = 8'b0;
    XRAM[58869] = 8'b0;
    XRAM[58870] = 8'b0;
    XRAM[58871] = 8'b0;
    XRAM[58872] = 8'b0;
    XRAM[58873] = 8'b0;
    XRAM[58874] = 8'b0;
    XRAM[58875] = 8'b0;
    XRAM[58876] = 8'b0;
    XRAM[58877] = 8'b0;
    XRAM[58878] = 8'b0;
    XRAM[58879] = 8'b0;
    XRAM[58880] = 8'b0;
    XRAM[58881] = 8'b0;
    XRAM[58882] = 8'b0;
    XRAM[58883] = 8'b0;
    XRAM[58884] = 8'b0;
    XRAM[58885] = 8'b0;
    XRAM[58886] = 8'b0;
    XRAM[58887] = 8'b0;
    XRAM[58888] = 8'b0;
    XRAM[58889] = 8'b0;
    XRAM[58890] = 8'b0;
    XRAM[58891] = 8'b0;
    XRAM[58892] = 8'b0;
    XRAM[58893] = 8'b0;
    XRAM[58894] = 8'b0;
    XRAM[58895] = 8'b0;
    XRAM[58896] = 8'b0;
    XRAM[58897] = 8'b0;
    XRAM[58898] = 8'b0;
    XRAM[58899] = 8'b0;
    XRAM[58900] = 8'b0;
    XRAM[58901] = 8'b0;
    XRAM[58902] = 8'b0;
    XRAM[58903] = 8'b0;
    XRAM[58904] = 8'b0;
    XRAM[58905] = 8'b0;
    XRAM[58906] = 8'b0;
    XRAM[58907] = 8'b0;
    XRAM[58908] = 8'b0;
    XRAM[58909] = 8'b0;
    XRAM[58910] = 8'b0;
    XRAM[58911] = 8'b0;
    XRAM[58912] = 8'b0;
    XRAM[58913] = 8'b0;
    XRAM[58914] = 8'b0;
    XRAM[58915] = 8'b0;
    XRAM[58916] = 8'b0;
    XRAM[58917] = 8'b0;
    XRAM[58918] = 8'b0;
    XRAM[58919] = 8'b0;
    XRAM[58920] = 8'b0;
    XRAM[58921] = 8'b0;
    XRAM[58922] = 8'b0;
    XRAM[58923] = 8'b0;
    XRAM[58924] = 8'b0;
    XRAM[58925] = 8'b0;
    XRAM[58926] = 8'b0;
    XRAM[58927] = 8'b0;
    XRAM[58928] = 8'b0;
    XRAM[58929] = 8'b0;
    XRAM[58930] = 8'b0;
    XRAM[58931] = 8'b0;
    XRAM[58932] = 8'b0;
    XRAM[58933] = 8'b0;
    XRAM[58934] = 8'b0;
    XRAM[58935] = 8'b0;
    XRAM[58936] = 8'b0;
    XRAM[58937] = 8'b0;
    XRAM[58938] = 8'b0;
    XRAM[58939] = 8'b0;
    XRAM[58940] = 8'b0;
    XRAM[58941] = 8'b0;
    XRAM[58942] = 8'b0;
    XRAM[58943] = 8'b0;
    XRAM[58944] = 8'b0;
    XRAM[58945] = 8'b0;
    XRAM[58946] = 8'b0;
    XRAM[58947] = 8'b0;
    XRAM[58948] = 8'b0;
    XRAM[58949] = 8'b0;
    XRAM[58950] = 8'b0;
    XRAM[58951] = 8'b0;
    XRAM[58952] = 8'b0;
    XRAM[58953] = 8'b0;
    XRAM[58954] = 8'b0;
    XRAM[58955] = 8'b0;
    XRAM[58956] = 8'b0;
    XRAM[58957] = 8'b0;
    XRAM[58958] = 8'b0;
    XRAM[58959] = 8'b0;
    XRAM[58960] = 8'b0;
    XRAM[58961] = 8'b0;
    XRAM[58962] = 8'b0;
    XRAM[58963] = 8'b0;
    XRAM[58964] = 8'b0;
    XRAM[58965] = 8'b0;
    XRAM[58966] = 8'b0;
    XRAM[58967] = 8'b0;
    XRAM[58968] = 8'b0;
    XRAM[58969] = 8'b0;
    XRAM[58970] = 8'b0;
    XRAM[58971] = 8'b0;
    XRAM[58972] = 8'b0;
    XRAM[58973] = 8'b0;
    XRAM[58974] = 8'b0;
    XRAM[58975] = 8'b0;
    XRAM[58976] = 8'b0;
    XRAM[58977] = 8'b0;
    XRAM[58978] = 8'b0;
    XRAM[58979] = 8'b0;
    XRAM[58980] = 8'b0;
    XRAM[58981] = 8'b0;
    XRAM[58982] = 8'b0;
    XRAM[58983] = 8'b0;
    XRAM[58984] = 8'b0;
    XRAM[58985] = 8'b0;
    XRAM[58986] = 8'b0;
    XRAM[58987] = 8'b0;
    XRAM[58988] = 8'b0;
    XRAM[58989] = 8'b0;
    XRAM[58990] = 8'b0;
    XRAM[58991] = 8'b0;
    XRAM[58992] = 8'b0;
    XRAM[58993] = 8'b0;
    XRAM[58994] = 8'b0;
    XRAM[58995] = 8'b0;
    XRAM[58996] = 8'b0;
    XRAM[58997] = 8'b0;
    XRAM[58998] = 8'b0;
    XRAM[58999] = 8'b0;
    XRAM[59000] = 8'b0;
    XRAM[59001] = 8'b0;
    XRAM[59002] = 8'b0;
    XRAM[59003] = 8'b0;
    XRAM[59004] = 8'b0;
    XRAM[59005] = 8'b0;
    XRAM[59006] = 8'b0;
    XRAM[59007] = 8'b0;
    XRAM[59008] = 8'b0;
    XRAM[59009] = 8'b0;
    XRAM[59010] = 8'b0;
    XRAM[59011] = 8'b0;
    XRAM[59012] = 8'b0;
    XRAM[59013] = 8'b0;
    XRAM[59014] = 8'b0;
    XRAM[59015] = 8'b0;
    XRAM[59016] = 8'b0;
    XRAM[59017] = 8'b0;
    XRAM[59018] = 8'b0;
    XRAM[59019] = 8'b0;
    XRAM[59020] = 8'b0;
    XRAM[59021] = 8'b0;
    XRAM[59022] = 8'b0;
    XRAM[59023] = 8'b0;
    XRAM[59024] = 8'b0;
    XRAM[59025] = 8'b0;
    XRAM[59026] = 8'b0;
    XRAM[59027] = 8'b0;
    XRAM[59028] = 8'b0;
    XRAM[59029] = 8'b0;
    XRAM[59030] = 8'b0;
    XRAM[59031] = 8'b0;
    XRAM[59032] = 8'b0;
    XRAM[59033] = 8'b0;
    XRAM[59034] = 8'b0;
    XRAM[59035] = 8'b0;
    XRAM[59036] = 8'b0;
    XRAM[59037] = 8'b0;
    XRAM[59038] = 8'b0;
    XRAM[59039] = 8'b0;
    XRAM[59040] = 8'b0;
    XRAM[59041] = 8'b0;
    XRAM[59042] = 8'b0;
    XRAM[59043] = 8'b0;
    XRAM[59044] = 8'b0;
    XRAM[59045] = 8'b0;
    XRAM[59046] = 8'b0;
    XRAM[59047] = 8'b0;
    XRAM[59048] = 8'b0;
    XRAM[59049] = 8'b0;
    XRAM[59050] = 8'b0;
    XRAM[59051] = 8'b0;
    XRAM[59052] = 8'b0;
    XRAM[59053] = 8'b0;
    XRAM[59054] = 8'b0;
    XRAM[59055] = 8'b0;
    XRAM[59056] = 8'b0;
    XRAM[59057] = 8'b0;
    XRAM[59058] = 8'b0;
    XRAM[59059] = 8'b0;
    XRAM[59060] = 8'b0;
    XRAM[59061] = 8'b0;
    XRAM[59062] = 8'b0;
    XRAM[59063] = 8'b0;
    XRAM[59064] = 8'b0;
    XRAM[59065] = 8'b0;
    XRAM[59066] = 8'b0;
    XRAM[59067] = 8'b0;
    XRAM[59068] = 8'b0;
    XRAM[59069] = 8'b0;
    XRAM[59070] = 8'b0;
    XRAM[59071] = 8'b0;
    XRAM[59072] = 8'b0;
    XRAM[59073] = 8'b0;
    XRAM[59074] = 8'b0;
    XRAM[59075] = 8'b0;
    XRAM[59076] = 8'b0;
    XRAM[59077] = 8'b0;
    XRAM[59078] = 8'b0;
    XRAM[59079] = 8'b0;
    XRAM[59080] = 8'b0;
    XRAM[59081] = 8'b0;
    XRAM[59082] = 8'b0;
    XRAM[59083] = 8'b0;
    XRAM[59084] = 8'b0;
    XRAM[59085] = 8'b0;
    XRAM[59086] = 8'b0;
    XRAM[59087] = 8'b0;
    XRAM[59088] = 8'b0;
    XRAM[59089] = 8'b0;
    XRAM[59090] = 8'b0;
    XRAM[59091] = 8'b0;
    XRAM[59092] = 8'b0;
    XRAM[59093] = 8'b0;
    XRAM[59094] = 8'b0;
    XRAM[59095] = 8'b0;
    XRAM[59096] = 8'b0;
    XRAM[59097] = 8'b0;
    XRAM[59098] = 8'b0;
    XRAM[59099] = 8'b0;
    XRAM[59100] = 8'b0;
    XRAM[59101] = 8'b0;
    XRAM[59102] = 8'b0;
    XRAM[59103] = 8'b0;
    XRAM[59104] = 8'b0;
    XRAM[59105] = 8'b0;
    XRAM[59106] = 8'b0;
    XRAM[59107] = 8'b0;
    XRAM[59108] = 8'b0;
    XRAM[59109] = 8'b0;
    XRAM[59110] = 8'b0;
    XRAM[59111] = 8'b0;
    XRAM[59112] = 8'b0;
    XRAM[59113] = 8'b0;
    XRAM[59114] = 8'b0;
    XRAM[59115] = 8'b0;
    XRAM[59116] = 8'b0;
    XRAM[59117] = 8'b0;
    XRAM[59118] = 8'b0;
    XRAM[59119] = 8'b0;
    XRAM[59120] = 8'b0;
    XRAM[59121] = 8'b0;
    XRAM[59122] = 8'b0;
    XRAM[59123] = 8'b0;
    XRAM[59124] = 8'b0;
    XRAM[59125] = 8'b0;
    XRAM[59126] = 8'b0;
    XRAM[59127] = 8'b0;
    XRAM[59128] = 8'b0;
    XRAM[59129] = 8'b0;
    XRAM[59130] = 8'b0;
    XRAM[59131] = 8'b0;
    XRAM[59132] = 8'b0;
    XRAM[59133] = 8'b0;
    XRAM[59134] = 8'b0;
    XRAM[59135] = 8'b0;
    XRAM[59136] = 8'b0;
    XRAM[59137] = 8'b0;
    XRAM[59138] = 8'b0;
    XRAM[59139] = 8'b0;
    XRAM[59140] = 8'b0;
    XRAM[59141] = 8'b0;
    XRAM[59142] = 8'b0;
    XRAM[59143] = 8'b0;
    XRAM[59144] = 8'b0;
    XRAM[59145] = 8'b0;
    XRAM[59146] = 8'b0;
    XRAM[59147] = 8'b0;
    XRAM[59148] = 8'b0;
    XRAM[59149] = 8'b0;
    XRAM[59150] = 8'b0;
    XRAM[59151] = 8'b0;
    XRAM[59152] = 8'b0;
    XRAM[59153] = 8'b0;
    XRAM[59154] = 8'b0;
    XRAM[59155] = 8'b0;
    XRAM[59156] = 8'b0;
    XRAM[59157] = 8'b0;
    XRAM[59158] = 8'b0;
    XRAM[59159] = 8'b0;
    XRAM[59160] = 8'b0;
    XRAM[59161] = 8'b0;
    XRAM[59162] = 8'b0;
    XRAM[59163] = 8'b0;
    XRAM[59164] = 8'b0;
    XRAM[59165] = 8'b0;
    XRAM[59166] = 8'b0;
    XRAM[59167] = 8'b0;
    XRAM[59168] = 8'b0;
    XRAM[59169] = 8'b0;
    XRAM[59170] = 8'b0;
    XRAM[59171] = 8'b0;
    XRAM[59172] = 8'b0;
    XRAM[59173] = 8'b0;
    XRAM[59174] = 8'b0;
    XRAM[59175] = 8'b0;
    XRAM[59176] = 8'b0;
    XRAM[59177] = 8'b0;
    XRAM[59178] = 8'b0;
    XRAM[59179] = 8'b0;
    XRAM[59180] = 8'b0;
    XRAM[59181] = 8'b0;
    XRAM[59182] = 8'b0;
    XRAM[59183] = 8'b0;
    XRAM[59184] = 8'b0;
    XRAM[59185] = 8'b0;
    XRAM[59186] = 8'b0;
    XRAM[59187] = 8'b0;
    XRAM[59188] = 8'b0;
    XRAM[59189] = 8'b0;
    XRAM[59190] = 8'b0;
    XRAM[59191] = 8'b0;
    XRAM[59192] = 8'b0;
    XRAM[59193] = 8'b0;
    XRAM[59194] = 8'b0;
    XRAM[59195] = 8'b0;
    XRAM[59196] = 8'b0;
    XRAM[59197] = 8'b0;
    XRAM[59198] = 8'b0;
    XRAM[59199] = 8'b0;
    XRAM[59200] = 8'b0;
    XRAM[59201] = 8'b0;
    XRAM[59202] = 8'b0;
    XRAM[59203] = 8'b0;
    XRAM[59204] = 8'b0;
    XRAM[59205] = 8'b0;
    XRAM[59206] = 8'b0;
    XRAM[59207] = 8'b0;
    XRAM[59208] = 8'b0;
    XRAM[59209] = 8'b0;
    XRAM[59210] = 8'b0;
    XRAM[59211] = 8'b0;
    XRAM[59212] = 8'b0;
    XRAM[59213] = 8'b0;
    XRAM[59214] = 8'b0;
    XRAM[59215] = 8'b0;
    XRAM[59216] = 8'b0;
    XRAM[59217] = 8'b0;
    XRAM[59218] = 8'b0;
    XRAM[59219] = 8'b0;
    XRAM[59220] = 8'b0;
    XRAM[59221] = 8'b0;
    XRAM[59222] = 8'b0;
    XRAM[59223] = 8'b0;
    XRAM[59224] = 8'b0;
    XRAM[59225] = 8'b0;
    XRAM[59226] = 8'b0;
    XRAM[59227] = 8'b0;
    XRAM[59228] = 8'b0;
    XRAM[59229] = 8'b0;
    XRAM[59230] = 8'b0;
    XRAM[59231] = 8'b0;
    XRAM[59232] = 8'b0;
    XRAM[59233] = 8'b0;
    XRAM[59234] = 8'b0;
    XRAM[59235] = 8'b0;
    XRAM[59236] = 8'b0;
    XRAM[59237] = 8'b0;
    XRAM[59238] = 8'b0;
    XRAM[59239] = 8'b0;
    XRAM[59240] = 8'b0;
    XRAM[59241] = 8'b0;
    XRAM[59242] = 8'b0;
    XRAM[59243] = 8'b0;
    XRAM[59244] = 8'b0;
    XRAM[59245] = 8'b0;
    XRAM[59246] = 8'b0;
    XRAM[59247] = 8'b0;
    XRAM[59248] = 8'b0;
    XRAM[59249] = 8'b0;
    XRAM[59250] = 8'b0;
    XRAM[59251] = 8'b0;
    XRAM[59252] = 8'b0;
    XRAM[59253] = 8'b0;
    XRAM[59254] = 8'b0;
    XRAM[59255] = 8'b0;
    XRAM[59256] = 8'b0;
    XRAM[59257] = 8'b0;
    XRAM[59258] = 8'b0;
    XRAM[59259] = 8'b0;
    XRAM[59260] = 8'b0;
    XRAM[59261] = 8'b0;
    XRAM[59262] = 8'b0;
    XRAM[59263] = 8'b0;
    XRAM[59264] = 8'b0;
    XRAM[59265] = 8'b0;
    XRAM[59266] = 8'b0;
    XRAM[59267] = 8'b0;
    XRAM[59268] = 8'b0;
    XRAM[59269] = 8'b0;
    XRAM[59270] = 8'b0;
    XRAM[59271] = 8'b0;
    XRAM[59272] = 8'b0;
    XRAM[59273] = 8'b0;
    XRAM[59274] = 8'b0;
    XRAM[59275] = 8'b0;
    XRAM[59276] = 8'b0;
    XRAM[59277] = 8'b0;
    XRAM[59278] = 8'b0;
    XRAM[59279] = 8'b0;
    XRAM[59280] = 8'b0;
    XRAM[59281] = 8'b0;
    XRAM[59282] = 8'b0;
    XRAM[59283] = 8'b0;
    XRAM[59284] = 8'b0;
    XRAM[59285] = 8'b0;
    XRAM[59286] = 8'b0;
    XRAM[59287] = 8'b0;
    XRAM[59288] = 8'b0;
    XRAM[59289] = 8'b0;
    XRAM[59290] = 8'b0;
    XRAM[59291] = 8'b0;
    XRAM[59292] = 8'b0;
    XRAM[59293] = 8'b0;
    XRAM[59294] = 8'b0;
    XRAM[59295] = 8'b0;
    XRAM[59296] = 8'b0;
    XRAM[59297] = 8'b0;
    XRAM[59298] = 8'b0;
    XRAM[59299] = 8'b0;
    XRAM[59300] = 8'b0;
    XRAM[59301] = 8'b0;
    XRAM[59302] = 8'b0;
    XRAM[59303] = 8'b0;
    XRAM[59304] = 8'b0;
    XRAM[59305] = 8'b0;
    XRAM[59306] = 8'b0;
    XRAM[59307] = 8'b0;
    XRAM[59308] = 8'b0;
    XRAM[59309] = 8'b0;
    XRAM[59310] = 8'b0;
    XRAM[59311] = 8'b0;
    XRAM[59312] = 8'b0;
    XRAM[59313] = 8'b0;
    XRAM[59314] = 8'b0;
    XRAM[59315] = 8'b0;
    XRAM[59316] = 8'b0;
    XRAM[59317] = 8'b0;
    XRAM[59318] = 8'b0;
    XRAM[59319] = 8'b0;
    XRAM[59320] = 8'b0;
    XRAM[59321] = 8'b0;
    XRAM[59322] = 8'b0;
    XRAM[59323] = 8'b0;
    XRAM[59324] = 8'b0;
    XRAM[59325] = 8'b0;
    XRAM[59326] = 8'b0;
    XRAM[59327] = 8'b0;
    XRAM[59328] = 8'b0;
    XRAM[59329] = 8'b0;
    XRAM[59330] = 8'b0;
    XRAM[59331] = 8'b0;
    XRAM[59332] = 8'b0;
    XRAM[59333] = 8'b0;
    XRAM[59334] = 8'b0;
    XRAM[59335] = 8'b0;
    XRAM[59336] = 8'b0;
    XRAM[59337] = 8'b0;
    XRAM[59338] = 8'b0;
    XRAM[59339] = 8'b0;
    XRAM[59340] = 8'b0;
    XRAM[59341] = 8'b0;
    XRAM[59342] = 8'b0;
    XRAM[59343] = 8'b0;
    XRAM[59344] = 8'b0;
    XRAM[59345] = 8'b0;
    XRAM[59346] = 8'b0;
    XRAM[59347] = 8'b0;
    XRAM[59348] = 8'b0;
    XRAM[59349] = 8'b0;
    XRAM[59350] = 8'b0;
    XRAM[59351] = 8'b0;
    XRAM[59352] = 8'b0;
    XRAM[59353] = 8'b0;
    XRAM[59354] = 8'b0;
    XRAM[59355] = 8'b0;
    XRAM[59356] = 8'b0;
    XRAM[59357] = 8'b0;
    XRAM[59358] = 8'b0;
    XRAM[59359] = 8'b0;
    XRAM[59360] = 8'b0;
    XRAM[59361] = 8'b0;
    XRAM[59362] = 8'b0;
    XRAM[59363] = 8'b0;
    XRAM[59364] = 8'b0;
    XRAM[59365] = 8'b0;
    XRAM[59366] = 8'b0;
    XRAM[59367] = 8'b0;
    XRAM[59368] = 8'b0;
    XRAM[59369] = 8'b0;
    XRAM[59370] = 8'b0;
    XRAM[59371] = 8'b0;
    XRAM[59372] = 8'b0;
    XRAM[59373] = 8'b0;
    XRAM[59374] = 8'b0;
    XRAM[59375] = 8'b0;
    XRAM[59376] = 8'b0;
    XRAM[59377] = 8'b0;
    XRAM[59378] = 8'b0;
    XRAM[59379] = 8'b0;
    XRAM[59380] = 8'b0;
    XRAM[59381] = 8'b0;
    XRAM[59382] = 8'b0;
    XRAM[59383] = 8'b0;
    XRAM[59384] = 8'b0;
    XRAM[59385] = 8'b0;
    XRAM[59386] = 8'b0;
    XRAM[59387] = 8'b0;
    XRAM[59388] = 8'b0;
    XRAM[59389] = 8'b0;
    XRAM[59390] = 8'b0;
    XRAM[59391] = 8'b0;
    XRAM[59392] = 8'b0;
    XRAM[59393] = 8'b0;
    XRAM[59394] = 8'b0;
    XRAM[59395] = 8'b0;
    XRAM[59396] = 8'b0;
    XRAM[59397] = 8'b0;
    XRAM[59398] = 8'b0;
    XRAM[59399] = 8'b0;
    XRAM[59400] = 8'b0;
    XRAM[59401] = 8'b0;
    XRAM[59402] = 8'b0;
    XRAM[59403] = 8'b0;
    XRAM[59404] = 8'b0;
    XRAM[59405] = 8'b0;
    XRAM[59406] = 8'b0;
    XRAM[59407] = 8'b0;
    XRAM[59408] = 8'b0;
    XRAM[59409] = 8'b0;
    XRAM[59410] = 8'b0;
    XRAM[59411] = 8'b0;
    XRAM[59412] = 8'b0;
    XRAM[59413] = 8'b0;
    XRAM[59414] = 8'b0;
    XRAM[59415] = 8'b0;
    XRAM[59416] = 8'b0;
    XRAM[59417] = 8'b0;
    XRAM[59418] = 8'b0;
    XRAM[59419] = 8'b0;
    XRAM[59420] = 8'b0;
    XRAM[59421] = 8'b0;
    XRAM[59422] = 8'b0;
    XRAM[59423] = 8'b0;
    XRAM[59424] = 8'b0;
    XRAM[59425] = 8'b0;
    XRAM[59426] = 8'b0;
    XRAM[59427] = 8'b0;
    XRAM[59428] = 8'b0;
    XRAM[59429] = 8'b0;
    XRAM[59430] = 8'b0;
    XRAM[59431] = 8'b0;
    XRAM[59432] = 8'b0;
    XRAM[59433] = 8'b0;
    XRAM[59434] = 8'b0;
    XRAM[59435] = 8'b0;
    XRAM[59436] = 8'b0;
    XRAM[59437] = 8'b0;
    XRAM[59438] = 8'b0;
    XRAM[59439] = 8'b0;
    XRAM[59440] = 8'b0;
    XRAM[59441] = 8'b0;
    XRAM[59442] = 8'b0;
    XRAM[59443] = 8'b0;
    XRAM[59444] = 8'b0;
    XRAM[59445] = 8'b0;
    XRAM[59446] = 8'b0;
    XRAM[59447] = 8'b0;
    XRAM[59448] = 8'b0;
    XRAM[59449] = 8'b0;
    XRAM[59450] = 8'b0;
    XRAM[59451] = 8'b0;
    XRAM[59452] = 8'b0;
    XRAM[59453] = 8'b0;
    XRAM[59454] = 8'b0;
    XRAM[59455] = 8'b0;
    XRAM[59456] = 8'b0;
    XRAM[59457] = 8'b0;
    XRAM[59458] = 8'b0;
    XRAM[59459] = 8'b0;
    XRAM[59460] = 8'b0;
    XRAM[59461] = 8'b0;
    XRAM[59462] = 8'b0;
    XRAM[59463] = 8'b0;
    XRAM[59464] = 8'b0;
    XRAM[59465] = 8'b0;
    XRAM[59466] = 8'b0;
    XRAM[59467] = 8'b0;
    XRAM[59468] = 8'b0;
    XRAM[59469] = 8'b0;
    XRAM[59470] = 8'b0;
    XRAM[59471] = 8'b0;
    XRAM[59472] = 8'b0;
    XRAM[59473] = 8'b0;
    XRAM[59474] = 8'b0;
    XRAM[59475] = 8'b0;
    XRAM[59476] = 8'b0;
    XRAM[59477] = 8'b0;
    XRAM[59478] = 8'b0;
    XRAM[59479] = 8'b0;
    XRAM[59480] = 8'b0;
    XRAM[59481] = 8'b0;
    XRAM[59482] = 8'b0;
    XRAM[59483] = 8'b0;
    XRAM[59484] = 8'b0;
    XRAM[59485] = 8'b0;
    XRAM[59486] = 8'b0;
    XRAM[59487] = 8'b0;
    XRAM[59488] = 8'b0;
    XRAM[59489] = 8'b0;
    XRAM[59490] = 8'b0;
    XRAM[59491] = 8'b0;
    XRAM[59492] = 8'b0;
    XRAM[59493] = 8'b0;
    XRAM[59494] = 8'b0;
    XRAM[59495] = 8'b0;
    XRAM[59496] = 8'b0;
    XRAM[59497] = 8'b0;
    XRAM[59498] = 8'b0;
    XRAM[59499] = 8'b0;
    XRAM[59500] = 8'b0;
    XRAM[59501] = 8'b0;
    XRAM[59502] = 8'b0;
    XRAM[59503] = 8'b0;
    XRAM[59504] = 8'b0;
    XRAM[59505] = 8'b0;
    XRAM[59506] = 8'b0;
    XRAM[59507] = 8'b0;
    XRAM[59508] = 8'b0;
    XRAM[59509] = 8'b0;
    XRAM[59510] = 8'b0;
    XRAM[59511] = 8'b0;
    XRAM[59512] = 8'b0;
    XRAM[59513] = 8'b0;
    XRAM[59514] = 8'b0;
    XRAM[59515] = 8'b0;
    XRAM[59516] = 8'b0;
    XRAM[59517] = 8'b0;
    XRAM[59518] = 8'b0;
    XRAM[59519] = 8'b0;
    XRAM[59520] = 8'b0;
    XRAM[59521] = 8'b0;
    XRAM[59522] = 8'b0;
    XRAM[59523] = 8'b0;
    XRAM[59524] = 8'b0;
    XRAM[59525] = 8'b0;
    XRAM[59526] = 8'b0;
    XRAM[59527] = 8'b0;
    XRAM[59528] = 8'b0;
    XRAM[59529] = 8'b0;
    XRAM[59530] = 8'b0;
    XRAM[59531] = 8'b0;
    XRAM[59532] = 8'b0;
    XRAM[59533] = 8'b0;
    XRAM[59534] = 8'b0;
    XRAM[59535] = 8'b0;
    XRAM[59536] = 8'b0;
    XRAM[59537] = 8'b0;
    XRAM[59538] = 8'b0;
    XRAM[59539] = 8'b0;
    XRAM[59540] = 8'b0;
    XRAM[59541] = 8'b0;
    XRAM[59542] = 8'b0;
    XRAM[59543] = 8'b0;
    XRAM[59544] = 8'b0;
    XRAM[59545] = 8'b0;
    XRAM[59546] = 8'b0;
    XRAM[59547] = 8'b0;
    XRAM[59548] = 8'b0;
    XRAM[59549] = 8'b0;
    XRAM[59550] = 8'b0;
    XRAM[59551] = 8'b0;
    XRAM[59552] = 8'b0;
    XRAM[59553] = 8'b0;
    XRAM[59554] = 8'b0;
    XRAM[59555] = 8'b0;
    XRAM[59556] = 8'b0;
    XRAM[59557] = 8'b0;
    XRAM[59558] = 8'b0;
    XRAM[59559] = 8'b0;
    XRAM[59560] = 8'b0;
    XRAM[59561] = 8'b0;
    XRAM[59562] = 8'b0;
    XRAM[59563] = 8'b0;
    XRAM[59564] = 8'b0;
    XRAM[59565] = 8'b0;
    XRAM[59566] = 8'b0;
    XRAM[59567] = 8'b0;
    XRAM[59568] = 8'b0;
    XRAM[59569] = 8'b0;
    XRAM[59570] = 8'b0;
    XRAM[59571] = 8'b0;
    XRAM[59572] = 8'b0;
    XRAM[59573] = 8'b0;
    XRAM[59574] = 8'b0;
    XRAM[59575] = 8'b0;
    XRAM[59576] = 8'b0;
    XRAM[59577] = 8'b0;
    XRAM[59578] = 8'b0;
    XRAM[59579] = 8'b0;
    XRAM[59580] = 8'b0;
    XRAM[59581] = 8'b0;
    XRAM[59582] = 8'b0;
    XRAM[59583] = 8'b0;
    XRAM[59584] = 8'b0;
    XRAM[59585] = 8'b0;
    XRAM[59586] = 8'b0;
    XRAM[59587] = 8'b0;
    XRAM[59588] = 8'b0;
    XRAM[59589] = 8'b0;
    XRAM[59590] = 8'b0;
    XRAM[59591] = 8'b0;
    XRAM[59592] = 8'b0;
    XRAM[59593] = 8'b0;
    XRAM[59594] = 8'b0;
    XRAM[59595] = 8'b0;
    XRAM[59596] = 8'b0;
    XRAM[59597] = 8'b0;
    XRAM[59598] = 8'b0;
    XRAM[59599] = 8'b0;
    XRAM[59600] = 8'b0;
    XRAM[59601] = 8'b0;
    XRAM[59602] = 8'b0;
    XRAM[59603] = 8'b0;
    XRAM[59604] = 8'b0;
    XRAM[59605] = 8'b0;
    XRAM[59606] = 8'b0;
    XRAM[59607] = 8'b0;
    XRAM[59608] = 8'b0;
    XRAM[59609] = 8'b0;
    XRAM[59610] = 8'b0;
    XRAM[59611] = 8'b0;
    XRAM[59612] = 8'b0;
    XRAM[59613] = 8'b0;
    XRAM[59614] = 8'b0;
    XRAM[59615] = 8'b0;
    XRAM[59616] = 8'b0;
    XRAM[59617] = 8'b0;
    XRAM[59618] = 8'b0;
    XRAM[59619] = 8'b0;
    XRAM[59620] = 8'b0;
    XRAM[59621] = 8'b0;
    XRAM[59622] = 8'b0;
    XRAM[59623] = 8'b0;
    XRAM[59624] = 8'b0;
    XRAM[59625] = 8'b0;
    XRAM[59626] = 8'b0;
    XRAM[59627] = 8'b0;
    XRAM[59628] = 8'b0;
    XRAM[59629] = 8'b0;
    XRAM[59630] = 8'b0;
    XRAM[59631] = 8'b0;
    XRAM[59632] = 8'b0;
    XRAM[59633] = 8'b0;
    XRAM[59634] = 8'b0;
    XRAM[59635] = 8'b0;
    XRAM[59636] = 8'b0;
    XRAM[59637] = 8'b0;
    XRAM[59638] = 8'b0;
    XRAM[59639] = 8'b0;
    XRAM[59640] = 8'b0;
    XRAM[59641] = 8'b0;
    XRAM[59642] = 8'b0;
    XRAM[59643] = 8'b0;
    XRAM[59644] = 8'b0;
    XRAM[59645] = 8'b0;
    XRAM[59646] = 8'b0;
    XRAM[59647] = 8'b0;
    XRAM[59648] = 8'b0;
    XRAM[59649] = 8'b0;
    XRAM[59650] = 8'b0;
    XRAM[59651] = 8'b0;
    XRAM[59652] = 8'b0;
    XRAM[59653] = 8'b0;
    XRAM[59654] = 8'b0;
    XRAM[59655] = 8'b0;
    XRAM[59656] = 8'b0;
    XRAM[59657] = 8'b0;
    XRAM[59658] = 8'b0;
    XRAM[59659] = 8'b0;
    XRAM[59660] = 8'b0;
    XRAM[59661] = 8'b0;
    XRAM[59662] = 8'b0;
    XRAM[59663] = 8'b0;
    XRAM[59664] = 8'b0;
    XRAM[59665] = 8'b0;
    XRAM[59666] = 8'b0;
    XRAM[59667] = 8'b0;
    XRAM[59668] = 8'b0;
    XRAM[59669] = 8'b0;
    XRAM[59670] = 8'b0;
    XRAM[59671] = 8'b0;
    XRAM[59672] = 8'b0;
    XRAM[59673] = 8'b0;
    XRAM[59674] = 8'b0;
    XRAM[59675] = 8'b0;
    XRAM[59676] = 8'b0;
    XRAM[59677] = 8'b0;
    XRAM[59678] = 8'b0;
    XRAM[59679] = 8'b0;
    XRAM[59680] = 8'b0;
    XRAM[59681] = 8'b0;
    XRAM[59682] = 8'b0;
    XRAM[59683] = 8'b0;
    XRAM[59684] = 8'b0;
    XRAM[59685] = 8'b0;
    XRAM[59686] = 8'b0;
    XRAM[59687] = 8'b0;
    XRAM[59688] = 8'b0;
    XRAM[59689] = 8'b0;
    XRAM[59690] = 8'b0;
    XRAM[59691] = 8'b0;
    XRAM[59692] = 8'b0;
    XRAM[59693] = 8'b0;
    XRAM[59694] = 8'b0;
    XRAM[59695] = 8'b0;
    XRAM[59696] = 8'b0;
    XRAM[59697] = 8'b0;
    XRAM[59698] = 8'b0;
    XRAM[59699] = 8'b0;
    XRAM[59700] = 8'b0;
    XRAM[59701] = 8'b0;
    XRAM[59702] = 8'b0;
    XRAM[59703] = 8'b0;
    XRAM[59704] = 8'b0;
    XRAM[59705] = 8'b0;
    XRAM[59706] = 8'b0;
    XRAM[59707] = 8'b0;
    XRAM[59708] = 8'b0;
    XRAM[59709] = 8'b0;
    XRAM[59710] = 8'b0;
    XRAM[59711] = 8'b0;
    XRAM[59712] = 8'b0;
    XRAM[59713] = 8'b0;
    XRAM[59714] = 8'b0;
    XRAM[59715] = 8'b0;
    XRAM[59716] = 8'b0;
    XRAM[59717] = 8'b0;
    XRAM[59718] = 8'b0;
    XRAM[59719] = 8'b0;
    XRAM[59720] = 8'b0;
    XRAM[59721] = 8'b0;
    XRAM[59722] = 8'b0;
    XRAM[59723] = 8'b0;
    XRAM[59724] = 8'b0;
    XRAM[59725] = 8'b0;
    XRAM[59726] = 8'b0;
    XRAM[59727] = 8'b0;
    XRAM[59728] = 8'b0;
    XRAM[59729] = 8'b0;
    XRAM[59730] = 8'b0;
    XRAM[59731] = 8'b0;
    XRAM[59732] = 8'b0;
    XRAM[59733] = 8'b0;
    XRAM[59734] = 8'b0;
    XRAM[59735] = 8'b0;
    XRAM[59736] = 8'b0;
    XRAM[59737] = 8'b0;
    XRAM[59738] = 8'b0;
    XRAM[59739] = 8'b0;
    XRAM[59740] = 8'b0;
    XRAM[59741] = 8'b0;
    XRAM[59742] = 8'b0;
    XRAM[59743] = 8'b0;
    XRAM[59744] = 8'b0;
    XRAM[59745] = 8'b0;
    XRAM[59746] = 8'b0;
    XRAM[59747] = 8'b0;
    XRAM[59748] = 8'b0;
    XRAM[59749] = 8'b0;
    XRAM[59750] = 8'b0;
    XRAM[59751] = 8'b0;
    XRAM[59752] = 8'b0;
    XRAM[59753] = 8'b0;
    XRAM[59754] = 8'b0;
    XRAM[59755] = 8'b0;
    XRAM[59756] = 8'b0;
    XRAM[59757] = 8'b0;
    XRAM[59758] = 8'b0;
    XRAM[59759] = 8'b0;
    XRAM[59760] = 8'b0;
    XRAM[59761] = 8'b0;
    XRAM[59762] = 8'b0;
    XRAM[59763] = 8'b0;
    XRAM[59764] = 8'b0;
    XRAM[59765] = 8'b0;
    XRAM[59766] = 8'b0;
    XRAM[59767] = 8'b0;
    XRAM[59768] = 8'b0;
    XRAM[59769] = 8'b0;
    XRAM[59770] = 8'b0;
    XRAM[59771] = 8'b0;
    XRAM[59772] = 8'b0;
    XRAM[59773] = 8'b0;
    XRAM[59774] = 8'b0;
    XRAM[59775] = 8'b0;
    XRAM[59776] = 8'b0;
    XRAM[59777] = 8'b0;
    XRAM[59778] = 8'b0;
    XRAM[59779] = 8'b0;
    XRAM[59780] = 8'b0;
    XRAM[59781] = 8'b0;
    XRAM[59782] = 8'b0;
    XRAM[59783] = 8'b0;
    XRAM[59784] = 8'b0;
    XRAM[59785] = 8'b0;
    XRAM[59786] = 8'b0;
    XRAM[59787] = 8'b0;
    XRAM[59788] = 8'b0;
    XRAM[59789] = 8'b0;
    XRAM[59790] = 8'b0;
    XRAM[59791] = 8'b0;
    XRAM[59792] = 8'b0;
    XRAM[59793] = 8'b0;
    XRAM[59794] = 8'b0;
    XRAM[59795] = 8'b0;
    XRAM[59796] = 8'b0;
    XRAM[59797] = 8'b0;
    XRAM[59798] = 8'b0;
    XRAM[59799] = 8'b0;
    XRAM[59800] = 8'b0;
    XRAM[59801] = 8'b0;
    XRAM[59802] = 8'b0;
    XRAM[59803] = 8'b0;
    XRAM[59804] = 8'b0;
    XRAM[59805] = 8'b0;
    XRAM[59806] = 8'b0;
    XRAM[59807] = 8'b0;
    XRAM[59808] = 8'b0;
    XRAM[59809] = 8'b0;
    XRAM[59810] = 8'b0;
    XRAM[59811] = 8'b0;
    XRAM[59812] = 8'b0;
    XRAM[59813] = 8'b0;
    XRAM[59814] = 8'b0;
    XRAM[59815] = 8'b0;
    XRAM[59816] = 8'b0;
    XRAM[59817] = 8'b0;
    XRAM[59818] = 8'b0;
    XRAM[59819] = 8'b0;
    XRAM[59820] = 8'b0;
    XRAM[59821] = 8'b0;
    XRAM[59822] = 8'b0;
    XRAM[59823] = 8'b0;
    XRAM[59824] = 8'b0;
    XRAM[59825] = 8'b0;
    XRAM[59826] = 8'b0;
    XRAM[59827] = 8'b0;
    XRAM[59828] = 8'b0;
    XRAM[59829] = 8'b0;
    XRAM[59830] = 8'b0;
    XRAM[59831] = 8'b0;
    XRAM[59832] = 8'b0;
    XRAM[59833] = 8'b0;
    XRAM[59834] = 8'b0;
    XRAM[59835] = 8'b0;
    XRAM[59836] = 8'b0;
    XRAM[59837] = 8'b0;
    XRAM[59838] = 8'b0;
    XRAM[59839] = 8'b0;
    XRAM[59840] = 8'b0;
    XRAM[59841] = 8'b0;
    XRAM[59842] = 8'b0;
    XRAM[59843] = 8'b0;
    XRAM[59844] = 8'b0;
    XRAM[59845] = 8'b0;
    XRAM[59846] = 8'b0;
    XRAM[59847] = 8'b0;
    XRAM[59848] = 8'b0;
    XRAM[59849] = 8'b0;
    XRAM[59850] = 8'b0;
    XRAM[59851] = 8'b0;
    XRAM[59852] = 8'b0;
    XRAM[59853] = 8'b0;
    XRAM[59854] = 8'b0;
    XRAM[59855] = 8'b0;
    XRAM[59856] = 8'b0;
    XRAM[59857] = 8'b0;
    XRAM[59858] = 8'b0;
    XRAM[59859] = 8'b0;
    XRAM[59860] = 8'b0;
    XRAM[59861] = 8'b0;
    XRAM[59862] = 8'b0;
    XRAM[59863] = 8'b0;
    XRAM[59864] = 8'b0;
    XRAM[59865] = 8'b0;
    XRAM[59866] = 8'b0;
    XRAM[59867] = 8'b0;
    XRAM[59868] = 8'b0;
    XRAM[59869] = 8'b0;
    XRAM[59870] = 8'b0;
    XRAM[59871] = 8'b0;
    XRAM[59872] = 8'b0;
    XRAM[59873] = 8'b0;
    XRAM[59874] = 8'b0;
    XRAM[59875] = 8'b0;
    XRAM[59876] = 8'b0;
    XRAM[59877] = 8'b0;
    XRAM[59878] = 8'b0;
    XRAM[59879] = 8'b0;
    XRAM[59880] = 8'b0;
    XRAM[59881] = 8'b0;
    XRAM[59882] = 8'b0;
    XRAM[59883] = 8'b0;
    XRAM[59884] = 8'b0;
    XRAM[59885] = 8'b0;
    XRAM[59886] = 8'b0;
    XRAM[59887] = 8'b0;
    XRAM[59888] = 8'b0;
    XRAM[59889] = 8'b0;
    XRAM[59890] = 8'b0;
    XRAM[59891] = 8'b0;
    XRAM[59892] = 8'b0;
    XRAM[59893] = 8'b0;
    XRAM[59894] = 8'b0;
    XRAM[59895] = 8'b0;
    XRAM[59896] = 8'b0;
    XRAM[59897] = 8'b0;
    XRAM[59898] = 8'b0;
    XRAM[59899] = 8'b0;
    XRAM[59900] = 8'b0;
    XRAM[59901] = 8'b0;
    XRAM[59902] = 8'b0;
    XRAM[59903] = 8'b0;
    XRAM[59904] = 8'b0;
    XRAM[59905] = 8'b0;
    XRAM[59906] = 8'b0;
    XRAM[59907] = 8'b0;
    XRAM[59908] = 8'b0;
    XRAM[59909] = 8'b0;
    XRAM[59910] = 8'b0;
    XRAM[59911] = 8'b0;
    XRAM[59912] = 8'b0;
    XRAM[59913] = 8'b0;
    XRAM[59914] = 8'b0;
    XRAM[59915] = 8'b0;
    XRAM[59916] = 8'b0;
    XRAM[59917] = 8'b0;
    XRAM[59918] = 8'b0;
    XRAM[59919] = 8'b0;
    XRAM[59920] = 8'b0;
    XRAM[59921] = 8'b0;
    XRAM[59922] = 8'b0;
    XRAM[59923] = 8'b0;
    XRAM[59924] = 8'b0;
    XRAM[59925] = 8'b0;
    XRAM[59926] = 8'b0;
    XRAM[59927] = 8'b0;
    XRAM[59928] = 8'b0;
    XRAM[59929] = 8'b0;
    XRAM[59930] = 8'b0;
    XRAM[59931] = 8'b0;
    XRAM[59932] = 8'b0;
    XRAM[59933] = 8'b0;
    XRAM[59934] = 8'b0;
    XRAM[59935] = 8'b0;
    XRAM[59936] = 8'b0;
    XRAM[59937] = 8'b0;
    XRAM[59938] = 8'b0;
    XRAM[59939] = 8'b0;
    XRAM[59940] = 8'b0;
    XRAM[59941] = 8'b0;
    XRAM[59942] = 8'b0;
    XRAM[59943] = 8'b0;
    XRAM[59944] = 8'b0;
    XRAM[59945] = 8'b0;
    XRAM[59946] = 8'b0;
    XRAM[59947] = 8'b0;
    XRAM[59948] = 8'b0;
    XRAM[59949] = 8'b0;
    XRAM[59950] = 8'b0;
    XRAM[59951] = 8'b0;
    XRAM[59952] = 8'b0;
    XRAM[59953] = 8'b0;
    XRAM[59954] = 8'b0;
    XRAM[59955] = 8'b0;
    XRAM[59956] = 8'b0;
    XRAM[59957] = 8'b0;
    XRAM[59958] = 8'b0;
    XRAM[59959] = 8'b0;
    XRAM[59960] = 8'b0;
    XRAM[59961] = 8'b0;
    XRAM[59962] = 8'b0;
    XRAM[59963] = 8'b0;
    XRAM[59964] = 8'b0;
    XRAM[59965] = 8'b0;
    XRAM[59966] = 8'b0;
    XRAM[59967] = 8'b0;
    XRAM[59968] = 8'b0;
    XRAM[59969] = 8'b0;
    XRAM[59970] = 8'b0;
    XRAM[59971] = 8'b0;
    XRAM[59972] = 8'b0;
    XRAM[59973] = 8'b0;
    XRAM[59974] = 8'b0;
    XRAM[59975] = 8'b0;
    XRAM[59976] = 8'b0;
    XRAM[59977] = 8'b0;
    XRAM[59978] = 8'b0;
    XRAM[59979] = 8'b0;
    XRAM[59980] = 8'b0;
    XRAM[59981] = 8'b0;
    XRAM[59982] = 8'b0;
    XRAM[59983] = 8'b0;
    XRAM[59984] = 8'b0;
    XRAM[59985] = 8'b0;
    XRAM[59986] = 8'b0;
    XRAM[59987] = 8'b0;
    XRAM[59988] = 8'b0;
    XRAM[59989] = 8'b0;
    XRAM[59990] = 8'b0;
    XRAM[59991] = 8'b0;
    XRAM[59992] = 8'b0;
    XRAM[59993] = 8'b0;
    XRAM[59994] = 8'b0;
    XRAM[59995] = 8'b0;
    XRAM[59996] = 8'b0;
    XRAM[59997] = 8'b0;
    XRAM[59998] = 8'b0;
    XRAM[59999] = 8'b0;
    XRAM[60000] = 8'b0;
    XRAM[60001] = 8'b0;
    XRAM[60002] = 8'b0;
    XRAM[60003] = 8'b0;
    XRAM[60004] = 8'b0;
    XRAM[60005] = 8'b0;
    XRAM[60006] = 8'b0;
    XRAM[60007] = 8'b0;
    XRAM[60008] = 8'b0;
    XRAM[60009] = 8'b0;
    XRAM[60010] = 8'b0;
    XRAM[60011] = 8'b0;
    XRAM[60012] = 8'b0;
    XRAM[60013] = 8'b0;
    XRAM[60014] = 8'b0;
    XRAM[60015] = 8'b0;
    XRAM[60016] = 8'b0;
    XRAM[60017] = 8'b0;
    XRAM[60018] = 8'b0;
    XRAM[60019] = 8'b0;
    XRAM[60020] = 8'b0;
    XRAM[60021] = 8'b0;
    XRAM[60022] = 8'b0;
    XRAM[60023] = 8'b0;
    XRAM[60024] = 8'b0;
    XRAM[60025] = 8'b0;
    XRAM[60026] = 8'b0;
    XRAM[60027] = 8'b0;
    XRAM[60028] = 8'b0;
    XRAM[60029] = 8'b0;
    XRAM[60030] = 8'b0;
    XRAM[60031] = 8'b0;
    XRAM[60032] = 8'b0;
    XRAM[60033] = 8'b0;
    XRAM[60034] = 8'b0;
    XRAM[60035] = 8'b0;
    XRAM[60036] = 8'b0;
    XRAM[60037] = 8'b0;
    XRAM[60038] = 8'b0;
    XRAM[60039] = 8'b0;
    XRAM[60040] = 8'b0;
    XRAM[60041] = 8'b0;
    XRAM[60042] = 8'b0;
    XRAM[60043] = 8'b0;
    XRAM[60044] = 8'b0;
    XRAM[60045] = 8'b0;
    XRAM[60046] = 8'b0;
    XRAM[60047] = 8'b0;
    XRAM[60048] = 8'b0;
    XRAM[60049] = 8'b0;
    XRAM[60050] = 8'b0;
    XRAM[60051] = 8'b0;
    XRAM[60052] = 8'b0;
    XRAM[60053] = 8'b0;
    XRAM[60054] = 8'b0;
    XRAM[60055] = 8'b0;
    XRAM[60056] = 8'b0;
    XRAM[60057] = 8'b0;
    XRAM[60058] = 8'b0;
    XRAM[60059] = 8'b0;
    XRAM[60060] = 8'b0;
    XRAM[60061] = 8'b0;
    XRAM[60062] = 8'b0;
    XRAM[60063] = 8'b0;
    XRAM[60064] = 8'b0;
    XRAM[60065] = 8'b0;
    XRAM[60066] = 8'b0;
    XRAM[60067] = 8'b0;
    XRAM[60068] = 8'b0;
    XRAM[60069] = 8'b0;
    XRAM[60070] = 8'b0;
    XRAM[60071] = 8'b0;
    XRAM[60072] = 8'b0;
    XRAM[60073] = 8'b0;
    XRAM[60074] = 8'b0;
    XRAM[60075] = 8'b0;
    XRAM[60076] = 8'b0;
    XRAM[60077] = 8'b0;
    XRAM[60078] = 8'b0;
    XRAM[60079] = 8'b0;
    XRAM[60080] = 8'b0;
    XRAM[60081] = 8'b0;
    XRAM[60082] = 8'b0;
    XRAM[60083] = 8'b0;
    XRAM[60084] = 8'b0;
    XRAM[60085] = 8'b0;
    XRAM[60086] = 8'b0;
    XRAM[60087] = 8'b0;
    XRAM[60088] = 8'b0;
    XRAM[60089] = 8'b0;
    XRAM[60090] = 8'b0;
    XRAM[60091] = 8'b0;
    XRAM[60092] = 8'b0;
    XRAM[60093] = 8'b0;
    XRAM[60094] = 8'b0;
    XRAM[60095] = 8'b0;
    XRAM[60096] = 8'b0;
    XRAM[60097] = 8'b0;
    XRAM[60098] = 8'b0;
    XRAM[60099] = 8'b0;
    XRAM[60100] = 8'b0;
    XRAM[60101] = 8'b0;
    XRAM[60102] = 8'b0;
    XRAM[60103] = 8'b0;
    XRAM[60104] = 8'b0;
    XRAM[60105] = 8'b0;
    XRAM[60106] = 8'b0;
    XRAM[60107] = 8'b0;
    XRAM[60108] = 8'b0;
    XRAM[60109] = 8'b0;
    XRAM[60110] = 8'b0;
    XRAM[60111] = 8'b0;
    XRAM[60112] = 8'b0;
    XRAM[60113] = 8'b0;
    XRAM[60114] = 8'b0;
    XRAM[60115] = 8'b0;
    XRAM[60116] = 8'b0;
    XRAM[60117] = 8'b0;
    XRAM[60118] = 8'b0;
    XRAM[60119] = 8'b0;
    XRAM[60120] = 8'b0;
    XRAM[60121] = 8'b0;
    XRAM[60122] = 8'b0;
    XRAM[60123] = 8'b0;
    XRAM[60124] = 8'b0;
    XRAM[60125] = 8'b0;
    XRAM[60126] = 8'b0;
    XRAM[60127] = 8'b0;
    XRAM[60128] = 8'b0;
    XRAM[60129] = 8'b0;
    XRAM[60130] = 8'b0;
    XRAM[60131] = 8'b0;
    XRAM[60132] = 8'b0;
    XRAM[60133] = 8'b0;
    XRAM[60134] = 8'b0;
    XRAM[60135] = 8'b0;
    XRAM[60136] = 8'b0;
    XRAM[60137] = 8'b0;
    XRAM[60138] = 8'b0;
    XRAM[60139] = 8'b0;
    XRAM[60140] = 8'b0;
    XRAM[60141] = 8'b0;
    XRAM[60142] = 8'b0;
    XRAM[60143] = 8'b0;
    XRAM[60144] = 8'b0;
    XRAM[60145] = 8'b0;
    XRAM[60146] = 8'b0;
    XRAM[60147] = 8'b0;
    XRAM[60148] = 8'b0;
    XRAM[60149] = 8'b0;
    XRAM[60150] = 8'b0;
    XRAM[60151] = 8'b0;
    XRAM[60152] = 8'b0;
    XRAM[60153] = 8'b0;
    XRAM[60154] = 8'b0;
    XRAM[60155] = 8'b0;
    XRAM[60156] = 8'b0;
    XRAM[60157] = 8'b0;
    XRAM[60158] = 8'b0;
    XRAM[60159] = 8'b0;
    XRAM[60160] = 8'b0;
    XRAM[60161] = 8'b0;
    XRAM[60162] = 8'b0;
    XRAM[60163] = 8'b0;
    XRAM[60164] = 8'b0;
    XRAM[60165] = 8'b0;
    XRAM[60166] = 8'b0;
    XRAM[60167] = 8'b0;
    XRAM[60168] = 8'b0;
    XRAM[60169] = 8'b0;
    XRAM[60170] = 8'b0;
    XRAM[60171] = 8'b0;
    XRAM[60172] = 8'b0;
    XRAM[60173] = 8'b0;
    XRAM[60174] = 8'b0;
    XRAM[60175] = 8'b0;
    XRAM[60176] = 8'b0;
    XRAM[60177] = 8'b0;
    XRAM[60178] = 8'b0;
    XRAM[60179] = 8'b0;
    XRAM[60180] = 8'b0;
    XRAM[60181] = 8'b0;
    XRAM[60182] = 8'b0;
    XRAM[60183] = 8'b0;
    XRAM[60184] = 8'b0;
    XRAM[60185] = 8'b0;
    XRAM[60186] = 8'b0;
    XRAM[60187] = 8'b0;
    XRAM[60188] = 8'b0;
    XRAM[60189] = 8'b0;
    XRAM[60190] = 8'b0;
    XRAM[60191] = 8'b0;
    XRAM[60192] = 8'b0;
    XRAM[60193] = 8'b0;
    XRAM[60194] = 8'b0;
    XRAM[60195] = 8'b0;
    XRAM[60196] = 8'b0;
    XRAM[60197] = 8'b0;
    XRAM[60198] = 8'b0;
    XRAM[60199] = 8'b0;
    XRAM[60200] = 8'b0;
    XRAM[60201] = 8'b0;
    XRAM[60202] = 8'b0;
    XRAM[60203] = 8'b0;
    XRAM[60204] = 8'b0;
    XRAM[60205] = 8'b0;
    XRAM[60206] = 8'b0;
    XRAM[60207] = 8'b0;
    XRAM[60208] = 8'b0;
    XRAM[60209] = 8'b0;
    XRAM[60210] = 8'b0;
    XRAM[60211] = 8'b0;
    XRAM[60212] = 8'b0;
    XRAM[60213] = 8'b0;
    XRAM[60214] = 8'b0;
    XRAM[60215] = 8'b0;
    XRAM[60216] = 8'b0;
    XRAM[60217] = 8'b0;
    XRAM[60218] = 8'b0;
    XRAM[60219] = 8'b0;
    XRAM[60220] = 8'b0;
    XRAM[60221] = 8'b0;
    XRAM[60222] = 8'b0;
    XRAM[60223] = 8'b0;
    XRAM[60224] = 8'b0;
    XRAM[60225] = 8'b0;
    XRAM[60226] = 8'b0;
    XRAM[60227] = 8'b0;
    XRAM[60228] = 8'b0;
    XRAM[60229] = 8'b0;
    XRAM[60230] = 8'b0;
    XRAM[60231] = 8'b0;
    XRAM[60232] = 8'b0;
    XRAM[60233] = 8'b0;
    XRAM[60234] = 8'b0;
    XRAM[60235] = 8'b0;
    XRAM[60236] = 8'b0;
    XRAM[60237] = 8'b0;
    XRAM[60238] = 8'b0;
    XRAM[60239] = 8'b0;
    XRAM[60240] = 8'b0;
    XRAM[60241] = 8'b0;
    XRAM[60242] = 8'b0;
    XRAM[60243] = 8'b0;
    XRAM[60244] = 8'b0;
    XRAM[60245] = 8'b0;
    XRAM[60246] = 8'b0;
    XRAM[60247] = 8'b0;
    XRAM[60248] = 8'b0;
    XRAM[60249] = 8'b0;
    XRAM[60250] = 8'b0;
    XRAM[60251] = 8'b0;
    XRAM[60252] = 8'b0;
    XRAM[60253] = 8'b0;
    XRAM[60254] = 8'b0;
    XRAM[60255] = 8'b0;
    XRAM[60256] = 8'b0;
    XRAM[60257] = 8'b0;
    XRAM[60258] = 8'b0;
    XRAM[60259] = 8'b0;
    XRAM[60260] = 8'b0;
    XRAM[60261] = 8'b0;
    XRAM[60262] = 8'b0;
    XRAM[60263] = 8'b0;
    XRAM[60264] = 8'b0;
    XRAM[60265] = 8'b0;
    XRAM[60266] = 8'b0;
    XRAM[60267] = 8'b0;
    XRAM[60268] = 8'b0;
    XRAM[60269] = 8'b0;
    XRAM[60270] = 8'b0;
    XRAM[60271] = 8'b0;
    XRAM[60272] = 8'b0;
    XRAM[60273] = 8'b0;
    XRAM[60274] = 8'b0;
    XRAM[60275] = 8'b0;
    XRAM[60276] = 8'b0;
    XRAM[60277] = 8'b0;
    XRAM[60278] = 8'b0;
    XRAM[60279] = 8'b0;
    XRAM[60280] = 8'b0;
    XRAM[60281] = 8'b0;
    XRAM[60282] = 8'b0;
    XRAM[60283] = 8'b0;
    XRAM[60284] = 8'b0;
    XRAM[60285] = 8'b0;
    XRAM[60286] = 8'b0;
    XRAM[60287] = 8'b0;
    XRAM[60288] = 8'b0;
    XRAM[60289] = 8'b0;
    XRAM[60290] = 8'b0;
    XRAM[60291] = 8'b0;
    XRAM[60292] = 8'b0;
    XRAM[60293] = 8'b0;
    XRAM[60294] = 8'b0;
    XRAM[60295] = 8'b0;
    XRAM[60296] = 8'b0;
    XRAM[60297] = 8'b0;
    XRAM[60298] = 8'b0;
    XRAM[60299] = 8'b0;
    XRAM[60300] = 8'b0;
    XRAM[60301] = 8'b0;
    XRAM[60302] = 8'b0;
    XRAM[60303] = 8'b0;
    XRAM[60304] = 8'b0;
    XRAM[60305] = 8'b0;
    XRAM[60306] = 8'b0;
    XRAM[60307] = 8'b0;
    XRAM[60308] = 8'b0;
    XRAM[60309] = 8'b0;
    XRAM[60310] = 8'b0;
    XRAM[60311] = 8'b0;
    XRAM[60312] = 8'b0;
    XRAM[60313] = 8'b0;
    XRAM[60314] = 8'b0;
    XRAM[60315] = 8'b0;
    XRAM[60316] = 8'b0;
    XRAM[60317] = 8'b0;
    XRAM[60318] = 8'b0;
    XRAM[60319] = 8'b0;
    XRAM[60320] = 8'b0;
    XRAM[60321] = 8'b0;
    XRAM[60322] = 8'b0;
    XRAM[60323] = 8'b0;
    XRAM[60324] = 8'b0;
    XRAM[60325] = 8'b0;
    XRAM[60326] = 8'b0;
    XRAM[60327] = 8'b0;
    XRAM[60328] = 8'b0;
    XRAM[60329] = 8'b0;
    XRAM[60330] = 8'b0;
    XRAM[60331] = 8'b0;
    XRAM[60332] = 8'b0;
    XRAM[60333] = 8'b0;
    XRAM[60334] = 8'b0;
    XRAM[60335] = 8'b0;
    XRAM[60336] = 8'b0;
    XRAM[60337] = 8'b0;
    XRAM[60338] = 8'b0;
    XRAM[60339] = 8'b0;
    XRAM[60340] = 8'b0;
    XRAM[60341] = 8'b0;
    XRAM[60342] = 8'b0;
    XRAM[60343] = 8'b0;
    XRAM[60344] = 8'b0;
    XRAM[60345] = 8'b0;
    XRAM[60346] = 8'b0;
    XRAM[60347] = 8'b0;
    XRAM[60348] = 8'b0;
    XRAM[60349] = 8'b0;
    XRAM[60350] = 8'b0;
    XRAM[60351] = 8'b0;
    XRAM[60352] = 8'b0;
    XRAM[60353] = 8'b0;
    XRAM[60354] = 8'b0;
    XRAM[60355] = 8'b0;
    XRAM[60356] = 8'b0;
    XRAM[60357] = 8'b0;
    XRAM[60358] = 8'b0;
    XRAM[60359] = 8'b0;
    XRAM[60360] = 8'b0;
    XRAM[60361] = 8'b0;
    XRAM[60362] = 8'b0;
    XRAM[60363] = 8'b0;
    XRAM[60364] = 8'b0;
    XRAM[60365] = 8'b0;
    XRAM[60366] = 8'b0;
    XRAM[60367] = 8'b0;
    XRAM[60368] = 8'b0;
    XRAM[60369] = 8'b0;
    XRAM[60370] = 8'b0;
    XRAM[60371] = 8'b0;
    XRAM[60372] = 8'b0;
    XRAM[60373] = 8'b0;
    XRAM[60374] = 8'b0;
    XRAM[60375] = 8'b0;
    XRAM[60376] = 8'b0;
    XRAM[60377] = 8'b0;
    XRAM[60378] = 8'b0;
    XRAM[60379] = 8'b0;
    XRAM[60380] = 8'b0;
    XRAM[60381] = 8'b0;
    XRAM[60382] = 8'b0;
    XRAM[60383] = 8'b0;
    XRAM[60384] = 8'b0;
    XRAM[60385] = 8'b0;
    XRAM[60386] = 8'b0;
    XRAM[60387] = 8'b0;
    XRAM[60388] = 8'b0;
    XRAM[60389] = 8'b0;
    XRAM[60390] = 8'b0;
    XRAM[60391] = 8'b0;
    XRAM[60392] = 8'b0;
    XRAM[60393] = 8'b0;
    XRAM[60394] = 8'b0;
    XRAM[60395] = 8'b0;
    XRAM[60396] = 8'b0;
    XRAM[60397] = 8'b0;
    XRAM[60398] = 8'b0;
    XRAM[60399] = 8'b0;
    XRAM[60400] = 8'b0;
    XRAM[60401] = 8'b0;
    XRAM[60402] = 8'b0;
    XRAM[60403] = 8'b0;
    XRAM[60404] = 8'b0;
    XRAM[60405] = 8'b0;
    XRAM[60406] = 8'b0;
    XRAM[60407] = 8'b0;
    XRAM[60408] = 8'b0;
    XRAM[60409] = 8'b0;
    XRAM[60410] = 8'b0;
    XRAM[60411] = 8'b0;
    XRAM[60412] = 8'b0;
    XRAM[60413] = 8'b0;
    XRAM[60414] = 8'b0;
    XRAM[60415] = 8'b0;
    XRAM[60416] = 8'b0;
    XRAM[60417] = 8'b0;
    XRAM[60418] = 8'b0;
    XRAM[60419] = 8'b0;
    XRAM[60420] = 8'b0;
    XRAM[60421] = 8'b0;
    XRAM[60422] = 8'b0;
    XRAM[60423] = 8'b0;
    XRAM[60424] = 8'b0;
    XRAM[60425] = 8'b0;
    XRAM[60426] = 8'b0;
    XRAM[60427] = 8'b0;
    XRAM[60428] = 8'b0;
    XRAM[60429] = 8'b0;
    XRAM[60430] = 8'b0;
    XRAM[60431] = 8'b0;
    XRAM[60432] = 8'b0;
    XRAM[60433] = 8'b0;
    XRAM[60434] = 8'b0;
    XRAM[60435] = 8'b0;
    XRAM[60436] = 8'b0;
    XRAM[60437] = 8'b0;
    XRAM[60438] = 8'b0;
    XRAM[60439] = 8'b0;
    XRAM[60440] = 8'b0;
    XRAM[60441] = 8'b0;
    XRAM[60442] = 8'b0;
    XRAM[60443] = 8'b0;
    XRAM[60444] = 8'b0;
    XRAM[60445] = 8'b0;
    XRAM[60446] = 8'b0;
    XRAM[60447] = 8'b0;
    XRAM[60448] = 8'b0;
    XRAM[60449] = 8'b0;
    XRAM[60450] = 8'b0;
    XRAM[60451] = 8'b0;
    XRAM[60452] = 8'b0;
    XRAM[60453] = 8'b0;
    XRAM[60454] = 8'b0;
    XRAM[60455] = 8'b0;
    XRAM[60456] = 8'b0;
    XRAM[60457] = 8'b0;
    XRAM[60458] = 8'b0;
    XRAM[60459] = 8'b0;
    XRAM[60460] = 8'b0;
    XRAM[60461] = 8'b0;
    XRAM[60462] = 8'b0;
    XRAM[60463] = 8'b0;
    XRAM[60464] = 8'b0;
    XRAM[60465] = 8'b0;
    XRAM[60466] = 8'b0;
    XRAM[60467] = 8'b0;
    XRAM[60468] = 8'b0;
    XRAM[60469] = 8'b0;
    XRAM[60470] = 8'b0;
    XRAM[60471] = 8'b0;
    XRAM[60472] = 8'b0;
    XRAM[60473] = 8'b0;
    XRAM[60474] = 8'b0;
    XRAM[60475] = 8'b0;
    XRAM[60476] = 8'b0;
    XRAM[60477] = 8'b0;
    XRAM[60478] = 8'b0;
    XRAM[60479] = 8'b0;
    XRAM[60480] = 8'b0;
    XRAM[60481] = 8'b0;
    XRAM[60482] = 8'b0;
    XRAM[60483] = 8'b0;
    XRAM[60484] = 8'b0;
    XRAM[60485] = 8'b0;
    XRAM[60486] = 8'b0;
    XRAM[60487] = 8'b0;
    XRAM[60488] = 8'b0;
    XRAM[60489] = 8'b0;
    XRAM[60490] = 8'b0;
    XRAM[60491] = 8'b0;
    XRAM[60492] = 8'b0;
    XRAM[60493] = 8'b0;
    XRAM[60494] = 8'b0;
    XRAM[60495] = 8'b0;
    XRAM[60496] = 8'b0;
    XRAM[60497] = 8'b0;
    XRAM[60498] = 8'b0;
    XRAM[60499] = 8'b0;
    XRAM[60500] = 8'b0;
    XRAM[60501] = 8'b0;
    XRAM[60502] = 8'b0;
    XRAM[60503] = 8'b0;
    XRAM[60504] = 8'b0;
    XRAM[60505] = 8'b0;
    XRAM[60506] = 8'b0;
    XRAM[60507] = 8'b0;
    XRAM[60508] = 8'b0;
    XRAM[60509] = 8'b0;
    XRAM[60510] = 8'b0;
    XRAM[60511] = 8'b0;
    XRAM[60512] = 8'b0;
    XRAM[60513] = 8'b0;
    XRAM[60514] = 8'b0;
    XRAM[60515] = 8'b0;
    XRAM[60516] = 8'b0;
    XRAM[60517] = 8'b0;
    XRAM[60518] = 8'b0;
    XRAM[60519] = 8'b0;
    XRAM[60520] = 8'b0;
    XRAM[60521] = 8'b0;
    XRAM[60522] = 8'b0;
    XRAM[60523] = 8'b0;
    XRAM[60524] = 8'b0;
    XRAM[60525] = 8'b0;
    XRAM[60526] = 8'b0;
    XRAM[60527] = 8'b0;
    XRAM[60528] = 8'b0;
    XRAM[60529] = 8'b0;
    XRAM[60530] = 8'b0;
    XRAM[60531] = 8'b0;
    XRAM[60532] = 8'b0;
    XRAM[60533] = 8'b0;
    XRAM[60534] = 8'b0;
    XRAM[60535] = 8'b0;
    XRAM[60536] = 8'b0;
    XRAM[60537] = 8'b0;
    XRAM[60538] = 8'b0;
    XRAM[60539] = 8'b0;
    XRAM[60540] = 8'b0;
    XRAM[60541] = 8'b0;
    XRAM[60542] = 8'b0;
    XRAM[60543] = 8'b0;
    XRAM[60544] = 8'b0;
    XRAM[60545] = 8'b0;
    XRAM[60546] = 8'b0;
    XRAM[60547] = 8'b0;
    XRAM[60548] = 8'b0;
    XRAM[60549] = 8'b0;
    XRAM[60550] = 8'b0;
    XRAM[60551] = 8'b0;
    XRAM[60552] = 8'b0;
    XRAM[60553] = 8'b0;
    XRAM[60554] = 8'b0;
    XRAM[60555] = 8'b0;
    XRAM[60556] = 8'b0;
    XRAM[60557] = 8'b0;
    XRAM[60558] = 8'b0;
    XRAM[60559] = 8'b0;
    XRAM[60560] = 8'b0;
    XRAM[60561] = 8'b0;
    XRAM[60562] = 8'b0;
    XRAM[60563] = 8'b0;
    XRAM[60564] = 8'b0;
    XRAM[60565] = 8'b0;
    XRAM[60566] = 8'b0;
    XRAM[60567] = 8'b0;
    XRAM[60568] = 8'b0;
    XRAM[60569] = 8'b0;
    XRAM[60570] = 8'b0;
    XRAM[60571] = 8'b0;
    XRAM[60572] = 8'b0;
    XRAM[60573] = 8'b0;
    XRAM[60574] = 8'b0;
    XRAM[60575] = 8'b0;
    XRAM[60576] = 8'b0;
    XRAM[60577] = 8'b0;
    XRAM[60578] = 8'b0;
    XRAM[60579] = 8'b0;
    XRAM[60580] = 8'b0;
    XRAM[60581] = 8'b0;
    XRAM[60582] = 8'b0;
    XRAM[60583] = 8'b0;
    XRAM[60584] = 8'b0;
    XRAM[60585] = 8'b0;
    XRAM[60586] = 8'b0;
    XRAM[60587] = 8'b0;
    XRAM[60588] = 8'b0;
    XRAM[60589] = 8'b0;
    XRAM[60590] = 8'b0;
    XRAM[60591] = 8'b0;
    XRAM[60592] = 8'b0;
    XRAM[60593] = 8'b0;
    XRAM[60594] = 8'b0;
    XRAM[60595] = 8'b0;
    XRAM[60596] = 8'b0;
    XRAM[60597] = 8'b0;
    XRAM[60598] = 8'b0;
    XRAM[60599] = 8'b0;
    XRAM[60600] = 8'b0;
    XRAM[60601] = 8'b0;
    XRAM[60602] = 8'b0;
    XRAM[60603] = 8'b0;
    XRAM[60604] = 8'b0;
    XRAM[60605] = 8'b0;
    XRAM[60606] = 8'b0;
    XRAM[60607] = 8'b0;
    XRAM[60608] = 8'b0;
    XRAM[60609] = 8'b0;
    XRAM[60610] = 8'b0;
    XRAM[60611] = 8'b0;
    XRAM[60612] = 8'b0;
    XRAM[60613] = 8'b0;
    XRAM[60614] = 8'b0;
    XRAM[60615] = 8'b0;
    XRAM[60616] = 8'b0;
    XRAM[60617] = 8'b0;
    XRAM[60618] = 8'b0;
    XRAM[60619] = 8'b0;
    XRAM[60620] = 8'b0;
    XRAM[60621] = 8'b0;
    XRAM[60622] = 8'b0;
    XRAM[60623] = 8'b0;
    XRAM[60624] = 8'b0;
    XRAM[60625] = 8'b0;
    XRAM[60626] = 8'b0;
    XRAM[60627] = 8'b0;
    XRAM[60628] = 8'b0;
    XRAM[60629] = 8'b0;
    XRAM[60630] = 8'b0;
    XRAM[60631] = 8'b0;
    XRAM[60632] = 8'b0;
    XRAM[60633] = 8'b0;
    XRAM[60634] = 8'b0;
    XRAM[60635] = 8'b0;
    XRAM[60636] = 8'b0;
    XRAM[60637] = 8'b0;
    XRAM[60638] = 8'b0;
    XRAM[60639] = 8'b0;
    XRAM[60640] = 8'b0;
    XRAM[60641] = 8'b0;
    XRAM[60642] = 8'b0;
    XRAM[60643] = 8'b0;
    XRAM[60644] = 8'b0;
    XRAM[60645] = 8'b0;
    XRAM[60646] = 8'b0;
    XRAM[60647] = 8'b0;
    XRAM[60648] = 8'b0;
    XRAM[60649] = 8'b0;
    XRAM[60650] = 8'b0;
    XRAM[60651] = 8'b0;
    XRAM[60652] = 8'b0;
    XRAM[60653] = 8'b0;
    XRAM[60654] = 8'b0;
    XRAM[60655] = 8'b0;
    XRAM[60656] = 8'b0;
    XRAM[60657] = 8'b0;
    XRAM[60658] = 8'b0;
    XRAM[60659] = 8'b0;
    XRAM[60660] = 8'b0;
    XRAM[60661] = 8'b0;
    XRAM[60662] = 8'b0;
    XRAM[60663] = 8'b0;
    XRAM[60664] = 8'b0;
    XRAM[60665] = 8'b0;
    XRAM[60666] = 8'b0;
    XRAM[60667] = 8'b0;
    XRAM[60668] = 8'b0;
    XRAM[60669] = 8'b0;
    XRAM[60670] = 8'b0;
    XRAM[60671] = 8'b0;
    XRAM[60672] = 8'b0;
    XRAM[60673] = 8'b0;
    XRAM[60674] = 8'b0;
    XRAM[60675] = 8'b0;
    XRAM[60676] = 8'b0;
    XRAM[60677] = 8'b0;
    XRAM[60678] = 8'b0;
    XRAM[60679] = 8'b0;
    XRAM[60680] = 8'b0;
    XRAM[60681] = 8'b0;
    XRAM[60682] = 8'b0;
    XRAM[60683] = 8'b0;
    XRAM[60684] = 8'b0;
    XRAM[60685] = 8'b0;
    XRAM[60686] = 8'b0;
    XRAM[60687] = 8'b0;
    XRAM[60688] = 8'b0;
    XRAM[60689] = 8'b0;
    XRAM[60690] = 8'b0;
    XRAM[60691] = 8'b0;
    XRAM[60692] = 8'b0;
    XRAM[60693] = 8'b0;
    XRAM[60694] = 8'b0;
    XRAM[60695] = 8'b0;
    XRAM[60696] = 8'b0;
    XRAM[60697] = 8'b0;
    XRAM[60698] = 8'b0;
    XRAM[60699] = 8'b0;
    XRAM[60700] = 8'b0;
    XRAM[60701] = 8'b0;
    XRAM[60702] = 8'b0;
    XRAM[60703] = 8'b0;
    XRAM[60704] = 8'b0;
    XRAM[60705] = 8'b0;
    XRAM[60706] = 8'b0;
    XRAM[60707] = 8'b0;
    XRAM[60708] = 8'b0;
    XRAM[60709] = 8'b0;
    XRAM[60710] = 8'b0;
    XRAM[60711] = 8'b0;
    XRAM[60712] = 8'b0;
    XRAM[60713] = 8'b0;
    XRAM[60714] = 8'b0;
    XRAM[60715] = 8'b0;
    XRAM[60716] = 8'b0;
    XRAM[60717] = 8'b0;
    XRAM[60718] = 8'b0;
    XRAM[60719] = 8'b0;
    XRAM[60720] = 8'b0;
    XRAM[60721] = 8'b0;
    XRAM[60722] = 8'b0;
    XRAM[60723] = 8'b0;
    XRAM[60724] = 8'b0;
    XRAM[60725] = 8'b0;
    XRAM[60726] = 8'b0;
    XRAM[60727] = 8'b0;
    XRAM[60728] = 8'b0;
    XRAM[60729] = 8'b0;
    XRAM[60730] = 8'b0;
    XRAM[60731] = 8'b0;
    XRAM[60732] = 8'b0;
    XRAM[60733] = 8'b0;
    XRAM[60734] = 8'b0;
    XRAM[60735] = 8'b0;
    XRAM[60736] = 8'b0;
    XRAM[60737] = 8'b0;
    XRAM[60738] = 8'b0;
    XRAM[60739] = 8'b0;
    XRAM[60740] = 8'b0;
    XRAM[60741] = 8'b0;
    XRAM[60742] = 8'b0;
    XRAM[60743] = 8'b0;
    XRAM[60744] = 8'b0;
    XRAM[60745] = 8'b0;
    XRAM[60746] = 8'b0;
    XRAM[60747] = 8'b0;
    XRAM[60748] = 8'b0;
    XRAM[60749] = 8'b0;
    XRAM[60750] = 8'b0;
    XRAM[60751] = 8'b0;
    XRAM[60752] = 8'b0;
    XRAM[60753] = 8'b0;
    XRAM[60754] = 8'b0;
    XRAM[60755] = 8'b0;
    XRAM[60756] = 8'b0;
    XRAM[60757] = 8'b0;
    XRAM[60758] = 8'b0;
    XRAM[60759] = 8'b0;
    XRAM[60760] = 8'b0;
    XRAM[60761] = 8'b0;
    XRAM[60762] = 8'b0;
    XRAM[60763] = 8'b0;
    XRAM[60764] = 8'b0;
    XRAM[60765] = 8'b0;
    XRAM[60766] = 8'b0;
    XRAM[60767] = 8'b0;
    XRAM[60768] = 8'b0;
    XRAM[60769] = 8'b0;
    XRAM[60770] = 8'b0;
    XRAM[60771] = 8'b0;
    XRAM[60772] = 8'b0;
    XRAM[60773] = 8'b0;
    XRAM[60774] = 8'b0;
    XRAM[60775] = 8'b0;
    XRAM[60776] = 8'b0;
    XRAM[60777] = 8'b0;
    XRAM[60778] = 8'b0;
    XRAM[60779] = 8'b0;
    XRAM[60780] = 8'b0;
    XRAM[60781] = 8'b0;
    XRAM[60782] = 8'b0;
    XRAM[60783] = 8'b0;
    XRAM[60784] = 8'b0;
    XRAM[60785] = 8'b0;
    XRAM[60786] = 8'b0;
    XRAM[60787] = 8'b0;
    XRAM[60788] = 8'b0;
    XRAM[60789] = 8'b0;
    XRAM[60790] = 8'b0;
    XRAM[60791] = 8'b0;
    XRAM[60792] = 8'b0;
    XRAM[60793] = 8'b0;
    XRAM[60794] = 8'b0;
    XRAM[60795] = 8'b0;
    XRAM[60796] = 8'b0;
    XRAM[60797] = 8'b0;
    XRAM[60798] = 8'b0;
    XRAM[60799] = 8'b0;
    XRAM[60800] = 8'b0;
    XRAM[60801] = 8'b0;
    XRAM[60802] = 8'b0;
    XRAM[60803] = 8'b0;
    XRAM[60804] = 8'b0;
    XRAM[60805] = 8'b0;
    XRAM[60806] = 8'b0;
    XRAM[60807] = 8'b0;
    XRAM[60808] = 8'b0;
    XRAM[60809] = 8'b0;
    XRAM[60810] = 8'b0;
    XRAM[60811] = 8'b0;
    XRAM[60812] = 8'b0;
    XRAM[60813] = 8'b0;
    XRAM[60814] = 8'b0;
    XRAM[60815] = 8'b0;
    XRAM[60816] = 8'b0;
    XRAM[60817] = 8'b0;
    XRAM[60818] = 8'b0;
    XRAM[60819] = 8'b0;
    XRAM[60820] = 8'b0;
    XRAM[60821] = 8'b0;
    XRAM[60822] = 8'b0;
    XRAM[60823] = 8'b0;
    XRAM[60824] = 8'b0;
    XRAM[60825] = 8'b0;
    XRAM[60826] = 8'b0;
    XRAM[60827] = 8'b0;
    XRAM[60828] = 8'b0;
    XRAM[60829] = 8'b0;
    XRAM[60830] = 8'b0;
    XRAM[60831] = 8'b0;
    XRAM[60832] = 8'b0;
    XRAM[60833] = 8'b0;
    XRAM[60834] = 8'b0;
    XRAM[60835] = 8'b0;
    XRAM[60836] = 8'b0;
    XRAM[60837] = 8'b0;
    XRAM[60838] = 8'b0;
    XRAM[60839] = 8'b0;
    XRAM[60840] = 8'b0;
    XRAM[60841] = 8'b0;
    XRAM[60842] = 8'b0;
    XRAM[60843] = 8'b0;
    XRAM[60844] = 8'b0;
    XRAM[60845] = 8'b0;
    XRAM[60846] = 8'b0;
    XRAM[60847] = 8'b0;
    XRAM[60848] = 8'b0;
    XRAM[60849] = 8'b0;
    XRAM[60850] = 8'b0;
    XRAM[60851] = 8'b0;
    XRAM[60852] = 8'b0;
    XRAM[60853] = 8'b0;
    XRAM[60854] = 8'b0;
    XRAM[60855] = 8'b0;
    XRAM[60856] = 8'b0;
    XRAM[60857] = 8'b0;
    XRAM[60858] = 8'b0;
    XRAM[60859] = 8'b0;
    XRAM[60860] = 8'b0;
    XRAM[60861] = 8'b0;
    XRAM[60862] = 8'b0;
    XRAM[60863] = 8'b0;
    XRAM[60864] = 8'b0;
    XRAM[60865] = 8'b0;
    XRAM[60866] = 8'b0;
    XRAM[60867] = 8'b0;
    XRAM[60868] = 8'b0;
    XRAM[60869] = 8'b0;
    XRAM[60870] = 8'b0;
    XRAM[60871] = 8'b0;
    XRAM[60872] = 8'b0;
    XRAM[60873] = 8'b0;
    XRAM[60874] = 8'b0;
    XRAM[60875] = 8'b0;
    XRAM[60876] = 8'b0;
    XRAM[60877] = 8'b0;
    XRAM[60878] = 8'b0;
    XRAM[60879] = 8'b0;
    XRAM[60880] = 8'b0;
    XRAM[60881] = 8'b0;
    XRAM[60882] = 8'b0;
    XRAM[60883] = 8'b0;
    XRAM[60884] = 8'b0;
    XRAM[60885] = 8'b0;
    XRAM[60886] = 8'b0;
    XRAM[60887] = 8'b0;
    XRAM[60888] = 8'b0;
    XRAM[60889] = 8'b0;
    XRAM[60890] = 8'b0;
    XRAM[60891] = 8'b0;
    XRAM[60892] = 8'b0;
    XRAM[60893] = 8'b0;
    XRAM[60894] = 8'b0;
    XRAM[60895] = 8'b0;
    XRAM[60896] = 8'b0;
    XRAM[60897] = 8'b0;
    XRAM[60898] = 8'b0;
    XRAM[60899] = 8'b0;
    XRAM[60900] = 8'b0;
    XRAM[60901] = 8'b0;
    XRAM[60902] = 8'b0;
    XRAM[60903] = 8'b0;
    XRAM[60904] = 8'b0;
    XRAM[60905] = 8'b0;
    XRAM[60906] = 8'b0;
    XRAM[60907] = 8'b0;
    XRAM[60908] = 8'b0;
    XRAM[60909] = 8'b0;
    XRAM[60910] = 8'b0;
    XRAM[60911] = 8'b0;
    XRAM[60912] = 8'b0;
    XRAM[60913] = 8'b0;
    XRAM[60914] = 8'b0;
    XRAM[60915] = 8'b0;
    XRAM[60916] = 8'b0;
    XRAM[60917] = 8'b0;
    XRAM[60918] = 8'b0;
    XRAM[60919] = 8'b0;
    XRAM[60920] = 8'b0;
    XRAM[60921] = 8'b0;
    XRAM[60922] = 8'b0;
    XRAM[60923] = 8'b0;
    XRAM[60924] = 8'b0;
    XRAM[60925] = 8'b0;
    XRAM[60926] = 8'b0;
    XRAM[60927] = 8'b0;
    XRAM[60928] = 8'b0;
    XRAM[60929] = 8'b0;
    XRAM[60930] = 8'b0;
    XRAM[60931] = 8'b0;
    XRAM[60932] = 8'b0;
    XRAM[60933] = 8'b0;
    XRAM[60934] = 8'b0;
    XRAM[60935] = 8'b0;
    XRAM[60936] = 8'b0;
    XRAM[60937] = 8'b0;
    XRAM[60938] = 8'b0;
    XRAM[60939] = 8'b0;
    XRAM[60940] = 8'b0;
    XRAM[60941] = 8'b0;
    XRAM[60942] = 8'b0;
    XRAM[60943] = 8'b0;
    XRAM[60944] = 8'b0;
    XRAM[60945] = 8'b0;
    XRAM[60946] = 8'b0;
    XRAM[60947] = 8'b0;
    XRAM[60948] = 8'b0;
    XRAM[60949] = 8'b0;
    XRAM[60950] = 8'b0;
    XRAM[60951] = 8'b0;
    XRAM[60952] = 8'b0;
    XRAM[60953] = 8'b0;
    XRAM[60954] = 8'b0;
    XRAM[60955] = 8'b0;
    XRAM[60956] = 8'b0;
    XRAM[60957] = 8'b0;
    XRAM[60958] = 8'b0;
    XRAM[60959] = 8'b0;
    XRAM[60960] = 8'b0;
    XRAM[60961] = 8'b0;
    XRAM[60962] = 8'b0;
    XRAM[60963] = 8'b0;
    XRAM[60964] = 8'b0;
    XRAM[60965] = 8'b0;
    XRAM[60966] = 8'b0;
    XRAM[60967] = 8'b0;
    XRAM[60968] = 8'b0;
    XRAM[60969] = 8'b0;
    XRAM[60970] = 8'b0;
    XRAM[60971] = 8'b0;
    XRAM[60972] = 8'b0;
    XRAM[60973] = 8'b0;
    XRAM[60974] = 8'b0;
    XRAM[60975] = 8'b0;
    XRAM[60976] = 8'b0;
    XRAM[60977] = 8'b0;
    XRAM[60978] = 8'b0;
    XRAM[60979] = 8'b0;
    XRAM[60980] = 8'b0;
    XRAM[60981] = 8'b0;
    XRAM[60982] = 8'b0;
    XRAM[60983] = 8'b0;
    XRAM[60984] = 8'b0;
    XRAM[60985] = 8'b0;
    XRAM[60986] = 8'b0;
    XRAM[60987] = 8'b0;
    XRAM[60988] = 8'b0;
    XRAM[60989] = 8'b0;
    XRAM[60990] = 8'b0;
    XRAM[60991] = 8'b0;
    XRAM[60992] = 8'b0;
    XRAM[60993] = 8'b0;
    XRAM[60994] = 8'b0;
    XRAM[60995] = 8'b0;
    XRAM[60996] = 8'b0;
    XRAM[60997] = 8'b0;
    XRAM[60998] = 8'b0;
    XRAM[60999] = 8'b0;
    XRAM[61000] = 8'b0;
    XRAM[61001] = 8'b0;
    XRAM[61002] = 8'b0;
    XRAM[61003] = 8'b0;
    XRAM[61004] = 8'b0;
    XRAM[61005] = 8'b0;
    XRAM[61006] = 8'b0;
    XRAM[61007] = 8'b0;
    XRAM[61008] = 8'b0;
    XRAM[61009] = 8'b0;
    XRAM[61010] = 8'b0;
    XRAM[61011] = 8'b0;
    XRAM[61012] = 8'b0;
    XRAM[61013] = 8'b0;
    XRAM[61014] = 8'b0;
    XRAM[61015] = 8'b0;
    XRAM[61016] = 8'b0;
    XRAM[61017] = 8'b0;
    XRAM[61018] = 8'b0;
    XRAM[61019] = 8'b0;
    XRAM[61020] = 8'b0;
    XRAM[61021] = 8'b0;
    XRAM[61022] = 8'b0;
    XRAM[61023] = 8'b0;
    XRAM[61024] = 8'b0;
    XRAM[61025] = 8'b0;
    XRAM[61026] = 8'b0;
    XRAM[61027] = 8'b0;
    XRAM[61028] = 8'b0;
    XRAM[61029] = 8'b0;
    XRAM[61030] = 8'b0;
    XRAM[61031] = 8'b0;
    XRAM[61032] = 8'b0;
    XRAM[61033] = 8'b0;
    XRAM[61034] = 8'b0;
    XRAM[61035] = 8'b0;
    XRAM[61036] = 8'b0;
    XRAM[61037] = 8'b0;
    XRAM[61038] = 8'b0;
    XRAM[61039] = 8'b0;
    XRAM[61040] = 8'b0;
    XRAM[61041] = 8'b0;
    XRAM[61042] = 8'b0;
    XRAM[61043] = 8'b0;
    XRAM[61044] = 8'b0;
    XRAM[61045] = 8'b0;
    XRAM[61046] = 8'b0;
    XRAM[61047] = 8'b0;
    XRAM[61048] = 8'b0;
    XRAM[61049] = 8'b0;
    XRAM[61050] = 8'b0;
    XRAM[61051] = 8'b0;
    XRAM[61052] = 8'b0;
    XRAM[61053] = 8'b0;
    XRAM[61054] = 8'b0;
    XRAM[61055] = 8'b0;
    XRAM[61056] = 8'b0;
    XRAM[61057] = 8'b0;
    XRAM[61058] = 8'b0;
    XRAM[61059] = 8'b0;
    XRAM[61060] = 8'b0;
    XRAM[61061] = 8'b0;
    XRAM[61062] = 8'b0;
    XRAM[61063] = 8'b0;
    XRAM[61064] = 8'b0;
    XRAM[61065] = 8'b0;
    XRAM[61066] = 8'b0;
    XRAM[61067] = 8'b0;
    XRAM[61068] = 8'b0;
    XRAM[61069] = 8'b0;
    XRAM[61070] = 8'b0;
    XRAM[61071] = 8'b0;
    XRAM[61072] = 8'b0;
    XRAM[61073] = 8'b0;
    XRAM[61074] = 8'b0;
    XRAM[61075] = 8'b0;
    XRAM[61076] = 8'b0;
    XRAM[61077] = 8'b0;
    XRAM[61078] = 8'b0;
    XRAM[61079] = 8'b0;
    XRAM[61080] = 8'b0;
    XRAM[61081] = 8'b0;
    XRAM[61082] = 8'b0;
    XRAM[61083] = 8'b0;
    XRAM[61084] = 8'b0;
    XRAM[61085] = 8'b0;
    XRAM[61086] = 8'b0;
    XRAM[61087] = 8'b0;
    XRAM[61088] = 8'b0;
    XRAM[61089] = 8'b0;
    XRAM[61090] = 8'b0;
    XRAM[61091] = 8'b0;
    XRAM[61092] = 8'b0;
    XRAM[61093] = 8'b0;
    XRAM[61094] = 8'b0;
    XRAM[61095] = 8'b0;
    XRAM[61096] = 8'b0;
    XRAM[61097] = 8'b0;
    XRAM[61098] = 8'b0;
    XRAM[61099] = 8'b0;
    XRAM[61100] = 8'b0;
    XRAM[61101] = 8'b0;
    XRAM[61102] = 8'b0;
    XRAM[61103] = 8'b0;
    XRAM[61104] = 8'b0;
    XRAM[61105] = 8'b0;
    XRAM[61106] = 8'b0;
    XRAM[61107] = 8'b0;
    XRAM[61108] = 8'b0;
    XRAM[61109] = 8'b0;
    XRAM[61110] = 8'b0;
    XRAM[61111] = 8'b0;
    XRAM[61112] = 8'b0;
    XRAM[61113] = 8'b0;
    XRAM[61114] = 8'b0;
    XRAM[61115] = 8'b0;
    XRAM[61116] = 8'b0;
    XRAM[61117] = 8'b0;
    XRAM[61118] = 8'b0;
    XRAM[61119] = 8'b0;
    XRAM[61120] = 8'b0;
    XRAM[61121] = 8'b0;
    XRAM[61122] = 8'b0;
    XRAM[61123] = 8'b0;
    XRAM[61124] = 8'b0;
    XRAM[61125] = 8'b0;
    XRAM[61126] = 8'b0;
    XRAM[61127] = 8'b0;
    XRAM[61128] = 8'b0;
    XRAM[61129] = 8'b0;
    XRAM[61130] = 8'b0;
    XRAM[61131] = 8'b0;
    XRAM[61132] = 8'b0;
    XRAM[61133] = 8'b0;
    XRAM[61134] = 8'b0;
    XRAM[61135] = 8'b0;
    XRAM[61136] = 8'b0;
    XRAM[61137] = 8'b0;
    XRAM[61138] = 8'b0;
    XRAM[61139] = 8'b0;
    XRAM[61140] = 8'b0;
    XRAM[61141] = 8'b0;
    XRAM[61142] = 8'b0;
    XRAM[61143] = 8'b0;
    XRAM[61144] = 8'b0;
    XRAM[61145] = 8'b0;
    XRAM[61146] = 8'b0;
    XRAM[61147] = 8'b0;
    XRAM[61148] = 8'b0;
    XRAM[61149] = 8'b0;
    XRAM[61150] = 8'b0;
    XRAM[61151] = 8'b0;
    XRAM[61152] = 8'b0;
    XRAM[61153] = 8'b0;
    XRAM[61154] = 8'b0;
    XRAM[61155] = 8'b0;
    XRAM[61156] = 8'b0;
    XRAM[61157] = 8'b0;
    XRAM[61158] = 8'b0;
    XRAM[61159] = 8'b0;
    XRAM[61160] = 8'b0;
    XRAM[61161] = 8'b0;
    XRAM[61162] = 8'b0;
    XRAM[61163] = 8'b0;
    XRAM[61164] = 8'b0;
    XRAM[61165] = 8'b0;
    XRAM[61166] = 8'b0;
    XRAM[61167] = 8'b0;
    XRAM[61168] = 8'b0;
    XRAM[61169] = 8'b0;
    XRAM[61170] = 8'b0;
    XRAM[61171] = 8'b0;
    XRAM[61172] = 8'b0;
    XRAM[61173] = 8'b0;
    XRAM[61174] = 8'b0;
    XRAM[61175] = 8'b0;
    XRAM[61176] = 8'b0;
    XRAM[61177] = 8'b0;
    XRAM[61178] = 8'b0;
    XRAM[61179] = 8'b0;
    XRAM[61180] = 8'b0;
    XRAM[61181] = 8'b0;
    XRAM[61182] = 8'b0;
    XRAM[61183] = 8'b0;
    XRAM[61184] = 8'b0;
    XRAM[61185] = 8'b0;
    XRAM[61186] = 8'b0;
    XRAM[61187] = 8'b0;
    XRAM[61188] = 8'b0;
    XRAM[61189] = 8'b0;
    XRAM[61190] = 8'b0;
    XRAM[61191] = 8'b0;
    XRAM[61192] = 8'b0;
    XRAM[61193] = 8'b0;
    XRAM[61194] = 8'b0;
    XRAM[61195] = 8'b0;
    XRAM[61196] = 8'b0;
    XRAM[61197] = 8'b0;
    XRAM[61198] = 8'b0;
    XRAM[61199] = 8'b0;
    XRAM[61200] = 8'b0;
    XRAM[61201] = 8'b0;
    XRAM[61202] = 8'b0;
    XRAM[61203] = 8'b0;
    XRAM[61204] = 8'b0;
    XRAM[61205] = 8'b0;
    XRAM[61206] = 8'b0;
    XRAM[61207] = 8'b0;
    XRAM[61208] = 8'b0;
    XRAM[61209] = 8'b0;
    XRAM[61210] = 8'b0;
    XRAM[61211] = 8'b0;
    XRAM[61212] = 8'b0;
    XRAM[61213] = 8'b0;
    XRAM[61214] = 8'b0;
    XRAM[61215] = 8'b0;
    XRAM[61216] = 8'b0;
    XRAM[61217] = 8'b0;
    XRAM[61218] = 8'b0;
    XRAM[61219] = 8'b0;
    XRAM[61220] = 8'b0;
    XRAM[61221] = 8'b0;
    XRAM[61222] = 8'b0;
    XRAM[61223] = 8'b0;
    XRAM[61224] = 8'b0;
    XRAM[61225] = 8'b0;
    XRAM[61226] = 8'b0;
    XRAM[61227] = 8'b0;
    XRAM[61228] = 8'b0;
    XRAM[61229] = 8'b0;
    XRAM[61230] = 8'b0;
    XRAM[61231] = 8'b0;
    XRAM[61232] = 8'b0;
    XRAM[61233] = 8'b0;
    XRAM[61234] = 8'b0;
    XRAM[61235] = 8'b0;
    XRAM[61236] = 8'b0;
    XRAM[61237] = 8'b0;
    XRAM[61238] = 8'b0;
    XRAM[61239] = 8'b0;
    XRAM[61240] = 8'b0;
    XRAM[61241] = 8'b0;
    XRAM[61242] = 8'b0;
    XRAM[61243] = 8'b0;
    XRAM[61244] = 8'b0;
    XRAM[61245] = 8'b0;
    XRAM[61246] = 8'b0;
    XRAM[61247] = 8'b0;
    XRAM[61248] = 8'b0;
    XRAM[61249] = 8'b0;
    XRAM[61250] = 8'b0;
    XRAM[61251] = 8'b0;
    XRAM[61252] = 8'b0;
    XRAM[61253] = 8'b0;
    XRAM[61254] = 8'b0;
    XRAM[61255] = 8'b0;
    XRAM[61256] = 8'b0;
    XRAM[61257] = 8'b0;
    XRAM[61258] = 8'b0;
    XRAM[61259] = 8'b0;
    XRAM[61260] = 8'b0;
    XRAM[61261] = 8'b0;
    XRAM[61262] = 8'b0;
    XRAM[61263] = 8'b0;
    XRAM[61264] = 8'b0;
    XRAM[61265] = 8'b0;
    XRAM[61266] = 8'b0;
    XRAM[61267] = 8'b0;
    XRAM[61268] = 8'b0;
    XRAM[61269] = 8'b0;
    XRAM[61270] = 8'b0;
    XRAM[61271] = 8'b0;
    XRAM[61272] = 8'b0;
    XRAM[61273] = 8'b0;
    XRAM[61274] = 8'b0;
    XRAM[61275] = 8'b0;
    XRAM[61276] = 8'b0;
    XRAM[61277] = 8'b0;
    XRAM[61278] = 8'b0;
    XRAM[61279] = 8'b0;
    XRAM[61280] = 8'b0;
    XRAM[61281] = 8'b0;
    XRAM[61282] = 8'b0;
    XRAM[61283] = 8'b0;
    XRAM[61284] = 8'b0;
    XRAM[61285] = 8'b0;
    XRAM[61286] = 8'b0;
    XRAM[61287] = 8'b0;
    XRAM[61288] = 8'b0;
    XRAM[61289] = 8'b0;
    XRAM[61290] = 8'b0;
    XRAM[61291] = 8'b0;
    XRAM[61292] = 8'b0;
    XRAM[61293] = 8'b0;
    XRAM[61294] = 8'b0;
    XRAM[61295] = 8'b0;
    XRAM[61296] = 8'b0;
    XRAM[61297] = 8'b0;
    XRAM[61298] = 8'b0;
    XRAM[61299] = 8'b0;
    XRAM[61300] = 8'b0;
    XRAM[61301] = 8'b0;
    XRAM[61302] = 8'b0;
    XRAM[61303] = 8'b0;
    XRAM[61304] = 8'b0;
    XRAM[61305] = 8'b0;
    XRAM[61306] = 8'b0;
    XRAM[61307] = 8'b0;
    XRAM[61308] = 8'b0;
    XRAM[61309] = 8'b0;
    XRAM[61310] = 8'b0;
    XRAM[61311] = 8'b0;
    XRAM[61312] = 8'b0;
    XRAM[61313] = 8'b0;
    XRAM[61314] = 8'b0;
    XRAM[61315] = 8'b0;
    XRAM[61316] = 8'b0;
    XRAM[61317] = 8'b0;
    XRAM[61318] = 8'b0;
    XRAM[61319] = 8'b0;
    XRAM[61320] = 8'b0;
    XRAM[61321] = 8'b0;
    XRAM[61322] = 8'b0;
    XRAM[61323] = 8'b0;
    XRAM[61324] = 8'b0;
    XRAM[61325] = 8'b0;
    XRAM[61326] = 8'b0;
    XRAM[61327] = 8'b0;
    XRAM[61328] = 8'b0;
    XRAM[61329] = 8'b0;
    XRAM[61330] = 8'b0;
    XRAM[61331] = 8'b0;
    XRAM[61332] = 8'b0;
    XRAM[61333] = 8'b0;
    XRAM[61334] = 8'b0;
    XRAM[61335] = 8'b0;
    XRAM[61336] = 8'b0;
    XRAM[61337] = 8'b0;
    XRAM[61338] = 8'b0;
    XRAM[61339] = 8'b0;
    XRAM[61340] = 8'b0;
    XRAM[61341] = 8'b0;
    XRAM[61342] = 8'b0;
    XRAM[61343] = 8'b0;
    XRAM[61344] = 8'b0;
    XRAM[61345] = 8'b0;
    XRAM[61346] = 8'b0;
    XRAM[61347] = 8'b0;
    XRAM[61348] = 8'b0;
    XRAM[61349] = 8'b0;
    XRAM[61350] = 8'b0;
    XRAM[61351] = 8'b0;
    XRAM[61352] = 8'b0;
    XRAM[61353] = 8'b0;
    XRAM[61354] = 8'b0;
    XRAM[61355] = 8'b0;
    XRAM[61356] = 8'b0;
    XRAM[61357] = 8'b0;
    XRAM[61358] = 8'b0;
    XRAM[61359] = 8'b0;
    XRAM[61360] = 8'b0;
    XRAM[61361] = 8'b0;
    XRAM[61362] = 8'b0;
    XRAM[61363] = 8'b0;
    XRAM[61364] = 8'b0;
    XRAM[61365] = 8'b0;
    XRAM[61366] = 8'b0;
    XRAM[61367] = 8'b0;
    XRAM[61368] = 8'b0;
    XRAM[61369] = 8'b0;
    XRAM[61370] = 8'b0;
    XRAM[61371] = 8'b0;
    XRAM[61372] = 8'b0;
    XRAM[61373] = 8'b0;
    XRAM[61374] = 8'b0;
    XRAM[61375] = 8'b0;
    XRAM[61376] = 8'b0;
    XRAM[61377] = 8'b0;
    XRAM[61378] = 8'b0;
    XRAM[61379] = 8'b0;
    XRAM[61380] = 8'b0;
    XRAM[61381] = 8'b0;
    XRAM[61382] = 8'b0;
    XRAM[61383] = 8'b0;
    XRAM[61384] = 8'b0;
    XRAM[61385] = 8'b0;
    XRAM[61386] = 8'b0;
    XRAM[61387] = 8'b0;
    XRAM[61388] = 8'b0;
    XRAM[61389] = 8'b0;
    XRAM[61390] = 8'b0;
    XRAM[61391] = 8'b0;
    XRAM[61392] = 8'b0;
    XRAM[61393] = 8'b0;
    XRAM[61394] = 8'b0;
    XRAM[61395] = 8'b0;
    XRAM[61396] = 8'b0;
    XRAM[61397] = 8'b0;
    XRAM[61398] = 8'b0;
    XRAM[61399] = 8'b0;
    XRAM[61400] = 8'b0;
    XRAM[61401] = 8'b0;
    XRAM[61402] = 8'b0;
    XRAM[61403] = 8'b0;
    XRAM[61404] = 8'b0;
    XRAM[61405] = 8'b0;
    XRAM[61406] = 8'b0;
    XRAM[61407] = 8'b0;
    XRAM[61408] = 8'b0;
    XRAM[61409] = 8'b0;
    XRAM[61410] = 8'b0;
    XRAM[61411] = 8'b0;
    XRAM[61412] = 8'b0;
    XRAM[61413] = 8'b0;
    XRAM[61414] = 8'b0;
    XRAM[61415] = 8'b0;
    XRAM[61416] = 8'b0;
    XRAM[61417] = 8'b0;
    XRAM[61418] = 8'b0;
    XRAM[61419] = 8'b0;
    XRAM[61420] = 8'b0;
    XRAM[61421] = 8'b0;
    XRAM[61422] = 8'b0;
    XRAM[61423] = 8'b0;
    XRAM[61424] = 8'b0;
    XRAM[61425] = 8'b0;
    XRAM[61426] = 8'b0;
    XRAM[61427] = 8'b0;
    XRAM[61428] = 8'b0;
    XRAM[61429] = 8'b0;
    XRAM[61430] = 8'b0;
    XRAM[61431] = 8'b0;
    XRAM[61432] = 8'b0;
    XRAM[61433] = 8'b0;
    XRAM[61434] = 8'b0;
    XRAM[61435] = 8'b0;
    XRAM[61436] = 8'b0;
    XRAM[61437] = 8'b0;
    XRAM[61438] = 8'b0;
    XRAM[61439] = 8'b0;
    XRAM[61440] = 8'b0;
    XRAM[61441] = 8'b0;
    XRAM[61442] = 8'b0;
    XRAM[61443] = 8'b0;
    XRAM[61444] = 8'b0;
    XRAM[61445] = 8'b0;
    XRAM[61446] = 8'b0;
    XRAM[61447] = 8'b0;
    XRAM[61448] = 8'b0;
    XRAM[61449] = 8'b0;
    XRAM[61450] = 8'b0;
    XRAM[61451] = 8'b0;
    XRAM[61452] = 8'b0;
    XRAM[61453] = 8'b0;
    XRAM[61454] = 8'b0;
    XRAM[61455] = 8'b0;
    XRAM[61456] = 8'b0;
    XRAM[61457] = 8'b0;
    XRAM[61458] = 8'b0;
    XRAM[61459] = 8'b0;
    XRAM[61460] = 8'b0;
    XRAM[61461] = 8'b0;
    XRAM[61462] = 8'b0;
    XRAM[61463] = 8'b0;
    XRAM[61464] = 8'b0;
    XRAM[61465] = 8'b0;
    XRAM[61466] = 8'b0;
    XRAM[61467] = 8'b0;
    XRAM[61468] = 8'b0;
    XRAM[61469] = 8'b0;
    XRAM[61470] = 8'b0;
    XRAM[61471] = 8'b0;
    XRAM[61472] = 8'b0;
    XRAM[61473] = 8'b0;
    XRAM[61474] = 8'b0;
    XRAM[61475] = 8'b0;
    XRAM[61476] = 8'b0;
    XRAM[61477] = 8'b0;
    XRAM[61478] = 8'b0;
    XRAM[61479] = 8'b0;
    XRAM[61480] = 8'b0;
    XRAM[61481] = 8'b0;
    XRAM[61482] = 8'b0;
    XRAM[61483] = 8'b0;
    XRAM[61484] = 8'b0;
    XRAM[61485] = 8'b0;
    XRAM[61486] = 8'b0;
    XRAM[61487] = 8'b0;
    XRAM[61488] = 8'b0;
    XRAM[61489] = 8'b0;
    XRAM[61490] = 8'b0;
    XRAM[61491] = 8'b0;
    XRAM[61492] = 8'b0;
    XRAM[61493] = 8'b0;
    XRAM[61494] = 8'b0;
    XRAM[61495] = 8'b0;
    XRAM[61496] = 8'b0;
    XRAM[61497] = 8'b0;
    XRAM[61498] = 8'b0;
    XRAM[61499] = 8'b0;
    XRAM[61500] = 8'b0;
    XRAM[61501] = 8'b0;
    XRAM[61502] = 8'b0;
    XRAM[61503] = 8'b0;
    XRAM[61504] = 8'b0;
    XRAM[61505] = 8'b0;
    XRAM[61506] = 8'b0;
    XRAM[61507] = 8'b0;
    XRAM[61508] = 8'b0;
    XRAM[61509] = 8'b0;
    XRAM[61510] = 8'b0;
    XRAM[61511] = 8'b0;
    XRAM[61512] = 8'b0;
    XRAM[61513] = 8'b0;
    XRAM[61514] = 8'b0;
    XRAM[61515] = 8'b0;
    XRAM[61516] = 8'b0;
    XRAM[61517] = 8'b0;
    XRAM[61518] = 8'b0;
    XRAM[61519] = 8'b0;
    XRAM[61520] = 8'b0;
    XRAM[61521] = 8'b0;
    XRAM[61522] = 8'b0;
    XRAM[61523] = 8'b0;
    XRAM[61524] = 8'b0;
    XRAM[61525] = 8'b0;
    XRAM[61526] = 8'b0;
    XRAM[61527] = 8'b0;
    XRAM[61528] = 8'b0;
    XRAM[61529] = 8'b0;
    XRAM[61530] = 8'b0;
    XRAM[61531] = 8'b0;
    XRAM[61532] = 8'b0;
    XRAM[61533] = 8'b0;
    XRAM[61534] = 8'b0;
    XRAM[61535] = 8'b0;
    XRAM[61536] = 8'b0;
    XRAM[61537] = 8'b0;
    XRAM[61538] = 8'b0;
    XRAM[61539] = 8'b0;
    XRAM[61540] = 8'b0;
    XRAM[61541] = 8'b0;
    XRAM[61542] = 8'b0;
    XRAM[61543] = 8'b0;
    XRAM[61544] = 8'b0;
    XRAM[61545] = 8'b0;
    XRAM[61546] = 8'b0;
    XRAM[61547] = 8'b0;
    XRAM[61548] = 8'b0;
    XRAM[61549] = 8'b0;
    XRAM[61550] = 8'b0;
    XRAM[61551] = 8'b0;
    XRAM[61552] = 8'b0;
    XRAM[61553] = 8'b0;
    XRAM[61554] = 8'b0;
    XRAM[61555] = 8'b0;
    XRAM[61556] = 8'b0;
    XRAM[61557] = 8'b0;
    XRAM[61558] = 8'b0;
    XRAM[61559] = 8'b0;
    XRAM[61560] = 8'b0;
    XRAM[61561] = 8'b0;
    XRAM[61562] = 8'b0;
    XRAM[61563] = 8'b0;
    XRAM[61564] = 8'b0;
    XRAM[61565] = 8'b0;
    XRAM[61566] = 8'b0;
    XRAM[61567] = 8'b0;
    XRAM[61568] = 8'b0;
    XRAM[61569] = 8'b0;
    XRAM[61570] = 8'b0;
    XRAM[61571] = 8'b0;
    XRAM[61572] = 8'b0;
    XRAM[61573] = 8'b0;
    XRAM[61574] = 8'b0;
    XRAM[61575] = 8'b0;
    XRAM[61576] = 8'b0;
    XRAM[61577] = 8'b0;
    XRAM[61578] = 8'b0;
    XRAM[61579] = 8'b0;
    XRAM[61580] = 8'b0;
    XRAM[61581] = 8'b0;
    XRAM[61582] = 8'b0;
    XRAM[61583] = 8'b0;
    XRAM[61584] = 8'b0;
    XRAM[61585] = 8'b0;
    XRAM[61586] = 8'b0;
    XRAM[61587] = 8'b0;
    XRAM[61588] = 8'b0;
    XRAM[61589] = 8'b0;
    XRAM[61590] = 8'b0;
    XRAM[61591] = 8'b0;
    XRAM[61592] = 8'b0;
    XRAM[61593] = 8'b0;
    XRAM[61594] = 8'b0;
    XRAM[61595] = 8'b0;
    XRAM[61596] = 8'b0;
    XRAM[61597] = 8'b0;
    XRAM[61598] = 8'b0;
    XRAM[61599] = 8'b0;
    XRAM[61600] = 8'b0;
    XRAM[61601] = 8'b0;
    XRAM[61602] = 8'b0;
    XRAM[61603] = 8'b0;
    XRAM[61604] = 8'b0;
    XRAM[61605] = 8'b0;
    XRAM[61606] = 8'b0;
    XRAM[61607] = 8'b0;
    XRAM[61608] = 8'b0;
    XRAM[61609] = 8'b0;
    XRAM[61610] = 8'b0;
    XRAM[61611] = 8'b0;
    XRAM[61612] = 8'b0;
    XRAM[61613] = 8'b0;
    XRAM[61614] = 8'b0;
    XRAM[61615] = 8'b0;
    XRAM[61616] = 8'b0;
    XRAM[61617] = 8'b0;
    XRAM[61618] = 8'b0;
    XRAM[61619] = 8'b0;
    XRAM[61620] = 8'b0;
    XRAM[61621] = 8'b0;
    XRAM[61622] = 8'b0;
    XRAM[61623] = 8'b0;
    XRAM[61624] = 8'b0;
    XRAM[61625] = 8'b0;
    XRAM[61626] = 8'b0;
    XRAM[61627] = 8'b0;
    XRAM[61628] = 8'b0;
    XRAM[61629] = 8'b0;
    XRAM[61630] = 8'b0;
    XRAM[61631] = 8'b0;
    XRAM[61632] = 8'b0;
    XRAM[61633] = 8'b0;
    XRAM[61634] = 8'b0;
    XRAM[61635] = 8'b0;
    XRAM[61636] = 8'b0;
    XRAM[61637] = 8'b0;
    XRAM[61638] = 8'b0;
    XRAM[61639] = 8'b0;
    XRAM[61640] = 8'b0;
    XRAM[61641] = 8'b0;
    XRAM[61642] = 8'b0;
    XRAM[61643] = 8'b0;
    XRAM[61644] = 8'b0;
    XRAM[61645] = 8'b0;
    XRAM[61646] = 8'b0;
    XRAM[61647] = 8'b0;
    XRAM[61648] = 8'b0;
    XRAM[61649] = 8'b0;
    XRAM[61650] = 8'b0;
    XRAM[61651] = 8'b0;
    XRAM[61652] = 8'b0;
    XRAM[61653] = 8'b0;
    XRAM[61654] = 8'b0;
    XRAM[61655] = 8'b0;
    XRAM[61656] = 8'b0;
    XRAM[61657] = 8'b0;
    XRAM[61658] = 8'b0;
    XRAM[61659] = 8'b0;
    XRAM[61660] = 8'b0;
    XRAM[61661] = 8'b0;
    XRAM[61662] = 8'b0;
    XRAM[61663] = 8'b0;
    XRAM[61664] = 8'b0;
    XRAM[61665] = 8'b0;
    XRAM[61666] = 8'b0;
    XRAM[61667] = 8'b0;
    XRAM[61668] = 8'b0;
    XRAM[61669] = 8'b0;
    XRAM[61670] = 8'b0;
    XRAM[61671] = 8'b0;
    XRAM[61672] = 8'b0;
    XRAM[61673] = 8'b0;
    XRAM[61674] = 8'b0;
    XRAM[61675] = 8'b0;
    XRAM[61676] = 8'b0;
    XRAM[61677] = 8'b0;
    XRAM[61678] = 8'b0;
    XRAM[61679] = 8'b0;
    XRAM[61680] = 8'b0;
    XRAM[61681] = 8'b0;
    XRAM[61682] = 8'b0;
    XRAM[61683] = 8'b0;
    XRAM[61684] = 8'b0;
    XRAM[61685] = 8'b0;
    XRAM[61686] = 8'b0;
    XRAM[61687] = 8'b0;
    XRAM[61688] = 8'b0;
    XRAM[61689] = 8'b0;
    XRAM[61690] = 8'b0;
    XRAM[61691] = 8'b0;
    XRAM[61692] = 8'b0;
    XRAM[61693] = 8'b0;
    XRAM[61694] = 8'b0;
    XRAM[61695] = 8'b0;
    XRAM[61696] = 8'b0;
    XRAM[61697] = 8'b0;
    XRAM[61698] = 8'b0;
    XRAM[61699] = 8'b0;
    XRAM[61700] = 8'b0;
    XRAM[61701] = 8'b0;
    XRAM[61702] = 8'b0;
    XRAM[61703] = 8'b0;
    XRAM[61704] = 8'b0;
    XRAM[61705] = 8'b0;
    XRAM[61706] = 8'b0;
    XRAM[61707] = 8'b0;
    XRAM[61708] = 8'b0;
    XRAM[61709] = 8'b0;
    XRAM[61710] = 8'b0;
    XRAM[61711] = 8'b0;
    XRAM[61712] = 8'b0;
    XRAM[61713] = 8'b0;
    XRAM[61714] = 8'b0;
    XRAM[61715] = 8'b0;
    XRAM[61716] = 8'b0;
    XRAM[61717] = 8'b0;
    XRAM[61718] = 8'b0;
    XRAM[61719] = 8'b0;
    XRAM[61720] = 8'b0;
    XRAM[61721] = 8'b0;
    XRAM[61722] = 8'b0;
    XRAM[61723] = 8'b0;
    XRAM[61724] = 8'b0;
    XRAM[61725] = 8'b0;
    XRAM[61726] = 8'b0;
    XRAM[61727] = 8'b0;
    XRAM[61728] = 8'b0;
    XRAM[61729] = 8'b0;
    XRAM[61730] = 8'b0;
    XRAM[61731] = 8'b0;
    XRAM[61732] = 8'b0;
    XRAM[61733] = 8'b0;
    XRAM[61734] = 8'b0;
    XRAM[61735] = 8'b0;
    XRAM[61736] = 8'b0;
    XRAM[61737] = 8'b0;
    XRAM[61738] = 8'b0;
    XRAM[61739] = 8'b0;
    XRAM[61740] = 8'b0;
    XRAM[61741] = 8'b0;
    XRAM[61742] = 8'b0;
    XRAM[61743] = 8'b0;
    XRAM[61744] = 8'b0;
    XRAM[61745] = 8'b0;
    XRAM[61746] = 8'b0;
    XRAM[61747] = 8'b0;
    XRAM[61748] = 8'b0;
    XRAM[61749] = 8'b0;
    XRAM[61750] = 8'b0;
    XRAM[61751] = 8'b0;
    XRAM[61752] = 8'b0;
    XRAM[61753] = 8'b0;
    XRAM[61754] = 8'b0;
    XRAM[61755] = 8'b0;
    XRAM[61756] = 8'b0;
    XRAM[61757] = 8'b0;
    XRAM[61758] = 8'b0;
    XRAM[61759] = 8'b0;
    XRAM[61760] = 8'b0;
    XRAM[61761] = 8'b0;
    XRAM[61762] = 8'b0;
    XRAM[61763] = 8'b0;
    XRAM[61764] = 8'b0;
    XRAM[61765] = 8'b0;
    XRAM[61766] = 8'b0;
    XRAM[61767] = 8'b0;
    XRAM[61768] = 8'b0;
    XRAM[61769] = 8'b0;
    XRAM[61770] = 8'b0;
    XRAM[61771] = 8'b0;
    XRAM[61772] = 8'b0;
    XRAM[61773] = 8'b0;
    XRAM[61774] = 8'b0;
    XRAM[61775] = 8'b0;
    XRAM[61776] = 8'b0;
    XRAM[61777] = 8'b0;
    XRAM[61778] = 8'b0;
    XRAM[61779] = 8'b0;
    XRAM[61780] = 8'b0;
    XRAM[61781] = 8'b0;
    XRAM[61782] = 8'b0;
    XRAM[61783] = 8'b0;
    XRAM[61784] = 8'b0;
    XRAM[61785] = 8'b0;
    XRAM[61786] = 8'b0;
    XRAM[61787] = 8'b0;
    XRAM[61788] = 8'b0;
    XRAM[61789] = 8'b0;
    XRAM[61790] = 8'b0;
    XRAM[61791] = 8'b0;
    XRAM[61792] = 8'b0;
    XRAM[61793] = 8'b0;
    XRAM[61794] = 8'b0;
    XRAM[61795] = 8'b0;
    XRAM[61796] = 8'b0;
    XRAM[61797] = 8'b0;
    XRAM[61798] = 8'b0;
    XRAM[61799] = 8'b0;
    XRAM[61800] = 8'b0;
    XRAM[61801] = 8'b0;
    XRAM[61802] = 8'b0;
    XRAM[61803] = 8'b0;
    XRAM[61804] = 8'b0;
    XRAM[61805] = 8'b0;
    XRAM[61806] = 8'b0;
    XRAM[61807] = 8'b0;
    XRAM[61808] = 8'b0;
    XRAM[61809] = 8'b0;
    XRAM[61810] = 8'b0;
    XRAM[61811] = 8'b0;
    XRAM[61812] = 8'b0;
    XRAM[61813] = 8'b0;
    XRAM[61814] = 8'b0;
    XRAM[61815] = 8'b0;
    XRAM[61816] = 8'b0;
    XRAM[61817] = 8'b0;
    XRAM[61818] = 8'b0;
    XRAM[61819] = 8'b0;
    XRAM[61820] = 8'b0;
    XRAM[61821] = 8'b0;
    XRAM[61822] = 8'b0;
    XRAM[61823] = 8'b0;
    XRAM[61824] = 8'b0;
    XRAM[61825] = 8'b0;
    XRAM[61826] = 8'b0;
    XRAM[61827] = 8'b0;
    XRAM[61828] = 8'b0;
    XRAM[61829] = 8'b0;
    XRAM[61830] = 8'b0;
    XRAM[61831] = 8'b0;
    XRAM[61832] = 8'b0;
    XRAM[61833] = 8'b0;
    XRAM[61834] = 8'b0;
    XRAM[61835] = 8'b0;
    XRAM[61836] = 8'b0;
    XRAM[61837] = 8'b0;
    XRAM[61838] = 8'b0;
    XRAM[61839] = 8'b0;
    XRAM[61840] = 8'b0;
    XRAM[61841] = 8'b0;
    XRAM[61842] = 8'b0;
    XRAM[61843] = 8'b0;
    XRAM[61844] = 8'b0;
    XRAM[61845] = 8'b0;
    XRAM[61846] = 8'b0;
    XRAM[61847] = 8'b0;
    XRAM[61848] = 8'b0;
    XRAM[61849] = 8'b0;
    XRAM[61850] = 8'b0;
    XRAM[61851] = 8'b0;
    XRAM[61852] = 8'b0;
    XRAM[61853] = 8'b0;
    XRAM[61854] = 8'b0;
    XRAM[61855] = 8'b0;
    XRAM[61856] = 8'b0;
    XRAM[61857] = 8'b0;
    XRAM[61858] = 8'b0;
    XRAM[61859] = 8'b0;
    XRAM[61860] = 8'b0;
    XRAM[61861] = 8'b0;
    XRAM[61862] = 8'b0;
    XRAM[61863] = 8'b0;
    XRAM[61864] = 8'b0;
    XRAM[61865] = 8'b0;
    XRAM[61866] = 8'b0;
    XRAM[61867] = 8'b0;
    XRAM[61868] = 8'b0;
    XRAM[61869] = 8'b0;
    XRAM[61870] = 8'b0;
    XRAM[61871] = 8'b0;
    XRAM[61872] = 8'b0;
    XRAM[61873] = 8'b0;
    XRAM[61874] = 8'b0;
    XRAM[61875] = 8'b0;
    XRAM[61876] = 8'b0;
    XRAM[61877] = 8'b0;
    XRAM[61878] = 8'b0;
    XRAM[61879] = 8'b0;
    XRAM[61880] = 8'b0;
    XRAM[61881] = 8'b0;
    XRAM[61882] = 8'b0;
    XRAM[61883] = 8'b0;
    XRAM[61884] = 8'b0;
    XRAM[61885] = 8'b0;
    XRAM[61886] = 8'b0;
    XRAM[61887] = 8'b0;
    XRAM[61888] = 8'b0;
    XRAM[61889] = 8'b0;
    XRAM[61890] = 8'b0;
    XRAM[61891] = 8'b0;
    XRAM[61892] = 8'b0;
    XRAM[61893] = 8'b0;
    XRAM[61894] = 8'b0;
    XRAM[61895] = 8'b0;
    XRAM[61896] = 8'b0;
    XRAM[61897] = 8'b0;
    XRAM[61898] = 8'b0;
    XRAM[61899] = 8'b0;
    XRAM[61900] = 8'b0;
    XRAM[61901] = 8'b0;
    XRAM[61902] = 8'b0;
    XRAM[61903] = 8'b0;
    XRAM[61904] = 8'b0;
    XRAM[61905] = 8'b0;
    XRAM[61906] = 8'b0;
    XRAM[61907] = 8'b0;
    XRAM[61908] = 8'b0;
    XRAM[61909] = 8'b0;
    XRAM[61910] = 8'b0;
    XRAM[61911] = 8'b0;
    XRAM[61912] = 8'b0;
    XRAM[61913] = 8'b0;
    XRAM[61914] = 8'b0;
    XRAM[61915] = 8'b0;
    XRAM[61916] = 8'b0;
    XRAM[61917] = 8'b0;
    XRAM[61918] = 8'b0;
    XRAM[61919] = 8'b0;
    XRAM[61920] = 8'b0;
    XRAM[61921] = 8'b0;
    XRAM[61922] = 8'b0;
    XRAM[61923] = 8'b0;
    XRAM[61924] = 8'b0;
    XRAM[61925] = 8'b0;
    XRAM[61926] = 8'b0;
    XRAM[61927] = 8'b0;
    XRAM[61928] = 8'b0;
    XRAM[61929] = 8'b0;
    XRAM[61930] = 8'b0;
    XRAM[61931] = 8'b0;
    XRAM[61932] = 8'b0;
    XRAM[61933] = 8'b0;
    XRAM[61934] = 8'b0;
    XRAM[61935] = 8'b0;
    XRAM[61936] = 8'b0;
    XRAM[61937] = 8'b0;
    XRAM[61938] = 8'b0;
    XRAM[61939] = 8'b0;
    XRAM[61940] = 8'b0;
    XRAM[61941] = 8'b0;
    XRAM[61942] = 8'b0;
    XRAM[61943] = 8'b0;
    XRAM[61944] = 8'b0;
    XRAM[61945] = 8'b0;
    XRAM[61946] = 8'b0;
    XRAM[61947] = 8'b0;
    XRAM[61948] = 8'b0;
    XRAM[61949] = 8'b0;
    XRAM[61950] = 8'b0;
    XRAM[61951] = 8'b0;
    XRAM[61952] = 8'b0;
    XRAM[61953] = 8'b0;
    XRAM[61954] = 8'b0;
    XRAM[61955] = 8'b0;
    XRAM[61956] = 8'b0;
    XRAM[61957] = 8'b0;
    XRAM[61958] = 8'b0;
    XRAM[61959] = 8'b0;
    XRAM[61960] = 8'b0;
    XRAM[61961] = 8'b0;
    XRAM[61962] = 8'b0;
    XRAM[61963] = 8'b0;
    XRAM[61964] = 8'b0;
    XRAM[61965] = 8'b0;
    XRAM[61966] = 8'b0;
    XRAM[61967] = 8'b0;
    XRAM[61968] = 8'b0;
    XRAM[61969] = 8'b0;
    XRAM[61970] = 8'b0;
    XRAM[61971] = 8'b0;
    XRAM[61972] = 8'b0;
    XRAM[61973] = 8'b0;
    XRAM[61974] = 8'b0;
    XRAM[61975] = 8'b0;
    XRAM[61976] = 8'b0;
    XRAM[61977] = 8'b0;
    XRAM[61978] = 8'b0;
    XRAM[61979] = 8'b0;
    XRAM[61980] = 8'b0;
    XRAM[61981] = 8'b0;
    XRAM[61982] = 8'b0;
    XRAM[61983] = 8'b0;
    XRAM[61984] = 8'b0;
    XRAM[61985] = 8'b0;
    XRAM[61986] = 8'b0;
    XRAM[61987] = 8'b0;
    XRAM[61988] = 8'b0;
    XRAM[61989] = 8'b0;
    XRAM[61990] = 8'b0;
    XRAM[61991] = 8'b0;
    XRAM[61992] = 8'b0;
    XRAM[61993] = 8'b0;
    XRAM[61994] = 8'b0;
    XRAM[61995] = 8'b0;
    XRAM[61996] = 8'b0;
    XRAM[61997] = 8'b0;
    XRAM[61998] = 8'b0;
    XRAM[61999] = 8'b0;
    XRAM[62000] = 8'b0;
    XRAM[62001] = 8'b0;
    XRAM[62002] = 8'b0;
    XRAM[62003] = 8'b0;
    XRAM[62004] = 8'b0;
    XRAM[62005] = 8'b0;
    XRAM[62006] = 8'b0;
    XRAM[62007] = 8'b0;
    XRAM[62008] = 8'b0;
    XRAM[62009] = 8'b0;
    XRAM[62010] = 8'b0;
    XRAM[62011] = 8'b0;
    XRAM[62012] = 8'b0;
    XRAM[62013] = 8'b0;
    XRAM[62014] = 8'b0;
    XRAM[62015] = 8'b0;
    XRAM[62016] = 8'b0;
    XRAM[62017] = 8'b0;
    XRAM[62018] = 8'b0;
    XRAM[62019] = 8'b0;
    XRAM[62020] = 8'b0;
    XRAM[62021] = 8'b0;
    XRAM[62022] = 8'b0;
    XRAM[62023] = 8'b0;
    XRAM[62024] = 8'b0;
    XRAM[62025] = 8'b0;
    XRAM[62026] = 8'b0;
    XRAM[62027] = 8'b0;
    XRAM[62028] = 8'b0;
    XRAM[62029] = 8'b0;
    XRAM[62030] = 8'b0;
    XRAM[62031] = 8'b0;
    XRAM[62032] = 8'b0;
    XRAM[62033] = 8'b0;
    XRAM[62034] = 8'b0;
    XRAM[62035] = 8'b0;
    XRAM[62036] = 8'b0;
    XRAM[62037] = 8'b0;
    XRAM[62038] = 8'b0;
    XRAM[62039] = 8'b0;
    XRAM[62040] = 8'b0;
    XRAM[62041] = 8'b0;
    XRAM[62042] = 8'b0;
    XRAM[62043] = 8'b0;
    XRAM[62044] = 8'b0;
    XRAM[62045] = 8'b0;
    XRAM[62046] = 8'b0;
    XRAM[62047] = 8'b0;
    XRAM[62048] = 8'b0;
    XRAM[62049] = 8'b0;
    XRAM[62050] = 8'b0;
    XRAM[62051] = 8'b0;
    XRAM[62052] = 8'b0;
    XRAM[62053] = 8'b0;
    XRAM[62054] = 8'b0;
    XRAM[62055] = 8'b0;
    XRAM[62056] = 8'b0;
    XRAM[62057] = 8'b0;
    XRAM[62058] = 8'b0;
    XRAM[62059] = 8'b0;
    XRAM[62060] = 8'b0;
    XRAM[62061] = 8'b0;
    XRAM[62062] = 8'b0;
    XRAM[62063] = 8'b0;
    XRAM[62064] = 8'b0;
    XRAM[62065] = 8'b0;
    XRAM[62066] = 8'b0;
    XRAM[62067] = 8'b0;
    XRAM[62068] = 8'b0;
    XRAM[62069] = 8'b0;
    XRAM[62070] = 8'b0;
    XRAM[62071] = 8'b0;
    XRAM[62072] = 8'b0;
    XRAM[62073] = 8'b0;
    XRAM[62074] = 8'b0;
    XRAM[62075] = 8'b0;
    XRAM[62076] = 8'b0;
    XRAM[62077] = 8'b0;
    XRAM[62078] = 8'b0;
    XRAM[62079] = 8'b0;
    XRAM[62080] = 8'b0;
    XRAM[62081] = 8'b0;
    XRAM[62082] = 8'b0;
    XRAM[62083] = 8'b0;
    XRAM[62084] = 8'b0;
    XRAM[62085] = 8'b0;
    XRAM[62086] = 8'b0;
    XRAM[62087] = 8'b0;
    XRAM[62088] = 8'b0;
    XRAM[62089] = 8'b0;
    XRAM[62090] = 8'b0;
    XRAM[62091] = 8'b0;
    XRAM[62092] = 8'b0;
    XRAM[62093] = 8'b0;
    XRAM[62094] = 8'b0;
    XRAM[62095] = 8'b0;
    XRAM[62096] = 8'b0;
    XRAM[62097] = 8'b0;
    XRAM[62098] = 8'b0;
    XRAM[62099] = 8'b0;
    XRAM[62100] = 8'b0;
    XRAM[62101] = 8'b0;
    XRAM[62102] = 8'b0;
    XRAM[62103] = 8'b0;
    XRAM[62104] = 8'b0;
    XRAM[62105] = 8'b0;
    XRAM[62106] = 8'b0;
    XRAM[62107] = 8'b0;
    XRAM[62108] = 8'b0;
    XRAM[62109] = 8'b0;
    XRAM[62110] = 8'b0;
    XRAM[62111] = 8'b0;
    XRAM[62112] = 8'b0;
    XRAM[62113] = 8'b0;
    XRAM[62114] = 8'b0;
    XRAM[62115] = 8'b0;
    XRAM[62116] = 8'b0;
    XRAM[62117] = 8'b0;
    XRAM[62118] = 8'b0;
    XRAM[62119] = 8'b0;
    XRAM[62120] = 8'b0;
    XRAM[62121] = 8'b0;
    XRAM[62122] = 8'b0;
    XRAM[62123] = 8'b0;
    XRAM[62124] = 8'b0;
    XRAM[62125] = 8'b0;
    XRAM[62126] = 8'b0;
    XRAM[62127] = 8'b0;
    XRAM[62128] = 8'b0;
    XRAM[62129] = 8'b0;
    XRAM[62130] = 8'b0;
    XRAM[62131] = 8'b0;
    XRAM[62132] = 8'b0;
    XRAM[62133] = 8'b0;
    XRAM[62134] = 8'b0;
    XRAM[62135] = 8'b0;
    XRAM[62136] = 8'b0;
    XRAM[62137] = 8'b0;
    XRAM[62138] = 8'b0;
    XRAM[62139] = 8'b0;
    XRAM[62140] = 8'b0;
    XRAM[62141] = 8'b0;
    XRAM[62142] = 8'b0;
    XRAM[62143] = 8'b0;
    XRAM[62144] = 8'b0;
    XRAM[62145] = 8'b0;
    XRAM[62146] = 8'b0;
    XRAM[62147] = 8'b0;
    XRAM[62148] = 8'b0;
    XRAM[62149] = 8'b0;
    XRAM[62150] = 8'b0;
    XRAM[62151] = 8'b0;
    XRAM[62152] = 8'b0;
    XRAM[62153] = 8'b0;
    XRAM[62154] = 8'b0;
    XRAM[62155] = 8'b0;
    XRAM[62156] = 8'b0;
    XRAM[62157] = 8'b0;
    XRAM[62158] = 8'b0;
    XRAM[62159] = 8'b0;
    XRAM[62160] = 8'b0;
    XRAM[62161] = 8'b0;
    XRAM[62162] = 8'b0;
    XRAM[62163] = 8'b0;
    XRAM[62164] = 8'b0;
    XRAM[62165] = 8'b0;
    XRAM[62166] = 8'b0;
    XRAM[62167] = 8'b0;
    XRAM[62168] = 8'b0;
    XRAM[62169] = 8'b0;
    XRAM[62170] = 8'b0;
    XRAM[62171] = 8'b0;
    XRAM[62172] = 8'b0;
    XRAM[62173] = 8'b0;
    XRAM[62174] = 8'b0;
    XRAM[62175] = 8'b0;
    XRAM[62176] = 8'b0;
    XRAM[62177] = 8'b0;
    XRAM[62178] = 8'b0;
    XRAM[62179] = 8'b0;
    XRAM[62180] = 8'b0;
    XRAM[62181] = 8'b0;
    XRAM[62182] = 8'b0;
    XRAM[62183] = 8'b0;
    XRAM[62184] = 8'b0;
    XRAM[62185] = 8'b0;
    XRAM[62186] = 8'b0;
    XRAM[62187] = 8'b0;
    XRAM[62188] = 8'b0;
    XRAM[62189] = 8'b0;
    XRAM[62190] = 8'b0;
    XRAM[62191] = 8'b0;
    XRAM[62192] = 8'b0;
    XRAM[62193] = 8'b0;
    XRAM[62194] = 8'b0;
    XRAM[62195] = 8'b0;
    XRAM[62196] = 8'b0;
    XRAM[62197] = 8'b0;
    XRAM[62198] = 8'b0;
    XRAM[62199] = 8'b0;
    XRAM[62200] = 8'b0;
    XRAM[62201] = 8'b0;
    XRAM[62202] = 8'b0;
    XRAM[62203] = 8'b0;
    XRAM[62204] = 8'b0;
    XRAM[62205] = 8'b0;
    XRAM[62206] = 8'b0;
    XRAM[62207] = 8'b0;
    XRAM[62208] = 8'b0;
    XRAM[62209] = 8'b0;
    XRAM[62210] = 8'b0;
    XRAM[62211] = 8'b0;
    XRAM[62212] = 8'b0;
    XRAM[62213] = 8'b0;
    XRAM[62214] = 8'b0;
    XRAM[62215] = 8'b0;
    XRAM[62216] = 8'b0;
    XRAM[62217] = 8'b0;
    XRAM[62218] = 8'b0;
    XRAM[62219] = 8'b0;
    XRAM[62220] = 8'b0;
    XRAM[62221] = 8'b0;
    XRAM[62222] = 8'b0;
    XRAM[62223] = 8'b0;
    XRAM[62224] = 8'b0;
    XRAM[62225] = 8'b0;
    XRAM[62226] = 8'b0;
    XRAM[62227] = 8'b0;
    XRAM[62228] = 8'b0;
    XRAM[62229] = 8'b0;
    XRAM[62230] = 8'b0;
    XRAM[62231] = 8'b0;
    XRAM[62232] = 8'b0;
    XRAM[62233] = 8'b0;
    XRAM[62234] = 8'b0;
    XRAM[62235] = 8'b0;
    XRAM[62236] = 8'b0;
    XRAM[62237] = 8'b0;
    XRAM[62238] = 8'b0;
    XRAM[62239] = 8'b0;
    XRAM[62240] = 8'b0;
    XRAM[62241] = 8'b0;
    XRAM[62242] = 8'b0;
    XRAM[62243] = 8'b0;
    XRAM[62244] = 8'b0;
    XRAM[62245] = 8'b0;
    XRAM[62246] = 8'b0;
    XRAM[62247] = 8'b0;
    XRAM[62248] = 8'b0;
    XRAM[62249] = 8'b0;
    XRAM[62250] = 8'b0;
    XRAM[62251] = 8'b0;
    XRAM[62252] = 8'b0;
    XRAM[62253] = 8'b0;
    XRAM[62254] = 8'b0;
    XRAM[62255] = 8'b0;
    XRAM[62256] = 8'b0;
    XRAM[62257] = 8'b0;
    XRAM[62258] = 8'b0;
    XRAM[62259] = 8'b0;
    XRAM[62260] = 8'b0;
    XRAM[62261] = 8'b0;
    XRAM[62262] = 8'b0;
    XRAM[62263] = 8'b0;
    XRAM[62264] = 8'b0;
    XRAM[62265] = 8'b0;
    XRAM[62266] = 8'b0;
    XRAM[62267] = 8'b0;
    XRAM[62268] = 8'b0;
    XRAM[62269] = 8'b0;
    XRAM[62270] = 8'b0;
    XRAM[62271] = 8'b0;
    XRAM[62272] = 8'b0;
    XRAM[62273] = 8'b0;
    XRAM[62274] = 8'b0;
    XRAM[62275] = 8'b0;
    XRAM[62276] = 8'b0;
    XRAM[62277] = 8'b0;
    XRAM[62278] = 8'b0;
    XRAM[62279] = 8'b0;
    XRAM[62280] = 8'b0;
    XRAM[62281] = 8'b0;
    XRAM[62282] = 8'b0;
    XRAM[62283] = 8'b0;
    XRAM[62284] = 8'b0;
    XRAM[62285] = 8'b0;
    XRAM[62286] = 8'b0;
    XRAM[62287] = 8'b0;
    XRAM[62288] = 8'b0;
    XRAM[62289] = 8'b0;
    XRAM[62290] = 8'b0;
    XRAM[62291] = 8'b0;
    XRAM[62292] = 8'b0;
    XRAM[62293] = 8'b0;
    XRAM[62294] = 8'b0;
    XRAM[62295] = 8'b0;
    XRAM[62296] = 8'b0;
    XRAM[62297] = 8'b0;
    XRAM[62298] = 8'b0;
    XRAM[62299] = 8'b0;
    XRAM[62300] = 8'b0;
    XRAM[62301] = 8'b0;
    XRAM[62302] = 8'b0;
    XRAM[62303] = 8'b0;
    XRAM[62304] = 8'b0;
    XRAM[62305] = 8'b0;
    XRAM[62306] = 8'b0;
    XRAM[62307] = 8'b0;
    XRAM[62308] = 8'b0;
    XRAM[62309] = 8'b0;
    XRAM[62310] = 8'b0;
    XRAM[62311] = 8'b0;
    XRAM[62312] = 8'b0;
    XRAM[62313] = 8'b0;
    XRAM[62314] = 8'b0;
    XRAM[62315] = 8'b0;
    XRAM[62316] = 8'b0;
    XRAM[62317] = 8'b0;
    XRAM[62318] = 8'b0;
    XRAM[62319] = 8'b0;
    XRAM[62320] = 8'b0;
    XRAM[62321] = 8'b0;
    XRAM[62322] = 8'b0;
    XRAM[62323] = 8'b0;
    XRAM[62324] = 8'b0;
    XRAM[62325] = 8'b0;
    XRAM[62326] = 8'b0;
    XRAM[62327] = 8'b0;
    XRAM[62328] = 8'b0;
    XRAM[62329] = 8'b0;
    XRAM[62330] = 8'b0;
    XRAM[62331] = 8'b0;
    XRAM[62332] = 8'b0;
    XRAM[62333] = 8'b0;
    XRAM[62334] = 8'b0;
    XRAM[62335] = 8'b0;
    XRAM[62336] = 8'b0;
    XRAM[62337] = 8'b0;
    XRAM[62338] = 8'b0;
    XRAM[62339] = 8'b0;
    XRAM[62340] = 8'b0;
    XRAM[62341] = 8'b0;
    XRAM[62342] = 8'b0;
    XRAM[62343] = 8'b0;
    XRAM[62344] = 8'b0;
    XRAM[62345] = 8'b0;
    XRAM[62346] = 8'b0;
    XRAM[62347] = 8'b0;
    XRAM[62348] = 8'b0;
    XRAM[62349] = 8'b0;
    XRAM[62350] = 8'b0;
    XRAM[62351] = 8'b0;
    XRAM[62352] = 8'b0;
    XRAM[62353] = 8'b0;
    XRAM[62354] = 8'b0;
    XRAM[62355] = 8'b0;
    XRAM[62356] = 8'b0;
    XRAM[62357] = 8'b0;
    XRAM[62358] = 8'b0;
    XRAM[62359] = 8'b0;
    XRAM[62360] = 8'b0;
    XRAM[62361] = 8'b0;
    XRAM[62362] = 8'b0;
    XRAM[62363] = 8'b0;
    XRAM[62364] = 8'b0;
    XRAM[62365] = 8'b0;
    XRAM[62366] = 8'b0;
    XRAM[62367] = 8'b0;
    XRAM[62368] = 8'b0;
    XRAM[62369] = 8'b0;
    XRAM[62370] = 8'b0;
    XRAM[62371] = 8'b0;
    XRAM[62372] = 8'b0;
    XRAM[62373] = 8'b0;
    XRAM[62374] = 8'b0;
    XRAM[62375] = 8'b0;
    XRAM[62376] = 8'b0;
    XRAM[62377] = 8'b0;
    XRAM[62378] = 8'b0;
    XRAM[62379] = 8'b0;
    XRAM[62380] = 8'b0;
    XRAM[62381] = 8'b0;
    XRAM[62382] = 8'b0;
    XRAM[62383] = 8'b0;
    XRAM[62384] = 8'b0;
    XRAM[62385] = 8'b0;
    XRAM[62386] = 8'b0;
    XRAM[62387] = 8'b0;
    XRAM[62388] = 8'b0;
    XRAM[62389] = 8'b0;
    XRAM[62390] = 8'b0;
    XRAM[62391] = 8'b0;
    XRAM[62392] = 8'b0;
    XRAM[62393] = 8'b0;
    XRAM[62394] = 8'b0;
    XRAM[62395] = 8'b0;
    XRAM[62396] = 8'b0;
    XRAM[62397] = 8'b0;
    XRAM[62398] = 8'b0;
    XRAM[62399] = 8'b0;
    XRAM[62400] = 8'b0;
    XRAM[62401] = 8'b0;
    XRAM[62402] = 8'b0;
    XRAM[62403] = 8'b0;
    XRAM[62404] = 8'b0;
    XRAM[62405] = 8'b0;
    XRAM[62406] = 8'b0;
    XRAM[62407] = 8'b0;
    XRAM[62408] = 8'b0;
    XRAM[62409] = 8'b0;
    XRAM[62410] = 8'b0;
    XRAM[62411] = 8'b0;
    XRAM[62412] = 8'b0;
    XRAM[62413] = 8'b0;
    XRAM[62414] = 8'b0;
    XRAM[62415] = 8'b0;
    XRAM[62416] = 8'b0;
    XRAM[62417] = 8'b0;
    XRAM[62418] = 8'b0;
    XRAM[62419] = 8'b0;
    XRAM[62420] = 8'b0;
    XRAM[62421] = 8'b0;
    XRAM[62422] = 8'b0;
    XRAM[62423] = 8'b0;
    XRAM[62424] = 8'b0;
    XRAM[62425] = 8'b0;
    XRAM[62426] = 8'b0;
    XRAM[62427] = 8'b0;
    XRAM[62428] = 8'b0;
    XRAM[62429] = 8'b0;
    XRAM[62430] = 8'b0;
    XRAM[62431] = 8'b0;
    XRAM[62432] = 8'b0;
    XRAM[62433] = 8'b0;
    XRAM[62434] = 8'b0;
    XRAM[62435] = 8'b0;
    XRAM[62436] = 8'b0;
    XRAM[62437] = 8'b0;
    XRAM[62438] = 8'b0;
    XRAM[62439] = 8'b0;
    XRAM[62440] = 8'b0;
    XRAM[62441] = 8'b0;
    XRAM[62442] = 8'b0;
    XRAM[62443] = 8'b0;
    XRAM[62444] = 8'b0;
    XRAM[62445] = 8'b0;
    XRAM[62446] = 8'b0;
    XRAM[62447] = 8'b0;
    XRAM[62448] = 8'b0;
    XRAM[62449] = 8'b0;
    XRAM[62450] = 8'b0;
    XRAM[62451] = 8'b0;
    XRAM[62452] = 8'b0;
    XRAM[62453] = 8'b0;
    XRAM[62454] = 8'b0;
    XRAM[62455] = 8'b0;
    XRAM[62456] = 8'b0;
    XRAM[62457] = 8'b0;
    XRAM[62458] = 8'b0;
    XRAM[62459] = 8'b0;
    XRAM[62460] = 8'b0;
    XRAM[62461] = 8'b0;
    XRAM[62462] = 8'b0;
    XRAM[62463] = 8'b0;
    XRAM[62464] = 8'b0;
    XRAM[62465] = 8'b0;
    XRAM[62466] = 8'b0;
    XRAM[62467] = 8'b0;
    XRAM[62468] = 8'b0;
    XRAM[62469] = 8'b0;
    XRAM[62470] = 8'b0;
    XRAM[62471] = 8'b0;
    XRAM[62472] = 8'b0;
    XRAM[62473] = 8'b0;
    XRAM[62474] = 8'b0;
    XRAM[62475] = 8'b0;
    XRAM[62476] = 8'b0;
    XRAM[62477] = 8'b0;
    XRAM[62478] = 8'b0;
    XRAM[62479] = 8'b0;
    XRAM[62480] = 8'b0;
    XRAM[62481] = 8'b0;
    XRAM[62482] = 8'b0;
    XRAM[62483] = 8'b0;
    XRAM[62484] = 8'b0;
    XRAM[62485] = 8'b0;
    XRAM[62486] = 8'b0;
    XRAM[62487] = 8'b0;
    XRAM[62488] = 8'b0;
    XRAM[62489] = 8'b0;
    XRAM[62490] = 8'b0;
    XRAM[62491] = 8'b0;
    XRAM[62492] = 8'b0;
    XRAM[62493] = 8'b0;
    XRAM[62494] = 8'b0;
    XRAM[62495] = 8'b0;
    XRAM[62496] = 8'b0;
    XRAM[62497] = 8'b0;
    XRAM[62498] = 8'b0;
    XRAM[62499] = 8'b0;
    XRAM[62500] = 8'b0;
    XRAM[62501] = 8'b0;
    XRAM[62502] = 8'b0;
    XRAM[62503] = 8'b0;
    XRAM[62504] = 8'b0;
    XRAM[62505] = 8'b0;
    XRAM[62506] = 8'b0;
    XRAM[62507] = 8'b0;
    XRAM[62508] = 8'b0;
    XRAM[62509] = 8'b0;
    XRAM[62510] = 8'b0;
    XRAM[62511] = 8'b0;
    XRAM[62512] = 8'b0;
    XRAM[62513] = 8'b0;
    XRAM[62514] = 8'b0;
    XRAM[62515] = 8'b0;
    XRAM[62516] = 8'b0;
    XRAM[62517] = 8'b0;
    XRAM[62518] = 8'b0;
    XRAM[62519] = 8'b0;
    XRAM[62520] = 8'b0;
    XRAM[62521] = 8'b0;
    XRAM[62522] = 8'b0;
    XRAM[62523] = 8'b0;
    XRAM[62524] = 8'b0;
    XRAM[62525] = 8'b0;
    XRAM[62526] = 8'b0;
    XRAM[62527] = 8'b0;
    XRAM[62528] = 8'b0;
    XRAM[62529] = 8'b0;
    XRAM[62530] = 8'b0;
    XRAM[62531] = 8'b0;
    XRAM[62532] = 8'b0;
    XRAM[62533] = 8'b0;
    XRAM[62534] = 8'b0;
    XRAM[62535] = 8'b0;
    XRAM[62536] = 8'b0;
    XRAM[62537] = 8'b0;
    XRAM[62538] = 8'b0;
    XRAM[62539] = 8'b0;
    XRAM[62540] = 8'b0;
    XRAM[62541] = 8'b0;
    XRAM[62542] = 8'b0;
    XRAM[62543] = 8'b0;
    XRAM[62544] = 8'b0;
    XRAM[62545] = 8'b0;
    XRAM[62546] = 8'b0;
    XRAM[62547] = 8'b0;
    XRAM[62548] = 8'b0;
    XRAM[62549] = 8'b0;
    XRAM[62550] = 8'b0;
    XRAM[62551] = 8'b0;
    XRAM[62552] = 8'b0;
    XRAM[62553] = 8'b0;
    XRAM[62554] = 8'b0;
    XRAM[62555] = 8'b0;
    XRAM[62556] = 8'b0;
    XRAM[62557] = 8'b0;
    XRAM[62558] = 8'b0;
    XRAM[62559] = 8'b0;
    XRAM[62560] = 8'b0;
    XRAM[62561] = 8'b0;
    XRAM[62562] = 8'b0;
    XRAM[62563] = 8'b0;
    XRAM[62564] = 8'b0;
    XRAM[62565] = 8'b0;
    XRAM[62566] = 8'b0;
    XRAM[62567] = 8'b0;
    XRAM[62568] = 8'b0;
    XRAM[62569] = 8'b0;
    XRAM[62570] = 8'b0;
    XRAM[62571] = 8'b0;
    XRAM[62572] = 8'b0;
    XRAM[62573] = 8'b0;
    XRAM[62574] = 8'b0;
    XRAM[62575] = 8'b0;
    XRAM[62576] = 8'b0;
    XRAM[62577] = 8'b0;
    XRAM[62578] = 8'b0;
    XRAM[62579] = 8'b0;
    XRAM[62580] = 8'b0;
    XRAM[62581] = 8'b0;
    XRAM[62582] = 8'b0;
    XRAM[62583] = 8'b0;
    XRAM[62584] = 8'b0;
    XRAM[62585] = 8'b0;
    XRAM[62586] = 8'b0;
    XRAM[62587] = 8'b0;
    XRAM[62588] = 8'b0;
    XRAM[62589] = 8'b0;
    XRAM[62590] = 8'b0;
    XRAM[62591] = 8'b0;
    XRAM[62592] = 8'b0;
    XRAM[62593] = 8'b0;
    XRAM[62594] = 8'b0;
    XRAM[62595] = 8'b0;
    XRAM[62596] = 8'b0;
    XRAM[62597] = 8'b0;
    XRAM[62598] = 8'b0;
    XRAM[62599] = 8'b0;
    XRAM[62600] = 8'b0;
    XRAM[62601] = 8'b0;
    XRAM[62602] = 8'b0;
    XRAM[62603] = 8'b0;
    XRAM[62604] = 8'b0;
    XRAM[62605] = 8'b0;
    XRAM[62606] = 8'b0;
    XRAM[62607] = 8'b0;
    XRAM[62608] = 8'b0;
    XRAM[62609] = 8'b0;
    XRAM[62610] = 8'b0;
    XRAM[62611] = 8'b0;
    XRAM[62612] = 8'b0;
    XRAM[62613] = 8'b0;
    XRAM[62614] = 8'b0;
    XRAM[62615] = 8'b0;
    XRAM[62616] = 8'b0;
    XRAM[62617] = 8'b0;
    XRAM[62618] = 8'b0;
    XRAM[62619] = 8'b0;
    XRAM[62620] = 8'b0;
    XRAM[62621] = 8'b0;
    XRAM[62622] = 8'b0;
    XRAM[62623] = 8'b0;
    XRAM[62624] = 8'b0;
    XRAM[62625] = 8'b0;
    XRAM[62626] = 8'b0;
    XRAM[62627] = 8'b0;
    XRAM[62628] = 8'b0;
    XRAM[62629] = 8'b0;
    XRAM[62630] = 8'b0;
    XRAM[62631] = 8'b0;
    XRAM[62632] = 8'b0;
    XRAM[62633] = 8'b0;
    XRAM[62634] = 8'b0;
    XRAM[62635] = 8'b0;
    XRAM[62636] = 8'b0;
    XRAM[62637] = 8'b0;
    XRAM[62638] = 8'b0;
    XRAM[62639] = 8'b0;
    XRAM[62640] = 8'b0;
    XRAM[62641] = 8'b0;
    XRAM[62642] = 8'b0;
    XRAM[62643] = 8'b0;
    XRAM[62644] = 8'b0;
    XRAM[62645] = 8'b0;
    XRAM[62646] = 8'b0;
    XRAM[62647] = 8'b0;
    XRAM[62648] = 8'b0;
    XRAM[62649] = 8'b0;
    XRAM[62650] = 8'b0;
    XRAM[62651] = 8'b0;
    XRAM[62652] = 8'b0;
    XRAM[62653] = 8'b0;
    XRAM[62654] = 8'b0;
    XRAM[62655] = 8'b0;
    XRAM[62656] = 8'b0;
    XRAM[62657] = 8'b0;
    XRAM[62658] = 8'b0;
    XRAM[62659] = 8'b0;
    XRAM[62660] = 8'b0;
    XRAM[62661] = 8'b0;
    XRAM[62662] = 8'b0;
    XRAM[62663] = 8'b0;
    XRAM[62664] = 8'b0;
    XRAM[62665] = 8'b0;
    XRAM[62666] = 8'b0;
    XRAM[62667] = 8'b0;
    XRAM[62668] = 8'b0;
    XRAM[62669] = 8'b0;
    XRAM[62670] = 8'b0;
    XRAM[62671] = 8'b0;
    XRAM[62672] = 8'b0;
    XRAM[62673] = 8'b0;
    XRAM[62674] = 8'b0;
    XRAM[62675] = 8'b0;
    XRAM[62676] = 8'b0;
    XRAM[62677] = 8'b0;
    XRAM[62678] = 8'b0;
    XRAM[62679] = 8'b0;
    XRAM[62680] = 8'b0;
    XRAM[62681] = 8'b0;
    XRAM[62682] = 8'b0;
    XRAM[62683] = 8'b0;
    XRAM[62684] = 8'b0;
    XRAM[62685] = 8'b0;
    XRAM[62686] = 8'b0;
    XRAM[62687] = 8'b0;
    XRAM[62688] = 8'b0;
    XRAM[62689] = 8'b0;
    XRAM[62690] = 8'b0;
    XRAM[62691] = 8'b0;
    XRAM[62692] = 8'b0;
    XRAM[62693] = 8'b0;
    XRAM[62694] = 8'b0;
    XRAM[62695] = 8'b0;
    XRAM[62696] = 8'b0;
    XRAM[62697] = 8'b0;
    XRAM[62698] = 8'b0;
    XRAM[62699] = 8'b0;
    XRAM[62700] = 8'b0;
    XRAM[62701] = 8'b0;
    XRAM[62702] = 8'b0;
    XRAM[62703] = 8'b0;
    XRAM[62704] = 8'b0;
    XRAM[62705] = 8'b0;
    XRAM[62706] = 8'b0;
    XRAM[62707] = 8'b0;
    XRAM[62708] = 8'b0;
    XRAM[62709] = 8'b0;
    XRAM[62710] = 8'b0;
    XRAM[62711] = 8'b0;
    XRAM[62712] = 8'b0;
    XRAM[62713] = 8'b0;
    XRAM[62714] = 8'b0;
    XRAM[62715] = 8'b0;
    XRAM[62716] = 8'b0;
    XRAM[62717] = 8'b0;
    XRAM[62718] = 8'b0;
    XRAM[62719] = 8'b0;
    XRAM[62720] = 8'b0;
    XRAM[62721] = 8'b0;
    XRAM[62722] = 8'b0;
    XRAM[62723] = 8'b0;
    XRAM[62724] = 8'b0;
    XRAM[62725] = 8'b0;
    XRAM[62726] = 8'b0;
    XRAM[62727] = 8'b0;
    XRAM[62728] = 8'b0;
    XRAM[62729] = 8'b0;
    XRAM[62730] = 8'b0;
    XRAM[62731] = 8'b0;
    XRAM[62732] = 8'b0;
    XRAM[62733] = 8'b0;
    XRAM[62734] = 8'b0;
    XRAM[62735] = 8'b0;
    XRAM[62736] = 8'b0;
    XRAM[62737] = 8'b0;
    XRAM[62738] = 8'b0;
    XRAM[62739] = 8'b0;
    XRAM[62740] = 8'b0;
    XRAM[62741] = 8'b0;
    XRAM[62742] = 8'b0;
    XRAM[62743] = 8'b0;
    XRAM[62744] = 8'b0;
    XRAM[62745] = 8'b0;
    XRAM[62746] = 8'b0;
    XRAM[62747] = 8'b0;
    XRAM[62748] = 8'b0;
    XRAM[62749] = 8'b0;
    XRAM[62750] = 8'b0;
    XRAM[62751] = 8'b0;
    XRAM[62752] = 8'b0;
    XRAM[62753] = 8'b0;
    XRAM[62754] = 8'b0;
    XRAM[62755] = 8'b0;
    XRAM[62756] = 8'b0;
    XRAM[62757] = 8'b0;
    XRAM[62758] = 8'b0;
    XRAM[62759] = 8'b0;
    XRAM[62760] = 8'b0;
    XRAM[62761] = 8'b0;
    XRAM[62762] = 8'b0;
    XRAM[62763] = 8'b0;
    XRAM[62764] = 8'b0;
    XRAM[62765] = 8'b0;
    XRAM[62766] = 8'b0;
    XRAM[62767] = 8'b0;
    XRAM[62768] = 8'b0;
    XRAM[62769] = 8'b0;
    XRAM[62770] = 8'b0;
    XRAM[62771] = 8'b0;
    XRAM[62772] = 8'b0;
    XRAM[62773] = 8'b0;
    XRAM[62774] = 8'b0;
    XRAM[62775] = 8'b0;
    XRAM[62776] = 8'b0;
    XRAM[62777] = 8'b0;
    XRAM[62778] = 8'b0;
    XRAM[62779] = 8'b0;
    XRAM[62780] = 8'b0;
    XRAM[62781] = 8'b0;
    XRAM[62782] = 8'b0;
    XRAM[62783] = 8'b0;
    XRAM[62784] = 8'b0;
    XRAM[62785] = 8'b0;
    XRAM[62786] = 8'b0;
    XRAM[62787] = 8'b0;
    XRAM[62788] = 8'b0;
    XRAM[62789] = 8'b0;
    XRAM[62790] = 8'b0;
    XRAM[62791] = 8'b0;
    XRAM[62792] = 8'b0;
    XRAM[62793] = 8'b0;
    XRAM[62794] = 8'b0;
    XRAM[62795] = 8'b0;
    XRAM[62796] = 8'b0;
    XRAM[62797] = 8'b0;
    XRAM[62798] = 8'b0;
    XRAM[62799] = 8'b0;
    XRAM[62800] = 8'b0;
    XRAM[62801] = 8'b0;
    XRAM[62802] = 8'b0;
    XRAM[62803] = 8'b0;
    XRAM[62804] = 8'b0;
    XRAM[62805] = 8'b0;
    XRAM[62806] = 8'b0;
    XRAM[62807] = 8'b0;
    XRAM[62808] = 8'b0;
    XRAM[62809] = 8'b0;
    XRAM[62810] = 8'b0;
    XRAM[62811] = 8'b0;
    XRAM[62812] = 8'b0;
    XRAM[62813] = 8'b0;
    XRAM[62814] = 8'b0;
    XRAM[62815] = 8'b0;
    XRAM[62816] = 8'b0;
    XRAM[62817] = 8'b0;
    XRAM[62818] = 8'b0;
    XRAM[62819] = 8'b0;
    XRAM[62820] = 8'b0;
    XRAM[62821] = 8'b0;
    XRAM[62822] = 8'b0;
    XRAM[62823] = 8'b0;
    XRAM[62824] = 8'b0;
    XRAM[62825] = 8'b0;
    XRAM[62826] = 8'b0;
    XRAM[62827] = 8'b0;
    XRAM[62828] = 8'b0;
    XRAM[62829] = 8'b0;
    XRAM[62830] = 8'b0;
    XRAM[62831] = 8'b0;
    XRAM[62832] = 8'b0;
    XRAM[62833] = 8'b0;
    XRAM[62834] = 8'b0;
    XRAM[62835] = 8'b0;
    XRAM[62836] = 8'b0;
    XRAM[62837] = 8'b0;
    XRAM[62838] = 8'b0;
    XRAM[62839] = 8'b0;
    XRAM[62840] = 8'b0;
    XRAM[62841] = 8'b0;
    XRAM[62842] = 8'b0;
    XRAM[62843] = 8'b0;
    XRAM[62844] = 8'b0;
    XRAM[62845] = 8'b0;
    XRAM[62846] = 8'b0;
    XRAM[62847] = 8'b0;
    XRAM[62848] = 8'b0;
    XRAM[62849] = 8'b0;
    XRAM[62850] = 8'b0;
    XRAM[62851] = 8'b0;
    XRAM[62852] = 8'b0;
    XRAM[62853] = 8'b0;
    XRAM[62854] = 8'b0;
    XRAM[62855] = 8'b0;
    XRAM[62856] = 8'b0;
    XRAM[62857] = 8'b0;
    XRAM[62858] = 8'b0;
    XRAM[62859] = 8'b0;
    XRAM[62860] = 8'b0;
    XRAM[62861] = 8'b0;
    XRAM[62862] = 8'b0;
    XRAM[62863] = 8'b0;
    XRAM[62864] = 8'b0;
    XRAM[62865] = 8'b0;
    XRAM[62866] = 8'b0;
    XRAM[62867] = 8'b0;
    XRAM[62868] = 8'b0;
    XRAM[62869] = 8'b0;
    XRAM[62870] = 8'b0;
    XRAM[62871] = 8'b0;
    XRAM[62872] = 8'b0;
    XRAM[62873] = 8'b0;
    XRAM[62874] = 8'b0;
    XRAM[62875] = 8'b0;
    XRAM[62876] = 8'b0;
    XRAM[62877] = 8'b0;
    XRAM[62878] = 8'b0;
    XRAM[62879] = 8'b0;
    XRAM[62880] = 8'b0;
    XRAM[62881] = 8'b0;
    XRAM[62882] = 8'b0;
    XRAM[62883] = 8'b0;
    XRAM[62884] = 8'b0;
    XRAM[62885] = 8'b0;
    XRAM[62886] = 8'b0;
    XRAM[62887] = 8'b0;
    XRAM[62888] = 8'b0;
    XRAM[62889] = 8'b0;
    XRAM[62890] = 8'b0;
    XRAM[62891] = 8'b0;
    XRAM[62892] = 8'b0;
    XRAM[62893] = 8'b0;
    XRAM[62894] = 8'b0;
    XRAM[62895] = 8'b0;
    XRAM[62896] = 8'b0;
    XRAM[62897] = 8'b0;
    XRAM[62898] = 8'b0;
    XRAM[62899] = 8'b0;
    XRAM[62900] = 8'b0;
    XRAM[62901] = 8'b0;
    XRAM[62902] = 8'b0;
    XRAM[62903] = 8'b0;
    XRAM[62904] = 8'b0;
    XRAM[62905] = 8'b0;
    XRAM[62906] = 8'b0;
    XRAM[62907] = 8'b0;
    XRAM[62908] = 8'b0;
    XRAM[62909] = 8'b0;
    XRAM[62910] = 8'b0;
    XRAM[62911] = 8'b0;
    XRAM[62912] = 8'b0;
    XRAM[62913] = 8'b0;
    XRAM[62914] = 8'b0;
    XRAM[62915] = 8'b0;
    XRAM[62916] = 8'b0;
    XRAM[62917] = 8'b0;
    XRAM[62918] = 8'b0;
    XRAM[62919] = 8'b0;
    XRAM[62920] = 8'b0;
    XRAM[62921] = 8'b0;
    XRAM[62922] = 8'b0;
    XRAM[62923] = 8'b0;
    XRAM[62924] = 8'b0;
    XRAM[62925] = 8'b0;
    XRAM[62926] = 8'b0;
    XRAM[62927] = 8'b0;
    XRAM[62928] = 8'b0;
    XRAM[62929] = 8'b0;
    XRAM[62930] = 8'b0;
    XRAM[62931] = 8'b0;
    XRAM[62932] = 8'b0;
    XRAM[62933] = 8'b0;
    XRAM[62934] = 8'b0;
    XRAM[62935] = 8'b0;
    XRAM[62936] = 8'b0;
    XRAM[62937] = 8'b0;
    XRAM[62938] = 8'b0;
    XRAM[62939] = 8'b0;
    XRAM[62940] = 8'b0;
    XRAM[62941] = 8'b0;
    XRAM[62942] = 8'b0;
    XRAM[62943] = 8'b0;
    XRAM[62944] = 8'b0;
    XRAM[62945] = 8'b0;
    XRAM[62946] = 8'b0;
    XRAM[62947] = 8'b0;
    XRAM[62948] = 8'b0;
    XRAM[62949] = 8'b0;
    XRAM[62950] = 8'b0;
    XRAM[62951] = 8'b0;
    XRAM[62952] = 8'b0;
    XRAM[62953] = 8'b0;
    XRAM[62954] = 8'b0;
    XRAM[62955] = 8'b0;
    XRAM[62956] = 8'b0;
    XRAM[62957] = 8'b0;
    XRAM[62958] = 8'b0;
    XRAM[62959] = 8'b0;
    XRAM[62960] = 8'b0;
    XRAM[62961] = 8'b0;
    XRAM[62962] = 8'b0;
    XRAM[62963] = 8'b0;
    XRAM[62964] = 8'b0;
    XRAM[62965] = 8'b0;
    XRAM[62966] = 8'b0;
    XRAM[62967] = 8'b0;
    XRAM[62968] = 8'b0;
    XRAM[62969] = 8'b0;
    XRAM[62970] = 8'b0;
    XRAM[62971] = 8'b0;
    XRAM[62972] = 8'b0;
    XRAM[62973] = 8'b0;
    XRAM[62974] = 8'b0;
    XRAM[62975] = 8'b0;
    XRAM[62976] = 8'b0;
    XRAM[62977] = 8'b0;
    XRAM[62978] = 8'b0;
    XRAM[62979] = 8'b0;
    XRAM[62980] = 8'b0;
    XRAM[62981] = 8'b0;
    XRAM[62982] = 8'b0;
    XRAM[62983] = 8'b0;
    XRAM[62984] = 8'b0;
    XRAM[62985] = 8'b0;
    XRAM[62986] = 8'b0;
    XRAM[62987] = 8'b0;
    XRAM[62988] = 8'b0;
    XRAM[62989] = 8'b0;
    XRAM[62990] = 8'b0;
    XRAM[62991] = 8'b0;
    XRAM[62992] = 8'b0;
    XRAM[62993] = 8'b0;
    XRAM[62994] = 8'b0;
    XRAM[62995] = 8'b0;
    XRAM[62996] = 8'b0;
    XRAM[62997] = 8'b0;
    XRAM[62998] = 8'b0;
    XRAM[62999] = 8'b0;
    XRAM[63000] = 8'b0;
    XRAM[63001] = 8'b0;
    XRAM[63002] = 8'b0;
    XRAM[63003] = 8'b0;
    XRAM[63004] = 8'b0;
    XRAM[63005] = 8'b0;
    XRAM[63006] = 8'b0;
    XRAM[63007] = 8'b0;
    XRAM[63008] = 8'b0;
    XRAM[63009] = 8'b0;
    XRAM[63010] = 8'b0;
    XRAM[63011] = 8'b0;
    XRAM[63012] = 8'b0;
    XRAM[63013] = 8'b0;
    XRAM[63014] = 8'b0;
    XRAM[63015] = 8'b0;
    XRAM[63016] = 8'b0;
    XRAM[63017] = 8'b0;
    XRAM[63018] = 8'b0;
    XRAM[63019] = 8'b0;
    XRAM[63020] = 8'b0;
    XRAM[63021] = 8'b0;
    XRAM[63022] = 8'b0;
    XRAM[63023] = 8'b0;
    XRAM[63024] = 8'b0;
    XRAM[63025] = 8'b0;
    XRAM[63026] = 8'b0;
    XRAM[63027] = 8'b0;
    XRAM[63028] = 8'b0;
    XRAM[63029] = 8'b0;
    XRAM[63030] = 8'b0;
    XRAM[63031] = 8'b0;
    XRAM[63032] = 8'b0;
    XRAM[63033] = 8'b0;
    XRAM[63034] = 8'b0;
    XRAM[63035] = 8'b0;
    XRAM[63036] = 8'b0;
    XRAM[63037] = 8'b0;
    XRAM[63038] = 8'b0;
    XRAM[63039] = 8'b0;
    XRAM[63040] = 8'b0;
    XRAM[63041] = 8'b0;
    XRAM[63042] = 8'b0;
    XRAM[63043] = 8'b0;
    XRAM[63044] = 8'b0;
    XRAM[63045] = 8'b0;
    XRAM[63046] = 8'b0;
    XRAM[63047] = 8'b0;
    XRAM[63048] = 8'b0;
    XRAM[63049] = 8'b0;
    XRAM[63050] = 8'b0;
    XRAM[63051] = 8'b0;
    XRAM[63052] = 8'b0;
    XRAM[63053] = 8'b0;
    XRAM[63054] = 8'b0;
    XRAM[63055] = 8'b0;
    XRAM[63056] = 8'b0;
    XRAM[63057] = 8'b0;
    XRAM[63058] = 8'b0;
    XRAM[63059] = 8'b0;
    XRAM[63060] = 8'b0;
    XRAM[63061] = 8'b0;
    XRAM[63062] = 8'b0;
    XRAM[63063] = 8'b0;
    XRAM[63064] = 8'b0;
    XRAM[63065] = 8'b0;
    XRAM[63066] = 8'b0;
    XRAM[63067] = 8'b0;
    XRAM[63068] = 8'b0;
    XRAM[63069] = 8'b0;
    XRAM[63070] = 8'b0;
    XRAM[63071] = 8'b0;
    XRAM[63072] = 8'b0;
    XRAM[63073] = 8'b0;
    XRAM[63074] = 8'b0;
    XRAM[63075] = 8'b0;
    XRAM[63076] = 8'b0;
    XRAM[63077] = 8'b0;
    XRAM[63078] = 8'b0;
    XRAM[63079] = 8'b0;
    XRAM[63080] = 8'b0;
    XRAM[63081] = 8'b0;
    XRAM[63082] = 8'b0;
    XRAM[63083] = 8'b0;
    XRAM[63084] = 8'b0;
    XRAM[63085] = 8'b0;
    XRAM[63086] = 8'b0;
    XRAM[63087] = 8'b0;
    XRAM[63088] = 8'b0;
    XRAM[63089] = 8'b0;
    XRAM[63090] = 8'b0;
    XRAM[63091] = 8'b0;
    XRAM[63092] = 8'b0;
    XRAM[63093] = 8'b0;
    XRAM[63094] = 8'b0;
    XRAM[63095] = 8'b0;
    XRAM[63096] = 8'b0;
    XRAM[63097] = 8'b0;
    XRAM[63098] = 8'b0;
    XRAM[63099] = 8'b0;
    XRAM[63100] = 8'b0;
    XRAM[63101] = 8'b0;
    XRAM[63102] = 8'b0;
    XRAM[63103] = 8'b0;
    XRAM[63104] = 8'b0;
    XRAM[63105] = 8'b0;
    XRAM[63106] = 8'b0;
    XRAM[63107] = 8'b0;
    XRAM[63108] = 8'b0;
    XRAM[63109] = 8'b0;
    XRAM[63110] = 8'b0;
    XRAM[63111] = 8'b0;
    XRAM[63112] = 8'b0;
    XRAM[63113] = 8'b0;
    XRAM[63114] = 8'b0;
    XRAM[63115] = 8'b0;
    XRAM[63116] = 8'b0;
    XRAM[63117] = 8'b0;
    XRAM[63118] = 8'b0;
    XRAM[63119] = 8'b0;
    XRAM[63120] = 8'b0;
    XRAM[63121] = 8'b0;
    XRAM[63122] = 8'b0;
    XRAM[63123] = 8'b0;
    XRAM[63124] = 8'b0;
    XRAM[63125] = 8'b0;
    XRAM[63126] = 8'b0;
    XRAM[63127] = 8'b0;
    XRAM[63128] = 8'b0;
    XRAM[63129] = 8'b0;
    XRAM[63130] = 8'b0;
    XRAM[63131] = 8'b0;
    XRAM[63132] = 8'b0;
    XRAM[63133] = 8'b0;
    XRAM[63134] = 8'b0;
    XRAM[63135] = 8'b0;
    XRAM[63136] = 8'b0;
    XRAM[63137] = 8'b0;
    XRAM[63138] = 8'b0;
    XRAM[63139] = 8'b0;
    XRAM[63140] = 8'b0;
    XRAM[63141] = 8'b0;
    XRAM[63142] = 8'b0;
    XRAM[63143] = 8'b0;
    XRAM[63144] = 8'b0;
    XRAM[63145] = 8'b0;
    XRAM[63146] = 8'b0;
    XRAM[63147] = 8'b0;
    XRAM[63148] = 8'b0;
    XRAM[63149] = 8'b0;
    XRAM[63150] = 8'b0;
    XRAM[63151] = 8'b0;
    XRAM[63152] = 8'b0;
    XRAM[63153] = 8'b0;
    XRAM[63154] = 8'b0;
    XRAM[63155] = 8'b0;
    XRAM[63156] = 8'b0;
    XRAM[63157] = 8'b0;
    XRAM[63158] = 8'b0;
    XRAM[63159] = 8'b0;
    XRAM[63160] = 8'b0;
    XRAM[63161] = 8'b0;
    XRAM[63162] = 8'b0;
    XRAM[63163] = 8'b0;
    XRAM[63164] = 8'b0;
    XRAM[63165] = 8'b0;
    XRAM[63166] = 8'b0;
    XRAM[63167] = 8'b0;
    XRAM[63168] = 8'b0;
    XRAM[63169] = 8'b0;
    XRAM[63170] = 8'b0;
    XRAM[63171] = 8'b0;
    XRAM[63172] = 8'b0;
    XRAM[63173] = 8'b0;
    XRAM[63174] = 8'b0;
    XRAM[63175] = 8'b0;
    XRAM[63176] = 8'b0;
    XRAM[63177] = 8'b0;
    XRAM[63178] = 8'b0;
    XRAM[63179] = 8'b0;
    XRAM[63180] = 8'b0;
    XRAM[63181] = 8'b0;
    XRAM[63182] = 8'b0;
    XRAM[63183] = 8'b0;
    XRAM[63184] = 8'b0;
    XRAM[63185] = 8'b0;
    XRAM[63186] = 8'b0;
    XRAM[63187] = 8'b0;
    XRAM[63188] = 8'b0;
    XRAM[63189] = 8'b0;
    XRAM[63190] = 8'b0;
    XRAM[63191] = 8'b0;
    XRAM[63192] = 8'b0;
    XRAM[63193] = 8'b0;
    XRAM[63194] = 8'b0;
    XRAM[63195] = 8'b0;
    XRAM[63196] = 8'b0;
    XRAM[63197] = 8'b0;
    XRAM[63198] = 8'b0;
    XRAM[63199] = 8'b0;
    XRAM[63200] = 8'b0;
    XRAM[63201] = 8'b0;
    XRAM[63202] = 8'b0;
    XRAM[63203] = 8'b0;
    XRAM[63204] = 8'b0;
    XRAM[63205] = 8'b0;
    XRAM[63206] = 8'b0;
    XRAM[63207] = 8'b0;
    XRAM[63208] = 8'b0;
    XRAM[63209] = 8'b0;
    XRAM[63210] = 8'b0;
    XRAM[63211] = 8'b0;
    XRAM[63212] = 8'b0;
    XRAM[63213] = 8'b0;
    XRAM[63214] = 8'b0;
    XRAM[63215] = 8'b0;
    XRAM[63216] = 8'b0;
    XRAM[63217] = 8'b0;
    XRAM[63218] = 8'b0;
    XRAM[63219] = 8'b0;
    XRAM[63220] = 8'b0;
    XRAM[63221] = 8'b0;
    XRAM[63222] = 8'b0;
    XRAM[63223] = 8'b0;
    XRAM[63224] = 8'b0;
    XRAM[63225] = 8'b0;
    XRAM[63226] = 8'b0;
    XRAM[63227] = 8'b0;
    XRAM[63228] = 8'b0;
    XRAM[63229] = 8'b0;
    XRAM[63230] = 8'b0;
    XRAM[63231] = 8'b0;
    XRAM[63232] = 8'b0;
    XRAM[63233] = 8'b0;
    XRAM[63234] = 8'b0;
    XRAM[63235] = 8'b0;
    XRAM[63236] = 8'b0;
    XRAM[63237] = 8'b0;
    XRAM[63238] = 8'b0;
    XRAM[63239] = 8'b0;
    XRAM[63240] = 8'b0;
    XRAM[63241] = 8'b0;
    XRAM[63242] = 8'b0;
    XRAM[63243] = 8'b0;
    XRAM[63244] = 8'b0;
    XRAM[63245] = 8'b0;
    XRAM[63246] = 8'b0;
    XRAM[63247] = 8'b0;
    XRAM[63248] = 8'b0;
    XRAM[63249] = 8'b0;
    XRAM[63250] = 8'b0;
    XRAM[63251] = 8'b0;
    XRAM[63252] = 8'b0;
    XRAM[63253] = 8'b0;
    XRAM[63254] = 8'b0;
    XRAM[63255] = 8'b0;
    XRAM[63256] = 8'b0;
    XRAM[63257] = 8'b0;
    XRAM[63258] = 8'b0;
    XRAM[63259] = 8'b0;
    XRAM[63260] = 8'b0;
    XRAM[63261] = 8'b0;
    XRAM[63262] = 8'b0;
    XRAM[63263] = 8'b0;
    XRAM[63264] = 8'b0;
    XRAM[63265] = 8'b0;
    XRAM[63266] = 8'b0;
    XRAM[63267] = 8'b0;
    XRAM[63268] = 8'b0;
    XRAM[63269] = 8'b0;
    XRAM[63270] = 8'b0;
    XRAM[63271] = 8'b0;
    XRAM[63272] = 8'b0;
    XRAM[63273] = 8'b0;
    XRAM[63274] = 8'b0;
    XRAM[63275] = 8'b0;
    XRAM[63276] = 8'b0;
    XRAM[63277] = 8'b0;
    XRAM[63278] = 8'b0;
    XRAM[63279] = 8'b0;
    XRAM[63280] = 8'b0;
    XRAM[63281] = 8'b0;
    XRAM[63282] = 8'b0;
    XRAM[63283] = 8'b0;
    XRAM[63284] = 8'b0;
    XRAM[63285] = 8'b0;
    XRAM[63286] = 8'b0;
    XRAM[63287] = 8'b0;
    XRAM[63288] = 8'b0;
    XRAM[63289] = 8'b0;
    XRAM[63290] = 8'b0;
    XRAM[63291] = 8'b0;
    XRAM[63292] = 8'b0;
    XRAM[63293] = 8'b0;
    XRAM[63294] = 8'b0;
    XRAM[63295] = 8'b0;
    XRAM[63296] = 8'b0;
    XRAM[63297] = 8'b0;
    XRAM[63298] = 8'b0;
    XRAM[63299] = 8'b0;
    XRAM[63300] = 8'b0;
    XRAM[63301] = 8'b0;
    XRAM[63302] = 8'b0;
    XRAM[63303] = 8'b0;
    XRAM[63304] = 8'b0;
    XRAM[63305] = 8'b0;
    XRAM[63306] = 8'b0;
    XRAM[63307] = 8'b0;
    XRAM[63308] = 8'b0;
    XRAM[63309] = 8'b0;
    XRAM[63310] = 8'b0;
    XRAM[63311] = 8'b0;
    XRAM[63312] = 8'b0;
    XRAM[63313] = 8'b0;
    XRAM[63314] = 8'b0;
    XRAM[63315] = 8'b0;
    XRAM[63316] = 8'b0;
    XRAM[63317] = 8'b0;
    XRAM[63318] = 8'b0;
    XRAM[63319] = 8'b0;
    XRAM[63320] = 8'b0;
    XRAM[63321] = 8'b0;
    XRAM[63322] = 8'b0;
    XRAM[63323] = 8'b0;
    XRAM[63324] = 8'b0;
    XRAM[63325] = 8'b0;
    XRAM[63326] = 8'b0;
    XRAM[63327] = 8'b0;
    XRAM[63328] = 8'b0;
    XRAM[63329] = 8'b0;
    XRAM[63330] = 8'b0;
    XRAM[63331] = 8'b0;
    XRAM[63332] = 8'b0;
    XRAM[63333] = 8'b0;
    XRAM[63334] = 8'b0;
    XRAM[63335] = 8'b0;
    XRAM[63336] = 8'b0;
    XRAM[63337] = 8'b0;
    XRAM[63338] = 8'b0;
    XRAM[63339] = 8'b0;
    XRAM[63340] = 8'b0;
    XRAM[63341] = 8'b0;
    XRAM[63342] = 8'b0;
    XRAM[63343] = 8'b0;
    XRAM[63344] = 8'b0;
    XRAM[63345] = 8'b0;
    XRAM[63346] = 8'b0;
    XRAM[63347] = 8'b0;
    XRAM[63348] = 8'b0;
    XRAM[63349] = 8'b0;
    XRAM[63350] = 8'b0;
    XRAM[63351] = 8'b0;
    XRAM[63352] = 8'b0;
    XRAM[63353] = 8'b0;
    XRAM[63354] = 8'b0;
    XRAM[63355] = 8'b0;
    XRAM[63356] = 8'b0;
    XRAM[63357] = 8'b0;
    XRAM[63358] = 8'b0;
    XRAM[63359] = 8'b0;
    XRAM[63360] = 8'b0;
    XRAM[63361] = 8'b0;
    XRAM[63362] = 8'b0;
    XRAM[63363] = 8'b0;
    XRAM[63364] = 8'b0;
    XRAM[63365] = 8'b0;
    XRAM[63366] = 8'b0;
    XRAM[63367] = 8'b0;
    XRAM[63368] = 8'b0;
    XRAM[63369] = 8'b0;
    XRAM[63370] = 8'b0;
    XRAM[63371] = 8'b0;
    XRAM[63372] = 8'b0;
    XRAM[63373] = 8'b0;
    XRAM[63374] = 8'b0;
    XRAM[63375] = 8'b0;
    XRAM[63376] = 8'b0;
    XRAM[63377] = 8'b0;
    XRAM[63378] = 8'b0;
    XRAM[63379] = 8'b0;
    XRAM[63380] = 8'b0;
    XRAM[63381] = 8'b0;
    XRAM[63382] = 8'b0;
    XRAM[63383] = 8'b0;
    XRAM[63384] = 8'b0;
    XRAM[63385] = 8'b0;
    XRAM[63386] = 8'b0;
    XRAM[63387] = 8'b0;
    XRAM[63388] = 8'b0;
    XRAM[63389] = 8'b0;
    XRAM[63390] = 8'b0;
    XRAM[63391] = 8'b0;
    XRAM[63392] = 8'b0;
    XRAM[63393] = 8'b0;
    XRAM[63394] = 8'b0;
    XRAM[63395] = 8'b0;
    XRAM[63396] = 8'b0;
    XRAM[63397] = 8'b0;
    XRAM[63398] = 8'b0;
    XRAM[63399] = 8'b0;
    XRAM[63400] = 8'b0;
    XRAM[63401] = 8'b0;
    XRAM[63402] = 8'b0;
    XRAM[63403] = 8'b0;
    XRAM[63404] = 8'b0;
    XRAM[63405] = 8'b0;
    XRAM[63406] = 8'b0;
    XRAM[63407] = 8'b0;
    XRAM[63408] = 8'b0;
    XRAM[63409] = 8'b0;
    XRAM[63410] = 8'b0;
    XRAM[63411] = 8'b0;
    XRAM[63412] = 8'b0;
    XRAM[63413] = 8'b0;
    XRAM[63414] = 8'b0;
    XRAM[63415] = 8'b0;
    XRAM[63416] = 8'b0;
    XRAM[63417] = 8'b0;
    XRAM[63418] = 8'b0;
    XRAM[63419] = 8'b0;
    XRAM[63420] = 8'b0;
    XRAM[63421] = 8'b0;
    XRAM[63422] = 8'b0;
    XRAM[63423] = 8'b0;
    XRAM[63424] = 8'b0;
    XRAM[63425] = 8'b0;
    XRAM[63426] = 8'b0;
    XRAM[63427] = 8'b0;
    XRAM[63428] = 8'b0;
    XRAM[63429] = 8'b0;
    XRAM[63430] = 8'b0;
    XRAM[63431] = 8'b0;
    XRAM[63432] = 8'b0;
    XRAM[63433] = 8'b0;
    XRAM[63434] = 8'b0;
    XRAM[63435] = 8'b0;
    XRAM[63436] = 8'b0;
    XRAM[63437] = 8'b0;
    XRAM[63438] = 8'b0;
    XRAM[63439] = 8'b0;
    XRAM[63440] = 8'b0;
    XRAM[63441] = 8'b0;
    XRAM[63442] = 8'b0;
    XRAM[63443] = 8'b0;
    XRAM[63444] = 8'b0;
    XRAM[63445] = 8'b0;
    XRAM[63446] = 8'b0;
    XRAM[63447] = 8'b0;
    XRAM[63448] = 8'b0;
    XRAM[63449] = 8'b0;
    XRAM[63450] = 8'b0;
    XRAM[63451] = 8'b0;
    XRAM[63452] = 8'b0;
    XRAM[63453] = 8'b0;
    XRAM[63454] = 8'b0;
    XRAM[63455] = 8'b0;
    XRAM[63456] = 8'b0;
    XRAM[63457] = 8'b0;
    XRAM[63458] = 8'b0;
    XRAM[63459] = 8'b0;
    XRAM[63460] = 8'b0;
    XRAM[63461] = 8'b0;
    XRAM[63462] = 8'b0;
    XRAM[63463] = 8'b0;
    XRAM[63464] = 8'b0;
    XRAM[63465] = 8'b0;
    XRAM[63466] = 8'b0;
    XRAM[63467] = 8'b0;
    XRAM[63468] = 8'b0;
    XRAM[63469] = 8'b0;
    XRAM[63470] = 8'b0;
    XRAM[63471] = 8'b0;
    XRAM[63472] = 8'b0;
    XRAM[63473] = 8'b0;
    XRAM[63474] = 8'b0;
    XRAM[63475] = 8'b0;
    XRAM[63476] = 8'b0;
    XRAM[63477] = 8'b0;
    XRAM[63478] = 8'b0;
    XRAM[63479] = 8'b0;
    XRAM[63480] = 8'b0;
    XRAM[63481] = 8'b0;
    XRAM[63482] = 8'b0;
    XRAM[63483] = 8'b0;
    XRAM[63484] = 8'b0;
    XRAM[63485] = 8'b0;
    XRAM[63486] = 8'b0;
    XRAM[63487] = 8'b0;
    XRAM[63488] = 8'b0;
    XRAM[63489] = 8'b0;
    XRAM[63490] = 8'b0;
    XRAM[63491] = 8'b0;
    XRAM[63492] = 8'b0;
    XRAM[63493] = 8'b0;
    XRAM[63494] = 8'b0;
    XRAM[63495] = 8'b0;
    XRAM[63496] = 8'b0;
    XRAM[63497] = 8'b0;
    XRAM[63498] = 8'b0;
    XRAM[63499] = 8'b0;
    XRAM[63500] = 8'b0;
    XRAM[63501] = 8'b0;
    XRAM[63502] = 8'b0;
    XRAM[63503] = 8'b0;
    XRAM[63504] = 8'b0;
    XRAM[63505] = 8'b0;
    XRAM[63506] = 8'b0;
    XRAM[63507] = 8'b0;
    XRAM[63508] = 8'b0;
    XRAM[63509] = 8'b0;
    XRAM[63510] = 8'b0;
    XRAM[63511] = 8'b0;
    XRAM[63512] = 8'b0;
    XRAM[63513] = 8'b0;
    XRAM[63514] = 8'b0;
    XRAM[63515] = 8'b0;
    XRAM[63516] = 8'b0;
    XRAM[63517] = 8'b0;
    XRAM[63518] = 8'b0;
    XRAM[63519] = 8'b0;
    XRAM[63520] = 8'b0;
    XRAM[63521] = 8'b0;
    XRAM[63522] = 8'b0;
    XRAM[63523] = 8'b0;
    XRAM[63524] = 8'b0;
    XRAM[63525] = 8'b0;
    XRAM[63526] = 8'b0;
    XRAM[63527] = 8'b0;
    XRAM[63528] = 8'b0;
    XRAM[63529] = 8'b0;
    XRAM[63530] = 8'b0;
    XRAM[63531] = 8'b0;
    XRAM[63532] = 8'b0;
    XRAM[63533] = 8'b0;
    XRAM[63534] = 8'b0;
    XRAM[63535] = 8'b0;
    XRAM[63536] = 8'b0;
    XRAM[63537] = 8'b0;
    XRAM[63538] = 8'b0;
    XRAM[63539] = 8'b0;
    XRAM[63540] = 8'b0;
    XRAM[63541] = 8'b0;
    XRAM[63542] = 8'b0;
    XRAM[63543] = 8'b0;
    XRAM[63544] = 8'b0;
    XRAM[63545] = 8'b0;
    XRAM[63546] = 8'b0;
    XRAM[63547] = 8'b0;
    XRAM[63548] = 8'b0;
    XRAM[63549] = 8'b0;
    XRAM[63550] = 8'b0;
    XRAM[63551] = 8'b0;
    XRAM[63552] = 8'b0;
    XRAM[63553] = 8'b0;
    XRAM[63554] = 8'b0;
    XRAM[63555] = 8'b0;
    XRAM[63556] = 8'b0;
    XRAM[63557] = 8'b0;
    XRAM[63558] = 8'b0;
    XRAM[63559] = 8'b0;
    XRAM[63560] = 8'b0;
    XRAM[63561] = 8'b0;
    XRAM[63562] = 8'b0;
    XRAM[63563] = 8'b0;
    XRAM[63564] = 8'b0;
    XRAM[63565] = 8'b0;
    XRAM[63566] = 8'b0;
    XRAM[63567] = 8'b0;
    XRAM[63568] = 8'b0;
    XRAM[63569] = 8'b0;
    XRAM[63570] = 8'b0;
    XRAM[63571] = 8'b0;
    XRAM[63572] = 8'b0;
    XRAM[63573] = 8'b0;
    XRAM[63574] = 8'b0;
    XRAM[63575] = 8'b0;
    XRAM[63576] = 8'b0;
    XRAM[63577] = 8'b0;
    XRAM[63578] = 8'b0;
    XRAM[63579] = 8'b0;
    XRAM[63580] = 8'b0;
    XRAM[63581] = 8'b0;
    XRAM[63582] = 8'b0;
    XRAM[63583] = 8'b0;
    XRAM[63584] = 8'b0;
    XRAM[63585] = 8'b0;
    XRAM[63586] = 8'b0;
    XRAM[63587] = 8'b0;
    XRAM[63588] = 8'b0;
    XRAM[63589] = 8'b0;
    XRAM[63590] = 8'b0;
    XRAM[63591] = 8'b0;
    XRAM[63592] = 8'b0;
    XRAM[63593] = 8'b0;
    XRAM[63594] = 8'b0;
    XRAM[63595] = 8'b0;
    XRAM[63596] = 8'b0;
    XRAM[63597] = 8'b0;
    XRAM[63598] = 8'b0;
    XRAM[63599] = 8'b0;
    XRAM[63600] = 8'b0;
    XRAM[63601] = 8'b0;
    XRAM[63602] = 8'b0;
    XRAM[63603] = 8'b0;
    XRAM[63604] = 8'b0;
    XRAM[63605] = 8'b0;
    XRAM[63606] = 8'b0;
    XRAM[63607] = 8'b0;
    XRAM[63608] = 8'b0;
    XRAM[63609] = 8'b0;
    XRAM[63610] = 8'b0;
    XRAM[63611] = 8'b0;
    XRAM[63612] = 8'b0;
    XRAM[63613] = 8'b0;
    XRAM[63614] = 8'b0;
    XRAM[63615] = 8'b0;
    XRAM[63616] = 8'b0;
    XRAM[63617] = 8'b0;
    XRAM[63618] = 8'b0;
    XRAM[63619] = 8'b0;
    XRAM[63620] = 8'b0;
    XRAM[63621] = 8'b0;
    XRAM[63622] = 8'b0;
    XRAM[63623] = 8'b0;
    XRAM[63624] = 8'b0;
    XRAM[63625] = 8'b0;
    XRAM[63626] = 8'b0;
    XRAM[63627] = 8'b0;
    XRAM[63628] = 8'b0;
    XRAM[63629] = 8'b0;
    XRAM[63630] = 8'b0;
    XRAM[63631] = 8'b0;
    XRAM[63632] = 8'b0;
    XRAM[63633] = 8'b0;
    XRAM[63634] = 8'b0;
    XRAM[63635] = 8'b0;
    XRAM[63636] = 8'b0;
    XRAM[63637] = 8'b0;
    XRAM[63638] = 8'b0;
    XRAM[63639] = 8'b0;
    XRAM[63640] = 8'b0;
    XRAM[63641] = 8'b0;
    XRAM[63642] = 8'b0;
    XRAM[63643] = 8'b0;
    XRAM[63644] = 8'b0;
    XRAM[63645] = 8'b0;
    XRAM[63646] = 8'b0;
    XRAM[63647] = 8'b0;
    XRAM[63648] = 8'b0;
    XRAM[63649] = 8'b0;
    XRAM[63650] = 8'b0;
    XRAM[63651] = 8'b0;
    XRAM[63652] = 8'b0;
    XRAM[63653] = 8'b0;
    XRAM[63654] = 8'b0;
    XRAM[63655] = 8'b0;
    XRAM[63656] = 8'b0;
    XRAM[63657] = 8'b0;
    XRAM[63658] = 8'b0;
    XRAM[63659] = 8'b0;
    XRAM[63660] = 8'b0;
    XRAM[63661] = 8'b0;
    XRAM[63662] = 8'b0;
    XRAM[63663] = 8'b0;
    XRAM[63664] = 8'b0;
    XRAM[63665] = 8'b0;
    XRAM[63666] = 8'b0;
    XRAM[63667] = 8'b0;
    XRAM[63668] = 8'b0;
    XRAM[63669] = 8'b0;
    XRAM[63670] = 8'b0;
    XRAM[63671] = 8'b0;
    XRAM[63672] = 8'b0;
    XRAM[63673] = 8'b0;
    XRAM[63674] = 8'b0;
    XRAM[63675] = 8'b0;
    XRAM[63676] = 8'b0;
    XRAM[63677] = 8'b0;
    XRAM[63678] = 8'b0;
    XRAM[63679] = 8'b0;
    XRAM[63680] = 8'b0;
    XRAM[63681] = 8'b0;
    XRAM[63682] = 8'b0;
    XRAM[63683] = 8'b0;
    XRAM[63684] = 8'b0;
    XRAM[63685] = 8'b0;
    XRAM[63686] = 8'b0;
    XRAM[63687] = 8'b0;
    XRAM[63688] = 8'b0;
    XRAM[63689] = 8'b0;
    XRAM[63690] = 8'b0;
    XRAM[63691] = 8'b0;
    XRAM[63692] = 8'b0;
    XRAM[63693] = 8'b0;
    XRAM[63694] = 8'b0;
    XRAM[63695] = 8'b0;
    XRAM[63696] = 8'b0;
    XRAM[63697] = 8'b0;
    XRAM[63698] = 8'b0;
    XRAM[63699] = 8'b0;
    XRAM[63700] = 8'b0;
    XRAM[63701] = 8'b0;
    XRAM[63702] = 8'b0;
    XRAM[63703] = 8'b0;
    XRAM[63704] = 8'b0;
    XRAM[63705] = 8'b0;
    XRAM[63706] = 8'b0;
    XRAM[63707] = 8'b0;
    XRAM[63708] = 8'b0;
    XRAM[63709] = 8'b0;
    XRAM[63710] = 8'b0;
    XRAM[63711] = 8'b0;
    XRAM[63712] = 8'b0;
    XRAM[63713] = 8'b0;
    XRAM[63714] = 8'b0;
    XRAM[63715] = 8'b0;
    XRAM[63716] = 8'b0;
    XRAM[63717] = 8'b0;
    XRAM[63718] = 8'b0;
    XRAM[63719] = 8'b0;
    XRAM[63720] = 8'b0;
    XRAM[63721] = 8'b0;
    XRAM[63722] = 8'b0;
    XRAM[63723] = 8'b0;
    XRAM[63724] = 8'b0;
    XRAM[63725] = 8'b0;
    XRAM[63726] = 8'b0;
    XRAM[63727] = 8'b0;
    XRAM[63728] = 8'b0;
    XRAM[63729] = 8'b0;
    XRAM[63730] = 8'b0;
    XRAM[63731] = 8'b0;
    XRAM[63732] = 8'b0;
    XRAM[63733] = 8'b0;
    XRAM[63734] = 8'b0;
    XRAM[63735] = 8'b0;
    XRAM[63736] = 8'b0;
    XRAM[63737] = 8'b0;
    XRAM[63738] = 8'b0;
    XRAM[63739] = 8'b0;
    XRAM[63740] = 8'b0;
    XRAM[63741] = 8'b0;
    XRAM[63742] = 8'b0;
    XRAM[63743] = 8'b0;
    XRAM[63744] = 8'b0;
    XRAM[63745] = 8'b0;
    XRAM[63746] = 8'b0;
    XRAM[63747] = 8'b0;
    XRAM[63748] = 8'b0;
    XRAM[63749] = 8'b0;
    XRAM[63750] = 8'b0;
    XRAM[63751] = 8'b0;
    XRAM[63752] = 8'b0;
    XRAM[63753] = 8'b0;
    XRAM[63754] = 8'b0;
    XRAM[63755] = 8'b0;
    XRAM[63756] = 8'b0;
    XRAM[63757] = 8'b0;
    XRAM[63758] = 8'b0;
    XRAM[63759] = 8'b0;
    XRAM[63760] = 8'b0;
    XRAM[63761] = 8'b0;
    XRAM[63762] = 8'b0;
    XRAM[63763] = 8'b0;
    XRAM[63764] = 8'b0;
    XRAM[63765] = 8'b0;
    XRAM[63766] = 8'b0;
    XRAM[63767] = 8'b0;
    XRAM[63768] = 8'b0;
    XRAM[63769] = 8'b0;
    XRAM[63770] = 8'b0;
    XRAM[63771] = 8'b0;
    XRAM[63772] = 8'b0;
    XRAM[63773] = 8'b0;
    XRAM[63774] = 8'b0;
    XRAM[63775] = 8'b0;
    XRAM[63776] = 8'b0;
    XRAM[63777] = 8'b0;
    XRAM[63778] = 8'b0;
    XRAM[63779] = 8'b0;
    XRAM[63780] = 8'b0;
    XRAM[63781] = 8'b0;
    XRAM[63782] = 8'b0;
    XRAM[63783] = 8'b0;
    XRAM[63784] = 8'b0;
    XRAM[63785] = 8'b0;
    XRAM[63786] = 8'b0;
    XRAM[63787] = 8'b0;
    XRAM[63788] = 8'b0;
    XRAM[63789] = 8'b0;
    XRAM[63790] = 8'b0;
    XRAM[63791] = 8'b0;
    XRAM[63792] = 8'b0;
    XRAM[63793] = 8'b0;
    XRAM[63794] = 8'b0;
    XRAM[63795] = 8'b0;
    XRAM[63796] = 8'b0;
    XRAM[63797] = 8'b0;
    XRAM[63798] = 8'b0;
    XRAM[63799] = 8'b0;
    XRAM[63800] = 8'b0;
    XRAM[63801] = 8'b0;
    XRAM[63802] = 8'b0;
    XRAM[63803] = 8'b0;
    XRAM[63804] = 8'b0;
    XRAM[63805] = 8'b0;
    XRAM[63806] = 8'b0;
    XRAM[63807] = 8'b0;
    XRAM[63808] = 8'b0;
    XRAM[63809] = 8'b0;
    XRAM[63810] = 8'b0;
    XRAM[63811] = 8'b0;
    XRAM[63812] = 8'b0;
    XRAM[63813] = 8'b0;
    XRAM[63814] = 8'b0;
    XRAM[63815] = 8'b0;
    XRAM[63816] = 8'b0;
    XRAM[63817] = 8'b0;
    XRAM[63818] = 8'b0;
    XRAM[63819] = 8'b0;
    XRAM[63820] = 8'b0;
    XRAM[63821] = 8'b0;
    XRAM[63822] = 8'b0;
    XRAM[63823] = 8'b0;
    XRAM[63824] = 8'b0;
    XRAM[63825] = 8'b0;
    XRAM[63826] = 8'b0;
    XRAM[63827] = 8'b0;
    XRAM[63828] = 8'b0;
    XRAM[63829] = 8'b0;
    XRAM[63830] = 8'b0;
    XRAM[63831] = 8'b0;
    XRAM[63832] = 8'b0;
    XRAM[63833] = 8'b0;
    XRAM[63834] = 8'b0;
    XRAM[63835] = 8'b0;
    XRAM[63836] = 8'b0;
    XRAM[63837] = 8'b0;
    XRAM[63838] = 8'b0;
    XRAM[63839] = 8'b0;
    XRAM[63840] = 8'b0;
    XRAM[63841] = 8'b0;
    XRAM[63842] = 8'b0;
    XRAM[63843] = 8'b0;
    XRAM[63844] = 8'b0;
    XRAM[63845] = 8'b0;
    XRAM[63846] = 8'b0;
    XRAM[63847] = 8'b0;
    XRAM[63848] = 8'b0;
    XRAM[63849] = 8'b0;
    XRAM[63850] = 8'b0;
    XRAM[63851] = 8'b0;
    XRAM[63852] = 8'b0;
    XRAM[63853] = 8'b0;
    XRAM[63854] = 8'b0;
    XRAM[63855] = 8'b0;
    XRAM[63856] = 8'b0;
    XRAM[63857] = 8'b0;
    XRAM[63858] = 8'b0;
    XRAM[63859] = 8'b0;
    XRAM[63860] = 8'b0;
    XRAM[63861] = 8'b0;
    XRAM[63862] = 8'b0;
    XRAM[63863] = 8'b0;
    XRAM[63864] = 8'b0;
    XRAM[63865] = 8'b0;
    XRAM[63866] = 8'b0;
    XRAM[63867] = 8'b0;
    XRAM[63868] = 8'b0;
    XRAM[63869] = 8'b0;
    XRAM[63870] = 8'b0;
    XRAM[63871] = 8'b0;
    XRAM[63872] = 8'b0;
    XRAM[63873] = 8'b0;
    XRAM[63874] = 8'b0;
    XRAM[63875] = 8'b0;
    XRAM[63876] = 8'b0;
    XRAM[63877] = 8'b0;
    XRAM[63878] = 8'b0;
    XRAM[63879] = 8'b0;
    XRAM[63880] = 8'b0;
    XRAM[63881] = 8'b0;
    XRAM[63882] = 8'b0;
    XRAM[63883] = 8'b0;
    XRAM[63884] = 8'b0;
    XRAM[63885] = 8'b0;
    XRAM[63886] = 8'b0;
    XRAM[63887] = 8'b0;
    XRAM[63888] = 8'b0;
    XRAM[63889] = 8'b0;
    XRAM[63890] = 8'b0;
    XRAM[63891] = 8'b0;
    XRAM[63892] = 8'b0;
    XRAM[63893] = 8'b0;
    XRAM[63894] = 8'b0;
    XRAM[63895] = 8'b0;
    XRAM[63896] = 8'b0;
    XRAM[63897] = 8'b0;
    XRAM[63898] = 8'b0;
    XRAM[63899] = 8'b0;
    XRAM[63900] = 8'b0;
    XRAM[63901] = 8'b0;
    XRAM[63902] = 8'b0;
    XRAM[63903] = 8'b0;
    XRAM[63904] = 8'b0;
    XRAM[63905] = 8'b0;
    XRAM[63906] = 8'b0;
    XRAM[63907] = 8'b0;
    XRAM[63908] = 8'b0;
    XRAM[63909] = 8'b0;
    XRAM[63910] = 8'b0;
    XRAM[63911] = 8'b0;
    XRAM[63912] = 8'b0;
    XRAM[63913] = 8'b0;
    XRAM[63914] = 8'b0;
    XRAM[63915] = 8'b0;
    XRAM[63916] = 8'b0;
    XRAM[63917] = 8'b0;
    XRAM[63918] = 8'b0;
    XRAM[63919] = 8'b0;
    XRAM[63920] = 8'b0;
    XRAM[63921] = 8'b0;
    XRAM[63922] = 8'b0;
    XRAM[63923] = 8'b0;
    XRAM[63924] = 8'b0;
    XRAM[63925] = 8'b0;
    XRAM[63926] = 8'b0;
    XRAM[63927] = 8'b0;
    XRAM[63928] = 8'b0;
    XRAM[63929] = 8'b0;
    XRAM[63930] = 8'b0;
    XRAM[63931] = 8'b0;
    XRAM[63932] = 8'b0;
    XRAM[63933] = 8'b0;
    XRAM[63934] = 8'b0;
    XRAM[63935] = 8'b0;
    XRAM[63936] = 8'b0;
    XRAM[63937] = 8'b0;
    XRAM[63938] = 8'b0;
    XRAM[63939] = 8'b0;
    XRAM[63940] = 8'b0;
    XRAM[63941] = 8'b0;
    XRAM[63942] = 8'b0;
    XRAM[63943] = 8'b0;
    XRAM[63944] = 8'b0;
    XRAM[63945] = 8'b0;
    XRAM[63946] = 8'b0;
    XRAM[63947] = 8'b0;
    XRAM[63948] = 8'b0;
    XRAM[63949] = 8'b0;
    XRAM[63950] = 8'b0;
    XRAM[63951] = 8'b0;
    XRAM[63952] = 8'b0;
    XRAM[63953] = 8'b0;
    XRAM[63954] = 8'b0;
    XRAM[63955] = 8'b0;
    XRAM[63956] = 8'b0;
    XRAM[63957] = 8'b0;
    XRAM[63958] = 8'b0;
    XRAM[63959] = 8'b0;
    XRAM[63960] = 8'b0;
    XRAM[63961] = 8'b0;
    XRAM[63962] = 8'b0;
    XRAM[63963] = 8'b0;
    XRAM[63964] = 8'b0;
    XRAM[63965] = 8'b0;
    XRAM[63966] = 8'b0;
    XRAM[63967] = 8'b0;
    XRAM[63968] = 8'b0;
    XRAM[63969] = 8'b0;
    XRAM[63970] = 8'b0;
    XRAM[63971] = 8'b0;
    XRAM[63972] = 8'b0;
    XRAM[63973] = 8'b0;
    XRAM[63974] = 8'b0;
    XRAM[63975] = 8'b0;
    XRAM[63976] = 8'b0;
    XRAM[63977] = 8'b0;
    XRAM[63978] = 8'b0;
    XRAM[63979] = 8'b0;
    XRAM[63980] = 8'b0;
    XRAM[63981] = 8'b0;
    XRAM[63982] = 8'b0;
    XRAM[63983] = 8'b0;
    XRAM[63984] = 8'b0;
    XRAM[63985] = 8'b0;
    XRAM[63986] = 8'b0;
    XRAM[63987] = 8'b0;
    XRAM[63988] = 8'b0;
    XRAM[63989] = 8'b0;
    XRAM[63990] = 8'b0;
    XRAM[63991] = 8'b0;
    XRAM[63992] = 8'b0;
    XRAM[63993] = 8'b0;
    XRAM[63994] = 8'b0;
    XRAM[63995] = 8'b0;
    XRAM[63996] = 8'b0;
    XRAM[63997] = 8'b0;
    XRAM[63998] = 8'b0;
    XRAM[63999] = 8'b0;
    XRAM[64000] = 8'b0;
    XRAM[64001] = 8'b0;
    XRAM[64002] = 8'b0;
    XRAM[64003] = 8'b0;
    XRAM[64004] = 8'b0;
    XRAM[64005] = 8'b0;
    XRAM[64006] = 8'b0;
    XRAM[64007] = 8'b0;
    XRAM[64008] = 8'b0;
    XRAM[64009] = 8'b0;
    XRAM[64010] = 8'b0;
    XRAM[64011] = 8'b0;
    XRAM[64012] = 8'b0;
    XRAM[64013] = 8'b0;
    XRAM[64014] = 8'b0;
    XRAM[64015] = 8'b0;
    XRAM[64016] = 8'b0;
    XRAM[64017] = 8'b0;
    XRAM[64018] = 8'b0;
    XRAM[64019] = 8'b0;
    XRAM[64020] = 8'b0;
    XRAM[64021] = 8'b0;
    XRAM[64022] = 8'b0;
    XRAM[64023] = 8'b0;
    XRAM[64024] = 8'b0;
    XRAM[64025] = 8'b0;
    XRAM[64026] = 8'b0;
    XRAM[64027] = 8'b0;
    XRAM[64028] = 8'b0;
    XRAM[64029] = 8'b0;
    XRAM[64030] = 8'b0;
    XRAM[64031] = 8'b0;
    XRAM[64032] = 8'b0;
    XRAM[64033] = 8'b0;
    XRAM[64034] = 8'b0;
    XRAM[64035] = 8'b0;
    XRAM[64036] = 8'b0;
    XRAM[64037] = 8'b0;
    XRAM[64038] = 8'b0;
    XRAM[64039] = 8'b0;
    XRAM[64040] = 8'b0;
    XRAM[64041] = 8'b0;
    XRAM[64042] = 8'b0;
    XRAM[64043] = 8'b0;
    XRAM[64044] = 8'b0;
    XRAM[64045] = 8'b0;
    XRAM[64046] = 8'b0;
    XRAM[64047] = 8'b0;
    XRAM[64048] = 8'b0;
    XRAM[64049] = 8'b0;
    XRAM[64050] = 8'b0;
    XRAM[64051] = 8'b0;
    XRAM[64052] = 8'b0;
    XRAM[64053] = 8'b0;
    XRAM[64054] = 8'b0;
    XRAM[64055] = 8'b0;
    XRAM[64056] = 8'b0;
    XRAM[64057] = 8'b0;
    XRAM[64058] = 8'b0;
    XRAM[64059] = 8'b0;
    XRAM[64060] = 8'b0;
    XRAM[64061] = 8'b0;
    XRAM[64062] = 8'b0;
    XRAM[64063] = 8'b0;
    XRAM[64064] = 8'b0;
    XRAM[64065] = 8'b0;
    XRAM[64066] = 8'b0;
    XRAM[64067] = 8'b0;
    XRAM[64068] = 8'b0;
    XRAM[64069] = 8'b0;
    XRAM[64070] = 8'b0;
    XRAM[64071] = 8'b0;
    XRAM[64072] = 8'b0;
    XRAM[64073] = 8'b0;
    XRAM[64074] = 8'b0;
    XRAM[64075] = 8'b0;
    XRAM[64076] = 8'b0;
    XRAM[64077] = 8'b0;
    XRAM[64078] = 8'b0;
    XRAM[64079] = 8'b0;
    XRAM[64080] = 8'b0;
    XRAM[64081] = 8'b0;
    XRAM[64082] = 8'b0;
    XRAM[64083] = 8'b0;
    XRAM[64084] = 8'b0;
    XRAM[64085] = 8'b0;
    XRAM[64086] = 8'b0;
    XRAM[64087] = 8'b0;
    XRAM[64088] = 8'b0;
    XRAM[64089] = 8'b0;
    XRAM[64090] = 8'b0;
    XRAM[64091] = 8'b0;
    XRAM[64092] = 8'b0;
    XRAM[64093] = 8'b0;
    XRAM[64094] = 8'b0;
    XRAM[64095] = 8'b0;
    XRAM[64096] = 8'b0;
    XRAM[64097] = 8'b0;
    XRAM[64098] = 8'b0;
    XRAM[64099] = 8'b0;
    XRAM[64100] = 8'b0;
    XRAM[64101] = 8'b0;
    XRAM[64102] = 8'b0;
    XRAM[64103] = 8'b0;
    XRAM[64104] = 8'b0;
    XRAM[64105] = 8'b0;
    XRAM[64106] = 8'b0;
    XRAM[64107] = 8'b0;
    XRAM[64108] = 8'b0;
    XRAM[64109] = 8'b0;
    XRAM[64110] = 8'b0;
    XRAM[64111] = 8'b0;
    XRAM[64112] = 8'b0;
    XRAM[64113] = 8'b0;
    XRAM[64114] = 8'b0;
    XRAM[64115] = 8'b0;
    XRAM[64116] = 8'b0;
    XRAM[64117] = 8'b0;
    XRAM[64118] = 8'b0;
    XRAM[64119] = 8'b0;
    XRAM[64120] = 8'b0;
    XRAM[64121] = 8'b0;
    XRAM[64122] = 8'b0;
    XRAM[64123] = 8'b0;
    XRAM[64124] = 8'b0;
    XRAM[64125] = 8'b0;
    XRAM[64126] = 8'b0;
    XRAM[64127] = 8'b0;
    XRAM[64128] = 8'b0;
    XRAM[64129] = 8'b0;
    XRAM[64130] = 8'b0;
    XRAM[64131] = 8'b0;
    XRAM[64132] = 8'b0;
    XRAM[64133] = 8'b0;
    XRAM[64134] = 8'b0;
    XRAM[64135] = 8'b0;
    XRAM[64136] = 8'b0;
    XRAM[64137] = 8'b0;
    XRAM[64138] = 8'b0;
    XRAM[64139] = 8'b0;
    XRAM[64140] = 8'b0;
    XRAM[64141] = 8'b0;
    XRAM[64142] = 8'b0;
    XRAM[64143] = 8'b0;
    XRAM[64144] = 8'b0;
    XRAM[64145] = 8'b0;
    XRAM[64146] = 8'b0;
    XRAM[64147] = 8'b0;
    XRAM[64148] = 8'b0;
    XRAM[64149] = 8'b0;
    XRAM[64150] = 8'b0;
    XRAM[64151] = 8'b0;
    XRAM[64152] = 8'b0;
    XRAM[64153] = 8'b0;
    XRAM[64154] = 8'b0;
    XRAM[64155] = 8'b0;
    XRAM[64156] = 8'b0;
    XRAM[64157] = 8'b0;
    XRAM[64158] = 8'b0;
    XRAM[64159] = 8'b0;
    XRAM[64160] = 8'b0;
    XRAM[64161] = 8'b0;
    XRAM[64162] = 8'b0;
    XRAM[64163] = 8'b0;
    XRAM[64164] = 8'b0;
    XRAM[64165] = 8'b0;
    XRAM[64166] = 8'b0;
    XRAM[64167] = 8'b0;
    XRAM[64168] = 8'b0;
    XRAM[64169] = 8'b0;
    XRAM[64170] = 8'b0;
    XRAM[64171] = 8'b0;
    XRAM[64172] = 8'b0;
    XRAM[64173] = 8'b0;
    XRAM[64174] = 8'b0;
    XRAM[64175] = 8'b0;
    XRAM[64176] = 8'b0;
    XRAM[64177] = 8'b0;
    XRAM[64178] = 8'b0;
    XRAM[64179] = 8'b0;
    XRAM[64180] = 8'b0;
    XRAM[64181] = 8'b0;
    XRAM[64182] = 8'b0;
    XRAM[64183] = 8'b0;
    XRAM[64184] = 8'b0;
    XRAM[64185] = 8'b0;
    XRAM[64186] = 8'b0;
    XRAM[64187] = 8'b0;
    XRAM[64188] = 8'b0;
    XRAM[64189] = 8'b0;
    XRAM[64190] = 8'b0;
    XRAM[64191] = 8'b0;
    XRAM[64192] = 8'b0;
    XRAM[64193] = 8'b0;
    XRAM[64194] = 8'b0;
    XRAM[64195] = 8'b0;
    XRAM[64196] = 8'b0;
    XRAM[64197] = 8'b0;
    XRAM[64198] = 8'b0;
    XRAM[64199] = 8'b0;
    XRAM[64200] = 8'b0;
    XRAM[64201] = 8'b0;
    XRAM[64202] = 8'b0;
    XRAM[64203] = 8'b0;
    XRAM[64204] = 8'b0;
    XRAM[64205] = 8'b0;
    XRAM[64206] = 8'b0;
    XRAM[64207] = 8'b0;
    XRAM[64208] = 8'b0;
    XRAM[64209] = 8'b0;
    XRAM[64210] = 8'b0;
    XRAM[64211] = 8'b0;
    XRAM[64212] = 8'b0;
    XRAM[64213] = 8'b0;
    XRAM[64214] = 8'b0;
    XRAM[64215] = 8'b0;
    XRAM[64216] = 8'b0;
    XRAM[64217] = 8'b0;
    XRAM[64218] = 8'b0;
    XRAM[64219] = 8'b0;
    XRAM[64220] = 8'b0;
    XRAM[64221] = 8'b0;
    XRAM[64222] = 8'b0;
    XRAM[64223] = 8'b0;
    XRAM[64224] = 8'b0;
    XRAM[64225] = 8'b0;
    XRAM[64226] = 8'b0;
    XRAM[64227] = 8'b0;
    XRAM[64228] = 8'b0;
    XRAM[64229] = 8'b0;
    XRAM[64230] = 8'b0;
    XRAM[64231] = 8'b0;
    XRAM[64232] = 8'b0;
    XRAM[64233] = 8'b0;
    XRAM[64234] = 8'b0;
    XRAM[64235] = 8'b0;
    XRAM[64236] = 8'b0;
    XRAM[64237] = 8'b0;
    XRAM[64238] = 8'b0;
    XRAM[64239] = 8'b0;
    XRAM[64240] = 8'b0;
    XRAM[64241] = 8'b0;
    XRAM[64242] = 8'b0;
    XRAM[64243] = 8'b0;
    XRAM[64244] = 8'b0;
    XRAM[64245] = 8'b0;
    XRAM[64246] = 8'b0;
    XRAM[64247] = 8'b0;
    XRAM[64248] = 8'b0;
    XRAM[64249] = 8'b0;
    XRAM[64250] = 8'b0;
    XRAM[64251] = 8'b0;
    XRAM[64252] = 8'b0;
    XRAM[64253] = 8'b0;
    XRAM[64254] = 8'b0;
    XRAM[64255] = 8'b0;
    XRAM[64256] = 8'b0;
    XRAM[64257] = 8'b0;
    XRAM[64258] = 8'b0;
    XRAM[64259] = 8'b0;
    XRAM[64260] = 8'b0;
    XRAM[64261] = 8'b0;
    XRAM[64262] = 8'b0;
    XRAM[64263] = 8'b0;
    XRAM[64264] = 8'b0;
    XRAM[64265] = 8'b0;
    XRAM[64266] = 8'b0;
    XRAM[64267] = 8'b0;
    XRAM[64268] = 8'b0;
    XRAM[64269] = 8'b0;
    XRAM[64270] = 8'b0;
    XRAM[64271] = 8'b0;
    XRAM[64272] = 8'b0;
    XRAM[64273] = 8'b0;
    XRAM[64274] = 8'b0;
    XRAM[64275] = 8'b0;
    XRAM[64276] = 8'b0;
    XRAM[64277] = 8'b0;
    XRAM[64278] = 8'b0;
    XRAM[64279] = 8'b0;
    XRAM[64280] = 8'b0;
    XRAM[64281] = 8'b0;
    XRAM[64282] = 8'b0;
    XRAM[64283] = 8'b0;
    XRAM[64284] = 8'b0;
    XRAM[64285] = 8'b0;
    XRAM[64286] = 8'b0;
    XRAM[64287] = 8'b0;
    XRAM[64288] = 8'b0;
    XRAM[64289] = 8'b0;
    XRAM[64290] = 8'b0;
    XRAM[64291] = 8'b0;
    XRAM[64292] = 8'b0;
    XRAM[64293] = 8'b0;
    XRAM[64294] = 8'b0;
    XRAM[64295] = 8'b0;
    XRAM[64296] = 8'b0;
    XRAM[64297] = 8'b0;
    XRAM[64298] = 8'b0;
    XRAM[64299] = 8'b0;
    XRAM[64300] = 8'b0;
    XRAM[64301] = 8'b0;
    XRAM[64302] = 8'b0;
    XRAM[64303] = 8'b0;
    XRAM[64304] = 8'b0;
    XRAM[64305] = 8'b0;
    XRAM[64306] = 8'b0;
    XRAM[64307] = 8'b0;
    XRAM[64308] = 8'b0;
    XRAM[64309] = 8'b0;
    XRAM[64310] = 8'b0;
    XRAM[64311] = 8'b0;
    XRAM[64312] = 8'b0;
    XRAM[64313] = 8'b0;
    XRAM[64314] = 8'b0;
    XRAM[64315] = 8'b0;
    XRAM[64316] = 8'b0;
    XRAM[64317] = 8'b0;
    XRAM[64318] = 8'b0;
    XRAM[64319] = 8'b0;
    XRAM[64320] = 8'b0;
    XRAM[64321] = 8'b0;
    XRAM[64322] = 8'b0;
    XRAM[64323] = 8'b0;
    XRAM[64324] = 8'b0;
    XRAM[64325] = 8'b0;
    XRAM[64326] = 8'b0;
    XRAM[64327] = 8'b0;
    XRAM[64328] = 8'b0;
    XRAM[64329] = 8'b0;
    XRAM[64330] = 8'b0;
    XRAM[64331] = 8'b0;
    XRAM[64332] = 8'b0;
    XRAM[64333] = 8'b0;
    XRAM[64334] = 8'b0;
    XRAM[64335] = 8'b0;
    XRAM[64336] = 8'b0;
    XRAM[64337] = 8'b0;
    XRAM[64338] = 8'b0;
    XRAM[64339] = 8'b0;
    XRAM[64340] = 8'b0;
    XRAM[64341] = 8'b0;
    XRAM[64342] = 8'b0;
    XRAM[64343] = 8'b0;
    XRAM[64344] = 8'b0;
    XRAM[64345] = 8'b0;
    XRAM[64346] = 8'b0;
    XRAM[64347] = 8'b0;
    XRAM[64348] = 8'b0;
    XRAM[64349] = 8'b0;
    XRAM[64350] = 8'b0;
    XRAM[64351] = 8'b0;
    XRAM[64352] = 8'b0;
    XRAM[64353] = 8'b0;
    XRAM[64354] = 8'b0;
    XRAM[64355] = 8'b0;
    XRAM[64356] = 8'b0;
    XRAM[64357] = 8'b0;
    XRAM[64358] = 8'b0;
    XRAM[64359] = 8'b0;
    XRAM[64360] = 8'b0;
    XRAM[64361] = 8'b0;
    XRAM[64362] = 8'b0;
    XRAM[64363] = 8'b0;
    XRAM[64364] = 8'b0;
    XRAM[64365] = 8'b0;
    XRAM[64366] = 8'b0;
    XRAM[64367] = 8'b0;
    XRAM[64368] = 8'b0;
    XRAM[64369] = 8'b0;
    XRAM[64370] = 8'b0;
    XRAM[64371] = 8'b0;
    XRAM[64372] = 8'b0;
    XRAM[64373] = 8'b0;
    XRAM[64374] = 8'b0;
    XRAM[64375] = 8'b0;
    XRAM[64376] = 8'b0;
    XRAM[64377] = 8'b0;
    XRAM[64378] = 8'b0;
    XRAM[64379] = 8'b0;
    XRAM[64380] = 8'b0;
    XRAM[64381] = 8'b0;
    XRAM[64382] = 8'b0;
    XRAM[64383] = 8'b0;
    XRAM[64384] = 8'b0;
    XRAM[64385] = 8'b0;
    XRAM[64386] = 8'b0;
    XRAM[64387] = 8'b0;
    XRAM[64388] = 8'b0;
    XRAM[64389] = 8'b0;
    XRAM[64390] = 8'b0;
    XRAM[64391] = 8'b0;
    XRAM[64392] = 8'b0;
    XRAM[64393] = 8'b0;
    XRAM[64394] = 8'b0;
    XRAM[64395] = 8'b0;
    XRAM[64396] = 8'b0;
    XRAM[64397] = 8'b0;
    XRAM[64398] = 8'b0;
    XRAM[64399] = 8'b0;
    XRAM[64400] = 8'b0;
    XRAM[64401] = 8'b0;
    XRAM[64402] = 8'b0;
    XRAM[64403] = 8'b0;
    XRAM[64404] = 8'b0;
    XRAM[64405] = 8'b0;
    XRAM[64406] = 8'b0;
    XRAM[64407] = 8'b0;
    XRAM[64408] = 8'b0;
    XRAM[64409] = 8'b0;
    XRAM[64410] = 8'b0;
    XRAM[64411] = 8'b0;
    XRAM[64412] = 8'b0;
    XRAM[64413] = 8'b0;
    XRAM[64414] = 8'b0;
    XRAM[64415] = 8'b0;
    XRAM[64416] = 8'b0;
    XRAM[64417] = 8'b0;
    XRAM[64418] = 8'b0;
    XRAM[64419] = 8'b0;
    XRAM[64420] = 8'b0;
    XRAM[64421] = 8'b0;
    XRAM[64422] = 8'b0;
    XRAM[64423] = 8'b0;
    XRAM[64424] = 8'b0;
    XRAM[64425] = 8'b0;
    XRAM[64426] = 8'b0;
    XRAM[64427] = 8'b0;
    XRAM[64428] = 8'b0;
    XRAM[64429] = 8'b0;
    XRAM[64430] = 8'b0;
    XRAM[64431] = 8'b0;
    XRAM[64432] = 8'b0;
    XRAM[64433] = 8'b0;
    XRAM[64434] = 8'b0;
    XRAM[64435] = 8'b0;
    XRAM[64436] = 8'b0;
    XRAM[64437] = 8'b0;
    XRAM[64438] = 8'b0;
    XRAM[64439] = 8'b0;
    XRAM[64440] = 8'b0;
    XRAM[64441] = 8'b0;
    XRAM[64442] = 8'b0;
    XRAM[64443] = 8'b0;
    XRAM[64444] = 8'b0;
    XRAM[64445] = 8'b0;
    XRAM[64446] = 8'b0;
    XRAM[64447] = 8'b0;
    XRAM[64448] = 8'b0;
    XRAM[64449] = 8'b0;
    XRAM[64450] = 8'b0;
    XRAM[64451] = 8'b0;
    XRAM[64452] = 8'b0;
    XRAM[64453] = 8'b0;
    XRAM[64454] = 8'b0;
    XRAM[64455] = 8'b0;
    XRAM[64456] = 8'b0;
    XRAM[64457] = 8'b0;
    XRAM[64458] = 8'b0;
    XRAM[64459] = 8'b0;
    XRAM[64460] = 8'b0;
    XRAM[64461] = 8'b0;
    XRAM[64462] = 8'b0;
    XRAM[64463] = 8'b0;
    XRAM[64464] = 8'b0;
    XRAM[64465] = 8'b0;
    XRAM[64466] = 8'b0;
    XRAM[64467] = 8'b0;
    XRAM[64468] = 8'b0;
    XRAM[64469] = 8'b0;
    XRAM[64470] = 8'b0;
    XRAM[64471] = 8'b0;
    XRAM[64472] = 8'b0;
    XRAM[64473] = 8'b0;
    XRAM[64474] = 8'b0;
    XRAM[64475] = 8'b0;
    XRAM[64476] = 8'b0;
    XRAM[64477] = 8'b0;
    XRAM[64478] = 8'b0;
    XRAM[64479] = 8'b0;
    XRAM[64480] = 8'b0;
    XRAM[64481] = 8'b0;
    XRAM[64482] = 8'b0;
    XRAM[64483] = 8'b0;
    XRAM[64484] = 8'b0;
    XRAM[64485] = 8'b0;
    XRAM[64486] = 8'b0;
    XRAM[64487] = 8'b0;
    XRAM[64488] = 8'b0;
    XRAM[64489] = 8'b0;
    XRAM[64490] = 8'b0;
    XRAM[64491] = 8'b0;
    XRAM[64492] = 8'b0;
    XRAM[64493] = 8'b0;
    XRAM[64494] = 8'b0;
    XRAM[64495] = 8'b0;
    XRAM[64496] = 8'b0;
    XRAM[64497] = 8'b0;
    XRAM[64498] = 8'b0;
    XRAM[64499] = 8'b0;
    XRAM[64500] = 8'b0;
    XRAM[64501] = 8'b0;
    XRAM[64502] = 8'b0;
    XRAM[64503] = 8'b0;
    XRAM[64504] = 8'b0;
    XRAM[64505] = 8'b0;
    XRAM[64506] = 8'b0;
    XRAM[64507] = 8'b0;
    XRAM[64508] = 8'b0;
    XRAM[64509] = 8'b0;
    XRAM[64510] = 8'b0;
    XRAM[64511] = 8'b0;
    XRAM[64512] = 8'b0;
    XRAM[64513] = 8'b0;
    XRAM[64514] = 8'b0;
    XRAM[64515] = 8'b0;
    XRAM[64516] = 8'b0;
    XRAM[64517] = 8'b0;
    XRAM[64518] = 8'b0;
    XRAM[64519] = 8'b0;
    XRAM[64520] = 8'b0;
    XRAM[64521] = 8'b0;
    XRAM[64522] = 8'b0;
    XRAM[64523] = 8'b0;
    XRAM[64524] = 8'b0;
    XRAM[64525] = 8'b0;
    XRAM[64526] = 8'b0;
    XRAM[64527] = 8'b0;
    XRAM[64528] = 8'b0;
    XRAM[64529] = 8'b0;
    XRAM[64530] = 8'b0;
    XRAM[64531] = 8'b0;
    XRAM[64532] = 8'b0;
    XRAM[64533] = 8'b0;
    XRAM[64534] = 8'b0;
    XRAM[64535] = 8'b0;
    XRAM[64536] = 8'b0;
    XRAM[64537] = 8'b0;
    XRAM[64538] = 8'b0;
    XRAM[64539] = 8'b0;
    XRAM[64540] = 8'b0;
    XRAM[64541] = 8'b0;
    XRAM[64542] = 8'b0;
    XRAM[64543] = 8'b0;
    XRAM[64544] = 8'b0;
    XRAM[64545] = 8'b0;
    XRAM[64546] = 8'b0;
    XRAM[64547] = 8'b0;
    XRAM[64548] = 8'b0;
    XRAM[64549] = 8'b0;
    XRAM[64550] = 8'b0;
    XRAM[64551] = 8'b0;
    XRAM[64552] = 8'b0;
    XRAM[64553] = 8'b0;
    XRAM[64554] = 8'b0;
    XRAM[64555] = 8'b0;
    XRAM[64556] = 8'b0;
    XRAM[64557] = 8'b0;
    XRAM[64558] = 8'b0;
    XRAM[64559] = 8'b0;
    XRAM[64560] = 8'b0;
    XRAM[64561] = 8'b0;
    XRAM[64562] = 8'b0;
    XRAM[64563] = 8'b0;
    XRAM[64564] = 8'b0;
    XRAM[64565] = 8'b0;
    XRAM[64566] = 8'b0;
    XRAM[64567] = 8'b0;
    XRAM[64568] = 8'b0;
    XRAM[64569] = 8'b0;
    XRAM[64570] = 8'b0;
    XRAM[64571] = 8'b0;
    XRAM[64572] = 8'b0;
    XRAM[64573] = 8'b0;
    XRAM[64574] = 8'b0;
    XRAM[64575] = 8'b0;
    XRAM[64576] = 8'b0;
    XRAM[64577] = 8'b0;
    XRAM[64578] = 8'b0;
    XRAM[64579] = 8'b0;
    XRAM[64580] = 8'b0;
    XRAM[64581] = 8'b0;
    XRAM[64582] = 8'b0;
    XRAM[64583] = 8'b0;
    XRAM[64584] = 8'b0;
    XRAM[64585] = 8'b0;
    XRAM[64586] = 8'b0;
    XRAM[64587] = 8'b0;
    XRAM[64588] = 8'b0;
    XRAM[64589] = 8'b0;
    XRAM[64590] = 8'b0;
    XRAM[64591] = 8'b0;
    XRAM[64592] = 8'b0;
    XRAM[64593] = 8'b0;
    XRAM[64594] = 8'b0;
    XRAM[64595] = 8'b0;
    XRAM[64596] = 8'b0;
    XRAM[64597] = 8'b0;
    XRAM[64598] = 8'b0;
    XRAM[64599] = 8'b0;
    XRAM[64600] = 8'b0;
    XRAM[64601] = 8'b0;
    XRAM[64602] = 8'b0;
    XRAM[64603] = 8'b0;
    XRAM[64604] = 8'b0;
    XRAM[64605] = 8'b0;
    XRAM[64606] = 8'b0;
    XRAM[64607] = 8'b0;
    XRAM[64608] = 8'b0;
    XRAM[64609] = 8'b0;
    XRAM[64610] = 8'b0;
    XRAM[64611] = 8'b0;
    XRAM[64612] = 8'b0;
    XRAM[64613] = 8'b0;
    XRAM[64614] = 8'b0;
    XRAM[64615] = 8'b0;
    XRAM[64616] = 8'b0;
    XRAM[64617] = 8'b0;
    XRAM[64618] = 8'b0;
    XRAM[64619] = 8'b0;
    XRAM[64620] = 8'b0;
    XRAM[64621] = 8'b0;
    XRAM[64622] = 8'b0;
    XRAM[64623] = 8'b0;
    XRAM[64624] = 8'b0;
    XRAM[64625] = 8'b0;
    XRAM[64626] = 8'b0;
    XRAM[64627] = 8'b0;
    XRAM[64628] = 8'b0;
    XRAM[64629] = 8'b0;
    XRAM[64630] = 8'b0;
    XRAM[64631] = 8'b0;
    XRAM[64632] = 8'b0;
    XRAM[64633] = 8'b0;
    XRAM[64634] = 8'b0;
    XRAM[64635] = 8'b0;
    XRAM[64636] = 8'b0;
    XRAM[64637] = 8'b0;
    XRAM[64638] = 8'b0;
    XRAM[64639] = 8'b0;
    XRAM[64640] = 8'b0;
    XRAM[64641] = 8'b0;
    XRAM[64642] = 8'b0;
    XRAM[64643] = 8'b0;
    XRAM[64644] = 8'b0;
    XRAM[64645] = 8'b0;
    XRAM[64646] = 8'b0;
    XRAM[64647] = 8'b0;
    XRAM[64648] = 8'b0;
    XRAM[64649] = 8'b0;
    XRAM[64650] = 8'b0;
    XRAM[64651] = 8'b0;
    XRAM[64652] = 8'b0;
    XRAM[64653] = 8'b0;
    XRAM[64654] = 8'b0;
    XRAM[64655] = 8'b0;
    XRAM[64656] = 8'b0;
    XRAM[64657] = 8'b0;
    XRAM[64658] = 8'b0;
    XRAM[64659] = 8'b0;
    XRAM[64660] = 8'b0;
    XRAM[64661] = 8'b0;
    XRAM[64662] = 8'b0;
    XRAM[64663] = 8'b0;
    XRAM[64664] = 8'b0;
    XRAM[64665] = 8'b0;
    XRAM[64666] = 8'b0;
    XRAM[64667] = 8'b0;
    XRAM[64668] = 8'b0;
    XRAM[64669] = 8'b0;
    XRAM[64670] = 8'b0;
    XRAM[64671] = 8'b0;
    XRAM[64672] = 8'b0;
    XRAM[64673] = 8'b0;
    XRAM[64674] = 8'b0;
    XRAM[64675] = 8'b0;
    XRAM[64676] = 8'b0;
    XRAM[64677] = 8'b0;
    XRAM[64678] = 8'b0;
    XRAM[64679] = 8'b0;
    XRAM[64680] = 8'b0;
    XRAM[64681] = 8'b0;
    XRAM[64682] = 8'b0;
    XRAM[64683] = 8'b0;
    XRAM[64684] = 8'b0;
    XRAM[64685] = 8'b0;
    XRAM[64686] = 8'b0;
    XRAM[64687] = 8'b0;
    XRAM[64688] = 8'b0;
    XRAM[64689] = 8'b0;
    XRAM[64690] = 8'b0;
    XRAM[64691] = 8'b0;
    XRAM[64692] = 8'b0;
    XRAM[64693] = 8'b0;
    XRAM[64694] = 8'b0;
    XRAM[64695] = 8'b0;
    XRAM[64696] = 8'b0;
    XRAM[64697] = 8'b0;
    XRAM[64698] = 8'b0;
    XRAM[64699] = 8'b0;
    XRAM[64700] = 8'b0;
    XRAM[64701] = 8'b0;
    XRAM[64702] = 8'b0;
    XRAM[64703] = 8'b0;
    XRAM[64704] = 8'b0;
    XRAM[64705] = 8'b0;
    XRAM[64706] = 8'b0;
    XRAM[64707] = 8'b0;
    XRAM[64708] = 8'b0;
    XRAM[64709] = 8'b0;
    XRAM[64710] = 8'b0;
    XRAM[64711] = 8'b0;
    XRAM[64712] = 8'b0;
    XRAM[64713] = 8'b0;
    XRAM[64714] = 8'b0;
    XRAM[64715] = 8'b0;
    XRAM[64716] = 8'b0;
    XRAM[64717] = 8'b0;
    XRAM[64718] = 8'b0;
    XRAM[64719] = 8'b0;
    XRAM[64720] = 8'b0;
    XRAM[64721] = 8'b0;
    XRAM[64722] = 8'b0;
    XRAM[64723] = 8'b0;
    XRAM[64724] = 8'b0;
    XRAM[64725] = 8'b0;
    XRAM[64726] = 8'b0;
    XRAM[64727] = 8'b0;
    XRAM[64728] = 8'b0;
    XRAM[64729] = 8'b0;
    XRAM[64730] = 8'b0;
    XRAM[64731] = 8'b0;
    XRAM[64732] = 8'b0;
    XRAM[64733] = 8'b0;
    XRAM[64734] = 8'b0;
    XRAM[64735] = 8'b0;
    XRAM[64736] = 8'b0;
    XRAM[64737] = 8'b0;
    XRAM[64738] = 8'b0;
    XRAM[64739] = 8'b0;
    XRAM[64740] = 8'b0;
    XRAM[64741] = 8'b0;
    XRAM[64742] = 8'b0;
    XRAM[64743] = 8'b0;
    XRAM[64744] = 8'b0;
    XRAM[64745] = 8'b0;
    XRAM[64746] = 8'b0;
    XRAM[64747] = 8'b0;
    XRAM[64748] = 8'b0;
    XRAM[64749] = 8'b0;
    XRAM[64750] = 8'b0;
    XRAM[64751] = 8'b0;
    XRAM[64752] = 8'b0;
    XRAM[64753] = 8'b0;
    XRAM[64754] = 8'b0;
    XRAM[64755] = 8'b0;
    XRAM[64756] = 8'b0;
    XRAM[64757] = 8'b0;
    XRAM[64758] = 8'b0;
    XRAM[64759] = 8'b0;
    XRAM[64760] = 8'b0;
    XRAM[64761] = 8'b0;
    XRAM[64762] = 8'b0;
    XRAM[64763] = 8'b0;
    XRAM[64764] = 8'b0;
    XRAM[64765] = 8'b0;
    XRAM[64766] = 8'b0;
    XRAM[64767] = 8'b0;
    XRAM[64768] = 8'b0;
    XRAM[64769] = 8'b0;
    XRAM[64770] = 8'b0;
    XRAM[64771] = 8'b0;
    XRAM[64772] = 8'b0;
    XRAM[64773] = 8'b0;
    XRAM[64774] = 8'b0;
    XRAM[64775] = 8'b0;
    XRAM[64776] = 8'b0;
    XRAM[64777] = 8'b0;
    XRAM[64778] = 8'b0;
    XRAM[64779] = 8'b0;
    XRAM[64780] = 8'b0;
    XRAM[64781] = 8'b0;
    XRAM[64782] = 8'b0;
    XRAM[64783] = 8'b0;
    XRAM[64784] = 8'b0;
    XRAM[64785] = 8'b0;
    XRAM[64786] = 8'b0;
    XRAM[64787] = 8'b0;
    XRAM[64788] = 8'b0;
    XRAM[64789] = 8'b0;
    XRAM[64790] = 8'b0;
    XRAM[64791] = 8'b0;
    XRAM[64792] = 8'b0;
    XRAM[64793] = 8'b0;
    XRAM[64794] = 8'b0;
    XRAM[64795] = 8'b0;
    XRAM[64796] = 8'b0;
    XRAM[64797] = 8'b0;
    XRAM[64798] = 8'b0;
    XRAM[64799] = 8'b0;
    XRAM[64800] = 8'b0;
    XRAM[64801] = 8'b0;
    XRAM[64802] = 8'b0;
    XRAM[64803] = 8'b0;
    XRAM[64804] = 8'b0;
    XRAM[64805] = 8'b0;
    XRAM[64806] = 8'b0;
    XRAM[64807] = 8'b0;
    XRAM[64808] = 8'b0;
    XRAM[64809] = 8'b0;
    XRAM[64810] = 8'b0;
    XRAM[64811] = 8'b0;
    XRAM[64812] = 8'b0;
    XRAM[64813] = 8'b0;
    XRAM[64814] = 8'b0;
    XRAM[64815] = 8'b0;
    XRAM[64816] = 8'b0;
    XRAM[64817] = 8'b0;
    XRAM[64818] = 8'b0;
    XRAM[64819] = 8'b0;
    XRAM[64820] = 8'b0;
    XRAM[64821] = 8'b0;
    XRAM[64822] = 8'b0;
    XRAM[64823] = 8'b0;
    XRAM[64824] = 8'b0;
    XRAM[64825] = 8'b0;
    XRAM[64826] = 8'b0;
    XRAM[64827] = 8'b0;
    XRAM[64828] = 8'b0;
    XRAM[64829] = 8'b0;
    XRAM[64830] = 8'b0;
    XRAM[64831] = 8'b0;
    XRAM[64832] = 8'b0;
    XRAM[64833] = 8'b0;
    XRAM[64834] = 8'b0;
    XRAM[64835] = 8'b0;
    XRAM[64836] = 8'b0;
    XRAM[64837] = 8'b0;
    XRAM[64838] = 8'b0;
    XRAM[64839] = 8'b0;
    XRAM[64840] = 8'b0;
    XRAM[64841] = 8'b0;
    XRAM[64842] = 8'b0;
    XRAM[64843] = 8'b0;
    XRAM[64844] = 8'b0;
    XRAM[64845] = 8'b0;
    XRAM[64846] = 8'b0;
    XRAM[64847] = 8'b0;
    XRAM[64848] = 8'b0;
    XRAM[64849] = 8'b0;
    XRAM[64850] = 8'b0;
    XRAM[64851] = 8'b0;
    XRAM[64852] = 8'b0;
    XRAM[64853] = 8'b0;
    XRAM[64854] = 8'b0;
    XRAM[64855] = 8'b0;
    XRAM[64856] = 8'b0;
    XRAM[64857] = 8'b0;
    XRAM[64858] = 8'b0;
    XRAM[64859] = 8'b0;
    XRAM[64860] = 8'b0;
    XRAM[64861] = 8'b0;
    XRAM[64862] = 8'b0;
    XRAM[64863] = 8'b0;
    XRAM[64864] = 8'b0;
    XRAM[64865] = 8'b0;
    XRAM[64866] = 8'b0;
    XRAM[64867] = 8'b0;
    XRAM[64868] = 8'b0;
    XRAM[64869] = 8'b0;
    XRAM[64870] = 8'b0;
    XRAM[64871] = 8'b0;
    XRAM[64872] = 8'b0;
    XRAM[64873] = 8'b0;
    XRAM[64874] = 8'b0;
    XRAM[64875] = 8'b0;
    XRAM[64876] = 8'b0;
    XRAM[64877] = 8'b0;
    XRAM[64878] = 8'b0;
    XRAM[64879] = 8'b0;
    XRAM[64880] = 8'b0;
    XRAM[64881] = 8'b0;
    XRAM[64882] = 8'b0;
    XRAM[64883] = 8'b0;
    XRAM[64884] = 8'b0;
    XRAM[64885] = 8'b0;
    XRAM[64886] = 8'b0;
    XRAM[64887] = 8'b0;
    XRAM[64888] = 8'b0;
    XRAM[64889] = 8'b0;
    XRAM[64890] = 8'b0;
    XRAM[64891] = 8'b0;
    XRAM[64892] = 8'b0;
    XRAM[64893] = 8'b0;
    XRAM[64894] = 8'b0;
    XRAM[64895] = 8'b0;
    XRAM[64896] = 8'b0;
    XRAM[64897] = 8'b0;
    XRAM[64898] = 8'b0;
    XRAM[64899] = 8'b0;
    XRAM[64900] = 8'b0;
    XRAM[64901] = 8'b0;
    XRAM[64902] = 8'b0;
    XRAM[64903] = 8'b0;
    XRAM[64904] = 8'b0;
    XRAM[64905] = 8'b0;
    XRAM[64906] = 8'b0;
    XRAM[64907] = 8'b0;
    XRAM[64908] = 8'b0;
    XRAM[64909] = 8'b0;
    XRAM[64910] = 8'b0;
    XRAM[64911] = 8'b0;
    XRAM[64912] = 8'b0;
    XRAM[64913] = 8'b0;
    XRAM[64914] = 8'b0;
    XRAM[64915] = 8'b0;
    XRAM[64916] = 8'b0;
    XRAM[64917] = 8'b0;
    XRAM[64918] = 8'b0;
    XRAM[64919] = 8'b0;
    XRAM[64920] = 8'b0;
    XRAM[64921] = 8'b0;
    XRAM[64922] = 8'b0;
    XRAM[64923] = 8'b0;
    XRAM[64924] = 8'b0;
    XRAM[64925] = 8'b0;
    XRAM[64926] = 8'b0;
    XRAM[64927] = 8'b0;
    XRAM[64928] = 8'b0;
    XRAM[64929] = 8'b0;
    XRAM[64930] = 8'b0;
    XRAM[64931] = 8'b0;
    XRAM[64932] = 8'b0;
    XRAM[64933] = 8'b0;
    XRAM[64934] = 8'b0;
    XRAM[64935] = 8'b0;
    XRAM[64936] = 8'b0;
    XRAM[64937] = 8'b0;
    XRAM[64938] = 8'b0;
    XRAM[64939] = 8'b0;
    XRAM[64940] = 8'b0;
    XRAM[64941] = 8'b0;
    XRAM[64942] = 8'b0;
    XRAM[64943] = 8'b0;
    XRAM[64944] = 8'b0;
    XRAM[64945] = 8'b0;
    XRAM[64946] = 8'b0;
    XRAM[64947] = 8'b0;
    XRAM[64948] = 8'b0;
    XRAM[64949] = 8'b0;
    XRAM[64950] = 8'b0;
    XRAM[64951] = 8'b0;
    XRAM[64952] = 8'b0;
    XRAM[64953] = 8'b0;
    XRAM[64954] = 8'b0;
    XRAM[64955] = 8'b0;
    XRAM[64956] = 8'b0;
    XRAM[64957] = 8'b0;
    XRAM[64958] = 8'b0;
    XRAM[64959] = 8'b0;
    XRAM[64960] = 8'b0;
    XRAM[64961] = 8'b0;
    XRAM[64962] = 8'b0;
    XRAM[64963] = 8'b0;
    XRAM[64964] = 8'b0;
    XRAM[64965] = 8'b0;
    XRAM[64966] = 8'b0;
    XRAM[64967] = 8'b0;
    XRAM[64968] = 8'b0;
    XRAM[64969] = 8'b0;
    XRAM[64970] = 8'b0;
    XRAM[64971] = 8'b0;
    XRAM[64972] = 8'b0;
    XRAM[64973] = 8'b0;
    XRAM[64974] = 8'b0;
    XRAM[64975] = 8'b0;
    XRAM[64976] = 8'b0;
    XRAM[64977] = 8'b0;
    XRAM[64978] = 8'b0;
    XRAM[64979] = 8'b0;
    XRAM[64980] = 8'b0;
    XRAM[64981] = 8'b0;
    XRAM[64982] = 8'b0;
    XRAM[64983] = 8'b0;
    XRAM[64984] = 8'b0;
    XRAM[64985] = 8'b0;
    XRAM[64986] = 8'b0;
    XRAM[64987] = 8'b0;
    XRAM[64988] = 8'b0;
    XRAM[64989] = 8'b0;
    XRAM[64990] = 8'b0;
    XRAM[64991] = 8'b0;
    XRAM[64992] = 8'b0;
    XRAM[64993] = 8'b0;
    XRAM[64994] = 8'b0;
    XRAM[64995] = 8'b0;
    XRAM[64996] = 8'b0;
    XRAM[64997] = 8'b0;
    XRAM[64998] = 8'b0;
    XRAM[64999] = 8'b0;
    XRAM[65000] = 8'b0;
    XRAM[65001] = 8'b0;
    XRAM[65002] = 8'b0;
    XRAM[65003] = 8'b0;
    XRAM[65004] = 8'b0;
    XRAM[65005] = 8'b0;
    XRAM[65006] = 8'b0;
    XRAM[65007] = 8'b0;
    XRAM[65008] = 8'b0;
    XRAM[65009] = 8'b0;
    XRAM[65010] = 8'b0;
    XRAM[65011] = 8'b0;
    XRAM[65012] = 8'b0;
    XRAM[65013] = 8'b0;
    XRAM[65014] = 8'b0;
    XRAM[65015] = 8'b0;
    XRAM[65016] = 8'b0;
    XRAM[65017] = 8'b0;
    XRAM[65018] = 8'b0;
    XRAM[65019] = 8'b0;
    XRAM[65020] = 8'b0;
    XRAM[65021] = 8'b0;
    XRAM[65022] = 8'b0;
    XRAM[65023] = 8'b0;
    XRAM[65024] = 8'b0;
    XRAM[65025] = 8'b0;
    XRAM[65026] = 8'b0;
    XRAM[65027] = 8'b0;
    XRAM[65028] = 8'b0;
    XRAM[65029] = 8'b0;
    XRAM[65030] = 8'b0;
    XRAM[65031] = 8'b0;
    XRAM[65032] = 8'b0;
    XRAM[65033] = 8'b0;
    XRAM[65034] = 8'b0;
    XRAM[65035] = 8'b0;
    XRAM[65036] = 8'b0;
    XRAM[65037] = 8'b0;
    XRAM[65038] = 8'b0;
    XRAM[65039] = 8'b0;
    XRAM[65040] = 8'b0;
    XRAM[65041] = 8'b0;
    XRAM[65042] = 8'b0;
    XRAM[65043] = 8'b0;
    XRAM[65044] = 8'b0;
    XRAM[65045] = 8'b0;
    XRAM[65046] = 8'b0;
    XRAM[65047] = 8'b0;
    XRAM[65048] = 8'b0;
    XRAM[65049] = 8'b0;
    XRAM[65050] = 8'b0;
    XRAM[65051] = 8'b0;
    XRAM[65052] = 8'b0;
    XRAM[65053] = 8'b0;
    XRAM[65054] = 8'b0;
    XRAM[65055] = 8'b0;
    XRAM[65056] = 8'b0;
    XRAM[65057] = 8'b0;
    XRAM[65058] = 8'b0;
    XRAM[65059] = 8'b0;
    XRAM[65060] = 8'b0;
    XRAM[65061] = 8'b0;
    XRAM[65062] = 8'b0;
    XRAM[65063] = 8'b0;
    XRAM[65064] = 8'b0;
    XRAM[65065] = 8'b0;
    XRAM[65066] = 8'b0;
    XRAM[65067] = 8'b0;
    XRAM[65068] = 8'b0;
    XRAM[65069] = 8'b0;
    XRAM[65070] = 8'b0;
    XRAM[65071] = 8'b0;
    XRAM[65072] = 8'b0;
    XRAM[65073] = 8'b0;
    XRAM[65074] = 8'b0;
    XRAM[65075] = 8'b0;
    XRAM[65076] = 8'b0;
    XRAM[65077] = 8'b0;
    XRAM[65078] = 8'b0;
    XRAM[65079] = 8'b0;
    XRAM[65080] = 8'b0;
    XRAM[65081] = 8'b0;
    XRAM[65082] = 8'b0;
    XRAM[65083] = 8'b0;
    XRAM[65084] = 8'b0;
    XRAM[65085] = 8'b0;
    XRAM[65086] = 8'b0;
    XRAM[65087] = 8'b0;
    XRAM[65088] = 8'b0;
    XRAM[65089] = 8'b0;
    XRAM[65090] = 8'b0;
    XRAM[65091] = 8'b0;
    XRAM[65092] = 8'b0;
    XRAM[65093] = 8'b0;
    XRAM[65094] = 8'b0;
    XRAM[65095] = 8'b0;
    XRAM[65096] = 8'b0;
    XRAM[65097] = 8'b0;
    XRAM[65098] = 8'b0;
    XRAM[65099] = 8'b0;
    XRAM[65100] = 8'b0;
    XRAM[65101] = 8'b0;
    XRAM[65102] = 8'b0;
    XRAM[65103] = 8'b0;
    XRAM[65104] = 8'b0;
    XRAM[65105] = 8'b0;
    XRAM[65106] = 8'b0;
    XRAM[65107] = 8'b0;
    XRAM[65108] = 8'b0;
    XRAM[65109] = 8'b0;
    XRAM[65110] = 8'b0;
    XRAM[65111] = 8'b0;
    XRAM[65112] = 8'b0;
    XRAM[65113] = 8'b0;
    XRAM[65114] = 8'b0;
    XRAM[65115] = 8'b0;
    XRAM[65116] = 8'b0;
    XRAM[65117] = 8'b0;
    XRAM[65118] = 8'b0;
    XRAM[65119] = 8'b0;
    XRAM[65120] = 8'b0;
    XRAM[65121] = 8'b0;
    XRAM[65122] = 8'b0;
    XRAM[65123] = 8'b0;
    XRAM[65124] = 8'b0;
    XRAM[65125] = 8'b0;
    XRAM[65126] = 8'b0;
    XRAM[65127] = 8'b0;
    XRAM[65128] = 8'b0;
    XRAM[65129] = 8'b0;
    XRAM[65130] = 8'b0;
    XRAM[65131] = 8'b0;
    XRAM[65132] = 8'b0;
    XRAM[65133] = 8'b0;
    XRAM[65134] = 8'b0;
    XRAM[65135] = 8'b0;
    XRAM[65136] = 8'b0;
    XRAM[65137] = 8'b0;
    XRAM[65138] = 8'b0;
    XRAM[65139] = 8'b0;
    XRAM[65140] = 8'b0;
    XRAM[65141] = 8'b0;
    XRAM[65142] = 8'b0;
    XRAM[65143] = 8'b0;
    XRAM[65144] = 8'b0;
    XRAM[65145] = 8'b0;
    XRAM[65146] = 8'b0;
    XRAM[65147] = 8'b0;
    XRAM[65148] = 8'b0;
    XRAM[65149] = 8'b0;
    XRAM[65150] = 8'b0;
    XRAM[65151] = 8'b0;
    XRAM[65152] = 8'b0;
    XRAM[65153] = 8'b0;
    XRAM[65154] = 8'b0;
    XRAM[65155] = 8'b0;
    XRAM[65156] = 8'b0;
    XRAM[65157] = 8'b0;
    XRAM[65158] = 8'b0;
    XRAM[65159] = 8'b0;
    XRAM[65160] = 8'b0;
    XRAM[65161] = 8'b0;
    XRAM[65162] = 8'b0;
    XRAM[65163] = 8'b0;
    XRAM[65164] = 8'b0;
    XRAM[65165] = 8'b0;
    XRAM[65166] = 8'b0;
    XRAM[65167] = 8'b0;
    XRAM[65168] = 8'b0;
    XRAM[65169] = 8'b0;
    XRAM[65170] = 8'b0;
    XRAM[65171] = 8'b0;
    XRAM[65172] = 8'b0;
    XRAM[65173] = 8'b0;
    XRAM[65174] = 8'b0;
    XRAM[65175] = 8'b0;
    XRAM[65176] = 8'b0;
    XRAM[65177] = 8'b0;
    XRAM[65178] = 8'b0;
    XRAM[65179] = 8'b0;
    XRAM[65180] = 8'b0;
    XRAM[65181] = 8'b0;
    XRAM[65182] = 8'b0;
    XRAM[65183] = 8'b0;
    XRAM[65184] = 8'b0;
    XRAM[65185] = 8'b0;
    XRAM[65186] = 8'b0;
    XRAM[65187] = 8'b0;
    XRAM[65188] = 8'b0;
    XRAM[65189] = 8'b0;
    XRAM[65190] = 8'b0;
    XRAM[65191] = 8'b0;
    XRAM[65192] = 8'b0;
    XRAM[65193] = 8'b0;
    XRAM[65194] = 8'b0;
    XRAM[65195] = 8'b0;
    XRAM[65196] = 8'b0;
    XRAM[65197] = 8'b0;
    XRAM[65198] = 8'b0;
    XRAM[65199] = 8'b0;
    XRAM[65200] = 8'b0;
    XRAM[65201] = 8'b0;
    XRAM[65202] = 8'b0;
    XRAM[65203] = 8'b0;
    XRAM[65204] = 8'b0;
    XRAM[65205] = 8'b0;
    XRAM[65206] = 8'b0;
    XRAM[65207] = 8'b0;
    XRAM[65208] = 8'b0;
    XRAM[65209] = 8'b0;
    XRAM[65210] = 8'b0;
    XRAM[65211] = 8'b0;
    XRAM[65212] = 8'b0;
    XRAM[65213] = 8'b0;
    XRAM[65214] = 8'b0;
    XRAM[65215] = 8'b0;
    XRAM[65216] = 8'b0;
    XRAM[65217] = 8'b0;
    XRAM[65218] = 8'b0;
    XRAM[65219] = 8'b0;
    XRAM[65220] = 8'b0;
    XRAM[65221] = 8'b0;
    XRAM[65222] = 8'b0;
    XRAM[65223] = 8'b0;
    XRAM[65224] = 8'b0;
    XRAM[65225] = 8'b0;
    XRAM[65226] = 8'b0;
    XRAM[65227] = 8'b0;
    XRAM[65228] = 8'b0;
    XRAM[65229] = 8'b0;
    XRAM[65230] = 8'b0;
    XRAM[65231] = 8'b0;
    XRAM[65232] = 8'b0;
    XRAM[65233] = 8'b0;
    XRAM[65234] = 8'b0;
    XRAM[65235] = 8'b0;
    XRAM[65236] = 8'b0;
    XRAM[65237] = 8'b0;
    XRAM[65238] = 8'b0;
    XRAM[65239] = 8'b0;
    XRAM[65240] = 8'b0;
    XRAM[65241] = 8'b0;
    XRAM[65242] = 8'b0;
    XRAM[65243] = 8'b0;
    XRAM[65244] = 8'b0;
    XRAM[65245] = 8'b0;
    XRAM[65246] = 8'b0;
    XRAM[65247] = 8'b0;
    XRAM[65248] = 8'b0;
    XRAM[65249] = 8'b0;
    XRAM[65250] = 8'b0;
    XRAM[65251] = 8'b0;
    XRAM[65252] = 8'b0;
    XRAM[65253] = 8'b0;
    XRAM[65254] = 8'b0;
    XRAM[65255] = 8'b0;
    XRAM[65256] = 8'b0;
    XRAM[65257] = 8'b0;
    XRAM[65258] = 8'b0;
    XRAM[65259] = 8'b0;
    XRAM[65260] = 8'b0;
    XRAM[65261] = 8'b0;
    XRAM[65262] = 8'b0;
    XRAM[65263] = 8'b0;
    XRAM[65264] = 8'b0;
    XRAM[65265] = 8'b0;
    XRAM[65266] = 8'b0;
    XRAM[65267] = 8'b0;
    XRAM[65268] = 8'b0;
    XRAM[65269] = 8'b0;
    XRAM[65270] = 8'b0;
    XRAM[65271] = 8'b0;
    XRAM[65272] = 8'b0;
    XRAM[65273] = 8'b0;
    XRAM[65274] = 8'b0;
    XRAM[65275] = 8'b0;
    XRAM[65276] = 8'b0;
    XRAM[65277] = 8'b0;
    XRAM[65278] = 8'b0;
    XRAM[65279] = 8'b0;
    XRAM[65280] = 8'b0;
    XRAM[65281] = 8'b0;
    XRAM[65282] = 8'b0;
    XRAM[65283] = 8'b0;
    XRAM[65284] = 8'b0;
    XRAM[65285] = 8'b0;
    XRAM[65286] = 8'b0;
    XRAM[65287] = 8'b0;
    XRAM[65288] = 8'b0;
    XRAM[65289] = 8'b0;
    XRAM[65290] = 8'b0;
    XRAM[65291] = 8'b0;
    XRAM[65292] = 8'b0;
    XRAM[65293] = 8'b0;
    XRAM[65294] = 8'b0;
    XRAM[65295] = 8'b0;
    XRAM[65296] = 8'b0;
    XRAM[65297] = 8'b0;
    XRAM[65298] = 8'b0;
    XRAM[65299] = 8'b0;
    XRAM[65300] = 8'b0;
    XRAM[65301] = 8'b0;
    XRAM[65302] = 8'b0;
    XRAM[65303] = 8'b0;
    XRAM[65304] = 8'b0;
    XRAM[65305] = 8'b0;
    XRAM[65306] = 8'b0;
    XRAM[65307] = 8'b0;
    XRAM[65308] = 8'b0;
    XRAM[65309] = 8'b0;
    XRAM[65310] = 8'b0;
    XRAM[65311] = 8'b0;
    XRAM[65312] = 8'b0;
    XRAM[65313] = 8'b0;
    XRAM[65314] = 8'b0;
    XRAM[65315] = 8'b0;
    XRAM[65316] = 8'b0;
    XRAM[65317] = 8'b0;
    XRAM[65318] = 8'b0;
    XRAM[65319] = 8'b0;
    XRAM[65320] = 8'b0;
    XRAM[65321] = 8'b0;
    XRAM[65322] = 8'b0;
    XRAM[65323] = 8'b0;
    XRAM[65324] = 8'b0;
    XRAM[65325] = 8'b0;
    XRAM[65326] = 8'b0;
    XRAM[65327] = 8'b0;
    XRAM[65328] = 8'b0;
    XRAM[65329] = 8'b0;
    XRAM[65330] = 8'b0;
    XRAM[65331] = 8'b0;
    XRAM[65332] = 8'b0;
    XRAM[65333] = 8'b0;
    XRAM[65334] = 8'b0;
    XRAM[65335] = 8'b0;
    XRAM[65336] = 8'b0;
    XRAM[65337] = 8'b0;
    XRAM[65338] = 8'b0;
    XRAM[65339] = 8'b0;
    XRAM[65340] = 8'b0;
    XRAM[65341] = 8'b0;
    XRAM[65342] = 8'b0;
    XRAM[65343] = 8'b0;
    XRAM[65344] = 8'b0;
    XRAM[65345] = 8'b0;
    XRAM[65346] = 8'b0;
    XRAM[65347] = 8'b0;
    XRAM[65348] = 8'b0;
    XRAM[65349] = 8'b0;
    XRAM[65350] = 8'b0;
    XRAM[65351] = 8'b0;
    XRAM[65352] = 8'b0;
    XRAM[65353] = 8'b0;
    XRAM[65354] = 8'b0;
    XRAM[65355] = 8'b0;
    XRAM[65356] = 8'b0;
    XRAM[65357] = 8'b0;
    XRAM[65358] = 8'b0;
    XRAM[65359] = 8'b0;
    XRAM[65360] = 8'b0;
    XRAM[65361] = 8'b0;
    XRAM[65362] = 8'b0;
    XRAM[65363] = 8'b0;
    XRAM[65364] = 8'b0;
    XRAM[65365] = 8'b0;
    XRAM[65366] = 8'b0;
    XRAM[65367] = 8'b0;
    XRAM[65368] = 8'b0;
    XRAM[65369] = 8'b0;
    XRAM[65370] = 8'b0;
    XRAM[65371] = 8'b0;
    XRAM[65372] = 8'b0;
    XRAM[65373] = 8'b0;
    XRAM[65374] = 8'b0;
    XRAM[65375] = 8'b0;
    XRAM[65376] = 8'b0;
    XRAM[65377] = 8'b0;
    XRAM[65378] = 8'b0;
    XRAM[65379] = 8'b0;
    XRAM[65380] = 8'b0;
    XRAM[65381] = 8'b0;
    XRAM[65382] = 8'b0;
    XRAM[65383] = 8'b0;
    XRAM[65384] = 8'b0;
    XRAM[65385] = 8'b0;
    XRAM[65386] = 8'b0;
    XRAM[65387] = 8'b0;
    XRAM[65388] = 8'b0;
    XRAM[65389] = 8'b0;
    XRAM[65390] = 8'b0;
    XRAM[65391] = 8'b0;
    XRAM[65392] = 8'b0;
    XRAM[65393] = 8'b0;
    XRAM[65394] = 8'b0;
    XRAM[65395] = 8'b0;
    XRAM[65396] = 8'b0;
    XRAM[65397] = 8'b0;
    XRAM[65398] = 8'b0;
    XRAM[65399] = 8'b0;
    XRAM[65400] = 8'b0;
    XRAM[65401] = 8'b0;
    XRAM[65402] = 8'b0;
    XRAM[65403] = 8'b0;
    XRAM[65404] = 8'b0;
    XRAM[65405] = 8'b0;
    XRAM[65406] = 8'b0;
    XRAM[65407] = 8'b0;
    XRAM[65408] = 8'b0;
    XRAM[65409] = 8'b0;
    XRAM[65410] = 8'b0;
    XRAM[65411] = 8'b0;
    XRAM[65412] = 8'b0;
    XRAM[65413] = 8'b0;
    XRAM[65414] = 8'b0;
    XRAM[65415] = 8'b0;
    XRAM[65416] = 8'b0;
    XRAM[65417] = 8'b0;
    XRAM[65418] = 8'b0;
    XRAM[65419] = 8'b0;
    XRAM[65420] = 8'b0;
    XRAM[65421] = 8'b0;
    XRAM[65422] = 8'b0;
    XRAM[65423] = 8'b0;
    XRAM[65424] = 8'b0;
    XRAM[65425] = 8'b0;
    XRAM[65426] = 8'b0;
    XRAM[65427] = 8'b0;
    XRAM[65428] = 8'b0;
    XRAM[65429] = 8'b0;
    XRAM[65430] = 8'b0;
    XRAM[65431] = 8'b0;
    XRAM[65432] = 8'b0;
    XRAM[65433] = 8'b0;
    XRAM[65434] = 8'b0;
    XRAM[65435] = 8'b0;
    XRAM[65436] = 8'b0;
    XRAM[65437] = 8'b0;
    XRAM[65438] = 8'b0;
    XRAM[65439] = 8'b0;
    XRAM[65440] = 8'b0;
    XRAM[65441] = 8'b0;
    XRAM[65442] = 8'b0;
    XRAM[65443] = 8'b0;
    XRAM[65444] = 8'b0;
    XRAM[65445] = 8'b0;
    XRAM[65446] = 8'b0;
    XRAM[65447] = 8'b0;
    XRAM[65448] = 8'b0;
    XRAM[65449] = 8'b0;
    XRAM[65450] = 8'b0;
    XRAM[65451] = 8'b0;
    XRAM[65452] = 8'b0;
    XRAM[65453] = 8'b0;
    XRAM[65454] = 8'b0;
    XRAM[65455] = 8'b0;
    XRAM[65456] = 8'b0;
    XRAM[65457] = 8'b0;
    XRAM[65458] = 8'b0;
    XRAM[65459] = 8'b0;
    XRAM[65460] = 8'b0;
    XRAM[65461] = 8'b0;
    XRAM[65462] = 8'b0;
    XRAM[65463] = 8'b0;
    XRAM[65464] = 8'b0;
    XRAM[65465] = 8'b0;
    XRAM[65466] = 8'b0;
    XRAM[65467] = 8'b0;
    XRAM[65468] = 8'b0;
    XRAM[65469] = 8'b0;
    XRAM[65470] = 8'b0;
    XRAM[65471] = 8'b0;
    XRAM[65472] = 8'b0;
    XRAM[65473] = 8'b0;
    XRAM[65474] = 8'b0;
    XRAM[65475] = 8'b0;
    XRAM[65476] = 8'b0;
    XRAM[65477] = 8'b0;
    XRAM[65478] = 8'b0;
    XRAM[65479] = 8'b0;
    XRAM[65480] = 8'b0;
    XRAM[65481] = 8'b0;
    XRAM[65482] = 8'b0;
    XRAM[65483] = 8'b0;
    XRAM[65484] = 8'b0;
    XRAM[65485] = 8'b0;
    XRAM[65486] = 8'b0;
    XRAM[65487] = 8'b0;
    XRAM[65488] = 8'b0;
    XRAM[65489] = 8'b0;
    XRAM[65490] = 8'b0;
    XRAM[65491] = 8'b0;
    XRAM[65492] = 8'b0;
    XRAM[65493] = 8'b0;
    XRAM[65494] = 8'b0;
    XRAM[65495] = 8'b0;
    XRAM[65496] = 8'b0;
    XRAM[65497] = 8'b0;
    XRAM[65498] = 8'b0;
    XRAM[65499] = 8'b0;
    XRAM[65500] = 8'b0;
    XRAM[65501] = 8'b0;
    XRAM[65502] = 8'b0;
    XRAM[65503] = 8'b0;
    XRAM[65504] = 8'b0;
    XRAM[65505] = 8'b0;
    XRAM[65506] = 8'b0;
    XRAM[65507] = 8'b0;
    XRAM[65508] = 8'b0;
    XRAM[65509] = 8'b0;
    XRAM[65510] = 8'b0;
    XRAM[65511] = 8'b0;
    XRAM[65512] = 8'b0;
    XRAM[65513] = 8'b0;
    XRAM[65514] = 8'b0;
    XRAM[65515] = 8'b0;
    XRAM[65516] = 8'b0;
    XRAM[65517] = 8'b0;
    XRAM[65518] = 8'b0;
    XRAM[65519] = 8'b0;
    XRAM[65520] = 8'b0;
    XRAM[65521] = 8'b0;
    XRAM[65522] = 8'b0;
    XRAM[65523] = 8'b0;
    XRAM[65524] = 8'b0;
    XRAM[65525] = 8'b0;
    XRAM[65526] = 8'b0;
    XRAM[65527] = 8'b0;
    XRAM[65528] = 8'b0;
    XRAM[65529] = 8'b0;
    XRAM[65530] = 8'b0;
    XRAM[65531] = 8'b0;
    XRAM[65532] = 8'b0;
    XRAM[65533] = 8'b0;
    XRAM[65534] = 8'b0;
    XRAM[65535] = 8'b0;
`endif
  end
  else begin
    if (step) begin
      P0INREG <= P0IN;
      P1INREG <= P1IN;
      P2INREG <= P2IN;
      P3INREG <= P3IN;
      ACC <= ACC_next;
      P2 <= P2_next;
      P0 <= P0_next;
      P1 <= P1_next;
      P3 <= P3_next;
      SP <= SP_next;
      PC <= PC_next;
      B <= B_next;
      DPL <= DPL_next;
      PSW <= PSW_next;
      DPH <= DPH_next;
      if (WR_COND_0_IRAM) IRAM[WR_ADDR_0_IRAM] <= WR_DATA_0_IRAM;
      if (WR_COND_1_IRAM) IRAM[WR_ADDR_1_IRAM] <= WR_DATA_1_IRAM;
    end
  end
end

endmodule
