
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire [7:0] _00003_;
  wire _00004_;
  wire [7:0] _00005_;
  wire [7:0] _00006_;
  wire [7:0] _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire _44107_;
  wire _44108_;
  wire _44109_;
  wire _44110_;
  wire _44111_;
  wire _44112_;
  wire _44113_;
  wire _44114_;
  wire _44115_;
  wire _44116_;
  wire _44117_;
  wire _44118_;
  wire _44119_;
  wire _44120_;
  wire _44121_;
  wire _44122_;
  wire _44123_;
  wire _44124_;
  wire _44125_;
  wire _44126_;
  wire _44127_;
  wire _44128_;
  wire _44129_;
  wire _44130_;
  wire _44131_;
  wire _44132_;
  wire _44133_;
  wire _44134_;
  wire _44135_;
  wire _44136_;
  wire _44137_;
  wire _44138_;
  wire _44139_;
  wire _44140_;
  wire _44141_;
  wire _44142_;
  wire _44143_;
  wire _44144_;
  wire _44145_;
  wire _44146_;
  wire _44147_;
  wire _44148_;
  wire _44149_;
  wire _44150_;
  wire _44151_;
  wire _44152_;
  wire _44153_;
  wire _44154_;
  wire _44155_;
  wire _44156_;
  wire _44157_;
  wire _44158_;
  wire _44159_;
  wire _44160_;
  wire _44161_;
  wire _44162_;
  wire _44163_;
  wire _44164_;
  wire _44165_;
  wire _44166_;
  wire _44167_;
  wire _44168_;
  wire _44169_;
  wire _44170_;
  wire _44171_;
  wire _44172_;
  wire _44173_;
  wire _44174_;
  wire _44175_;
  wire _44176_;
  wire _44177_;
  wire _44178_;
  wire _44179_;
  wire _44180_;
  wire _44181_;
  wire _44182_;
  wire _44183_;
  wire _44184_;
  wire _44185_;
  wire _44186_;
  wire _44187_;
  wire _44188_;
  wire _44189_;
  wire _44190_;
  wire _44191_;
  wire _44192_;
  wire _44193_;
  wire _44194_;
  wire _44195_;
  wire _44196_;
  wire _44197_;
  wire _44198_;
  wire _44199_;
  wire _44200_;
  wire _44201_;
  wire _44202_;
  wire _44203_;
  wire _44204_;
  wire _44205_;
  wire _44206_;
  wire _44207_;
  wire _44208_;
  wire _44209_;
  wire _44210_;
  wire _44211_;
  wire _44212_;
  wire _44213_;
  wire _44214_;
  wire _44215_;
  wire _44216_;
  wire _44217_;
  wire _44218_;
  wire _44219_;
  wire _44220_;
  wire _44221_;
  wire _44222_;
  wire _44223_;
  wire _44224_;
  wire _44225_;
  wire _44226_;
  wire _44227_;
  wire _44228_;
  wire _44229_;
  wire _44230_;
  wire _44231_;
  wire _44232_;
  wire _44233_;
  wire _44234_;
  wire _44235_;
  wire _44236_;
  wire _44237_;
  wire _44238_;
  wire _44239_;
  wire _44240_;
  wire _44241_;
  wire _44242_;
  wire _44243_;
  wire _44244_;
  wire _44245_;
  wire _44246_;
  wire _44247_;
  wire _44248_;
  wire _44249_;
  wire _44250_;
  wire _44251_;
  wire _44252_;
  wire _44253_;
  wire _44254_;
  wire _44255_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire \oc8051_golden_model_1.n1046 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire \oc8051_golden_model_1.n1063 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1214 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire \oc8051_golden_model_1.n1300 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1424 ;
  wire \oc8051_golden_model_1.n1425 ;
  wire [4:0] \oc8051_golden_model_1.n1430 ;
  wire \oc8051_golden_model_1.n1431 ;
  wire \oc8051_golden_model_1.n1439 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1456 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [8:0] \oc8051_golden_model_1.n1461 ;
  wire \oc8051_golden_model_1.n1462 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire \oc8051_golden_model_1.n1475 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [8:0] \oc8051_golden_model_1.n1496 ;
  wire \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [8:0] \oc8051_golden_model_1.n1593 ;
  wire \oc8051_golden_model_1.n1594 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [4:0] \oc8051_golden_model_1.n1597 ;
  wire \oc8051_golden_model_1.n1598 ;
  wire \oc8051_golden_model_1.n1605 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1622 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [8:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire [4:0] \oc8051_golden_model_1.n1630 ;
  wire \oc8051_golden_model_1.n1631 ;
  wire \oc8051_golden_model_1.n1638 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1655 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire [6:0] \oc8051_golden_model_1.n1748 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1879 ;
  wire [6:0] \oc8051_golden_model_1.n1880 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire \oc8051_golden_model_1.n1936 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire \oc8051_golden_model_1.n1953 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire \oc8051_golden_model_1.n2085 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire \oc8051_golden_model_1.n2102 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire \oc8051_golden_model_1.n2141 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire \oc8051_golden_model_1.n2200 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2444 ;
  wire \oc8051_golden_model_1.n2446 ;
  wire \oc8051_golden_model_1.n2452 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [7:0] \oc8051_golden_model_1.n2734 ;
  wire [6:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire \oc8051_golden_model_1.n2853 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire \oc8051_golden_model_1.n2875 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire [7:0] \oc8051_golden_model_1.n2914 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire p1_valid_r;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  output property_invalid_sp;
  wire property_valid_psw_1_r;
  wire property_valid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire regs_always_zero;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_42003_, rst);
  not (_15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_15704_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15715_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15704_);
  and (_15726_, _15715_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15737_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15704_);
  and (_15748_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15704_);
  nor (_15759_, _15748_, _15737_);
  and (_15770_, _15759_, _15726_);
  nor (_15781_, _15770_, _15693_);
  and (_15792_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15803_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_15813_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15803_);
  nor (_15824_, _15813_, _15792_);
  not (_15835_, _15824_);
  and (_15846_, _15835_, _15770_);
  or (_15857_, _15846_, _15781_);
  and (_22436_, _15857_, _42003_);
  nor (_15878_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15889_, _15878_);
  and (_15900_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_15911_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_15922_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_15933_, _15922_);
  not (_15944_, _15813_);
  nor (_15955_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_15966_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_15977_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15966_);
  nor (_15988_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_15999_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_16010_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15999_);
  nor (_16021_, _16010_, _15988_);
  nor (_16032_, _16021_, _15977_);
  not (_16043_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_16054_, _15977_, _16043_);
  nor (_16065_, _16054_, _16032_);
  and (_16076_, _16065_, _15955_);
  not (_16087_, _16076_);
  and (_16098_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16109_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_16120_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16131_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16120_);
  and (_16142_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_16152_, _16142_, _16109_);
  and (_16163_, _16152_, _16087_);
  nor (_16174_, _16163_, _15944_);
  not (_16185_, _15792_);
  nor (_16196_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_16207_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15999_);
  nor (_16218_, _16207_, _16196_);
  nor (_16229_, _16218_, _15977_);
  not (_16240_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_16251_, _15977_, _16240_);
  nor (_16262_, _16251_, _16229_);
  and (_16273_, _16262_, _15955_);
  not (_16284_, _16273_);
  and (_16295_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_16306_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_16317_, _16306_, _16295_);
  and (_16328_, _16317_, _16284_);
  nor (_16339_, _16328_, _16185_);
  nor (_16350_, _16339_, _16174_);
  nor (_16361_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_16372_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15999_);
  nor (_16383_, _16372_, _16361_);
  nor (_16394_, _16383_, _15977_);
  not (_16405_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_16416_, _15977_, _16405_);
  nor (_16427_, _16416_, _16394_);
  and (_16438_, _16427_, _15955_);
  not (_16449_, _16438_);
  and (_16460_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16471_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16481_, _16471_, _16460_);
  and (_16492_, _16481_, _16449_);
  nor (_16503_, _16492_, _15835_);
  nor (_16514_, _16503_, _15878_);
  and (_16525_, _16514_, _16350_);
  nor (_16536_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16558_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15999_);
  nor (_16559_, _16558_, _16536_);
  nor (_16570_, _16559_, _15977_);
  not (_16581_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16592_, _15977_, _16581_);
  nor (_16603_, _16592_, _16570_);
  and (_16614_, _16603_, _15955_);
  not (_16625_, _16614_);
  and (_16636_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_16647_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16658_, _16647_, _16636_);
  and (_16669_, _16658_, _16625_);
  and (_16680_, _16669_, _15878_);
  nor (_16691_, _16680_, _16525_);
  not (_16702_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16713_, _16702_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16724_, _16713_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16735_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16746_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16757_, _16746_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16768_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_16779_, _16768_, _16735_);
  nor (_16790_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16801_, _16790_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16811_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_16822_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16833_, _16713_, _16822_);
  and (_16844_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_16855_, _16844_, _16811_);
  and (_16866_, _16855_, _16779_);
  and (_16877_, _16790_, _16702_);
  and (_16888_, _16877_, _16603_);
  and (_16899_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16910_, _16899_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16921_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_16932_, _16899_, _16822_);
  and (_16943_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16954_, _16943_, _16921_);
  not (_16965_, _16954_);
  nor (_16976_, _16965_, _16888_);
  and (_16987_, _16976_, _16866_);
  not (_16998_, _16987_);
  and (_17009_, _16998_, _16691_);
  not (_17020_, _17009_);
  nor (_17031_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_17042_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15999_);
  nor (_17053_, _17042_, _17031_);
  nor (_17064_, _17053_, _15977_);
  not (_17075_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_17086_, _15977_, _17075_);
  nor (_17097_, _17086_, _17064_);
  and (_17108_, _17097_, _15955_);
  not (_17118_, _17108_);
  and (_17129_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_17140_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17151_, _17140_, _17129_);
  and (_17162_, _17151_, _17118_);
  nor (_17173_, _17162_, _15944_);
  nor (_17184_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_17195_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15999_);
  nor (_17205_, _17195_, _17184_);
  nor (_17216_, _17205_, _15977_);
  not (_17227_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_17238_, _15977_, _17227_);
  nor (_17249_, _17238_, _17216_);
  and (_17260_, _17249_, _15955_);
  not (_17281_, _17260_);
  and (_17282_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_17302_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17303_, _17302_, _17282_);
  and (_17314_, _17303_, _17281_);
  nor (_17325_, _17314_, _16185_);
  nor (_17336_, _17325_, _17173_);
  nor (_17347_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_17358_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15999_);
  nor (_17369_, _17358_, _17347_);
  nor (_17380_, _17369_, _15977_);
  not (_17391_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_17401_, _15977_, _17391_);
  nor (_17412_, _17401_, _17380_);
  and (_17423_, _17412_, _15955_);
  not (_17434_, _17423_);
  and (_17445_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_17456_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17467_, _17456_, _17445_);
  and (_17478_, _17467_, _17434_);
  nor (_17488_, _17478_, _15835_);
  nor (_17499_, _17488_, _15878_);
  and (_17510_, _17499_, _17336_);
  nor (_17521_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17532_, _15999_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17543_, _17532_, _17521_);
  nor (_17554_, _17543_, _15977_);
  not (_17565_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17576_, _15977_, _17565_);
  nor (_17586_, _17576_, _17554_);
  and (_17597_, _17586_, _15955_);
  not (_17608_, _17597_);
  and (_17619_, _16098_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17630_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_17641_, _17630_, _17619_);
  and (_17652_, _17641_, _17608_);
  and (_17663_, _17652_, _15878_);
  or (_17674_, _17663_, _17510_);
  and (_17684_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_17695_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_17706_, _17695_, _17684_);
  and (_17717_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17728_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_17739_, _17728_, _17717_);
  and (_17750_, _17739_, _17706_);
  and (_17761_, _17586_, _16877_);
  and (_17771_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17782_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_17793_, _17782_, _17771_);
  not (_17804_, _17793_);
  nor (_17815_, _17804_, _17761_);
  and (_17826_, _17815_, _17750_);
  nor (_17837_, _17826_, _17674_);
  and (_17848_, _17837_, _17020_);
  not (_17858_, _17848_);
  and (_17869_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17880_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_17891_, _17880_, _17869_);
  and (_17902_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_17913_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_17924_, _17913_, _17902_);
  and (_17935_, _17924_, _17891_);
  and (_17946_, _17249_, _16877_);
  and (_17956_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_17967_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17978_, _17967_, _17956_);
  not (_17989_, _17978_);
  nor (_18000_, _17989_, _17946_);
  and (_18011_, _18000_, _17935_);
  nor (_18022_, _18011_, _17674_);
  and (_18033_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_18044_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_18054_, _18044_, _18033_);
  and (_18065_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_18076_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_18087_, _18076_, _18065_);
  and (_18098_, _18087_, _18054_);
  and (_18109_, _16877_, _16262_);
  and (_18120_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_18131_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_18141_, _18131_, _18120_);
  not (_18152_, _18141_);
  nor (_18163_, _18152_, _18109_);
  and (_18174_, _18163_, _18098_);
  not (_18185_, _18174_);
  and (_18196_, _18185_, _16691_);
  and (_18207_, _18022_, _18196_);
  and (_18218_, _16998_, _18207_);
  nor (_18229_, _17009_, _18207_);
  nor (_18239_, _18229_, _18218_);
  and (_18250_, _18239_, _18022_);
  and (_18261_, _17837_, _17009_);
  nor (_18272_, _16987_, _17674_);
  not (_18283_, _17826_);
  and (_18294_, _18283_, _16691_);
  nor (_18305_, _18294_, _18272_);
  nor (_18316_, _18305_, _18261_);
  and (_18326_, _18316_, _18250_);
  nor (_18337_, _18316_, _18250_);
  nor (_18348_, _18337_, _18326_);
  and (_18359_, _18348_, _18218_);
  nor (_18370_, _18359_, _18326_);
  nor (_18381_, _18370_, _17858_);
  nor (_18392_, _17674_, _18174_);
  and (_18403_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_18414_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_18424_, _18414_, _18403_);
  and (_18435_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_18446_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_18457_, _18446_, _18435_);
  and (_18468_, _18457_, _18424_);
  and (_18479_, _17097_, _16877_);
  and (_18490_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_18501_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_18512_, _18501_, _18490_);
  not (_18523_, _18512_);
  nor (_18533_, _18523_, _18479_);
  and (_18544_, _18533_, _18468_);
  not (_18555_, _18544_);
  and (_18566_, _18555_, _16691_);
  and (_18577_, _18566_, _18392_);
  not (_18588_, _18011_);
  and (_18599_, _18588_, _16691_);
  nor (_18610_, _18599_, _18392_);
  nor (_18621_, _18610_, _18207_);
  and (_18632_, _18621_, _18577_);
  nor (_18642_, _17009_, _18022_);
  nor (_18653_, _18642_, _18250_);
  and (_18664_, _18653_, _18632_);
  nor (_18675_, _18348_, _18218_);
  nor (_18686_, _18675_, _18359_);
  and (_18697_, _18686_, _18664_);
  nor (_18708_, _18686_, _18664_);
  nor (_18719_, _18708_, _18697_);
  not (_18730_, _18719_);
  and (_18741_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_18752_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_18762_, _18752_, _18741_);
  and (_18773_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_18784_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor (_18795_, _18784_, _18773_);
  and (_18806_, _18795_, _18762_);
  and (_18817_, _17412_, _16877_);
  and (_18828_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_18839_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nor (_18850_, _18839_, _18828_);
  not (_18861_, _18850_);
  nor (_18871_, _18861_, _18817_);
  and (_18882_, _18871_, _18806_);
  nor (_18893_, _18882_, _17674_);
  and (_18904_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_18915_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_18926_, _18915_, _18904_);
  and (_18937_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_18948_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_18959_, _18948_, _18937_);
  and (_18970_, _18959_, _18926_);
  and (_18981_, _16877_, _16065_);
  and (_18991_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and (_19002_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19013_, _19002_, _18991_);
  not (_19024_, _19013_);
  nor (_19035_, _19024_, _18981_);
  and (_19046_, _19035_, _18970_);
  not (_19057_, _19046_);
  and (_19068_, _19057_, _16691_);
  and (_19079_, _19068_, _18893_);
  not (_19090_, _18882_);
  and (_19100_, _19090_, _16691_);
  not (_19111_, _19100_);
  nor (_19122_, _19046_, _17674_);
  and (_19133_, _19122_, _19111_);
  and (_19144_, _19133_, _18566_);
  nor (_19155_, _19144_, _19079_);
  nor (_19166_, _18544_, _17674_);
  nor (_19177_, _19166_, _18196_);
  nor (_19188_, _19177_, _18577_);
  not (_19199_, _19188_);
  nor (_19210_, _19199_, _19155_);
  nor (_19220_, _18621_, _18577_);
  nor (_19231_, _19220_, _18632_);
  and (_19242_, _19231_, _19210_);
  nor (_19253_, _18653_, _18632_);
  nor (_19264_, _19253_, _18664_);
  and (_19275_, _19264_, _19242_);
  and (_19286_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_19297_, _16757_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_19308_, _19297_, _19286_);
  and (_19319_, _16801_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_19329_, _16833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_19340_, _19329_, _19319_);
  and (_19351_, _19340_, _19308_);
  and (_19362_, _16877_, _16427_);
  and (_19373_, _16910_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_19384_, _16932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19395_, _19384_, _19373_);
  not (_19406_, _19395_);
  nor (_19417_, _19406_, _19362_);
  and (_19428_, _19417_, _19351_);
  nor (_19438_, _19428_, _17674_);
  and (_19449_, _19438_, _19100_);
  nor (_19460_, _19068_, _18893_);
  nor (_19471_, _19460_, _19079_);
  and (_19482_, _19471_, _19449_);
  nor (_19493_, _19133_, _18566_);
  nor (_19504_, _19493_, _19144_);
  and (_19515_, _19504_, _19482_);
  and (_19526_, _19199_, _19155_);
  nor (_19537_, _19526_, _19210_);
  and (_19548_, _19537_, _19515_);
  nor (_19558_, _19231_, _19210_);
  nor (_19569_, _19558_, _19242_);
  and (_19580_, _19569_, _19548_);
  nor (_19591_, _19264_, _19242_);
  nor (_19602_, _19591_, _19275_);
  and (_19613_, _19602_, _19580_);
  nor (_19624_, _19613_, _19275_);
  nor (_19635_, _19624_, _18730_);
  nor (_19646_, _19635_, _18697_);
  and (_19657_, _18370_, _17858_);
  nor (_19667_, _19657_, _18381_);
  not (_19678_, _19667_);
  nor (_19689_, _19678_, _19646_);
  or (_19700_, _19689_, _18261_);
  nor (_19711_, _19700_, _18381_);
  nor (_19722_, _19711_, _15933_);
  and (_19733_, _19711_, _15933_);
  nor (_19744_, _19733_, _19722_);
  not (_19755_, _19744_);
  and (_19766_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_19777_, _19678_, _19646_);
  nor (_19787_, _19777_, _19689_);
  and (_19798_, _19787_, _19766_);
  and (_19809_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_19820_, _19624_, _18730_);
  nor (_19831_, _19820_, _19635_);
  and (_19842_, _19831_, _19809_);
  nor (_19853_, _19831_, _19809_);
  nor (_19864_, _19853_, _19842_);
  not (_19875_, _19864_);
  and (_19886_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_19896_, _19602_, _19580_);
  nor (_19907_, _19896_, _19613_);
  and (_19918_, _19907_, _19886_);
  nor (_19929_, _19907_, _19886_);
  nor (_19940_, _19929_, _19918_);
  not (_19951_, _19940_);
  and (_19962_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_19973_, _19569_, _19548_);
  nor (_19984_, _19973_, _19580_);
  and (_19995_, _19984_, _19962_);
  nor (_20006_, _19984_, _19962_);
  nor (_20016_, _20006_, _19995_);
  not (_20027_, _20016_);
  and (_20038_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_20049_, _19537_, _19515_);
  nor (_20060_, _20049_, _19548_);
  and (_20071_, _20060_, _20038_);
  and (_20082_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_20093_, _19504_, _19482_);
  nor (_20104_, _20093_, _19515_);
  and (_20115_, _20104_, _20082_);
  and (_20126_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_20136_, _19471_, _19449_);
  nor (_20147_, _20136_, _19482_);
  and (_20158_, _20147_, _20126_);
  nor (_20169_, _20104_, _20082_);
  nor (_20180_, _20169_, _20115_);
  and (_20191_, _20180_, _20158_);
  nor (_20202_, _20191_, _20115_);
  not (_20213_, _20202_);
  nor (_20224_, _20060_, _20038_);
  nor (_20235_, _20224_, _20071_);
  and (_20246_, _20235_, _20213_);
  nor (_20256_, _20246_, _20071_);
  nor (_20267_, _20256_, _20027_);
  nor (_20278_, _20267_, _19995_);
  nor (_20289_, _20278_, _19951_);
  nor (_20300_, _20289_, _19918_);
  nor (_20311_, _20300_, _19875_);
  nor (_20322_, _20311_, _19842_);
  nor (_20333_, _19787_, _19766_);
  nor (_20344_, _20333_, _19798_);
  not (_20355_, _20344_);
  nor (_20366_, _20355_, _20322_);
  nor (_20376_, _20366_, _19798_);
  nor (_20387_, _20376_, _19755_);
  nor (_20398_, _20387_, _19722_);
  not (_20409_, _20398_);
  and (_20420_, _20409_, _15911_);
  and (_20431_, _20420_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_20442_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_20453_, _20442_, _20431_);
  and (_20464_, _20453_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20475_, _20464_, _15900_);
  and (_20486_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20497_, _20486_, _20475_);
  and (_20508_, _20475_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20518_, _20508_, _20497_);
  and (_24622_, _20518_, _42003_);
  nor (_20539_, _15770_, _15803_);
  and (_20550_, _15770_, _15803_);
  or (_20561_, _20550_, _20539_);
  and (_02472_, _20561_, _42003_);
  not (_20582_, _19428_);
  and (_20593_, _20582_, _16691_);
  and (_02667_, _20593_, _42003_);
  nor (_20614_, _19438_, _19100_);
  nor (_20625_, _20614_, _19449_);
  and (_02861_, _20625_, _42003_);
  nor (_20645_, _20147_, _20126_);
  nor (_20656_, _20645_, _20158_);
  and (_03065_, _20656_, _42003_);
  nor (_20677_, _20180_, _20158_);
  nor (_20688_, _20677_, _20191_);
  and (_03276_, _20688_, _42003_);
  nor (_20709_, _20235_, _20213_);
  nor (_20720_, _20709_, _20246_);
  and (_03477_, _20720_, _42003_);
  and (_20741_, _20256_, _20027_);
  nor (_20752_, _20741_, _20267_);
  and (_03678_, _20752_, _42003_);
  and (_20772_, _20278_, _19951_);
  nor (_20783_, _20772_, _20289_);
  and (_03879_, _20783_, _42003_);
  and (_20804_, _20300_, _19875_);
  nor (_20815_, _20804_, _20311_);
  and (_04080_, _20815_, _42003_);
  and (_20836_, _20355_, _20322_);
  nor (_20847_, _20836_, _20366_);
  and (_04181_, _20847_, _42003_);
  and (_20868_, _20376_, _19755_);
  nor (_20878_, _20868_, _20387_);
  and (_04282_, _20878_, _42003_);
  nor (_20899_, _20409_, _15911_);
  nor (_20910_, _20899_, _20420_);
  and (_04383_, _20910_, _42003_);
  and (_20931_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_20942_, _20931_, _20420_);
  nor (_20953_, _20942_, _20431_);
  and (_04484_, _20953_, _42003_);
  nor (_20974_, _20442_, _20431_);
  nor (_20984_, _20974_, _20453_);
  and (_04585_, _20984_, _42003_);
  and (_21005_, _15889_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_21016_, _21005_, _20453_);
  nor (_21027_, _21016_, _20464_);
  and (_04686_, _21027_, _42003_);
  nor (_21048_, _20464_, _15900_);
  nor (_21059_, _21048_, _20475_);
  and (_04787_, _21059_, _42003_);
  and (_21080_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15704_);
  nor (_21090_, _21080_, _15715_);
  not (_21101_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_21112_, _15737_, _21101_);
  and (_21123_, _21112_, _21090_);
  and (_21134_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_21145_, _21134_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21156_, _21134_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21167_, _21156_, _21145_);
  and (_00870_, _21167_, _42003_);
  and (_00901_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42003_);
  not (_21197_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_21208_, _17478_, _21197_);
  and (_21219_, _17162_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21230_, _21219_, _21208_);
  nor (_21241_, _21230_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21252_, _17314_, _21197_);
  and (_21263_, _17652_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_21274_, _21263_, _21252_);
  and (_21285_, _21274_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21296_, _21285_, _21241_);
  nor (_21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_21317_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_21328_, _21306_, _17826_);
  nor (_21339_, _21328_, _21317_);
  not (_21350_, _21339_);
  and (_21361_, _16492_, _21197_);
  and (_21372_, _16163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21383_, _21372_, _21361_);
  nor (_21394_, _21383_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21405_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21415_, _16328_, _21197_);
  and (_21426_, _16669_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21437_, _21426_, _21415_);
  nor (_21448_, _21437_, _21405_);
  nor (_21459_, _21448_, _21394_);
  nor (_21470_, _21459_, _21350_);
  and (_21492_, _21459_, _21350_);
  nor (_21504_, _21492_, _21470_);
  nor (_21516_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_21528_, _21306_, _16987_);
  nor (_21539_, _21528_, _21516_);
  not (_21551_, _21539_);
  nor (_21552_, _17478_, _21197_);
  nor (_21563_, _21552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21574_, _17162_, _21197_);
  and (_21585_, _17314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21596_, _21585_, _21574_);
  nor (_21607_, _21596_, _21405_);
  nor (_21618_, _21607_, _21563_);
  nor (_21629_, _21618_, _21551_);
  and (_21640_, _21618_, _21551_);
  nor (_21650_, _21640_, _21629_);
  not (_21661_, _21650_);
  nor (_21672_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_21683_, _21306_, _18011_);
  nor (_21694_, _21683_, _21672_);
  not (_21705_, _21694_);
  nor (_21716_, _16492_, _21197_);
  nor (_21727_, _21716_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21738_, _16163_, _21197_);
  and (_21748_, _16328_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21759_, _21748_, _21738_);
  nor (_21770_, _21759_, _21405_);
  nor (_21781_, _21770_, _21727_);
  nor (_21792_, _21781_, _21705_);
  and (_21803_, _21781_, _21705_);
  and (_21814_, _21230_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21825_, _21814_);
  nor (_21836_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_21847_, _21306_, _18174_);
  nor (_21857_, _21847_, _21836_);
  and (_21868_, _21857_, _21825_);
  and (_21879_, _21383_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21890_, _21879_);
  and (_21901_, _21306_, _18544_);
  nor (_21912_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_21923_, _21912_, _21901_);
  and (_21934_, _21923_, _21890_);
  nor (_21945_, _21923_, _21890_);
  nor (_21956_, _21945_, _21934_);
  not (_21967_, _21956_);
  and (_21977_, _21552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21988_, _21977_);
  and (_21999_, _21306_, _19046_);
  nor (_22010_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_22021_, _22010_, _21999_);
  and (_22032_, _22021_, _21988_);
  and (_22043_, _21716_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22064_, _22043_);
  nor (_22065_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_22076_, _21306_, _18882_);
  nor (_22086_, _22076_, _22065_);
  nor (_22097_, _22086_, _22064_);
  not (_22108_, _22097_);
  nor (_22119_, _22021_, _21988_);
  nor (_22130_, _22119_, _22032_);
  and (_22141_, _22130_, _22108_);
  nor (_22152_, _22141_, _22032_);
  nor (_22163_, _22152_, _21967_);
  nor (_22174_, _22163_, _21934_);
  nor (_22185_, _21857_, _21825_);
  nor (_22195_, _22185_, _21868_);
  not (_22206_, _22195_);
  nor (_22217_, _22206_, _22174_);
  nor (_22228_, _22217_, _21868_);
  nor (_22239_, _22228_, _21803_);
  nor (_22250_, _22239_, _21792_);
  nor (_22261_, _22250_, _21661_);
  nor (_22272_, _22261_, _21629_);
  not (_22283_, _22272_);
  and (_22294_, _22283_, _21504_);
  or (_22304_, _22294_, _21470_);
  and (_22326_, _17652_, _16669_);
  or (_22327_, _22326_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_22338_, _21596_);
  and (_22349_, _21274_, _22338_);
  nor (_22360_, _21759_, _21437_);
  and (_22371_, _22360_, _22349_);
  or (_22382_, _22371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22393_, _22382_, _22327_);
  and (_22404_, _22393_, _22304_);
  and (_22414_, _22404_, _21296_);
  nor (_22425_, _22283_, _21504_);
  or (_22437_, _22425_, _22294_);
  and (_22448_, _22437_, _22414_);
  nor (_22459_, _22414_, _21339_);
  nor (_22470_, _22459_, _22448_);
  not (_22481_, _22470_);
  and (_22492_, _22470_, _21296_);
  not (_22503_, _21459_);
  nor (_22514_, _22414_, _21551_);
  and (_22524_, _22250_, _21661_);
  nor (_22535_, _22524_, _22261_);
  and (_22546_, _22535_, _22414_);
  or (_22557_, _22546_, _22514_);
  and (_22568_, _22557_, _22503_);
  nor (_22579_, _22557_, _22503_);
  nor (_22590_, _22579_, _22568_);
  not (_22601_, _22590_);
  not (_22612_, _21618_);
  nor (_22623_, _22414_, _21705_);
  nor (_22633_, _21803_, _21792_);
  nor (_22644_, _22633_, _22228_);
  and (_22655_, _22633_, _22228_);
  or (_22666_, _22655_, _22644_);
  and (_22677_, _22666_, _22414_);
  or (_22688_, _22677_, _22623_);
  and (_22699_, _22688_, _22612_);
  nor (_22710_, _22688_, _22612_);
  not (_22721_, _21781_);
  and (_22732_, _22206_, _22174_);
  or (_22742_, _22732_, _22217_);
  and (_22753_, _22742_, _22414_);
  nor (_22764_, _22414_, _21857_);
  nor (_22775_, _22764_, _22753_);
  and (_22786_, _22775_, _22721_);
  and (_22797_, _22152_, _21967_);
  nor (_22808_, _22797_, _22163_);
  not (_22819_, _22808_);
  and (_22830_, _22819_, _22414_);
  nor (_22841_, _22414_, _21923_);
  nor (_22851_, _22841_, _22830_);
  and (_22862_, _22851_, _21825_);
  nor (_22873_, _22851_, _21825_);
  nor (_22884_, _22873_, _22862_);
  not (_22895_, _22884_);
  nor (_22906_, _22130_, _22108_);
  nor (_22917_, _22906_, _22141_);
  not (_22928_, _22917_);
  and (_22939_, _22928_, _22414_);
  nor (_22950_, _22414_, _22021_);
  nor (_22960_, _22950_, _22939_);
  and (_22971_, _22960_, _21890_);
  not (_22982_, _22086_);
  and (_23003_, _22414_, _22043_);
  or (_23004_, _23003_, _22982_);
  nand (_23015_, _22414_, _22043_);
  or (_23036_, _23015_, _22086_);
  and (_23037_, _23036_, _23004_);
  nor (_23048_, _23037_, _21977_);
  and (_23068_, _23037_, _21977_);
  nor (_23069_, _23068_, _23048_);
  and (_23080_, _21306_, _19428_);
  nor (_23101_, _21306_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_23102_, _23101_, _23080_);
  nor (_23113_, _23102_, _22064_);
  not (_23134_, _23113_);
  and (_23135_, _23134_, _23069_);
  nor (_23146_, _23135_, _23048_);
  nor (_23167_, _22960_, _21890_);
  nor (_23168_, _23167_, _22971_);
  not (_23178_, _23168_);
  nor (_23199_, _23178_, _23146_);
  nor (_23200_, _23199_, _22971_);
  nor (_23211_, _23200_, _22895_);
  nor (_23222_, _23211_, _22862_);
  nor (_23233_, _22775_, _22721_);
  nor (_23244_, _23233_, _22786_);
  not (_23255_, _23244_);
  nor (_23266_, _23255_, _23222_);
  nor (_23277_, _23266_, _22786_);
  nor (_23288_, _23277_, _22710_);
  nor (_23299_, _23288_, _22699_);
  nor (_23310_, _23299_, _22601_);
  or (_23321_, _23310_, _22568_);
  or (_23332_, _23321_, _22492_);
  and (_23343_, _23332_, _22393_);
  nor (_23354_, _23343_, _22481_);
  and (_23365_, _22492_, _22393_);
  and (_23376_, _23365_, _23321_);
  or (_23387_, _23376_, _23354_);
  and (_00922_, _23387_, _42003_);
  or (_23408_, _22470_, _21296_);
  and (_23419_, _23408_, _23343_);
  and (_03022_, _23419_, _42003_);
  and (_03033_, _22414_, _42003_);
  and (_03054_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42003_);
  and (_03076_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42003_);
  and (_03097_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42003_);
  or (_23480_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23491_, _21134_, rst);
  and (_03108_, _23491_, _23480_);
  not (_23512_, _23102_);
  and (_23523_, _23419_, _22043_);
  nor (_23534_, _23523_, _23512_);
  and (_23545_, _23523_, _23512_);
  or (_23556_, _23545_, _23534_);
  and (_03119_, _23556_, _42003_);
  nor (_23577_, _23419_, _23037_);
  nor (_23588_, _23134_, _23069_);
  nor (_23599_, _23588_, _23135_);
  and (_23610_, _23599_, _23419_);
  or (_23621_, _23610_, _23577_);
  and (_03130_, _23621_, _42003_);
  and (_23642_, _23178_, _23146_);
  or (_23653_, _23642_, _23199_);
  nand (_23664_, _23653_, _23419_);
  or (_23675_, _23419_, _22960_);
  and (_23686_, _23675_, _23664_);
  and (_03141_, _23686_, _42003_);
  and (_23707_, _23200_, _22895_);
  or (_23718_, _23707_, _23211_);
  nand (_23729_, _23718_, _23419_);
  or (_23740_, _23419_, _22851_);
  and (_23751_, _23740_, _23729_);
  and (_03152_, _23751_, _42003_);
  and (_23772_, _23255_, _23222_);
  or (_23783_, _23772_, _23266_);
  nand (_23794_, _23783_, _23419_);
  or (_23805_, _23419_, _22775_);
  and (_23816_, _23805_, _23794_);
  and (_03163_, _23816_, _42003_);
  or (_23837_, _22710_, _22699_);
  and (_23848_, _23837_, _23277_);
  nor (_23859_, _23837_, _23277_);
  or (_23870_, _23859_, _23848_);
  nand (_23881_, _23870_, _23419_);
  or (_23892_, _23419_, _22688_);
  and (_23903_, _23892_, _23881_);
  and (_03174_, _23903_, _42003_);
  and (_23924_, _23299_, _22601_);
  or (_23935_, _23924_, _23310_);
  nand (_23946_, _23935_, _23419_);
  or (_23957_, _23419_, _22557_);
  and (_23968_, _23957_, _23946_);
  and (_03185_, _23968_, _42003_);
  not (_23989_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24000_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15704_);
  and (_24011_, _24000_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24022_, _24011_, _23989_);
  and (_24033_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24044_, _24033_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24055_, _24033_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24066_, _24055_, _24044_);
  and (_24077_, _24066_, _24022_);
  not (_24088_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24099_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15704_);
  and (_24110_, _24099_, _23989_);
  and (_24121_, _24110_, _24088_);
  and (_24132_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24143_, _24132_, _24077_);
  not (_24154_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24165_, _24000_, _24154_);
  and (_24187_, _24165_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24199_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24211_, _24165_, _23989_);
  and (_24223_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_24235_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24247_, _24235_, _15704_);
  nor (_24259_, _24247_, _24000_);
  and (_24260_, _24259_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24271_, _24260_, _24223_);
  nor (_24282_, _24271_, _24199_);
  and (_24293_, _24282_, _24143_);
  nor (_24304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24315_, _24304_, _24033_);
  and (_24326_, _24315_, _24022_);
  and (_24337_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24348_, _24337_, _24326_);
  and (_24359_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24370_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_24381_, _24259_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_24392_, _24381_, _24370_);
  nor (_24403_, _24392_, _24359_);
  and (_24414_, _24403_, _24348_);
  and (_24425_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_24436_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_24447_, _24436_, _24425_);
  and (_24458_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_24469_, _24458_);
  not (_24480_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24491_, _24022_, _24480_);
  and (_24502_, _24259_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24513_, _24502_, _24491_);
  and (_24524_, _24513_, _24469_);
  and (_24535_, _24524_, _24447_);
  and (_24546_, _24535_, _24414_);
  and (_24557_, _24546_, _24293_);
  and (_24568_, _24044_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24579_, _24568_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_24590_, _24579_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24601_, _24590_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_24612_, _24601_);
  not (_24623_, _24022_);
  nor (_24634_, _24590_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_24645_, _24634_, _24623_);
  and (_24656_, _24645_, _24612_);
  not (_24667_, _24656_);
  and (_24678_, _24011_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24689_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_24700_, _24689_, _24678_);
  and (_24711_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_24722_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_24732_, _24722_, _24711_);
  and (_24743_, _24732_, _24700_);
  and (_24754_, _24743_, _24667_);
  nor (_24765_, _24579_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_24776_, _24765_);
  nor (_24787_, _24590_, _24623_);
  and (_24798_, _24787_, _24776_);
  not (_24809_, _24798_);
  and (_24820_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_24831_, _24820_, _24678_);
  and (_24842_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_24853_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_24864_, _24853_, _24842_);
  and (_24875_, _24864_, _24831_);
  and (_24886_, _24875_, _24809_);
  nor (_24897_, _24886_, _24754_);
  not (_24908_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_24919_, _24601_, _24908_);
  and (_24930_, _24601_, _24908_);
  nor (_24941_, _24930_, _24919_);
  nor (_24952_, _24941_, _24623_);
  not (_24963_, _24952_);
  and (_24973_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_24984_, _24973_);
  not (_24995_, _24678_);
  and (_25006_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_25017_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_25028_, _25017_, _25006_);
  and (_25039_, _25028_, _24995_);
  and (_25050_, _25039_, _24984_);
  and (_25061_, _25050_, _24963_);
  not (_25072_, _25061_);
  and (_25082_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_25093_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_25114_, _25093_, _25082_);
  not (_25115_, _24568_);
  nor (_25126_, _24044_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25137_, _25126_, _24623_);
  and (_25158_, _25137_, _25115_);
  and (_25159_, _24259_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_25170_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25191_, _25170_, _25159_);
  not (_25192_, _25191_);
  nor (_25202_, _25192_, _25158_);
  and (_25213_, _25202_, _25114_);
  nor (_25224_, _24568_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_25245_, _25224_, _24623_);
  nor (_25246_, _25245_, _24579_);
  and (_25257_, _24187_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_25268_, _25257_, _25246_);
  and (_25279_, _24211_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_25290_, _24259_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_25301_, _25290_, _25279_);
  and (_25312_, _24121_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25322_, _25312_, _24678_);
  and (_25333_, _25322_, _25301_);
  and (_25344_, _25333_, _25268_);
  not (_25355_, _25344_);
  and (_25376_, _25355_, _25213_);
  and (_25377_, _25376_, _25072_);
  and (_25388_, _25377_, _24897_);
  nand (_25399_, _25388_, _24557_);
  and (_25410_, _23387_, _21123_);
  not (_25421_, _25410_);
  and (_25432_, _20518_, _15770_);
  not (_25443_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_25454_, _21080_, _25443_);
  and (_25465_, _25454_, _15759_);
  nor (_25476_, _16987_, _16669_);
  and (_25486_, _16987_, _16669_);
  nor (_25497_, _25486_, _25476_);
  not (_25508_, _25497_);
  nor (_25519_, _18011_, _17314_);
  nor (_25530_, _18174_, _16328_);
  and (_25551_, _18011_, _17314_);
  nor (_25552_, _25551_, _25519_);
  and (_25563_, _25552_, _25530_);
  nor (_25573_, _25563_, _25519_);
  nor (_25584_, _25573_, _25508_);
  and (_25595_, _18174_, _16328_);
  nor (_25606_, _25595_, _25530_);
  nor (_25617_, _18544_, _17162_);
  and (_25628_, _18544_, _17162_);
  nor (_25639_, _25628_, _25617_);
  nor (_25650_, _19046_, _16163_);
  and (_25660_, _19046_, _16163_);
  nor (_25671_, _25660_, _25650_);
  not (_25682_, _25671_);
  nor (_25693_, _18882_, _17478_);
  nor (_25704_, _19428_, _16492_);
  and (_25715_, _18882_, _17478_);
  nor (_25726_, _25715_, _25693_);
  and (_25746_, _25726_, _25704_);
  nor (_25747_, _25746_, _25693_);
  nor (_25758_, _25747_, _25682_);
  nor (_25769_, _25758_, _25650_);
  nor (_25780_, _25769_, _25639_);
  and (_25791_, _25769_, _25639_);
  nor (_25802_, _25791_, _25780_);
  not (_25813_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_25824_, _15977_, _25813_);
  not (_25834_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25845_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25856_, _25845_, _17543_);
  nor (_25867_, _25856_, _25834_);
  nor (_25878_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25889_, _25878_, _16218_);
  not (_25900_, _25889_);
  not (_25911_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25921_, _25911_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25932_, _25921_, _16559_);
  not (_25943_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25954_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25943_);
  and (_25965_, _25954_, _17205_);
  nor (_25976_, _25965_, _25932_);
  and (_25987_, _25976_, _25900_);
  and (_25998_, _25987_, _25867_);
  and (_26008_, _25845_, _17053_);
  nor (_26019_, _26008_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26030_, _25954_, _17369_);
  not (_26041_, _26030_);
  and (_26052_, _25921_, _16021_);
  and (_26063_, _25878_, _16383_);
  nor (_26074_, _26063_, _26052_);
  and (_26094_, _26074_, _26041_);
  and (_26095_, _26094_, _26019_);
  nor (_26106_, _26095_, _25998_);
  nor (_26117_, _26106_, _15977_);
  nor (_26128_, _26117_, _25824_);
  and (_26139_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26150_, _26139_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_26161_, _26150_);
  and (_26172_, _26161_, _26128_);
  and (_26182_, _26161_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_26203_, _26182_, _26172_);
  and (_26204_, _19428_, _16492_);
  nor (_26215_, _26204_, _25704_);
  not (_26226_, _26215_);
  nor (_26237_, _26226_, _26203_);
  and (_26248_, _26237_, _25726_);
  and (_26259_, _25747_, _25682_);
  nor (_26269_, _26259_, _25758_);
  and (_26280_, _26269_, _26248_);
  not (_26291_, _26280_);
  nor (_26302_, _26291_, _25802_);
  nor (_26313_, _25769_, _25628_);
  or (_26324_, _26313_, _25617_);
  or (_26335_, _26324_, _26302_);
  and (_26346_, _26335_, _25606_);
  nor (_26356_, _25552_, _25530_);
  nor (_26367_, _26356_, _25563_);
  and (_26378_, _26367_, _26346_);
  and (_26389_, _25573_, _25508_);
  nor (_26400_, _26389_, _25584_);
  and (_26411_, _26400_, _26378_);
  or (_26422_, _26411_, _25584_);
  nor (_26433_, _26422_, _25476_);
  nor (_26443_, _17826_, _17652_);
  and (_26454_, _17826_, _17652_);
  nor (_26465_, _26454_, _26443_);
  not (_26476_, _26465_);
  nor (_26487_, _26476_, _26433_);
  and (_26498_, _26476_, _26433_);
  nor (_26509_, _26498_, _26487_);
  and (_26520_, _26509_, _25465_);
  not (_26531_, _26520_);
  not (_26541_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_26552_, _15715_, _26541_);
  and (_26563_, _26552_, _15759_);
  not (_26574_, _26563_);
  not (_26585_, _16669_);
  nor (_26596_, _16987_, _26585_);
  not (_26607_, _17314_);
  nor (_26618_, _18011_, _26607_);
  not (_26628_, _16328_);
  and (_26649_, _18174_, _26628_);
  nor (_26650_, _26649_, _25552_);
  nor (_26661_, _26650_, _26618_);
  nor (_26672_, _26661_, _25497_);
  nor (_26683_, _26672_, _26596_);
  and (_26694_, _26661_, _25497_);
  nor (_26705_, _26694_, _26672_);
  not (_26715_, _26705_);
  and (_26726_, _26649_, _25552_);
  nor (_26737_, _26726_, _26650_);
  not (_26748_, _26737_);
  not (_26759_, _25606_);
  not (_26770_, _16492_);
  and (_26781_, _19428_, _26770_);
  nor (_26792_, _26781_, _25726_);
  not (_26803_, _17478_);
  nor (_26814_, _18882_, _26803_);
  nor (_26824_, _26814_, _26792_);
  nor (_26835_, _26824_, _25671_);
  not (_26846_, _16163_);
  nor (_26857_, _19046_, _26846_);
  nor (_26868_, _26857_, _26835_);
  nor (_26879_, _26868_, _25639_);
  and (_26890_, _26868_, _25639_);
  nor (_26901_, _26890_, _26879_);
  not (_26912_, _26901_);
  and (_26923_, _26824_, _25671_);
  nor (_26943_, _26923_, _26835_);
  not (_26944_, _26943_);
  nor (_26955_, _26215_, _26203_);
  and (_26966_, _26781_, _25726_);
  nor (_26977_, _26966_, _26792_);
  not (_26988_, _26977_);
  and (_26999_, _26988_, _26955_);
  and (_27010_, _26999_, _26944_);
  and (_27021_, _27010_, _26912_);
  not (_27032_, _17162_);
  or (_27052_, _18544_, _27032_);
  and (_27053_, _18544_, _27032_);
  or (_27064_, _26868_, _27053_);
  and (_27075_, _27064_, _27052_);
  or (_27086_, _27075_, _27021_);
  and (_27097_, _27086_, _26759_);
  and (_27108_, _27097_, _26748_);
  and (_27119_, _27108_, _26715_);
  nor (_27130_, _27119_, _26683_);
  nor (_27141_, _27130_, _26465_);
  and (_27152_, _27130_, _26465_);
  nor (_27162_, _27152_, _27141_);
  nor (_27173_, _27162_, _26574_);
  not (_27184_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27195_, _15748_, _27184_);
  and (_27206_, _27195_, _25454_);
  not (_27217_, _27206_);
  nor (_27228_, _27217_, _26454_);
  and (_27239_, _27195_, _21090_);
  and (_27250_, _27239_, _26465_);
  nor (_27271_, _27250_, _27228_);
  and (_27272_, _15748_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27282_, _27272_, _21090_);
  not (_27293_, _27282_);
  nor (_27304_, _27293_, _19428_);
  and (_27315_, _27195_, _15715_);
  not (_27326_, _27315_);
  nor (_27337_, _27326_, _16987_);
  nor (_27348_, _27337_, _27304_);
  and (_27359_, _27272_, _25454_);
  not (_27370_, _27359_);
  nor (_27381_, _27370_, _26203_);
  and (_27391_, _21112_, _15726_);
  and (_27402_, _27391_, _26443_);
  and (_27413_, _26552_, _21112_);
  and (_27424_, _27413_, _17826_);
  nor (_27435_, _27424_, _27402_);
  and (_27446_, _21090_, _15759_);
  not (_27457_, _27446_);
  nor (_27468_, _27457_, _17826_);
  not (_27479_, _27468_);
  nand (_27490_, _27479_, _27435_);
  nor (_27501_, _27490_, _27381_);
  and (_27511_, _27501_, _27348_);
  and (_27532_, _27272_, _26552_);
  nor (_27533_, _19428_, _18882_);
  and (_27544_, _27533_, _19057_);
  and (_27555_, _27544_, _18555_);
  and (_27566_, _27555_, _18185_);
  and (_27577_, _27566_, _18588_);
  and (_27588_, _27577_, _16998_);
  and (_27598_, _27588_, _26203_);
  not (_27609_, _26203_);
  and (_27620_, _16987_, _18011_);
  and (_27631_, _19428_, _18882_);
  and (_27642_, _27631_, _19046_);
  and (_27653_, _27642_, _18544_);
  and (_27664_, _27653_, _18174_);
  and (_27675_, _27664_, _27620_);
  and (_27686_, _27675_, _27609_);
  nor (_27697_, _27686_, _27598_);
  and (_27708_, _27697_, _17826_);
  nor (_27718_, _27697_, _17826_);
  nor (_27729_, _27718_, _27708_);
  and (_27740_, _27729_, _27532_);
  not (_27751_, _17652_);
  nor (_27762_, _26203_, _27751_);
  not (_27773_, _27762_);
  and (_27784_, _26203_, _17826_);
  and (_27795_, _27272_, _15726_);
  not (_27816_, _27795_);
  nor (_27817_, _27816_, _27784_);
  and (_27828_, _27817_, _27773_);
  nor (_27838_, _27828_, _27740_);
  and (_27849_, _25454_, _21112_);
  not (_27860_, _27849_);
  and (_27871_, _19046_, _18882_);
  nor (_27882_, _27871_, _18544_);
  and (_27893_, _27882_, _27849_);
  and (_27904_, _27893_, _18185_);
  nor (_27915_, _27904_, _18588_);
  and (_27926_, _27915_, _16987_);
  nor (_27937_, _27620_, _17826_);
  nor (_27948_, _27937_, _27893_);
  and (_27958_, _27948_, _26203_);
  nor (_27969_, _27958_, _27926_);
  and (_27980_, _27969_, _17826_);
  nor (_27991_, _27969_, _17826_);
  nor (_28002_, _27991_, _27980_);
  nor (_28013_, _28002_, _27860_);
  not (_28024_, _28013_);
  and (_28035_, _28024_, _27838_);
  and (_28046_, _28035_, _27511_);
  and (_28057_, _28046_, _27271_);
  not (_28068_, _28057_);
  nor (_28079_, _28068_, _27173_);
  and (_28089_, _28079_, _26531_);
  not (_28100_, _28089_);
  nor (_28111_, _28100_, _25432_);
  and (_28122_, _28111_, _25421_);
  not (_28133_, _28122_);
  or (_28144_, _28133_, _25399_);
  not (_28155_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_28166_, \oc8051_top_1.oc8051_decoder1.wr , _15704_);
  not (_28177_, _28166_);
  nor (_28188_, _28177_, _24110_);
  and (_28199_, _28188_, _28155_);
  not (_28210_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_28221_, _25399_, _28210_);
  and (_28231_, _28221_, _28199_);
  and (_28252_, _28231_, _28144_);
  nor (_28253_, _28188_, _28210_);
  not (_28264_, _25465_);
  nor (_28275_, _26487_, _26443_);
  nor (_28286_, _28275_, _28264_);
  not (_28297_, _28286_);
  and (_28308_, _17826_, _27751_);
  nor (_28319_, _28308_, _27141_);
  nor (_28330_, _28319_, _26574_);
  and (_28341_, _26203_, _16987_);
  and (_28351_, _28341_, _27915_);
  nor (_28362_, _28351_, _27784_);
  nor (_28373_, _26203_, _17826_);
  not (_28384_, _28373_);
  nor (_28395_, _28384_, _27926_);
  nor (_28406_, _28395_, _27860_);
  and (_28417_, _28406_, _28362_);
  or (_28438_, _28417_, _27893_);
  nor (_28439_, _26182_, _26128_);
  not (_28450_, _27239_);
  nor (_28460_, _28450_, _26172_);
  not (_28471_, _28460_);
  nor (_28482_, _27293_, _26128_);
  nor (_28493_, _28482_, _27206_);
  and (_28504_, _28493_, _28471_);
  nor (_28515_, _28504_, _28439_);
  not (_28526_, _28515_);
  nor (_28537_, _27457_, _26203_);
  nor (_28548_, _27370_, _19428_);
  and (_28559_, _27195_, _15726_);
  not (_28569_, _28559_);
  nor (_28580_, _28569_, _17826_);
  nor (_28591_, _28580_, _28548_);
  not (_28602_, _28591_);
  nor (_28613_, _28602_, _28537_);
  and (_28624_, _27413_, _26203_);
  and (_28635_, _26150_, _26128_);
  and (_28646_, _27195_, _26552_);
  and (_28657_, _27391_, _26128_);
  nor (_28668_, _28657_, _28646_);
  nor (_28679_, _28668_, _28635_);
  nor (_28689_, _28679_, _28624_);
  and (_28700_, _28689_, _28613_);
  and (_28711_, _28700_, _28526_);
  not (_28722_, _28711_);
  nor (_28733_, _28722_, _28438_);
  not (_28744_, _28733_);
  nor (_28755_, _28744_, _28330_);
  and (_28766_, _28755_, _28297_);
  not (_28777_, _24293_);
  nor (_28788_, _24535_, _24414_);
  and (_28798_, _28788_, _28777_);
  and (_28809_, _28798_, _25388_);
  nand (_28820_, _28809_, _28766_);
  and (_28831_, _28188_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_28842_, _28809_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_28853_, _28842_, _28831_);
  and (_28864_, _28853_, _28820_);
  or (_28875_, _28864_, _28253_);
  or (_28886_, _28875_, _28252_);
  and (_06703_, _28886_, _42003_);
  and (_28907_, _23556_, _21123_);
  not (_28917_, _28907_);
  and (_28928_, _26226_, _26203_);
  nor (_28939_, _28928_, _26237_);
  and (_28950_, _28939_, _25465_);
  not (_28971_, _28950_);
  and (_28972_, _27272_, _25443_);
  not (_28983_, _28972_);
  nor (_28994_, _28983_, _18882_);
  and (_29005_, _28646_, _18283_);
  nor (_29016_, _29005_, _28994_);
  and (_29027_, _27391_, _25704_);
  and (_29037_, _27413_, _19428_);
  nor (_29048_, _29037_, _29027_);
  nor (_29059_, _27816_, _16492_);
  and (_29070_, _27532_, _19428_);
  nor (_29081_, _29070_, _29059_);
  nor (_29092_, _27446_, _27849_);
  nor (_29103_, _29092_, _19428_);
  not (_29114_, _29103_);
  and (_29125_, _29114_, _29081_);
  and (_29136_, _29125_, _29048_);
  and (_29146_, _29136_, _29016_);
  and (_29157_, _20847_, _15770_);
  and (_29168_, _28939_, _26563_);
  nor (_29179_, _28569_, _26203_);
  not (_29190_, _29179_);
  nor (_29201_, _28450_, _25704_);
  nor (_29212_, _29201_, _27206_);
  or (_29223_, _29212_, _26204_);
  nand (_29233_, _29223_, _29190_);
  or (_29244_, _29233_, _29168_);
  nor (_29255_, _29244_, _29157_);
  and (_29266_, _29255_, _29146_);
  and (_29277_, _29266_, _28971_);
  and (_29288_, _29277_, _28917_);
  not (_29299_, _29288_);
  or (_29310_, _29299_, _25399_);
  not (_29320_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_29331_, _25399_, _29320_);
  and (_29342_, _29331_, _28199_);
  and (_29353_, _29342_, _29310_);
  nor (_29364_, _28188_, _29320_);
  not (_29375_, _28766_);
  or (_29386_, _29375_, _25399_);
  and (_29397_, _29331_, _28831_);
  and (_29407_, _29397_, _29386_);
  or (_29418_, _29407_, _29364_);
  or (_29429_, _29418_, _29353_);
  and (_08941_, _29429_, _42003_);
  and (_29450_, _20878_, _15770_);
  not (_29461_, _29450_);
  and (_29472_, _23621_, _21123_);
  nor (_29483_, _27816_, _17478_);
  nor (_29493_, _27631_, _27533_);
  not (_29514_, _29493_);
  nor (_29515_, _29514_, _26203_);
  and (_29526_, _29514_, _26203_);
  nor (_29537_, _29526_, _29515_);
  and (_29548_, _29537_, _27532_);
  nor (_29559_, _29548_, _29483_);
  nor (_29570_, _27882_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29580_, _29570_, _19090_);
  nor (_29591_, _29570_, _19090_);
  nor (_29602_, _29591_, _29580_);
  nor (_29613_, _29602_, _27860_);
  not (_29624_, _29613_);
  and (_29635_, _27239_, _25726_);
  nor (_29646_, _27217_, _25715_);
  not (_29657_, _29646_);
  and (_29667_, _27391_, _25693_);
  and (_29678_, _27413_, _18882_);
  nor (_29689_, _29678_, _29667_);
  nand (_29700_, _29689_, _29657_);
  nor (_29711_, _29700_, _29635_);
  nor (_29722_, _28983_, _19046_);
  not (_29733_, _29722_);
  nor (_29744_, _27457_, _18882_);
  nor (_29754_, _27326_, _19428_);
  nor (_29775_, _29754_, _29744_);
  and (_29776_, _29775_, _29733_);
  and (_29787_, _29776_, _29711_);
  and (_29798_, _29787_, _29624_);
  and (_29809_, _29798_, _29559_);
  nor (_29820_, _25726_, _25704_);
  or (_29830_, _29820_, _25746_);
  and (_29841_, _29830_, _26237_);
  nor (_29852_, _29830_, _26237_);
  or (_29863_, _29852_, _29841_);
  and (_29874_, _29863_, _25465_);
  nor (_29885_, _26988_, _26955_);
  nor (_29896_, _29885_, _26999_);
  nor (_29907_, _29896_, _26574_);
  nor (_29918_, _29907_, _29874_);
  and (_29928_, _29918_, _29809_);
  not (_29939_, _29928_);
  nor (_29950_, _29939_, _29472_);
  and (_29961_, _29950_, _29461_);
  not (_29972_, _29961_);
  or (_29983_, _29972_, _25399_);
  not (_29994_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_30005_, _25399_, _29994_);
  and (_30015_, _30005_, _28199_);
  and (_30026_, _30015_, _29983_);
  nor (_30037_, _28188_, _29994_);
  not (_30048_, _24535_);
  and (_30059_, _30048_, _24414_);
  and (_30080_, _30059_, _24293_);
  and (_30081_, _30080_, _25388_);
  or (_30092_, _30081_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30102_, _30092_, _28831_);
  nand (_30113_, _30081_, _28766_);
  and (_30124_, _30113_, _30102_);
  or (_30135_, _30124_, _30037_);
  or (_30146_, _30135_, _30026_);
  and (_08952_, _30146_, _42003_);
  and (_30167_, _20910_, _15770_);
  not (_30178_, _30167_);
  and (_30188_, _23686_, _21123_);
  nor (_30199_, _27816_, _16163_);
  and (_30210_, _27533_, _26203_);
  and (_30221_, _27631_, _27609_);
  nor (_30232_, _30221_, _30210_);
  and (_30243_, _30232_, _19046_);
  nor (_30254_, _30232_, _19046_);
  nor (_30265_, _30254_, _30243_);
  and (_30275_, _30265_, _27532_);
  nor (_30286_, _30275_, _30199_);
  nor (_30297_, _26999_, _26944_);
  nor (_30308_, _30297_, _27010_);
  nor (_30319_, _30308_, _26574_);
  and (_30330_, _27239_, _25671_);
  nor (_30341_, _27217_, _25660_);
  not (_30352_, _30341_);
  and (_30362_, _27391_, _25650_);
  and (_30373_, _27413_, _19046_);
  nor (_30384_, _30373_, _30362_);
  nand (_30405_, _30384_, _30352_);
  nor (_30406_, _30405_, _30330_);
  nor (_30417_, _27326_, _18882_);
  not (_30428_, _30417_);
  nor (_30438_, _27457_, _19046_);
  nor (_30449_, _28983_, _18544_);
  nor (_30460_, _30449_, _30438_);
  and (_30472_, _30460_, _30428_);
  and (_30493_, _30472_, _30406_);
  not (_30504_, _30493_);
  nor (_30515_, _30504_, _30319_);
  nor (_30526_, _26269_, _26248_);
  nor (_30536_, _30526_, _28264_);
  and (_30547_, _30536_, _26291_);
  nor (_30558_, _29591_, _19046_);
  and (_30569_, _27871_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30580_, _30569_, _30558_);
  nor (_30591_, _30580_, _27860_);
  nor (_30602_, _30591_, _30547_);
  and (_30613_, _30602_, _30515_);
  and (_30624_, _30613_, _30286_);
  not (_30634_, _30624_);
  nor (_30645_, _30634_, _30188_);
  and (_30656_, _30645_, _30178_);
  not (_30667_, _30656_);
  or (_30678_, _30667_, _25399_);
  not (_30689_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_30700_, _25399_, _30689_);
  and (_30711_, _30700_, _28199_);
  and (_30721_, _30711_, _30678_);
  nor (_30732_, _28188_, _30689_);
  nand (_30743_, _25388_, _24293_);
  or (_30754_, _28788_, _30743_);
  and (_30765_, _30754_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_30776_, _24414_);
  and (_30787_, _24293_, _24535_);
  and (_30798_, _30787_, _30776_);
  and (_30808_, _30798_, _29375_);
  and (_30819_, _24293_, _24414_);
  and (_30830_, _30819_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_30841_, _30830_, _30808_);
  and (_30852_, _30841_, _25388_);
  or (_30863_, _30852_, _30765_);
  and (_30874_, _30863_, _28831_);
  or (_30894_, _30874_, _30732_);
  or (_30895_, _30894_, _30721_);
  and (_08963_, _30895_, _42003_);
  and (_30916_, _23751_, _21123_);
  not (_30927_, _30916_);
  and (_30938_, _20953_, _15770_);
  nor (_30949_, _27010_, _26912_);
  nor (_30960_, _30949_, _27021_);
  nor (_30971_, _30960_, _26574_);
  not (_30981_, _30971_);
  and (_30992_, _26291_, _25802_);
  or (_31003_, _30992_, _28264_);
  nor (_31014_, _31003_, _26302_);
  not (_31025_, _31014_);
  nor (_31036_, _27816_, _17162_);
  nor (_31047_, _27642_, _26203_);
  nor (_31057_, _27544_, _27609_);
  nor (_31068_, _31057_, _31047_);
  and (_31079_, _31068_, _18555_);
  not (_31090_, _27532_);
  nor (_31101_, _31068_, _18555_);
  or (_31122_, _31101_, _31090_);
  nor (_31123_, _31122_, _31079_);
  nor (_31134_, _31123_, _31036_);
  not (_31144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_31155_, _27871_, _31144_);
  nor (_31166_, _31155_, _18555_);
  nor (_31177_, _27457_, _18544_);
  nor (_31188_, _27882_, _27860_);
  nor (_31199_, _31188_, _31177_);
  nor (_31210_, _31199_, _31166_);
  not (_31221_, _31210_);
  nor (_31231_, _27217_, _25628_);
  and (_31242_, _27239_, _25639_);
  nor (_31253_, _31242_, _31231_);
  and (_31264_, _27391_, _25617_);
  and (_31275_, _27413_, _18544_);
  nor (_31286_, _31275_, _31264_);
  nor (_31297_, _28983_, _18174_);
  nor (_31308_, _27326_, _19046_);
  nor (_31318_, _31308_, _31297_);
  and (_31329_, _31318_, _31286_);
  and (_31340_, _31329_, _31253_);
  and (_31351_, _31340_, _31221_);
  and (_31362_, _31351_, _31134_);
  and (_31373_, _31362_, _31025_);
  and (_31384_, _31373_, _30981_);
  not (_31395_, _31384_);
  nor (_31405_, _31395_, _30938_);
  and (_31416_, _31405_, _30927_);
  not (_31427_, _31416_);
  or (_31438_, _31427_, _25399_);
  not (_31449_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_31460_, _25399_, _31449_);
  and (_31471_, _31460_, _28199_);
  and (_31482_, _31471_, _31438_);
  nor (_31492_, _28188_, _31449_);
  and (_31503_, _30743_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_31514_, _28788_, _24293_);
  not (_31525_, _31514_);
  nor (_31536_, _31525_, _28766_);
  nor (_31547_, _30819_, _30787_);
  nor (_31558_, _31547_, _31449_);
  or (_31569_, _31558_, _31536_);
  and (_31579_, _31569_, _25388_);
  or (_31590_, _31579_, _31503_);
  and (_31601_, _31590_, _28831_);
  or (_31612_, _31601_, _31492_);
  or (_31623_, _31612_, _31482_);
  and (_08974_, _31623_, _42003_);
  and (_31644_, _23816_, _21123_);
  not (_31655_, _31644_);
  and (_31665_, _20984_, _15770_);
  nor (_31676_, _27086_, _25606_);
  and (_31697_, _27086_, _25606_);
  nor (_31698_, _31697_, _31676_);
  and (_31709_, _31698_, _26563_);
  or (_31720_, _26335_, _25606_);
  nor (_31731_, _28264_, _26346_);
  and (_31742_, _31731_, _31720_);
  and (_31752_, _27555_, _26203_);
  and (_31763_, _27653_, _27609_);
  nor (_31774_, _31763_, _31752_);
  nor (_31785_, _31774_, _18174_);
  and (_31796_, _31774_, _18174_);
  or (_31807_, _31796_, _31090_);
  nor (_31818_, _31807_, _31785_);
  and (_31829_, _26203_, _18185_);
  nor (_31839_, _26203_, _16328_);
  or (_31850_, _31839_, _31829_);
  and (_31861_, _31850_, _27795_);
  and (_31872_, _27391_, _25530_);
  and (_31883_, _27413_, _18174_);
  nor (_31894_, _31883_, _31872_);
  not (_31905_, _31894_);
  and (_31916_, _27239_, _25606_);
  nor (_31926_, _27217_, _25595_);
  or (_31937_, _31926_, _31916_);
  nor (_31948_, _31937_, _31905_);
  not (_31959_, _31948_);
  or (_31970_, _31959_, _31861_);
  or (_31981_, _31970_, _31818_);
  or (_31992_, _27893_, _18185_);
  nor (_32003_, _27457_, _18174_);
  nor (_32013_, _27904_, _27860_);
  or (_32024_, _32013_, _32003_);
  and (_32035_, _32024_, _31992_);
  nor (_32046_, _28983_, _18011_);
  nor (_32057_, _27326_, _18544_);
  or (_32068_, _32057_, _32046_);
  or (_32079_, _32068_, _32035_);
  or (_32090_, _32079_, _31981_);
  or (_32100_, _32090_, _31742_);
  or (_32111_, _32100_, _31709_);
  nor (_32122_, _32111_, _31665_);
  and (_32133_, _32122_, _31655_);
  not (_32144_, _32133_);
  or (_32155_, _32144_, _25399_);
  not (_32166_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_32177_, _25399_, _32166_);
  and (_32187_, _32177_, _28199_);
  and (_32198_, _32187_, _32155_);
  nor (_32209_, _28188_, _32166_);
  not (_32220_, _25388_);
  and (_32231_, _24546_, _28777_);
  nor (_32242_, _24546_, _28777_);
  nor (_32253_, _32242_, _32231_);
  or (_32264_, _32253_, _32220_);
  and (_32275_, _32264_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_32286_, _32231_, _29375_);
  and (_32297_, _32242_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_32308_, _32297_, _32286_);
  and (_32329_, _32308_, _25388_);
  or (_32330_, _32329_, _32275_);
  and (_32341_, _32330_, _28831_);
  or (_32352_, _32341_, _32209_);
  or (_32363_, _32352_, _32198_);
  and (_08985_, _32363_, _42003_);
  and (_32384_, _21027_, _15770_);
  not (_32395_, _32384_);
  and (_32406_, _23903_, _21123_);
  nor (_32417_, _26367_, _26346_);
  not (_32428_, _32417_);
  nor (_32439_, _28264_, _26378_);
  and (_32449_, _32439_, _32428_);
  not (_32460_, _32449_);
  nor (_32471_, _27097_, _26748_);
  nor (_32482_, _32471_, _27108_);
  nor (_32493_, _32482_, _26574_);
  nor (_32504_, _26203_, _17314_);
  and (_32515_, _26203_, _18588_);
  nor (_32526_, _32515_, _32504_);
  nor (_32537_, _32526_, _27816_);
  nor (_32548_, _27566_, _27609_);
  nor (_32559_, _27664_, _26203_);
  nor (_32570_, _32559_, _32548_);
  and (_32581_, _32570_, _18588_);
  nor (_32592_, _32570_, _18588_);
  or (_32603_, _32592_, _31090_);
  nor (_32614_, _32603_, _32581_);
  nor (_32635_, _32614_, _32537_);
  not (_32636_, _27958_);
  and (_32647_, _32636_, _27915_);
  nor (_32658_, _27958_, _27904_);
  nor (_32669_, _32658_, _18011_);
  nor (_32680_, _32669_, _32647_);
  nor (_32691_, _32680_, _27860_);
  nor (_32702_, _27217_, _25551_);
  and (_32713_, _27239_, _25552_);
  nor (_32724_, _32713_, _32702_);
  and (_32735_, _27391_, _25519_);
  and (_32746_, _27413_, _18011_);
  nor (_32757_, _32746_, _32735_);
  nor (_32768_, _27326_, _18174_);
  not (_32779_, _32768_);
  nor (_32790_, _27457_, _18011_);
  nor (_32801_, _28983_, _16987_);
  nor (_32812_, _32801_, _32790_);
  and (_32823_, _32812_, _32779_);
  and (_32834_, _32823_, _32757_);
  and (_32845_, _32834_, _32724_);
  not (_32855_, _32845_);
  nor (_32866_, _32855_, _32691_);
  and (_32877_, _32866_, _32635_);
  not (_32888_, _32877_);
  nor (_32899_, _32888_, _32493_);
  and (_32910_, _32899_, _32460_);
  not (_32921_, _32910_);
  nor (_32932_, _32921_, _32406_);
  and (_32943_, _32932_, _32395_);
  not (_32954_, _32943_);
  or (_32965_, _32954_, _25399_);
  not (_32986_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_32987_, _25399_, _32986_);
  and (_32998_, _32987_, _28199_);
  and (_33009_, _32998_, _32965_);
  nor (_33020_, _28188_, _32986_);
  and (_33031_, _30059_, _28777_);
  and (_33042_, _33031_, _25388_);
  nand (_33053_, _33042_, _28766_);
  or (_33064_, _33042_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_33075_, _33064_, _28831_);
  and (_33086_, _33075_, _33053_);
  or (_33097_, _33086_, _33020_);
  or (_33108_, _33097_, _33009_);
  and (_08996_, _33108_, _42003_);
  and (_33129_, _23968_, _21123_);
  not (_33140_, _33129_);
  and (_33151_, _21059_, _15770_);
  nor (_33162_, _26400_, _26378_);
  not (_33173_, _33162_);
  nor (_33184_, _28264_, _26411_);
  and (_33195_, _33184_, _33173_);
  not (_33206_, _33195_);
  nor (_33217_, _27108_, _26715_);
  nor (_33227_, _33217_, _27119_);
  nor (_33238_, _33227_, _26574_);
  nor (_33249_, _26203_, _26585_);
  or (_33260_, _33249_, _27816_);
  nor (_33271_, _33260_, _28341_);
  nor (_33282_, _26203_, _18588_);
  nand (_33293_, _33282_, _27664_);
  nand (_33304_, _27577_, _26203_);
  and (_33315_, _33304_, _33293_);
  and (_33326_, _33315_, _16987_);
  nor (_33337_, _33315_, _16987_);
  or (_33358_, _33337_, _31090_);
  nor (_33359_, _33358_, _33326_);
  nor (_33370_, _33359_, _33271_);
  nor (_33381_, _32647_, _16987_);
  and (_33392_, _32647_, _16987_);
  nor (_33403_, _33392_, _33381_);
  nor (_33414_, _33403_, _27860_);
  and (_33425_, _27239_, _25497_);
  nor (_33436_, _27217_, _25486_);
  not (_33447_, _33436_);
  and (_33458_, _27391_, _25476_);
  and (_33469_, _27413_, _16987_);
  nor (_33480_, _33469_, _33458_);
  nand (_33491_, _33480_, _33447_);
  nor (_33502_, _33491_, _33425_);
  nor (_33513_, _28983_, _17826_);
  not (_33524_, _33513_);
  nor (_33535_, _27457_, _16987_);
  nor (_33546_, _27326_, _18011_);
  nor (_33557_, _33546_, _33535_);
  and (_33568_, _33557_, _33524_);
  and (_33579_, _33568_, _33502_);
  not (_33589_, _33579_);
  nor (_33600_, _33589_, _33414_);
  and (_33611_, _33600_, _33370_);
  not (_33622_, _33611_);
  nor (_33633_, _33622_, _33238_);
  and (_33644_, _33633_, _33206_);
  not (_33655_, _33644_);
  nor (_33666_, _33655_, _33151_);
  and (_33677_, _33666_, _33140_);
  not (_33688_, _33677_);
  or (_33699_, _33688_, _25399_);
  not (_33710_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_33721_, _25399_, _33710_);
  and (_33732_, _33721_, _28199_);
  and (_33743_, _33732_, _33699_);
  nor (_33754_, _28188_, _33710_);
  nor (_33765_, _24293_, _24414_);
  and (_33776_, _33765_, _24535_);
  and (_33787_, _33776_, _25388_);
  nand (_33798_, _33787_, _28766_);
  or (_33809_, _33787_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_33820_, _33809_, _28831_);
  and (_33831_, _33820_, _33798_);
  or (_33842_, _33831_, _33754_);
  or (_33853_, _33842_, _33743_);
  and (_09006_, _33853_, _42003_);
  and (_33884_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_33885_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_33896_, _33885_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33907_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_33918_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_33929_, _33918_, _33907_);
  and (_33939_, _33885_, _15704_);
  and (_33950_, _33939_, _33929_);
  not (_33961_, _33950_);
  and (_33972_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_33983_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_33994_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_34005_, _33994_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34016_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34027_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_34038_, _34027_, _34016_);
  and (_34049_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_34060_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_34071_, _34060_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34082_, _34071_, _34016_);
  and (_34093_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_34104_, _34093_, _34049_);
  and (_34115_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34126_, _34115_, _34016_);
  and (_34137_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_34158_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34159_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34158_);
  and (_34170_, _34159_, _34016_);
  and (_34181_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34192_, _34181_, _34137_);
  and (_34203_, _34027_, _34016_);
  and (_34214_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_34225_, _34027_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34236_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34247_, _34236_, _34214_);
  and (_34258_, _34247_, _34192_);
  and (_34269_, _34258_, _34104_);
  nor (_34280_, _34269_, _34005_);
  nor (_34291_, _34280_, _33983_);
  nor (_34302_, _34291_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34312_, _34302_, _33972_);
  nor (_34323_, _34312_, _33961_);
  and (_34334_, _33929_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34345_, _34334_, _33961_);
  nor (_34356_, _34345_, _34323_);
  and (_34367_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34378_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34389_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34400_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_34411_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34422_, _34411_, _34400_);
  and (_34433_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34444_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34455_, _34444_, _34433_);
  and (_34466_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_34477_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34488_, _34477_, _34466_);
  and (_34499_, _34488_, _34455_);
  and (_34510_, _34499_, _34422_);
  nor (_34521_, _34510_, _33994_);
  and (_34532_, _34521_, _34389_);
  nor (_34543_, _34532_, _34378_);
  nor (_34554_, _34543_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34565_, _34554_, _34367_);
  nor (_34576_, _34565_, _33961_);
  and (_34587_, _33929_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34598_, _34587_, _33961_);
  nor (_34609_, _34598_, _34576_);
  not (_34620_, _34609_);
  and (_34631_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34642_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34653_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34664_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_34674_, _34664_, _34653_);
  and (_34685_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_34696_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34707_, _34696_, _34685_);
  and (_34718_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_34729_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_34740_, _34729_, _34718_);
  and (_34751_, _34740_, _34707_);
  and (_34762_, _34751_, _34674_);
  nor (_34783_, _34762_, _34005_);
  nor (_34784_, _34783_, _34642_);
  nor (_34795_, _34784_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34806_, _34795_, _34631_);
  nor (_34817_, _34806_, _33961_);
  and (_34828_, _33929_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34839_, _34828_, _33961_);
  nor (_34850_, _34839_, _34817_);
  nor (_34861_, _34850_, _34620_);
  and (_34872_, _34861_, _34356_);
  and (_34883_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_34894_, _34883_);
  and (_34905_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_34916_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_34927_, _34916_, _34905_);
  and (_34938_, _34927_, _34894_);
  and (_34949_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_34960_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_34971_, _34960_, _34949_);
  and (_34982_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34993_, _33994_, _34982_);
  and (_35004_, _34993_, _34971_);
  and (_35015_, _35004_, _34938_);
  and (_35026_, _35015_, _34389_);
  nor (_35036_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34389_);
  nor (_35047_, _35036_, _35026_);
  nor (_35058_, _35047_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_35069_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35080_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _35069_);
  nor (_35091_, _35080_, _35058_);
  and (_35102_, _35091_, _33950_);
  and (_35113_, _33929_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_35124_, _35113_, _33961_);
  nor (_35135_, _35124_, _35102_);
  and (_35146_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35157_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35168_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_35179_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_35190_, _35179_, _35168_);
  and (_35201_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_35212_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_35223_, _35212_, _35201_);
  and (_35234_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_35245_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_35256_, _35245_, _35234_);
  and (_35267_, _35256_, _35223_);
  and (_35278_, _35267_, _35190_);
  nor (_35289_, _35278_, _34005_);
  nor (_35300_, _35289_, _35157_);
  nor (_35311_, _35300_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35322_, _35311_, _35146_);
  nor (_35333_, _35322_, _33961_);
  and (_35344_, _33929_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_35355_, _35344_, _33961_);
  nor (_35366_, _35355_, _35333_);
  nor (_35376_, _35366_, _35135_);
  and (_35387_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35398_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35409_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_35420_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_35431_, _35420_, _35409_);
  and (_35442_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_35453_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_35464_, _35453_, _35442_);
  and (_35475_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_35497_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_35498_, _35497_, _35475_);
  and (_35520_, _35498_, _35464_);
  and (_35521_, _35520_, _35431_);
  nor (_35543_, _35521_, _33994_);
  and (_35544_, _35543_, _34389_);
  or (_35566_, _35544_, _35398_);
  and (_35567_, _35566_, _35069_);
  nor (_35578_, _35567_, _35387_);
  nor (_35589_, _35578_, _33961_);
  and (_35600_, _33929_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_35611_, _35600_, _33961_);
  nor (_35622_, _35611_, _35589_);
  and (_35633_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_35644_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_35655_, _35644_, _35633_);
  and (_35666_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_35677_, _35666_, _33994_);
  and (_35688_, _35677_, _35655_);
  and (_35699_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_35709_, _35699_);
  and (_35720_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_35731_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_35742_, _35731_, _35720_);
  and (_35753_, _35742_, _35709_);
  and (_35764_, _35753_, _35688_);
  and (_35775_, _35764_, _34389_);
  nor (_35786_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34389_);
  or (_35797_, _35786_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35808_, _35797_, _35775_);
  and (_35819_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_35830_, _35819_, _35808_);
  and (_35841_, _35830_, _33950_);
  and (_35852_, _33929_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_35863_, _35852_, _33961_);
  nor (_35874_, _35863_, _35841_);
  not (_35885_, _35874_);
  and (_35896_, _35885_, _35622_);
  and (_35907_, _35896_, _35376_);
  and (_35918_, _35907_, _34872_);
  and (_35929_, _35376_, _35622_);
  and (_35940_, _34850_, _34356_);
  and (_35951_, _35940_, _34620_);
  and (_35962_, _35951_, _35929_);
  or (_35973_, _35962_, _35918_);
  not (_35984_, _35973_);
  and (_35995_, _35940_, _34609_);
  and (_36006_, _35995_, _35929_);
  not (_36016_, _34356_);
  and (_36027_, _34850_, _36016_);
  and (_36038_, _36027_, _34620_);
  and (_36049_, _36038_, _35907_);
  nor (_36060_, _36049_, _36006_);
  not (_36071_, _36060_);
  and (_36082_, _36027_, _34609_);
  and (_36093_, _36082_, _35874_);
  and (_36104_, _36093_, _35929_);
  nor (_36115_, _36104_, _36071_);
  and (_36126_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36137_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_36148_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_36159_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_36170_, _36159_, _36148_);
  and (_36181_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_36192_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_36203_, _36192_, _36181_);
  and (_36214_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_36225_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_36236_, _36225_, _36214_);
  and (_36247_, _36236_, _36203_);
  and (_36258_, _36247_, _36170_);
  nor (_36269_, _36258_, _33994_);
  and (_36280_, _36269_, _34389_);
  nor (_36291_, _36280_, _36137_);
  nor (_36302_, _36291_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36313_, _36302_, _36126_);
  nor (_36324_, _36313_, _33961_);
  and (_36334_, _33929_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_36345_, _36334_, _33961_);
  nor (_36356_, _36345_, _36324_);
  not (_36367_, _35135_);
  and (_36378_, _35622_, _35366_);
  and (_36389_, _36378_, _36367_);
  and (_36400_, _36389_, _36356_);
  and (_36411_, _36400_, _35951_);
  not (_36422_, _36411_);
  and (_36433_, _34861_, _36016_);
  and (_36444_, _36433_, _35929_);
  and (_36455_, _36082_, _35885_);
  and (_36466_, _36455_, _35929_);
  nor (_36477_, _36466_, _36444_);
  and (_36488_, _36477_, _36422_);
  and (_36499_, _36488_, _36115_);
  and (_36510_, _36499_, _35984_);
  not (_36521_, _36356_);
  and (_36532_, _36389_, _36521_);
  and (_36543_, _36038_, _35874_);
  and (_36554_, _36543_, _36532_);
  and (_36565_, _36532_, _36455_);
  nor (_36576_, _34850_, _34609_);
  and (_36587_, _36576_, _34356_);
  and (_36598_, _36587_, _35885_);
  and (_36609_, _36598_, _36532_);
  or (_36620_, _36609_, _36565_);
  nor (_36631_, _36620_, _36554_);
  and (_36641_, _36356_, _35135_);
  and (_36652_, _36641_, _36378_);
  and (_36663_, _36433_, _35885_);
  and (_36674_, _36663_, _36652_);
  not (_36685_, _36674_);
  and (_36696_, _35874_, _35929_);
  and (_36707_, _36576_, _36016_);
  or (_36718_, _36707_, _34872_);
  and (_36729_, _36718_, _36696_);
  and (_36740_, _36587_, _35874_);
  and (_36751_, _36740_, _35929_);
  nor (_36762_, _36751_, _36729_);
  and (_36773_, _36762_, _36685_);
  and (_36784_, _36773_, _36631_);
  and (_36795_, _36784_, _36510_);
  nor (_36806_, _36795_, _33896_);
  not (_36817_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_36828_, _15704_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_36839_, _36828_, _36817_);
  and (_36850_, _36839_, _36587_);
  and (_36861_, _36850_, _36652_);
  and (_36872_, _36411_, _36828_);
  and (_36883_, _36872_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_36894_, _36883_, _36861_);
  nor (_36905_, _36894_, _36806_);
  nor (_36916_, _36905_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36927_, _36916_, _33884_);
  and (_36938_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36949_, _33896_);
  not (_36959_, _35366_);
  and (_36970_, _35622_, _36959_);
  nor (_36981_, _36356_, _36367_);
  and (_36992_, _36981_, _36970_);
  and (_37003_, _36027_, _35885_);
  and (_37014_, _37003_, _36992_);
  and (_37025_, _36707_, _35874_);
  and (_37036_, _37025_, _36992_);
  and (_37047_, _36038_, _36696_);
  or (_37058_, _37047_, _37036_);
  or (_37069_, _37058_, _37014_);
  and (_37080_, _34872_, _35885_);
  or (_37091_, _37080_, _35951_);
  and (_37102_, _36992_, _37091_);
  nor (_37113_, _35885_, _35622_);
  and (_37124_, _37113_, _36038_);
  and (_37135_, _35995_, _35874_);
  and (_37146_, _37135_, _36992_);
  or (_37157_, _37146_, _37124_);
  or (_37168_, _37157_, _36411_);
  or (_37179_, _37168_, _37102_);
  and (_37190_, _36992_, _36740_);
  and (_37201_, _36433_, _35874_);
  and (_37212_, _37201_, _36992_);
  or (_37223_, _37212_, _37190_);
  and (_37234_, _36543_, _36400_);
  and (_37245_, _36663_, _36400_);
  nor (_37256_, _37245_, _37234_);
  not (_37264_, _37256_);
  or (_37271_, _37264_, _37223_);
  or (_37279_, _37271_, _37179_);
  or (_37287_, _37279_, _37069_);
  and (_37294_, _34872_, _35874_);
  and (_37302_, _37294_, _36389_);
  and (_37310_, _35995_, _35885_);
  and (_37317_, _37310_, _36992_);
  and (_37322_, _36038_, _35885_);
  and (_37323_, _36652_, _37322_);
  or (_37324_, _37323_, _37317_);
  nor (_37331_, _37324_, _37302_);
  and (_37342_, _36598_, _36400_);
  and (_37353_, _36992_, _36663_);
  nor (_37364_, _37353_, _37342_);
  and (_37375_, _37364_, _37331_);
  and (_37386_, _36652_, _36543_);
  and (_37397_, _37294_, _36992_);
  nor (_37408_, _37397_, _37386_);
  and (_37419_, _36400_, _37322_);
  and (_37430_, _37201_, _36400_);
  nor (_37441_, _37430_, _37419_);
  and (_37452_, _37441_, _37408_);
  and (_37463_, _37452_, _37375_);
  and (_37474_, _36455_, _36400_);
  and (_37485_, _36992_, _36093_);
  or (_37496_, _37485_, _37474_);
  and (_37507_, _36652_, _36433_);
  and (_37518_, _36740_, _36389_);
  or (_37529_, _37518_, _37507_);
  or (_37540_, _37529_, _37496_);
  and (_37551_, _36400_, _36093_);
  and (_37562_, _36389_, _37080_);
  or (_37573_, _37562_, _37551_);
  and (_37584_, _36652_, _35951_);
  and (_37595_, _37584_, _35874_);
  and (_37606_, _35885_, _35951_);
  or (_37617_, _37310_, _37606_);
  and (_37628_, _37617_, _36652_);
  nor (_37639_, _37628_, _37595_);
  not (_37650_, _37639_);
  or (_37661_, _37650_, _37573_);
  nor (_37672_, _37661_, _37540_);
  nand (_37683_, _37672_, _37463_);
  or (_37694_, _37683_, _37287_);
  and (_37705_, _37694_, _36949_);
  and (_37716_, _36828_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37727_, _37716_, _36411_);
  not (_37738_, _37727_);
  nor (_37749_, _34850_, _36016_);
  and (_37760_, _36652_, _37749_);
  and (_37771_, _37760_, _36839_);
  not (_37782_, _36839_);
  and (_37793_, _35874_, _35951_);
  and (_37804_, _37793_, _36652_);
  and (_37815_, _37310_, _36652_);
  nor (_37826_, _37815_, _37804_);
  nor (_37837_, _37826_, _37782_);
  nor (_37848_, _37837_, _37771_);
  and (_37859_, _37848_, _37738_);
  not (_37870_, _37859_);
  nor (_37881_, _37870_, _37705_);
  nor (_37892_, _37881_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37903_, _37892_, _36938_);
  nor (_37914_, _37903_, _36927_);
  and (_37925_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37936_, _36641_, _36970_);
  and (_37947_, _37936_, _36093_);
  and (_37958_, _37936_, _36543_);
  nor (_37969_, _37958_, _37947_);
  and (_37980_, _37969_, _36631_);
  nor (_37991_, _37980_, _33896_);
  not (_38002_, _33885_);
  and (_38013_, _37958_, _15704_);
  and (_38024_, _37947_, _15704_);
  or (_38035_, _38024_, _38013_);
  and (_38046_, _38035_, _38002_);
  or (_38057_, _38046_, _37771_);
  nor (_38068_, _38057_, _37991_);
  nor (_38079_, _38068_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38090_, _38079_, _37925_);
  and (_38101_, _38090_, _42003_);
  and (_09552_, _38101_, _37914_);
  and (_38122_, _28199_, _25213_);
  and (_38133_, _24886_, _24754_);
  and (_38144_, _38133_, _25344_);
  and (_38155_, _38144_, _25072_);
  and (_38166_, _38155_, _30080_);
  and (_38177_, _38166_, _38122_);
  not (_38188_, _38177_);
  and (_38199_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_38210_, _38155_, _25213_);
  and (_38221_, _38210_, _24293_);
  and (_38232_, _38221_, _30059_);
  and (_38243_, _38232_, _28199_);
  not (_38254_, _38243_);
  or (_38265_, _21123_, _15770_);
  and (_38276_, _25454_, _21101_);
  or (_38287_, _27315_, _27446_);
  or (_38298_, _38287_, _38276_);
  or (_38309_, _38298_, _38265_);
  nor (_38320_, _38309_, _28972_);
  nor (_38331_, _38320_, _16987_);
  not (_38342_, _38331_);
  and (_38353_, _38342_, _33502_);
  and (_38364_, _38353_, _33370_);
  nor (_38375_, _38364_, _38254_);
  nor (_38386_, _38375_, _38199_);
  and (_38397_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38408_, _38320_, _18011_);
  not (_38419_, _38408_);
  and (_38430_, _38419_, _32757_);
  and (_38441_, _38430_, _32724_);
  and (_38452_, _38441_, _32635_);
  nor (_38462_, _38452_, _38254_);
  nor (_38473_, _38462_, _38397_);
  and (_38484_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38495_, _38320_, _18174_);
  nor (_38506_, _38495_, _31981_);
  nor (_38517_, _38506_, _38254_);
  nor (_38528_, _38517_, _38484_);
  and (_38538_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38549_, _38320_, _18544_);
  not (_38560_, _38549_);
  and (_38570_, _38560_, _31286_);
  and (_38581_, _38570_, _31253_);
  and (_38592_, _38581_, _31134_);
  nor (_38596_, _38592_, _38254_);
  nor (_38602_, _38596_, _38538_);
  and (_38608_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38610_, _38320_, _19046_);
  not (_38611_, _38610_);
  and (_38612_, _38611_, _30406_);
  and (_38613_, _38612_, _30286_);
  nor (_38614_, _38613_, _38254_);
  nor (_38615_, _38614_, _38608_);
  and (_38616_, _38188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38617_, _38320_, _18882_);
  not (_38618_, _38617_);
  and (_38619_, _38618_, _29711_);
  and (_38620_, _38619_, _29559_);
  nor (_38621_, _38620_, _38188_);
  nor (_38622_, _38621_, _38616_);
  nor (_38623_, _38177_, _24480_);
  nor (_38624_, _38320_, _19428_);
  not (_38625_, _38624_);
  and (_38626_, _38625_, _29081_);
  and (_38627_, _38626_, _29048_);
  and (_38628_, _38627_, _29223_);
  not (_38629_, _38628_);
  and (_38630_, _38629_, _38177_);
  nor (_38631_, _38630_, _38623_);
  and (_38632_, _38631_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38633_, _38632_, _38622_);
  and (_38634_, _38633_, _38615_);
  and (_38635_, _38634_, _38602_);
  and (_38636_, _38635_, _38528_);
  and (_38637_, _38636_, _38473_);
  and (_38638_, _38637_, _38386_);
  nor (_38639_, _38177_, _24908_);
  and (_38640_, _38639_, _38638_);
  nor (_38641_, _38639_, _38638_);
  nor (_38642_, _38641_, _38640_);
  and (_38643_, _38642_, _24623_);
  nor (_38644_, _38177_, _24952_);
  not (_38645_, _38644_);
  nor (_38646_, _38645_, _38643_);
  nor (_38647_, _38320_, _17826_);
  not (_38648_, _38647_);
  and (_38649_, _38648_, _27435_);
  and (_38650_, _38649_, _27271_);
  and (_38651_, _38650_, _27838_);
  and (_38652_, _38651_, _38243_);
  nor (_38653_, _38652_, _38646_);
  and (_09573_, _38653_, _42003_);
  not (_38654_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38655_, _38631_, _38654_);
  nor (_38656_, _38631_, _38654_);
  nor (_38657_, _38656_, _38655_);
  and (_38658_, _38657_, _24623_);
  nor (_38659_, _38658_, _24491_);
  nor (_38660_, _38659_, _38243_);
  nor (_38661_, _38660_, _38630_);
  nand (_10699_, _38661_, _42003_);
  nor (_38662_, _38632_, _38622_);
  nor (_38663_, _38662_, _38633_);
  nor (_38664_, _38663_, _24022_);
  nor (_38665_, _38664_, _24326_);
  nor (_38666_, _38665_, _38243_);
  nor (_38667_, _38666_, _38621_);
  nand (_10710_, _38667_, _42003_);
  nor (_38668_, _38633_, _38615_);
  nor (_38669_, _38668_, _38634_);
  nor (_38670_, _38669_, _24022_);
  nor (_38671_, _38670_, _24077_);
  nor (_38672_, _38671_, _38243_);
  nor (_38673_, _38672_, _38614_);
  nand (_10721_, _38673_, _42003_);
  nor (_38674_, _38634_, _38602_);
  nor (_38675_, _38674_, _38635_);
  nor (_38676_, _38675_, _24022_);
  nor (_38677_, _38676_, _25158_);
  nor (_38678_, _38677_, _38243_);
  nor (_38679_, _38678_, _38596_);
  nor (_10731_, _38679_, rst);
  nor (_38680_, _38635_, _38528_);
  nor (_38681_, _38680_, _38636_);
  nor (_38682_, _38681_, _24022_);
  nor (_38683_, _38682_, _25246_);
  nor (_38684_, _38683_, _38243_);
  nor (_38685_, _38684_, _38517_);
  nor (_10742_, _38685_, rst);
  nor (_38686_, _38636_, _38473_);
  nor (_38687_, _38686_, _38637_);
  nor (_38688_, _38687_, _24022_);
  nor (_38689_, _38688_, _24798_);
  nor (_38690_, _38689_, _38243_);
  nor (_38691_, _38690_, _38462_);
  nor (_10753_, _38691_, rst);
  nor (_38692_, _38637_, _38386_);
  nor (_38693_, _38692_, _38638_);
  nor (_38694_, _38693_, _24022_);
  nor (_38695_, _38694_, _24656_);
  nor (_38696_, _38695_, _38243_);
  nor (_38697_, _38696_, _38375_);
  nor (_10764_, _38697_, rst);
  and (_38698_, _38122_, _31514_);
  nand (_38699_, _38698_, _38155_);
  nor (_38700_, _38699_, _28122_);
  and (_38701_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15704_);
  and (_38702_, _38701_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38703_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38704_, _38703_, _38702_);
  or (_38705_, _38704_, _38700_);
  nor (_38706_, _27457_, _17652_);
  nor (_38707_, _28569_, _18544_);
  and (_38708_, _26203_, _17314_);
  not (_38709_, _38708_);
  nor (_38710_, _17826_, _16492_);
  and (_38711_, _38710_, _27588_);
  and (_38712_, _38711_, _26803_);
  and (_38713_, _38712_, _26846_);
  and (_38714_, _38713_, _27032_);
  nor (_38715_, _38714_, _27609_);
  and (_38716_, _26203_, _16328_);
  nor (_38717_, _38716_, _38715_);
  and (_38718_, _38717_, _38709_);
  and (_38719_, _27675_, _17826_);
  and (_38720_, _17162_, _16163_);
  and (_38721_, _17478_, _16492_);
  and (_38722_, _38721_, _38720_);
  and (_38723_, _38722_, _38719_);
  and (_38724_, _17314_, _16328_);
  and (_38725_, _38724_, _38723_);
  nor (_38726_, _38725_, _26203_);
  not (_38727_, _38726_);
  and (_38728_, _38727_, _38718_);
  nor (_38729_, _26203_, _16669_);
  and (_38730_, _26203_, _16669_);
  nor (_38731_, _38730_, _38729_);
  and (_38732_, _38731_, _38728_);
  and (_38733_, _38732_, _27751_);
  nor (_38734_, _38732_, _27751_);
  nor (_38735_, _38734_, _38733_);
  and (_38736_, _38735_, _27532_);
  and (_38737_, _26203_, _27751_);
  nor (_38738_, _38737_, _28373_);
  nor (_38739_, _38738_, _27816_);
  or (_38740_, _38739_, _38736_);
  or (_38741_, _38740_, _38707_);
  and (_38742_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_38743_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38744_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38745_, _38744_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38746_, _38745_, _38743_);
  nor (_38747_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38748_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38749_, _38748_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38750_, _38749_, _38747_);
  nor (_38751_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38752_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38753_, _38752_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38754_, _38753_, _38751_);
  not (_38755_, _38754_);
  nor (_38756_, _38755_, _28275_);
  nor (_38757_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38758_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38759_, _38758_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38760_, _38759_, _38757_);
  and (_38761_, _38760_, _38756_);
  nor (_38762_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38763_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38764_, _38763_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38765_, _38764_, _38762_);
  and (_38766_, _38765_, _38761_);
  and (_38767_, _38766_, _38750_);
  nor (_38768_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38769_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38770_, _38769_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38771_, _38770_, _38768_);
  and (_38772_, _38771_, _38767_);
  and (_38773_, _38772_, _38746_);
  nor (_38774_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38775_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38776_, _38775_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38777_, _38776_, _38774_);
  and (_38778_, _38777_, _38773_);
  nor (_38779_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38780_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38781_, _38780_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38782_, _38781_, _38779_);
  or (_38783_, _38782_, _38778_);
  nand (_38784_, _38782_, _38778_);
  and (_38785_, _38784_, _25465_);
  and (_38786_, _38785_, _38783_);
  and (_38787_, _20815_, _15770_);
  or (_38788_, _38787_, _38786_);
  or (_38789_, _38788_, _38742_);
  or (_38790_, _38789_, _38741_);
  nor (_38791_, _38790_, _38706_);
  nand (_38792_, _38791_, _38702_);
  and (_38793_, _38792_, _42003_);
  and (_12710_, _38793_, _38705_);
  and (_38794_, _38122_, _30798_);
  and (_38795_, _38794_, _38155_);
  nor (_38796_, _38795_, _38702_);
  not (_38797_, _38796_);
  nand (_38798_, _38797_, _28122_);
  not (_38799_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_38800_, _38796_, _38799_);
  and (_38801_, _38800_, _42003_);
  and (_12731_, _38801_, _38798_);
  nor (_38802_, _38699_, _29288_);
  and (_38803_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38804_, _38803_, _38702_);
  or (_38805_, _38804_, _38802_);
  and (_38806_, _23419_, _21123_);
  and (_38807_, _38755_, _28275_);
  nor (_38808_, _38807_, _38756_);
  and (_38809_, _38808_, _25465_);
  nor (_38810_, _27457_, _16492_);
  and (_38811_, _20593_, _15770_);
  nor (_38812_, _28569_, _18174_);
  nor (_38813_, _27816_, _19428_);
  or (_38814_, _38813_, _38812_);
  or (_38815_, _38814_, _38811_);
  nor (_38816_, _38815_, _38810_);
  nor (_38817_, _28373_, _27784_);
  not (_38818_, _38817_);
  nor (_38819_, _38818_, _27697_);
  nor (_38820_, _38819_, _26770_);
  and (_38821_, _38819_, _26770_);
  or (_38822_, _38821_, _31090_);
  or (_38823_, _38822_, _38820_);
  and (_38824_, _38823_, _38816_);
  not (_38825_, _38824_);
  nor (_38826_, _38825_, _38809_);
  not (_38827_, _38826_);
  nor (_38828_, _38827_, _38806_);
  nand (_38829_, _38828_, _38702_);
  and (_38830_, _38829_, _42003_);
  and (_13625_, _38830_, _38805_);
  nor (_38831_, _38699_, _29961_);
  and (_38832_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38833_, _38832_, _38702_);
  or (_38834_, _38833_, _38831_);
  nor (_38835_, _27457_, _17478_);
  nor (_38836_, _28569_, _18011_);
  and (_38837_, _38711_, _26203_);
  and (_38838_, _38719_, _16492_);
  and (_38839_, _38838_, _27609_);
  nor (_38840_, _38839_, _38837_);
  and (_38841_, _38840_, _17478_);
  nor (_38842_, _38840_, _17478_);
  or (_38843_, _38842_, _31090_);
  nor (_38844_, _38843_, _38841_);
  nor (_38845_, _27816_, _18882_);
  or (_38846_, _38845_, _38844_);
  or (_38847_, _38846_, _38836_);
  and (_38848_, _22414_, _21123_);
  nor (_38849_, _38760_, _38756_);
  nor (_38850_, _38849_, _38761_);
  and (_38851_, _38850_, _25465_);
  and (_38852_, _20625_, _15770_);
  or (_38853_, _38852_, _38851_);
  or (_38854_, _38853_, _38848_);
  or (_38855_, _38854_, _38847_);
  nor (_38856_, _38855_, _38835_);
  nand (_38857_, _38856_, _38702_);
  and (_38858_, _38857_, _42003_);
  and (_13634_, _38858_, _38834_);
  nor (_38859_, _38699_, _30656_);
  and (_38860_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38861_, _38860_, _38702_);
  or (_38862_, _38861_, _38859_);
  nor (_38863_, _27457_, _16163_);
  nor (_38864_, _28569_, _16987_);
  and (_38865_, _38838_, _17478_);
  and (_38866_, _38865_, _27609_);
  and (_38867_, _38712_, _26203_);
  nor (_38868_, _38867_, _38866_);
  and (_38869_, _38868_, _16163_);
  nor (_38870_, _38868_, _16163_);
  nor (_38871_, _38870_, _38869_);
  and (_38872_, _38871_, _27532_);
  nor (_38873_, _27816_, _19046_);
  or (_38874_, _38873_, _38872_);
  or (_38875_, _38874_, _38864_);
  and (_38876_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38877_, _38765_, _38761_);
  nor (_38878_, _38877_, _38766_);
  and (_38879_, _38878_, _25465_);
  and (_38880_, _20656_, _15770_);
  or (_38881_, _38880_, _38879_);
  or (_38882_, _38881_, _38876_);
  or (_38883_, _38882_, _38875_);
  nor (_38884_, _38883_, _38863_);
  nand (_38885_, _38884_, _38702_);
  and (_38886_, _38885_, _42003_);
  and (_13644_, _38886_, _38862_);
  nor (_38887_, _38699_, _31416_);
  and (_38888_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38889_, _38888_, _38702_);
  or (_38890_, _38889_, _38887_);
  nor (_38891_, _27457_, _17162_);
  nor (_38892_, _38713_, _27032_);
  not (_38893_, _38892_);
  and (_38894_, _38893_, _38715_);
  and (_38895_, _38865_, _16163_);
  nor (_38896_, _38895_, _17162_);
  nor (_38897_, _38896_, _38723_);
  nor (_38898_, _38897_, _26203_);
  nor (_38899_, _38898_, _38894_);
  nor (_38900_, _38899_, _31090_);
  nor (_38901_, _27816_, _18544_);
  or (_38902_, _38901_, _38900_);
  or (_38903_, _38902_, _28580_);
  and (_38904_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_38905_, _38766_, _38750_);
  not (_38906_, _38905_);
  nor (_38907_, _38767_, _28264_);
  and (_38908_, _38907_, _38906_);
  and (_38909_, _20688_, _15770_);
  or (_38910_, _38909_, _38908_);
  or (_38911_, _38910_, _38904_);
  or (_38912_, _38911_, _38903_);
  nor (_38913_, _38912_, _38891_);
  nand (_38914_, _38913_, _38702_);
  and (_38915_, _38914_, _42003_);
  and (_13655_, _38915_, _38890_);
  nor (_38916_, _38699_, _32133_);
  and (_38917_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38918_, _38917_, _38702_);
  or (_38919_, _38918_, _38916_);
  nor (_38920_, _27457_, _16328_);
  nor (_38921_, _28569_, _19428_);
  nor (_38922_, _38723_, _26203_);
  nor (_38923_, _38922_, _38715_);
  nor (_38924_, _38923_, _26628_);
  and (_38925_, _38923_, _26628_);
  nor (_38926_, _38925_, _38924_);
  and (_38927_, _38926_, _27532_);
  nor (_38928_, _26203_, _18185_);
  or (_38929_, _38928_, _27816_);
  nor (_38930_, _38929_, _38716_);
  or (_38931_, _38930_, _38927_);
  or (_38932_, _38931_, _38921_);
  and (_38933_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38934_, _38771_, _38767_);
  nor (_38935_, _38934_, _38772_);
  and (_38936_, _38935_, _25465_);
  and (_38937_, _20720_, _15770_);
  or (_38938_, _38937_, _38936_);
  or (_38939_, _38938_, _38933_);
  or (_38940_, _38939_, _38932_);
  nor (_38941_, _38940_, _38920_);
  nand (_38942_, _38941_, _38702_);
  and (_38943_, _38942_, _42003_);
  and (_13664_, _38943_, _38919_);
  nor (_38944_, _38699_, _32943_);
  and (_38945_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38946_, _38945_, _38702_);
  or (_38947_, _38946_, _38944_);
  nor (_38948_, _27457_, _17314_);
  nor (_38949_, _28569_, _18882_);
  and (_38950_, _38723_, _16328_);
  nor (_38951_, _38950_, _26203_);
  not (_38952_, _38951_);
  and (_38953_, _38952_, _38717_);
  and (_38954_, _38953_, _17314_);
  nor (_38955_, _38953_, _17314_);
  or (_38956_, _38955_, _38954_);
  and (_38957_, _38956_, _27532_);
  nor (_38958_, _33282_, _27816_);
  and (_38959_, _38958_, _38709_);
  or (_38960_, _38959_, _38957_);
  or (_38961_, _38960_, _38949_);
  and (_38962_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38963_, _38772_, _38746_);
  nor (_38964_, _38963_, _38773_);
  and (_38965_, _38964_, _25465_);
  and (_38966_, _20752_, _15770_);
  or (_38967_, _38966_, _38965_);
  or (_38968_, _38967_, _38962_);
  or (_38969_, _38968_, _38961_);
  nor (_38970_, _38969_, _38948_);
  nand (_38971_, _38970_, _38702_);
  and (_38972_, _38971_, _42003_);
  and (_13673_, _38972_, _38947_);
  nor (_38973_, _38699_, _33677_);
  and (_38974_, _38699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38975_, _38974_, _38702_);
  or (_38976_, _38975_, _38973_);
  nor (_38977_, _27457_, _16669_);
  nor (_38978_, _28569_, _19046_);
  nor (_38979_, _38728_, _16669_);
  and (_38980_, _38728_, _16669_);
  nor (_38981_, _38980_, _38979_);
  nor (_38982_, _38981_, _31090_);
  nor (_38983_, _26203_, _16998_);
  or (_38984_, _38983_, _27816_);
  nor (_38985_, _38984_, _38730_);
  or (_38986_, _38985_, _38982_);
  or (_38987_, _38986_, _38978_);
  and (_38988_, _21123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38989_, _38777_, _38773_);
  nor (_38990_, _38989_, _38778_);
  and (_38991_, _38990_, _25465_);
  and (_38992_, _20783_, _15770_);
  or (_38993_, _38992_, _38991_);
  or (_38994_, _38993_, _38988_);
  or (_38995_, _38994_, _38987_);
  nor (_38996_, _38995_, _38977_);
  nand (_38997_, _38996_, _38702_);
  and (_38998_, _38997_, _42003_);
  and (_13683_, _38998_, _38976_);
  nand (_38999_, _38797_, _29288_);
  or (_39000_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_39001_, _39000_, _42003_);
  and (_13692_, _39001_, _38999_);
  nand (_39002_, _38797_, _29961_);
  or (_39003_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_39004_, _39003_, _42003_);
  and (_13702_, _39004_, _39002_);
  nand (_39005_, _38797_, _30656_);
  not (_39006_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_39007_, _38796_, _39006_);
  and (_39008_, _39007_, _42003_);
  and (_13712_, _39008_, _39005_);
  nand (_39009_, _38797_, _31416_);
  or (_39010_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_39011_, _39010_, _42003_);
  and (_13721_, _39011_, _39009_);
  nand (_39012_, _38797_, _32133_);
  or (_39014_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_39017_, _39014_, _42003_);
  and (_13731_, _39017_, _39012_);
  nand (_39018_, _38797_, _32943_);
  or (_39019_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_39020_, _39019_, _42003_);
  and (_13740_, _39020_, _39018_);
  nand (_39021_, _38797_, _33677_);
  or (_39022_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_39023_, _39022_, _42003_);
  and (_13750_, _39023_, _39021_);
  not (_39024_, _24754_);
  and (_39033_, _25376_, _24886_);
  and (_39039_, _39033_, _39024_);
  and (_39045_, _28831_, _25072_);
  and (_39049_, _39045_, _39039_);
  not (_39050_, _28798_);
  nor (_39051_, _39050_, _28766_);
  not (_39052_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_39053_, _28798_, _39052_);
  or (_39054_, _39053_, _39051_);
  and (_39055_, _39054_, _39049_);
  and (_39056_, _28199_, _24557_);
  nor (_39057_, _24754_, _25061_);
  and (_39058_, _39033_, _39057_);
  and (_39059_, _39058_, _39056_);
  nor (_39060_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_39061_, _39060_);
  nand (_39062_, _39061_, _28766_);
  and (_39063_, _39060_, _39052_);
  nor (_39064_, _39049_, _39063_);
  and (_39065_, _39064_, _39062_);
  or (_39066_, _39065_, _39059_);
  or (_39067_, _39066_, _39055_);
  nand (_39068_, _39059_, _38651_);
  and (_39069_, _39068_, _39067_);
  and (_16547_, _39069_, _42003_);
  not (_39070_, _39059_);
  nor (_39071_, _39070_, _38620_);
  not (_39072_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_39074_, _39058_, _28831_);
  nand (_39076_, _39074_, _30080_);
  nand (_39077_, _39076_, _39072_);
  and (_39078_, _39077_, _39070_);
  or (_39079_, _39076_, _29375_);
  and (_39080_, _39079_, _39078_);
  or (_39081_, _39080_, _39071_);
  and (_21481_, _39081_, _42003_);
  nor (_39082_, _39070_, _38613_);
  not (_39083_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39084_, _30798_, _39083_);
  or (_39085_, _39084_, _30808_);
  and (_39086_, _39085_, _39074_);
  or (_39087_, _20878_, _20847_);
  or (_39088_, _39087_, _20910_);
  or (_39089_, _39088_, _20953_);
  or (_39090_, _39089_, _21027_);
  or (_39091_, _39090_, _21059_);
  and (_39092_, _39091_, _15770_);
  and (_39093_, _28308_, _27130_);
  not (_39094_, _27130_);
  and (_39095_, _28319_, _39094_);
  or (_39096_, _39095_, _39093_);
  and (_39097_, _39096_, _26563_);
  not (_39098_, _26443_);
  nand (_39099_, _26433_, _39098_);
  or (_39100_, _26454_, _26433_);
  and (_39101_, _25465_, _39100_);
  and (_39102_, _39101_, _39099_);
  and (_39103_, _38724_, _22326_);
  and (_39104_, _38722_, _21123_);
  nand (_39105_, _39104_, _39103_);
  nand (_39106_, _39105_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39107_, _39106_, _39102_);
  or (_39108_, _39107_, _39097_);
  or (_39109_, _39108_, _31665_);
  or (_39110_, _39109_, _25432_);
  or (_39111_, _39110_, _39092_);
  nor (_39113_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39116_, _39113_, _39074_);
  and (_39122_, _39116_, _39111_);
  or (_39127_, _39122_, _39086_);
  and (_39134_, _39127_, _39070_);
  or (_39141_, _39134_, _39082_);
  and (_21493_, _39141_, _42003_);
  nor (_39151_, _39070_, _38592_);
  and (_39152_, _39074_, _31514_);
  nand (_39153_, _39152_, _28766_);
  or (_39154_, _39152_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_39155_, _39154_, _39070_);
  and (_39156_, _39155_, _39153_);
  or (_39157_, _39156_, _39151_);
  and (_21505_, _39157_, _42003_);
  nor (_39158_, _39070_, _38506_);
  not (_39159_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_39160_, _39059_, _39159_);
  or (_39161_, _39160_, _39158_);
  not (_39162_, _39074_);
  or (_39163_, _39162_, _32253_);
  and (_39164_, _39163_, _39161_);
  and (_39165_, _32242_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39166_, _39165_, _32286_);
  and (_39167_, _39166_, _39074_);
  or (_39168_, _39167_, _39164_);
  and (_21517_, _39168_, _42003_);
  nor (_39169_, _39070_, _38452_);
  not (_39170_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_39171_, _39074_, _33031_);
  nand (_39172_, _39171_, _39170_);
  and (_39173_, _39172_, _39070_);
  or (_39174_, _39171_, _29375_);
  and (_39175_, _39174_, _39173_);
  or (_39176_, _39175_, _39169_);
  and (_21529_, _39176_, _42003_);
  and (_39177_, _33776_, _29375_);
  nor (_39178_, _33776_, _31144_);
  or (_39179_, _39178_, _39177_);
  and (_39180_, _39179_, _39074_);
  and (_39181_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_39182_, _39181_, _27457_);
  and (_39183_, _39182_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_39184_, _25465_, _26335_);
  and (_39188_, _27086_, _26563_);
  or (_39199_, _39188_, _39184_);
  and (_39202_, _39199_, _39181_);
  or (_39203_, _39202_, _39183_);
  and (_39204_, _39203_, _39162_);
  or (_39213_, _39204_, _39180_);
  and (_39221_, _39213_, _39070_);
  nor (_39222_, _39070_, _38364_);
  or (_39223_, _39222_, _39221_);
  and (_21540_, _39223_, _42003_);
  not (_39224_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39225_, _38701_, _39224_);
  and (_39226_, _39225_, _38791_);
  nor (_39227_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39228_, _39227_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39229_, _24557_, _25213_);
  not (_39230_, _24886_);
  and (_39231_, _25344_, _39230_);
  and (_39232_, _39231_, _28199_);
  and (_39233_, _39232_, _39229_);
  and (_39234_, _39233_, _39057_);
  nor (_39235_, _39234_, _39228_);
  nor (_39236_, _39235_, _28122_);
  and (_39237_, _25344_, _25213_);
  and (_39238_, _39237_, _24897_);
  and (_39239_, _39238_, _39045_);
  and (_39240_, _39239_, _28798_);
  and (_39241_, _39240_, _28766_);
  nor (_39242_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_39243_, _39228_, _39225_);
  nor (_39244_, _39243_, _39234_);
  not (_39245_, _39244_);
  nor (_39246_, _39245_, _39242_);
  not (_39247_, _39246_);
  nor (_39248_, _39247_, _39241_);
  nor (_39249_, _39248_, _39225_);
  not (_39250_, _39249_);
  nor (_39251_, _39250_, _39236_);
  nor (_39252_, _39251_, _39226_);
  and (_22315_, _39252_, _42003_);
  not (_39253_, _39225_);
  nor (_39254_, _39235_, _29288_);
  and (_39255_, _39239_, _24557_);
  and (_39256_, _39255_, _28766_);
  nor (_39257_, _39255_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_39258_, _39257_, _39245_);
  not (_39259_, _39258_);
  nor (_39260_, _39259_, _39256_);
  or (_39261_, _39260_, _39254_);
  and (_39262_, _39261_, _39253_);
  nor (_39263_, _39253_, _38828_);
  or (_39264_, _39263_, _39262_);
  and (_24176_, _39264_, _42003_);
  and (_39265_, _39225_, _38856_);
  nor (_39266_, _39235_, _29961_);
  and (_39267_, _39239_, _30080_);
  and (_39268_, _39267_, _28766_);
  nor (_39269_, _39267_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_39270_, _39269_, _39245_);
  not (_39271_, _39270_);
  nor (_39272_, _39271_, _39268_);
  nor (_39273_, _39272_, _39225_);
  not (_39274_, _39273_);
  nor (_39275_, _39274_, _39266_);
  nor (_39276_, _39275_, _39265_);
  and (_24188_, _39276_, _42003_);
  nor (_39277_, _39235_, _30656_);
  and (_39278_, _39239_, _30798_);
  and (_39279_, _39278_, _28766_);
  nor (_39280_, _39278_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_39281_, _39280_, _39245_);
  not (_39282_, _39281_);
  nor (_39283_, _39282_, _39279_);
  or (_39284_, _39283_, _39277_);
  and (_39285_, _39284_, _39253_);
  nor (_39286_, _39253_, _38884_);
  or (_39287_, _39286_, _39285_);
  and (_24200_, _39287_, _42003_);
  nor (_39288_, _39235_, _31416_);
  not (_39289_, _39239_);
  and (_39290_, _39244_, _39289_);
  and (_39291_, _39290_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_39292_, _31525_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39293_, _39292_, _31536_);
  and (_39294_, _39239_, _39253_);
  not (_39295_, _39294_);
  nor (_39296_, _39295_, _39293_);
  and (_39297_, _39296_, _39244_);
  nor (_39298_, _39297_, _39291_);
  and (_39299_, _39298_, _39253_);
  not (_39300_, _39299_);
  nor (_39301_, _39300_, _39288_);
  and (_39302_, _39225_, _38913_);
  or (_39303_, _39302_, _39301_);
  nor (_24212_, _39303_, rst);
  nor (_39304_, _39235_, _32133_);
  and (_39305_, _39239_, _32231_);
  and (_39306_, _39305_, _28766_);
  nor (_39307_, _39305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_39308_, _39307_, _39245_);
  not (_39309_, _39308_);
  nor (_39310_, _39309_, _39306_);
  or (_39311_, _39310_, _39304_);
  and (_39312_, _39311_, _39253_);
  nor (_39313_, _39253_, _38941_);
  or (_39314_, _39313_, _39312_);
  and (_24224_, _39314_, _42003_);
  nor (_39315_, _39235_, _32943_);
  and (_39316_, _39239_, _33031_);
  and (_39317_, _39316_, _28766_);
  nor (_39318_, _39316_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_39319_, _39318_, _39245_);
  not (_39320_, _39319_);
  nor (_39321_, _39320_, _39317_);
  or (_39322_, _39321_, _39315_);
  and (_39323_, _39322_, _39253_);
  nor (_39324_, _39253_, _38970_);
  or (_39325_, _39324_, _39323_);
  and (_24236_, _39325_, _42003_);
  nor (_39326_, _39235_, _33677_);
  and (_39327_, _39239_, _33776_);
  and (_39328_, _39327_, _28766_);
  nor (_39329_, _39327_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_39330_, _39329_, _39245_);
  not (_39331_, _39330_);
  nor (_39332_, _39331_, _39328_);
  or (_39333_, _39332_, _39326_);
  and (_39334_, _39333_, _39253_);
  nor (_39335_, _39253_, _38996_);
  or (_39336_, _39335_, _39334_);
  and (_24248_, _39336_, _42003_);
  and (_39337_, _38210_, _28798_);
  nand (_39338_, _39337_, _28766_);
  or (_39339_, _39337_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39340_, _39339_, _28831_);
  and (_39341_, _39340_, _39338_);
  and (_39342_, _38155_, _39229_);
  nand (_39343_, _39342_, _38651_);
  or (_39344_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39345_, _39344_, _28199_);
  and (_39346_, _39345_, _39343_);
  not (_39347_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39348_, _28188_, _39347_);
  or (_39349_, _39348_, rst);
  or (_39350_, _39349_, _39346_);
  or (_35486_, _39350_, _39341_);
  nor (_39351_, _39024_, _25061_);
  and (_39352_, _39033_, _39351_);
  and (_39353_, _39352_, _28798_);
  nand (_39354_, _39353_, _28766_);
  or (_39355_, _39353_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39356_, _39355_, _28831_);
  and (_39357_, _39356_, _39354_);
  and (_39358_, _39352_, _24557_);
  not (_39359_, _39358_);
  nor (_39360_, _39359_, _38651_);
  not (_39361_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39362_, _39358_, _39361_);
  or (_39363_, _39362_, _39360_);
  and (_39364_, _39363_, _28199_);
  nor (_39365_, _28188_, _39361_);
  or (_39366_, _39365_, rst);
  or (_39367_, _39366_, _39364_);
  or (_35509_, _39367_, _39357_);
  and (_39368_, _39230_, _24754_);
  and (_39369_, _39368_, _39237_);
  and (_39370_, _39369_, _25072_);
  and (_39371_, _39370_, _28798_);
  nand (_39372_, _39371_, _28766_);
  or (_39373_, _39371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39374_, _39373_, _28831_);
  and (_39375_, _39374_, _39372_);
  and (_39376_, _39231_, _39351_);
  and (_39377_, _39376_, _39229_);
  not (_39378_, _39377_);
  nor (_39379_, _39378_, _38651_);
  not (_39380_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39381_, _39377_, _39380_);
  or (_39382_, _39381_, _39379_);
  and (_39383_, _39382_, _28199_);
  nor (_39384_, _28188_, _39380_);
  or (_39385_, _39384_, rst);
  or (_39386_, _39385_, _39383_);
  or (_35532_, _39386_, _39375_);
  and (_39387_, _39368_, _25377_);
  and (_39388_, _39387_, _28798_);
  nand (_39389_, _39388_, _28766_);
  or (_39390_, _39388_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39391_, _39390_, _28831_);
  and (_39392_, _39391_, _39389_);
  nor (_39393_, _25344_, _24886_);
  and (_39394_, _39351_, _39393_);
  and (_39395_, _39394_, _39229_);
  not (_39396_, _39395_);
  nor (_39403_, _39396_, _38651_);
  not (_39414_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_39425_, _39395_, _39414_);
  or (_39435_, _39425_, _39403_);
  and (_39441_, _39435_, _28199_);
  nor (_39451_, _28188_, _39414_);
  or (_39462_, _39451_, rst);
  or (_39473_, _39462_, _39441_);
  or (_35555_, _39473_, _39392_);
  not (_39494_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39505_, _39342_, _39494_);
  nand (_39516_, _38210_, _24557_);
  nor (_39527_, _39516_, _28766_);
  or (_39538_, _39527_, _39505_);
  and (_39549_, _39538_, _28831_);
  and (_39560_, _39342_, _38629_);
  or (_39571_, _39560_, _39505_);
  and (_39582_, _39571_, _28199_);
  nor (_39593_, _28188_, _39494_);
  or (_39604_, _39593_, rst);
  or (_39610_, _39604_, _39582_);
  or (_41403_, _39610_, _39549_);
  or (_39611_, _38232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39612_, _39611_, _28831_);
  nand (_39613_, _38232_, _28766_);
  and (_39614_, _39613_, _39612_);
  nand (_39615_, _39342_, _38620_);
  or (_39616_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39617_, _39616_, _28199_);
  and (_39618_, _39617_, _39615_);
  not (_39619_, _28188_);
  and (_39620_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39621_, _39620_, rst);
  or (_39622_, _39621_, _39618_);
  or (_41404_, _39622_, _39614_);
  not (_39623_, _31547_);
  nand (_39624_, _38210_, _39623_);
  and (_39625_, _39624_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39626_, _30819_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39627_, _39626_, _30808_);
  and (_39628_, _39627_, _38210_);
  or (_39629_, _39628_, _39625_);
  and (_39630_, _39629_, _28831_);
  nand (_39631_, _39342_, _38613_);
  or (_39632_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39633_, _39632_, _28199_);
  and (_39634_, _39633_, _39631_);
  not (_39635_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_39636_, _28188_, _39635_);
  or (_39637_, _39636_, rst);
  or (_39638_, _39637_, _39634_);
  or (_41406_, _39638_, _39630_);
  not (_39639_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_39640_, _38221_, _39639_);
  nor (_39641_, _31547_, _39639_);
  or (_39642_, _39641_, _31536_);
  and (_39643_, _39642_, _38210_);
  or (_39644_, _39643_, _39640_);
  and (_39645_, _39644_, _28831_);
  nand (_39646_, _39342_, _38592_);
  or (_39647_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39648_, _39647_, _28199_);
  and (_39649_, _39648_, _39646_);
  nor (_39650_, _28188_, _39639_);
  or (_39651_, _39650_, rst);
  or (_39652_, _39651_, _39649_);
  or (_41408_, _39652_, _39645_);
  not (_39653_, _38210_);
  or (_39654_, _39653_, _32253_);
  and (_39655_, _39654_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39656_, _32242_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39657_, _39656_, _32286_);
  and (_39658_, _39657_, _38210_);
  or (_39659_, _39658_, _39655_);
  and (_39660_, _39659_, _28831_);
  nand (_39661_, _39342_, _38506_);
  or (_39662_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39663_, _39662_, _28199_);
  and (_39664_, _39663_, _39661_);
  and (_39665_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39666_, _39665_, rst);
  or (_39667_, _39666_, _39664_);
  or (_41409_, _39667_, _39660_);
  and (_39668_, _38210_, _33031_);
  nand (_39669_, _39668_, _28766_);
  or (_39670_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39671_, _39670_, _28831_);
  and (_39672_, _39671_, _39669_);
  nand (_39673_, _39342_, _38452_);
  or (_39674_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39675_, _39674_, _28199_);
  and (_39676_, _39675_, _39673_);
  and (_39677_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39678_, _39677_, rst);
  or (_39679_, _39678_, _39676_);
  or (_41411_, _39679_, _39672_);
  and (_39680_, _38210_, _33776_);
  nand (_39681_, _39680_, _28766_);
  or (_39682_, _39680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39683_, _39682_, _28831_);
  and (_39684_, _39683_, _39681_);
  nand (_39685_, _39342_, _38364_);
  or (_39686_, _39342_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39687_, _39686_, _28199_);
  and (_39688_, _39687_, _39685_);
  and (_39689_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39690_, _39689_, rst);
  or (_39691_, _39690_, _39688_);
  or (_41413_, _39691_, _39684_);
  nand (_39692_, _39358_, _28766_);
  or (_39693_, _39358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39694_, _39693_, _28831_);
  and (_39695_, _39694_, _39692_);
  and (_39696_, _39358_, _38629_);
  and (_39697_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39698_, _39697_, _39696_);
  and (_39699_, _39698_, _28199_);
  and (_39700_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39701_, _39700_, rst);
  or (_39702_, _39701_, _39699_);
  or (_41415_, _39702_, _39695_);
  and (_39703_, _39352_, _30080_);
  nand (_39704_, _39703_, _28766_);
  or (_39705_, _39703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39706_, _39705_, _28831_);
  and (_39707_, _39706_, _39704_);
  nor (_39708_, _39359_, _38620_);
  and (_39709_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39710_, _39709_, _39708_);
  and (_39711_, _39710_, _28199_);
  and (_39712_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39713_, _39712_, rst);
  or (_39714_, _39713_, _39711_);
  or (_41416_, _39714_, _39707_);
  and (_39715_, _39352_, _30798_);
  nand (_39716_, _39715_, _28766_);
  or (_39717_, _39715_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39718_, _39717_, _28831_);
  and (_39719_, _39718_, _39716_);
  nor (_39720_, _39359_, _38613_);
  not (_39721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_39722_, _39358_, _39721_);
  or (_39723_, _39722_, _39720_);
  and (_39724_, _39723_, _28199_);
  nor (_39725_, _28188_, _39721_);
  or (_39726_, _39725_, rst);
  or (_39727_, _39726_, _39724_);
  or (_41418_, _39727_, _39719_);
  and (_39728_, _39352_, _31514_);
  nand (_39729_, _39728_, _28766_);
  or (_39730_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39731_, _39730_, _28831_);
  and (_39732_, _39731_, _39729_);
  nor (_39733_, _39359_, _38592_);
  and (_39734_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39735_, _39734_, _39733_);
  and (_39736_, _39735_, _28199_);
  and (_39737_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39738_, _39737_, rst);
  or (_39739_, _39738_, _39736_);
  or (_41420_, _39739_, _39732_);
  and (_39740_, _39352_, _32231_);
  nand (_39741_, _39740_, _28766_);
  or (_39742_, _39740_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39743_, _39742_, _28831_);
  and (_39744_, _39743_, _39741_);
  nor (_39745_, _39359_, _38506_);
  and (_39746_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39747_, _39746_, _39745_);
  and (_39748_, _39747_, _28199_);
  and (_39749_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39750_, _39749_, rst);
  or (_39751_, _39750_, _39748_);
  or (_41421_, _39751_, _39744_);
  and (_39752_, _39352_, _33031_);
  nand (_39753_, _39752_, _28766_);
  or (_39754_, _39752_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39755_, _39754_, _28831_);
  and (_39756_, _39755_, _39753_);
  nor (_39757_, _39359_, _38452_);
  and (_39758_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39759_, _39758_, _39757_);
  and (_39760_, _39759_, _28199_);
  and (_39761_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39762_, _39761_, rst);
  or (_39763_, _39762_, _39760_);
  or (_41423_, _39763_, _39756_);
  and (_39764_, _39352_, _33776_);
  nand (_39765_, _39764_, _28766_);
  or (_39766_, _39764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39767_, _39766_, _28831_);
  and (_39768_, _39767_, _39765_);
  nor (_39769_, _39359_, _38364_);
  and (_39770_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39771_, _39770_, _39769_);
  and (_39772_, _39771_, _28199_);
  and (_39773_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39774_, _39773_, rst);
  or (_39775_, _39774_, _39772_);
  or (_41425_, _39775_, _39768_);
  nand (_39776_, _39377_, _28766_);
  or (_39777_, _39377_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39778_, _39777_, _28831_);
  and (_39779_, _39778_, _39776_);
  and (_39780_, _39377_, _38629_);
  and (_39781_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39782_, _39781_, _39780_);
  and (_39783_, _39782_, _28199_);
  and (_39784_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39785_, _39784_, rst);
  or (_39786_, _39785_, _39783_);
  or (_41427_, _39786_, _39779_);
  and (_39787_, _39370_, _30080_);
  nand (_39788_, _39787_, _28766_);
  or (_39789_, _39787_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39790_, _39789_, _28831_);
  and (_39791_, _39790_, _39788_);
  nor (_39792_, _39378_, _38620_);
  and (_39793_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39794_, _39793_, _39792_);
  and (_39795_, _39794_, _28199_);
  and (_39796_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39797_, _39796_, rst);
  or (_39798_, _39797_, _39795_);
  or (_41429_, _39798_, _39791_);
  and (_39799_, _39370_, _30798_);
  nand (_39800_, _39799_, _28766_);
  or (_39801_, _39799_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39802_, _39801_, _28831_);
  and (_39803_, _39802_, _39800_);
  nor (_39804_, _39378_, _38613_);
  not (_39805_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_39806_, _39377_, _39805_);
  or (_39807_, _39806_, _39804_);
  and (_39808_, _39807_, _28199_);
  nor (_39809_, _28188_, _39805_);
  or (_39810_, _39809_, rst);
  or (_39811_, _39810_, _39808_);
  or (_41430_, _39811_, _39803_);
  and (_39812_, _39370_, _31514_);
  nand (_39813_, _39812_, _28766_);
  or (_39814_, _39812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39815_, _39814_, _28831_);
  and (_39817_, _39815_, _39813_);
  nor (_39818_, _39378_, _38592_);
  and (_39819_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39820_, _39819_, _39818_);
  and (_39821_, _39820_, _28199_);
  and (_39822_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39823_, _39822_, rst);
  or (_39824_, _39823_, _39821_);
  or (_41432_, _39824_, _39817_);
  and (_39825_, _39370_, _32231_);
  nand (_39826_, _39825_, _28766_);
  or (_39827_, _39825_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39828_, _39827_, _28831_);
  and (_39829_, _39828_, _39826_);
  nor (_39830_, _39378_, _38506_);
  and (_39831_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39832_, _39831_, _39830_);
  and (_39833_, _39832_, _28199_);
  and (_39834_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39835_, _39834_, rst);
  or (_39836_, _39835_, _39833_);
  or (_41434_, _39836_, _39829_);
  and (_39837_, _39370_, _33031_);
  nand (_39838_, _39837_, _28766_);
  or (_39839_, _39837_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39840_, _39839_, _28831_);
  and (_39841_, _39840_, _39838_);
  nor (_39842_, _39378_, _38452_);
  and (_39843_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39844_, _39843_, _39842_);
  and (_39845_, _39844_, _28199_);
  and (_39846_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39851_, _39846_, rst);
  or (_39852_, _39851_, _39845_);
  or (_41435_, _39852_, _39841_);
  and (_39853_, _39370_, _33776_);
  nand (_39854_, _39853_, _28766_);
  or (_39855_, _39853_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39856_, _39855_, _28831_);
  and (_39857_, _39856_, _39854_);
  nor (_39858_, _39378_, _38364_);
  and (_39859_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39860_, _39859_, _39858_);
  and (_39861_, _39860_, _28199_);
  and (_39862_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39863_, _39862_, rst);
  or (_39864_, _39863_, _39861_);
  or (_41437_, _39864_, _39857_);
  and (_39865_, _39387_, _24557_);
  nand (_39866_, _39865_, _28766_);
  or (_39867_, _39865_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39868_, _39867_, _28831_);
  and (_39869_, _39868_, _39866_);
  and (_39870_, _39395_, _38629_);
  and (_39871_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39872_, _39871_, _39870_);
  and (_39873_, _39872_, _28199_);
  and (_39874_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39875_, _39874_, rst);
  or (_39876_, _39875_, _39873_);
  or (_41439_, _39876_, _39869_);
  and (_39877_, _39387_, _30080_);
  nand (_39878_, _39877_, _28766_);
  or (_39879_, _39877_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39880_, _39879_, _28831_);
  and (_39881_, _39880_, _39878_);
  nor (_39882_, _39396_, _38620_);
  and (_39883_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39884_, _39883_, _39882_);
  and (_39885_, _39884_, _28199_);
  and (_39886_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39887_, _39886_, rst);
  or (_39888_, _39887_, _39885_);
  or (_41440_, _39888_, _39881_);
  and (_39889_, _39387_, _30798_);
  nand (_39890_, _39889_, _28766_);
  or (_39891_, _39889_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39892_, _39891_, _28831_);
  and (_39893_, _39892_, _39890_);
  nor (_39894_, _39396_, _38613_);
  not (_39895_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_39896_, _39395_, _39895_);
  or (_39897_, _39896_, _39894_);
  and (_39898_, _39897_, _28199_);
  nor (_39899_, _28188_, _39895_);
  or (_39900_, _39899_, rst);
  or (_39901_, _39900_, _39898_);
  or (_41442_, _39901_, _39893_);
  and (_39902_, _39387_, _31514_);
  nand (_39903_, _39902_, _28766_);
  or (_39904_, _39902_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39905_, _39904_, _28831_);
  and (_39906_, _39905_, _39903_);
  nor (_39907_, _39396_, _38592_);
  and (_39908_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39909_, _39908_, _39907_);
  and (_39910_, _39909_, _28199_);
  and (_39911_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39919_, _39911_, rst);
  or (_39920_, _39919_, _39910_);
  or (_41444_, _39920_, _39906_);
  and (_39921_, _39387_, _32231_);
  nand (_39922_, _39921_, _28766_);
  or (_39923_, _39921_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39924_, _39923_, _28831_);
  and (_39925_, _39924_, _39922_);
  nor (_39926_, _39396_, _38506_);
  and (_39927_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39928_, _39927_, _39926_);
  and (_39929_, _39928_, _28199_);
  and (_39930_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39931_, _39930_, rst);
  or (_39932_, _39931_, _39929_);
  or (_41445_, _39932_, _39925_);
  and (_39933_, _39387_, _33031_);
  nand (_39934_, _39933_, _28766_);
  or (_39935_, _39933_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39936_, _39935_, _28831_);
  and (_39937_, _39936_, _39934_);
  nor (_39938_, _39396_, _38452_);
  and (_39939_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39940_, _39939_, _39938_);
  and (_39941_, _39940_, _28199_);
  and (_39942_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39943_, _39942_, rst);
  or (_39944_, _39943_, _39941_);
  or (_41447_, _39944_, _39937_);
  and (_39945_, _39387_, _33776_);
  nand (_39946_, _39945_, _28766_);
  or (_39947_, _39945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39948_, _39947_, _28831_);
  and (_39949_, _39948_, _39946_);
  nor (_39950_, _39396_, _38364_);
  and (_39951_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39952_, _39951_, _39950_);
  and (_39953_, _39952_, _28199_);
  and (_39954_, _39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39955_, _39954_, rst);
  or (_39956_, _39955_, _39953_);
  or (_41449_, _39956_, _39949_);
  nor (_39957_, _25344_, _25213_);
  and (_39958_, _39957_, _39368_);
  and (_39959_, _39958_, _39045_);
  and (_39960_, _39959_, _28798_);
  nand (_39961_, _39960_, _28766_);
  not (_39966_, _25213_);
  and (_39967_, _39056_, _39966_);
  and (_39968_, _39967_, _39394_);
  not (_39969_, _39968_);
  or (_39970_, _39960_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39971_, _39970_, _39969_);
  and (_39972_, _39971_, _39961_);
  nor (_39973_, _39969_, _38651_);
  or (_39974_, _39973_, _39972_);
  and (_41945_, _39974_, _42003_);
  and (_39975_, _25344_, _39966_);
  and (_39976_, _39975_, _39045_);
  and (_39977_, _39976_, _39368_);
  and (_39978_, _39977_, _28798_);
  nand (_39979_, _39978_, _28766_);
  and (_39980_, _39967_, _39376_);
  not (_39990_, _39980_);
  or (_39991_, _39978_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39992_, _39991_, _39990_);
  and (_39993_, _39992_, _39979_);
  nor (_39994_, _39990_, _38651_);
  or (_39995_, _39994_, _39993_);
  and (_41948_, _39995_, _42003_);
  or (_39996_, _24546_, _30787_);
  and (_39997_, _39996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39998_, _39997_, _39177_);
  and (_39999_, _39976_, _38133_);
  and (_40000_, _39999_, _39998_);
  and (_40001_, _39967_, _38155_);
  nand (_40002_, _39999_, _24535_);
  and (_40003_, _40002_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40004_, _40003_, _40001_);
  or (_40005_, _40004_, _40000_);
  nand (_40006_, _40001_, _38364_);
  and (_40007_, _40006_, _42003_);
  and (_41950_, _40007_, _40005_);
  not (_40008_, _40001_);
  not (_40009_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40011_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40011_);
  and (_40013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40014_, _40013_, _40012_);
  nor (_40015_, _40014_, _40010_);
  or (_40016_, _40015_, _40009_);
  and (_40017_, _40011_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40018_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40019_, _40018_, _40017_);
  nor (_40020_, _40019_, _40010_);
  and (_40021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40011_);
  and (_40022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40023_, _40022_, _40021_);
  nand (_40024_, _40023_, _40020_);
  or (_40025_, _40024_, _40016_);
  and (_40026_, _40025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_40027_, _24293_, _25213_);
  and (_40028_, _28831_, _28788_);
  and (_40029_, _40028_, _38155_);
  and (_40030_, _40029_, _40027_);
  or (_40031_, _40030_, _40026_);
  and (_40032_, _40031_, _40008_);
  nand (_40033_, _40030_, _28766_);
  and (_40034_, _40033_, _40032_);
  nor (_40035_, _40008_, _38651_);
  or (_40036_, _40035_, _40034_);
  and (_41952_, _40036_, _42003_);
  nor (_40037_, _40023_, _40010_);
  nand (_40038_, _40037_, _40019_);
  or (_40039_, _40038_, _40016_);
  and (_40040_, _40039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_40041_, _28831_, _30059_);
  and (_40042_, _40041_, _38155_);
  and (_40043_, _40042_, _40027_);
  or (_40044_, _40043_, _40040_);
  and (_40045_, _40044_, _40008_);
  nand (_40046_, _40043_, _28766_);
  and (_40047_, _40046_, _40045_);
  nor (_40048_, _40008_, _38452_);
  or (_40049_, _40048_, _40047_);
  and (_41954_, _40049_, _42003_);
  not (_40050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40050_);
  nand (_40052_, _40015_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40053_, _40037_, _40020_);
  or (_40054_, _40053_, _40052_);
  and (_40055_, _40054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40056_, _40055_, _40051_);
  nor (_40057_, _28777_, _25213_);
  and (_40058_, _40042_, _40057_);
  or (_40059_, _40058_, _40056_);
  and (_40060_, _40059_, _40008_);
  nand (_40061_, _40058_, _28766_);
  and (_40062_, _40061_, _40060_);
  nor (_40063_, _40008_, _38620_);
  or (_40064_, _40063_, _40062_);
  and (_41956_, _40064_, _42003_);
  and (_40065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40066_, _40052_, _40038_);
  and (_40067_, _40066_, _40065_);
  and (_40068_, _40029_, _40057_);
  or (_40069_, _40068_, _40067_);
  and (_40070_, _40069_, _40008_);
  nand (_40071_, _40068_, _28766_);
  and (_40072_, _40071_, _40070_);
  nor (_40073_, _40008_, _38592_);
  or (_40074_, _40073_, _40072_);
  and (_41958_, _40074_, _42003_);
  and (_40075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40076_, _40075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40077_, _40076_);
  and (_40078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40079_, _40078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40081_, _40080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_40082_, _40081_, _40079_);
  and (_40083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40084_, _40083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not (_40085_, _40084_);
  and (_40086_, _40085_, _40082_);
  and (_40087_, _40086_, _40077_);
  not (_40088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40011_);
  or (_40091_, _40090_, _40089_);
  nor (_40092_, _40091_, _40088_);
  nor (_40093_, _40092_, _40010_);
  nor (_40094_, _40093_, _40087_);
  and (_40095_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40096_, _40095_, _40011_);
  and (_40097_, _40096_, _40094_);
  and (_40098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40010_);
  not (_40099_, _40098_);
  not (_40100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40101_, _40078_, _40100_);
  not (_40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40103_, _40080_, _40102_);
  nor (_40104_, _40103_, _40101_);
  not (_40105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40106_, _40083_, _40105_);
  not (_40107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40108_, _40075_, _40107_);
  nor (_40109_, _40108_, _40106_);
  and (_40110_, _40109_, _40104_);
  nor (_40111_, _40110_, _40099_);
  nand (_40112_, _40111_, _40096_);
  and (_40113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42003_);
  nand (_40114_, _40113_, _40112_);
  nor (_41990_, _40114_, _40097_);
  nor (_40115_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40116_, _40115_);
  nor (_40117_, _40111_, _40094_);
  nor (_40118_, _40117_, _40116_);
  nand (_40119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42003_);
  nor (_41992_, _40119_, _40118_);
  nor (_40120_, _40117_, _40095_);
  not (_40121_, _40120_);
  and (_40122_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40123_, _40095_);
  and (_40124_, _40076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40125_, _40082_);
  or (_40126_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40127_, _40126_, _40124_);
  or (_40128_, _40086_, _40017_);
  and (_40129_, _40128_, _40127_);
  and (_40130_, _40129_, _40094_);
  not (_40131_, _40094_);
  and (_40132_, _40111_, _40131_);
  and (_40133_, _40108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40134_, _40133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40135_, _40104_);
  and (_40136_, _40106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40137_, _40136_, _40135_);
  and (_40138_, _40137_, _40134_);
  and (_40139_, _40135_, _40017_);
  or (_40140_, _40139_, _40138_);
  and (_40141_, _40140_, _40132_);
  or (_40142_, _40141_, _40130_);
  and (_40143_, _40142_, _40123_);
  or (_40144_, _40143_, _40122_);
  and (_41994_, _40144_, _42003_);
  and (_40145_, _40076_, _40011_);
  or (_40146_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_40147_, _40146_, _40145_);
  or (_40148_, _40086_, _40018_);
  and (_40149_, _40148_, _40147_);
  and (_40150_, _40149_, _40094_);
  or (_40151_, _40150_, _40095_);
  and (_40152_, _40117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40153_, _40108_, _40011_);
  or (_40154_, _40153_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40155_, _40106_, _40011_);
  nor (_40156_, _40155_, _40135_);
  and (_40157_, _40156_, _40154_);
  and (_40158_, _40135_, _40018_);
  or (_40159_, _40158_, _40157_);
  and (_40160_, _40159_, _40132_);
  or (_40161_, _40160_, _40152_);
  or (_40162_, _40161_, _40151_);
  or (_40163_, _40123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40164_, _40163_, _42003_);
  and (_41995_, _40164_, _40162_);
  nand (_40165_, _40117_, _40010_);
  nor (_40166_, _40011_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40167_, _40166_, _40095_);
  and (_40168_, _40167_, _42003_);
  and (_41997_, _40168_, _40165_);
  and (_40169_, _40117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40170_, _40011_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40171_, _40170_, _40166_);
  nor (_40172_, _40171_, _40131_);
  or (_40173_, _40172_, _40095_);
  or (_40174_, _40173_, _40169_);
  or (_40175_, _40171_, _40123_);
  and (_40176_, _40175_, _42003_);
  and (_41999_, _40176_, _40174_);
  and (_40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42003_);
  and (_42001_, _40177_, _40095_);
  and (_40178_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40179_, _40178_, _40120_);
  and (_42928_, _40179_, _42003_);
  and (_40180_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40181_, _40180_, _40120_);
  and (_42930_, _40181_, _42003_);
  and (_40182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42003_);
  and (_42932_, _40182_, _40095_);
  not (_40183_, _40101_);
  nor (_40184_, _40108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40185_, _40184_, _40106_);
  or (_40186_, _40185_, _40103_);
  and (_40187_, _40186_, _40183_);
  and (_40188_, _40187_, _40132_);
  not (_40189_, _40079_);
  or (_40190_, _40076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40191_, _40190_, _40085_);
  or (_40192_, _40191_, _40081_);
  and (_40193_, _40192_, _40189_);
  and (_40194_, _40193_, _40094_);
  or (_40195_, _40194_, _40095_);
  or (_40196_, _40195_, _40188_);
  or (_40197_, _40123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40198_, _40197_, _42003_);
  and (_42934_, _40198_, _40196_);
  nand (_40199_, _40104_, _40098_);
  nor (_40200_, _40199_, _40109_);
  or (_40201_, _40200_, _40094_);
  nand (_40202_, _40094_, _40125_);
  and (_40203_, _40202_, _40201_);
  or (_40204_, _40203_, _40095_);
  or (_40205_, _40123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40206_, _40205_, _42003_);
  and (_42936_, _40206_, _40204_);
  and (_40207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42003_);
  and (_42938_, _40207_, _40095_);
  and (_40208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42003_);
  and (_42940_, _40208_, _40095_);
  nand (_40209_, _40117_, _40115_);
  nor (_40210_, _40095_, _40094_);
  or (_40211_, _40210_, _40011_);
  and (_40212_, _40211_, _42003_);
  and (_42942_, _40212_, _40209_);
  and (_40213_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40214_, _40145_);
  and (_40215_, _40214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40216_, _40084_, _40011_);
  or (_40217_, _40216_, _40081_);
  or (_40218_, _40217_, _40215_);
  not (_40219_, _40081_);
  or (_40220_, _40219_, _40013_);
  and (_40221_, _40220_, _40218_);
  or (_40222_, _40221_, _40079_);
  or (_40223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40011_);
  or (_40224_, _40223_, _40189_);
  and (_40225_, _40224_, _40094_);
  and (_40226_, _40225_, _40222_);
  not (_40227_, _40153_);
  and (_40228_, _40227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_40229_, _40155_, _40103_);
  or (_40230_, _40229_, _40228_);
  not (_40231_, _40103_);
  or (_40232_, _40231_, _40013_);
  and (_40233_, _40232_, _40183_);
  and (_40234_, _40233_, _40230_);
  and (_40235_, _40223_, _40101_);
  or (_40236_, _40235_, _40234_);
  and (_40237_, _40236_, _40132_);
  or (_40238_, _40237_, _40226_);
  and (_40239_, _40238_, _40123_);
  or (_40240_, _40239_, _40213_);
  and (_42944_, _40240_, _42003_);
  and (_40241_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40242_, _40214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40243_, _40242_, _40217_);
  or (_40244_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40011_);
  or (_40245_, _40244_, _40219_);
  and (_40246_, _40245_, _40189_);
  and (_40247_, _40246_, _40243_);
  and (_40248_, _40079_, _40022_);
  or (_40249_, _40248_, _40247_);
  and (_40250_, _40249_, _40094_);
  and (_40251_, _40227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40252_, _40251_, _40229_);
  or (_40253_, _40244_, _40231_);
  and (_40254_, _40253_, _40183_);
  and (_40255_, _40254_, _40252_);
  and (_40256_, _40101_, _40022_);
  or (_40257_, _40256_, _40255_);
  and (_40258_, _40257_, _40132_);
  or (_40259_, _40258_, _40250_);
  and (_40260_, _40259_, _40123_);
  or (_40261_, _40260_, _40241_);
  and (_42946_, _40261_, _42003_);
  and (_40262_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_40263_, _40124_);
  and (_40264_, _40263_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40265_, _40084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40266_, _40265_, _40081_);
  or (_40267_, _40266_, _40264_);
  or (_40268_, _40219_, _40012_);
  and (_40269_, _40268_, _40267_);
  or (_40270_, _40269_, _40079_);
  or (_40271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40272_, _40271_, _40189_);
  and (_40273_, _40272_, _40094_);
  and (_40274_, _40273_, _40270_);
  not (_40275_, _40133_);
  and (_40276_, _40275_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40277_, _40136_, _40103_);
  or (_40278_, _40277_, _40276_);
  or (_40279_, _40231_, _40012_);
  and (_40280_, _40279_, _40183_);
  and (_40281_, _40280_, _40278_);
  and (_40282_, _40271_, _40101_);
  or (_40283_, _40282_, _40281_);
  and (_40284_, _40283_, _40132_);
  or (_40285_, _40284_, _40274_);
  and (_40286_, _40285_, _40123_);
  or (_40287_, _40286_, _40262_);
  and (_42948_, _40287_, _42003_);
  and (_40288_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40289_, _40263_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40290_, _40289_, _40266_);
  or (_40291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40292_, _40291_, _40219_);
  and (_40293_, _40292_, _40189_);
  and (_40294_, _40293_, _40290_);
  and (_40295_, _40079_, _40021_);
  or (_40296_, _40295_, _40294_);
  and (_40297_, _40296_, _40094_);
  and (_40298_, _40275_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40299_, _40298_, _40277_);
  or (_40300_, _40291_, _40231_);
  and (_40301_, _40300_, _40183_);
  and (_40302_, _40301_, _40299_);
  and (_40303_, _40101_, _40021_);
  or (_40304_, _40303_, _40302_);
  and (_40305_, _40304_, _40132_);
  or (_40306_, _40305_, _40297_);
  and (_40307_, _40306_, _40123_);
  or (_40308_, _40307_, _40288_);
  and (_42950_, _40308_, _42003_);
  and (_40309_, _40115_, _40094_);
  nand (_40310_, _40115_, _40111_);
  and (_40311_, _40310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40312_, _40311_, _40309_);
  and (_42952_, _40312_, _42003_);
  and (_40313_, _40112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40314_, _40313_, _40097_);
  and (_42954_, _40314_, _42003_);
  and (_40315_, _39999_, _24557_);
  or (_40316_, _40315_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40317_, _40316_, _40008_);
  nand (_40318_, _40315_, _28766_);
  and (_40319_, _40318_, _40317_);
  and (_40320_, _40001_, _38629_);
  or (_40321_, _40320_, _40319_);
  and (_42956_, _40321_, _42003_);
  and (_40322_, _39999_, _30798_);
  nand (_40323_, _40322_, _28766_);
  or (_40324_, _40322_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40325_, _40324_, _40008_);
  and (_40326_, _40325_, _40323_);
  nor (_40327_, _40008_, _38613_);
  or (_40328_, _40327_, _40326_);
  and (_42958_, _40328_, _42003_);
  and (_40329_, _39999_, _32231_);
  nand (_40330_, _40329_, _28766_);
  or (_40331_, _40329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40332_, _40331_, _40008_);
  and (_40333_, _40332_, _40330_);
  nor (_40334_, _40008_, _38506_);
  or (_40335_, _40334_, _40333_);
  and (_42960_, _40335_, _42003_);
  and (_40336_, _39977_, _24557_);
  nand (_40337_, _40336_, _28766_);
  or (_40338_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40339_, _40338_, _39990_);
  and (_40340_, _40339_, _40337_);
  and (_40341_, _39980_, _38629_);
  or (_40342_, _40341_, _40340_);
  and (_42962_, _40342_, _42003_);
  and (_40343_, _39977_, _30080_);
  nand (_40344_, _40343_, _28766_);
  or (_40345_, _40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40346_, _40345_, _39990_);
  and (_40347_, _40346_, _40344_);
  nor (_40348_, _39990_, _38620_);
  or (_40349_, _40348_, _40347_);
  and (_42964_, _40349_, _42003_);
  and (_40350_, _30819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40351_, _40350_, _30808_);
  and (_40352_, _40351_, _39977_);
  nand (_40353_, _39977_, _39623_);
  and (_40354_, _40353_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40355_, _40354_, _39980_);
  or (_40356_, _40355_, _40352_);
  nand (_40357_, _39980_, _38613_);
  and (_40358_, _40357_, _42003_);
  and (_42966_, _40358_, _40356_);
  and (_40359_, _39977_, _31514_);
  nand (_40360_, _40359_, _28766_);
  or (_40361_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40362_, _40361_, _39990_);
  and (_40363_, _40362_, _40360_);
  nor (_40364_, _39990_, _38592_);
  or (_40365_, _40364_, _40363_);
  and (_42968_, _40365_, _42003_);
  and (_40366_, _39977_, _32231_);
  nand (_40367_, _40366_, _28766_);
  or (_40368_, _40366_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40369_, _40368_, _39990_);
  and (_40370_, _40369_, _40367_);
  nor (_40371_, _39990_, _38506_);
  or (_40372_, _40371_, _40370_);
  and (_42970_, _40372_, _42003_);
  and (_40373_, _39977_, _33031_);
  nand (_40374_, _40373_, _28766_);
  or (_40375_, _40373_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40376_, _40375_, _39990_);
  and (_40377_, _40376_, _40374_);
  nor (_40378_, _39990_, _38452_);
  or (_40379_, _40378_, _40377_);
  and (_42972_, _40379_, _42003_);
  and (_40380_, _39977_, _33776_);
  nand (_40381_, _40380_, _28766_);
  or (_40382_, _40380_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40383_, _40382_, _39990_);
  and (_40384_, _40383_, _40381_);
  nor (_40385_, _39990_, _38364_);
  or (_40386_, _40385_, _40384_);
  and (_42973_, _40386_, _42003_);
  and (_40387_, _39959_, _24557_);
  nand (_40388_, _40387_, _28766_);
  or (_40389_, _40387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40390_, _40389_, _39969_);
  and (_40391_, _40390_, _40388_);
  and (_40392_, _39968_, _38629_);
  or (_40393_, _40392_, _40391_);
  and (_42975_, _40393_, _42003_);
  and (_40394_, _39959_, _30080_);
  nand (_40395_, _40394_, _28766_);
  or (_40396_, _40394_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40397_, _40396_, _39969_);
  and (_40398_, _40397_, _40395_);
  nor (_40399_, _39969_, _38620_);
  or (_40400_, _40399_, _40398_);
  and (_42977_, _40400_, _42003_);
  and (_40401_, _30819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40402_, _40401_, _30808_);
  and (_40403_, _40402_, _39959_);
  nand (_40404_, _39959_, _39623_);
  and (_40405_, _40404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40406_, _40405_, _39968_);
  or (_40407_, _40406_, _40403_);
  nand (_40408_, _39968_, _38613_);
  and (_40409_, _40408_, _42003_);
  and (_42979_, _40409_, _40407_);
  and (_40410_, _39959_, _31514_);
  nand (_40411_, _40410_, _28766_);
  or (_40412_, _40410_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40413_, _40412_, _39969_);
  and (_40414_, _40413_, _40411_);
  nor (_40415_, _39969_, _38592_);
  or (_40416_, _40415_, _40414_);
  and (_42981_, _40416_, _42003_);
  and (_40417_, _39959_, _32231_);
  nand (_40418_, _40417_, _28766_);
  or (_40419_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40420_, _40419_, _40418_);
  or (_40421_, _40420_, _39968_);
  nand (_40422_, _39968_, _38506_);
  and (_40423_, _40422_, _42003_);
  and (_42983_, _40423_, _40421_);
  and (_40424_, _39959_, _33031_);
  nand (_40425_, _40424_, _28766_);
  or (_40426_, _40424_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40427_, _40426_, _39969_);
  and (_40428_, _40427_, _40425_);
  nor (_40429_, _39969_, _38452_);
  or (_40430_, _40429_, _40428_);
  and (_42985_, _40430_, _42003_);
  and (_40431_, _39959_, _33776_);
  nand (_40432_, _40431_, _28766_);
  or (_40433_, _40431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40434_, _40433_, _40432_);
  or (_40435_, _40434_, _39968_);
  nand (_40436_, _39968_, _38364_);
  and (_40437_, _40436_, _42003_);
  and (_42987_, _40437_, _40435_);
  and (_40438_, _28166_, _25039_);
  not (_40439_, _40438_);
  and (_40440_, _38090_, _37914_);
  and (_40441_, _38653_, _40440_);
  not (_40442_, _40441_);
  not (_40443_, _36927_);
  and (_40444_, _37903_, _40443_);
  not (_40445_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_40446_, _39059_, _40445_);
  nor (_40447_, _40446_, _39151_);
  and (_40448_, _40447_, _39966_);
  nor (_40449_, _40447_, _39966_);
  not (_40450_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_40451_, _30819_, _40450_);
  and (_40452_, _40451_, _40438_);
  and (_40453_, _36356_, _30048_);
  nor (_40454_, _36356_, _30048_);
  nor (_40455_, _40454_, _40453_);
  and (_40456_, _40455_, _40452_);
  not (_40457_, _40456_);
  or (_40458_, _40457_, _40449_);
  nor (_40459_, _40458_, _40448_);
  nor (_40460_, _40447_, _36521_);
  and (_40461_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_40462_, _40447_, _36521_);
  and (_40463_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40464_, _40463_, _40461_);
  nor (_40465_, _40447_, _36356_);
  and (_40466_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40467_, _40447_, _36356_);
  and (_40468_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_40469_, _40468_, _40466_);
  and (_40470_, _40469_, _40464_);
  nor (_40471_, _40470_, _40459_);
  not (_40472_, _38651_);
  and (_40473_, _40459_, _40472_);
  nor (_40474_, _40473_, _40471_);
  not (_40475_, _40474_);
  and (_40476_, _40475_, _40444_);
  not (_40477_, _40476_);
  not (_40478_, _38090_);
  nor (_40479_, _37903_, _40443_);
  not (_40480_, _33939_);
  and (_40481_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_40482_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_40483_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_40484_, _40483_, _40482_);
  and (_40485_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40486_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_40487_, _40486_, _40485_);
  and (_40488_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_40489_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_40490_, _40489_, _40488_);
  and (_40491_, _40490_, _40487_);
  and (_40492_, _40491_, _40484_);
  nor (_40493_, _33994_, _40480_);
  not (_40494_, _40493_);
  nor (_40495_, _40494_, _40492_);
  nor (_40496_, _40495_, _40481_);
  not (_40497_, _40496_);
  and (_40498_, _40497_, _40479_);
  nor (_40499_, _40498_, _40478_);
  and (_40500_, _40499_, _40477_);
  and (_40501_, _40500_, _40442_);
  nor (_40502_, _37474_, _37264_);
  nor (_40503_, _37386_, _37342_);
  nor (_40504_, _37551_, _37323_);
  and (_40505_, _40504_, _40503_);
  and (_40506_, _37639_, _37441_);
  and (_40507_, _40506_, _40505_);
  and (_40508_, _40507_, _40502_);
  nor (_40509_, _40508_, _33896_);
  and (_40510_, _37606_, _36652_);
  nor (_40511_, _37815_, _40510_);
  nor (_40512_, _40511_, _37782_);
  nor (_40513_, _40512_, _40509_);
  not (_40514_, _40513_);
  and (_40515_, _40514_, _40501_);
  not (_40516_, _40447_);
  and (_40517_, _38090_, _36927_);
  and (_40518_, _40517_, _37903_);
  and (_40519_, _40518_, _40516_);
  and (_40520_, _40479_, _38090_);
  and (_40521_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_40522_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_40523_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_40524_, _40523_, _40522_);
  and (_40525_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40526_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_40527_, _40526_, _40525_);
  and (_40528_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_40529_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_40530_, _40529_, _40528_);
  and (_40531_, _40530_, _40527_);
  and (_40532_, _40531_, _40524_);
  nor (_40533_, _40532_, _40494_);
  nor (_40534_, _40533_, _40521_);
  not (_40535_, _40534_);
  and (_40536_, _40535_, _40520_);
  nor (_40537_, _40536_, _40519_);
  not (_40538_, _38679_);
  and (_40539_, _40538_, _40440_);
  and (_40540_, _40444_, _38090_);
  and (_40541_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_40542_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_40543_, _40542_, _40541_);
  and (_40544_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_40545_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_40546_, _40545_, _40544_);
  and (_40547_, _40546_, _40543_);
  nor (_40548_, _40547_, _40459_);
  not (_40549_, _38592_);
  and (_40550_, _40459_, _40549_);
  nor (_40551_, _40550_, _40548_);
  not (_40552_, _40551_);
  and (_40553_, _40552_, _40540_);
  nor (_40554_, _40553_, _40539_);
  and (_40555_, _40554_, _40537_);
  not (_40556_, _40555_);
  and (_40557_, _40556_, _40515_);
  and (_40558_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_40559_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_40560_, _40559_, _40558_);
  and (_40561_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_40562_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_40563_, _40562_, _40561_);
  and (_40564_, _40563_, _40560_);
  nor (_40565_, _40564_, _40459_);
  and (_40566_, _40459_, _38629_);
  nor (_40567_, _40566_, _40565_);
  not (_40568_, _40567_);
  and (_40569_, _40568_, _40540_);
  and (_40570_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_40571_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_40572_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_40573_, _40572_, _40571_);
  and (_40574_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40575_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_40576_, _40575_, _40574_);
  and (_40577_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_40578_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_40579_, _40578_, _40577_);
  and (_40580_, _40579_, _40576_);
  and (_40581_, _40580_, _40573_);
  nor (_40582_, _40581_, _40494_);
  nor (_40583_, _40582_, _40570_);
  not (_40584_, _40583_);
  and (_40585_, _40584_, _40520_);
  nor (_40586_, _40585_, _40569_);
  not (_40587_, _38661_);
  and (_40588_, _40587_, _40440_);
  and (_40589_, _40518_, _36521_);
  nor (_40590_, _40589_, _40588_);
  and (_40591_, _40590_, _40586_);
  nor (_40592_, _40591_, _40514_);
  nor (_40593_, _40592_, _40557_);
  and (_40594_, _25061_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40595_, _40594_, _39966_);
  nor (_40596_, _24535_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40597_, _40596_, _40595_);
  not (_40598_, _40597_);
  and (_40599_, _40598_, _40593_);
  nor (_40600_, _40599_, _40439_);
  not (_40601_, _38452_);
  and (_40602_, _40459_, _40601_);
  and (_40603_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_40604_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40605_, _40604_, _40603_);
  and (_40606_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_40607_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_40608_, _40607_, _40606_);
  and (_40609_, _40608_, _40605_);
  nor (_40610_, _40609_, _40459_);
  nor (_40611_, _40610_, _40602_);
  not (_40612_, _40611_);
  and (_40613_, _40612_, _40540_);
  not (_40614_, _40613_);
  and (_40615_, _40478_, _36927_);
  and (_40616_, _40615_, _37903_);
  not (_40617_, _38691_);
  and (_40618_, _40617_, _40440_);
  nor (_40619_, _40618_, _40616_);
  and (_40620_, _40619_, _40614_);
  and (_40621_, _40478_, _37914_);
  and (_40622_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40623_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40624_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_40625_, _40624_, _40623_);
  and (_40626_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_40627_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40628_, _40627_, _40626_);
  and (_40629_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40630_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40631_, _40630_, _40629_);
  and (_40632_, _40631_, _40628_);
  and (_40633_, _40632_, _40625_);
  nor (_40634_, _40633_, _40494_);
  nor (_40635_, _40634_, _40622_);
  not (_40636_, _40635_);
  and (_40637_, _40636_, _40520_);
  nor (_40638_, _40637_, _40621_);
  and (_40639_, _40638_, _40620_);
  not (_40640_, _40639_);
  and (_40641_, _40640_, _40515_);
  and (_40642_, _40518_, _36959_);
  and (_40643_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40644_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40645_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_40646_, _40645_, _40644_);
  and (_40647_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_40648_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40649_, _40648_, _40647_);
  and (_40650_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_40651_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_40652_, _40651_, _40650_);
  and (_40653_, _40652_, _40649_);
  and (_40654_, _40653_, _40646_);
  nor (_40655_, _40654_, _40494_);
  nor (_40656_, _40655_, _40643_);
  not (_40657_, _40656_);
  and (_40658_, _40657_, _40520_);
  nor (_40659_, _40658_, _40642_);
  not (_40660_, _38673_);
  and (_40661_, _40660_, _40440_);
  and (_40662_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_40663_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_40664_, _40663_, _40662_);
  and (_40665_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_40666_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_40667_, _40666_, _40665_);
  and (_40668_, _40667_, _40664_);
  nor (_40669_, _40668_, _40459_);
  not (_40670_, _38613_);
  and (_40671_, _40459_, _40670_);
  nor (_40672_, _40671_, _40669_);
  not (_40673_, _40672_);
  and (_40674_, _40673_, _40540_);
  nor (_40675_, _40674_, _40661_);
  and (_40676_, _40675_, _40659_);
  nor (_40677_, _40676_, _40514_);
  nor (_40678_, _40677_, _40641_);
  and (_40679_, _40594_, _39230_);
  nor (_40680_, _24293_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40681_, _40680_, _40679_);
  not (_40682_, _40681_);
  and (_40683_, _40682_, _40678_);
  nor (_40684_, _40598_, _40593_);
  nor (_40685_, _40684_, _40683_);
  and (_40686_, _40685_, _40600_);
  and (_40687_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_40688_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_40689_, _40688_, _40687_);
  and (_40690_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_40691_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_40692_, _40691_, _40690_);
  and (_40693_, _40692_, _40689_);
  nor (_40694_, _40693_, _40459_);
  not (_40695_, _38506_);
  and (_40696_, _40459_, _40695_);
  nor (_40697_, _40696_, _40694_);
  not (_40698_, _40697_);
  and (_40699_, _40698_, _40540_);
  not (_40700_, _40699_);
  not (_40701_, _38685_);
  and (_40702_, _40701_, _40440_);
  nor (_40703_, _40702_, _40615_);
  and (_40704_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40705_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40706_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_40707_, _40706_, _40705_);
  and (_40708_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40709_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_40710_, _40709_, _40708_);
  and (_40711_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_40712_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40713_, _40712_, _40711_);
  and (_40714_, _40713_, _40710_);
  and (_40715_, _40714_, _40707_);
  nor (_40716_, _40715_, _40494_);
  nor (_40717_, _40716_, _40704_);
  not (_40718_, _40717_);
  and (_40719_, _40718_, _40520_);
  and (_40720_, _40518_, _39161_);
  nor (_40721_, _40720_, _40719_);
  and (_40722_, _40721_, _40703_);
  and (_40723_, _40722_, _40700_);
  not (_40724_, _40723_);
  and (_40725_, _40724_, _40515_);
  and (_40726_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40727_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40728_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40729_, _40728_, _40727_);
  and (_40730_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40731_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_40732_, _40731_, _40730_);
  and (_40733_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_40734_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_40735_, _40734_, _40733_);
  and (_40736_, _40735_, _40732_);
  and (_40737_, _40736_, _40729_);
  nor (_40738_, _40737_, _40494_);
  nor (_40739_, _40738_, _40726_);
  not (_40740_, _40739_);
  and (_40741_, _40740_, _40520_);
  and (_40742_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_40743_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_40744_, _40743_, _40742_);
  and (_40745_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_40746_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_40747_, _40746_, _40745_);
  and (_40748_, _40747_, _40744_);
  nor (_40749_, _40748_, _40459_);
  not (_40750_, _38620_);
  and (_40751_, _40459_, _40750_);
  nor (_40752_, _40751_, _40749_);
  not (_40753_, _40752_);
  and (_40754_, _40753_, _40540_);
  nor (_40755_, _40754_, _40741_);
  not (_40756_, _38667_);
  and (_40757_, _40756_, _40440_);
  not (_40758_, _40757_);
  and (_40759_, _40444_, _40478_);
  and (_40760_, _40518_, _36367_);
  nor (_40761_, _40760_, _40759_);
  and (_40762_, _40761_, _40758_);
  and (_40763_, _40762_, _40755_);
  nor (_40764_, _40763_, _40514_);
  nor (_40765_, _40764_, _40725_);
  and (_40766_, _40594_, _25355_);
  nor (_40767_, _24414_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40768_, _40767_, _40766_);
  nand (_40771_, _40768_, _40765_);
  or (_40777_, _40768_, _40765_);
  and (_40783_, _40777_, _40771_);
  not (_40789_, _40783_);
  nor (_40795_, _40682_, _40678_);
  not (_40801_, _40795_);
  not (_40802_, _38697_);
  and (_40803_, _40802_, _40440_);
  and (_40804_, _40460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_40805_, _40462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_40806_, _40805_, _40804_);
  and (_40807_, _40465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_40808_, _40467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_40809_, _40808_, _40807_);
  and (_40810_, _40809_, _40806_);
  nor (_40811_, _40810_, _40459_);
  not (_40812_, _38364_);
  and (_40813_, _40459_, _40812_);
  nor (_40814_, _40813_, _40811_);
  not (_40815_, _40814_);
  and (_40816_, _40815_, _40540_);
  or (_40817_, _40816_, _40615_);
  nor (_40818_, _40817_, _40803_);
  and (_40819_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40820_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40821_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_40822_, _40821_, _40820_);
  and (_40823_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_40824_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40825_, _40824_, _40823_);
  and (_40826_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_40827_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_40828_, _40827_, _40826_);
  and (_40829_, _40828_, _40825_);
  and (_40830_, _40829_, _40822_);
  nor (_40831_, _40830_, _40494_);
  nor (_40832_, _40831_, _40819_);
  not (_40833_, _40832_);
  and (_40834_, _40833_, _40479_);
  nor (_40835_, _40834_, _40621_);
  and (_40836_, _40835_, _40818_);
  and (_40837_, _40836_, _40515_);
  nor (_40838_, _40556_, _40515_);
  nor (_40842_, _40838_, _40837_);
  nor (_40845_, _40594_, _39966_);
  and (_40849_, _40594_, _24754_);
  nor (_40850_, _40849_, _40845_);
  not (_40851_, _40850_);
  and (_40852_, _40851_, _40842_);
  nor (_40858_, _40851_, _40842_);
  nor (_40862_, _40858_, _40852_);
  and (_40863_, _40862_, _40801_);
  and (_40864_, _40863_, _40789_);
  and (_40867_, _40864_, _40686_);
  not (_40873_, _40678_);
  and (_40875_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40876_, _40593_);
  and (_40877_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_40883_, _40877_, _40875_);
  and (_40887_, _40883_, _40765_);
  not (_40888_, _40765_);
  not (_40889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40892_, _40593_, _40889_);
  and (_40898_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40900_, _40898_, _40892_);
  and (_40901_, _40900_, _40888_);
  or (_40903_, _40901_, _40887_);
  or (_40909_, _40903_, _40873_);
  not (_40912_, _40842_);
  and (_40913_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_40915_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_40921_, _40915_, _40913_);
  and (_40924_, _40921_, _40765_);
  not (_40925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40926_, _40593_, _40925_);
  and (_40932_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40936_, _40932_, _40926_);
  and (_40937_, _40936_, _40888_);
  or (_40938_, _40937_, _40924_);
  or (_40941_, _40938_, _40678_);
  and (_40947_, _40941_, _40912_);
  and (_40949_, _40947_, _40909_);
  or (_40950_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_40952_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40958_, _40952_, _40950_);
  and (_40961_, _40958_, _40765_);
  or (_40962_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_40970_, _40593_, _40964_);
  and (_40973_, _40970_, _40962_);
  and (_40974_, _40973_, _40888_);
  or (_40975_, _40974_, _40961_);
  or (_40981_, _40975_, _40873_);
  or (_40985_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_40986_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_40987_, _40986_, _40985_);
  and (_40992_, _40987_, _40765_);
  or (_40997_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_40998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_40999_, _40593_, _40998_);
  and (_41003_, _40999_, _40997_);
  and (_41009_, _41003_, _40888_);
  or (_41010_, _41009_, _40992_);
  or (_41011_, _41010_, _40678_);
  and (_41015_, _41011_, _40842_);
  and (_41021_, _41015_, _40981_);
  or (_41022_, _41021_, _40949_);
  or (_41023_, _41022_, _40867_);
  not (_41027_, _40867_);
  or (_41032_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_41033_, _41032_, _42003_);
  and (_43063_, _41033_, _41023_);
  nor (_41034_, _40597_, _40439_);
  nor (_41035_, _40768_, _40439_);
  and (_41036_, _41035_, _41034_);
  and (_41037_, _40850_, _40438_);
  nor (_41038_, _40681_, _40439_);
  and (_41039_, _41038_, _41037_);
  and (_41040_, _41039_, _41036_);
  and (_41041_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_41042_, _41041_, _25845_);
  nor (_41043_, _41042_, _28766_);
  nand (_41044_, _25845_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41045_, _17543_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41046_, _41045_, _41044_);
  nor (_41047_, _38651_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_41048_, _41047_, _41046_);
  or (_41049_, _41048_, _41043_);
  and (_41050_, _41049_, _40438_);
  and (_41051_, _41050_, _41040_);
  not (_41052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_41053_, _41040_, _41052_);
  or (_43069_, _41053_, _41051_);
  nor (_41054_, _41038_, _41037_);
  nor (_41055_, _41035_, _41034_);
  and (_41056_, _41055_, _40438_);
  and (_41057_, _41056_, _41054_);
  and (_41058_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25834_);
  and (_41059_, _41058_, _25878_);
  not (_41060_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41061_, _38628_, _41060_);
  or (_41062_, _16383_, _41060_);
  and (_41063_, _41062_, _41061_);
  or (_41064_, _41063_, _41059_);
  nand (_41065_, _41059_, _28766_);
  and (_41066_, _41065_, _41064_);
  and (_41067_, _41066_, _41057_);
  not (_41068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_41069_, _41057_, _41068_);
  or (_43333_, _41069_, _41067_);
  nand (_41070_, _41058_, _25954_);
  nor (_41071_, _41070_, _28766_);
  nor (_41072_, _38620_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41073_, _41058_, _25911_);
  and (_41074_, _41058_, _25845_);
  or (_41075_, _41074_, _41041_);
  or (_41076_, _41075_, _41073_);
  and (_41077_, _41076_, _17369_);
  or (_41078_, _41077_, _41072_);
  or (_41079_, _41078_, _41071_);
  and (_41080_, _41079_, _41057_);
  not (_41081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_41082_, _41057_, _41081_);
  or (_43339_, _41082_, _41080_);
  not (_41083_, _41057_);
  and (_41084_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_41085_, _41058_, _25921_);
  nor (_41086_, _41085_, _28766_);
  nor (_41087_, _38613_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41088_, _41058_, _25943_);
  or (_41089_, _41088_, _41075_);
  and (_41090_, _41089_, _16021_);
  or (_41091_, _41090_, _41087_);
  or (_41092_, _41091_, _41086_);
  and (_41093_, _41092_, _41057_);
  or (_43345_, _41093_, _41084_);
  and (_41094_, _41074_, _29375_);
  nor (_41095_, _38592_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_41096_, _41073_, _41041_);
  or (_41097_, _41096_, _41088_);
  and (_41098_, _41097_, _17053_);
  or (_41099_, _41098_, _41095_);
  or (_41100_, _41099_, _41094_);
  and (_41101_, _41100_, _41057_);
  and (_41102_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_43351_, _41102_, _41101_);
  nand (_41103_, _41041_, _25878_);
  nor (_41104_, _41103_, _28766_);
  nor (_41105_, _38506_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41106_, _25878_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41107_, _16218_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41108_, _41107_, _41106_);
  or (_41109_, _41108_, _41105_);
  or (_41110_, _41109_, _41104_);
  and (_41111_, _41110_, _41057_);
  and (_41112_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_43357_, _41112_, _41111_);
  and (_41113_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_41114_, _41041_, _25954_);
  nor (_41115_, _41114_, _28766_);
  nor (_41116_, _38452_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41117_, _25954_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41118_, _17205_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41119_, _41118_, _41117_);
  or (_41120_, _41119_, _41116_);
  or (_41121_, _41120_, _41115_);
  and (_41122_, _41121_, _41057_);
  or (_43363_, _41122_, _41113_);
  nand (_41123_, _41041_, _25921_);
  nor (_41124_, _41123_, _28766_);
  nor (_41125_, _38364_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41126_, _25921_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41127_, _16559_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41128_, _41127_, _41126_);
  or (_41129_, _41128_, _41125_);
  or (_41130_, _41129_, _41124_);
  and (_41131_, _41130_, _41057_);
  and (_41132_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_43369_, _41132_, _41131_);
  and (_41133_, _41057_, _41049_);
  and (_41134_, _41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_43372_, _41134_, _41133_);
  and (_41135_, _41066_, _40438_);
  and (_41136_, _41034_, _40768_);
  and (_41137_, _41136_, _41054_);
  and (_41138_, _41137_, _41135_);
  not (_41139_, _41137_);
  and (_41140_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_43380_, _41140_, _41138_);
  and (_41141_, _41079_, _40438_);
  and (_41142_, _41137_, _41141_);
  and (_41143_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_43384_, _41143_, _41142_);
  and (_41144_, _41092_, _40438_);
  and (_41145_, _41137_, _41144_);
  and (_41146_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_43388_, _41146_, _41145_);
  and (_41147_, _41100_, _40438_);
  and (_41148_, _41137_, _41147_);
  and (_41149_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_43392_, _41149_, _41148_);
  and (_41150_, _41110_, _40438_);
  and (_41151_, _41137_, _41150_);
  not (_41152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_41153_, _41137_, _41152_);
  or (_43396_, _41153_, _41151_);
  and (_41154_, _41121_, _40438_);
  and (_41155_, _41137_, _41154_);
  not (_41156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_41157_, _41137_, _41156_);
  or (_43400_, _41157_, _41155_);
  and (_41158_, _41130_, _40438_);
  and (_41159_, _41137_, _41158_);
  and (_41160_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_43404_, _41160_, _41159_);
  and (_41161_, _41137_, _41050_);
  and (_41162_, _41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_43407_, _41162_, _41161_);
  and (_41163_, _41035_, _40597_);
  and (_41164_, _41163_, _41054_);
  and (_41165_, _41164_, _41135_);
  not (_41166_, _41164_);
  and (_41167_, _41166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43415_, _41167_, _41165_);
  and (_41168_, _41164_, _41141_);
  and (_41169_, _41166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43419_, _41169_, _41168_);
  and (_41170_, _41164_, _41144_);
  not (_41171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_41172_, _41164_, _41171_);
  or (_43423_, _41172_, _41170_);
  and (_41173_, _41164_, _41147_);
  not (_41174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_41175_, _41164_, _41174_);
  or (_43427_, _41175_, _41173_);
  and (_41176_, _41164_, _41150_);
  not (_41177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_41178_, _41164_, _41177_);
  or (_43431_, _41178_, _41176_);
  and (_41179_, _41164_, _41154_);
  not (_41180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_41181_, _41164_, _41180_);
  or (_43435_, _41181_, _41179_);
  and (_41182_, _41164_, _41158_);
  and (_41183_, _41166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43439_, _41183_, _41182_);
  and (_41184_, _41164_, _41050_);
  not (_41185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_41186_, _41164_, _41185_);
  or (_43442_, _41186_, _41184_);
  and (_41187_, _41054_, _41036_);
  and (_41188_, _41187_, _41135_);
  not (_41189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_41190_, _41187_, _41189_);
  or (_43448_, _41190_, _41188_);
  and (_41191_, _41187_, _41141_);
  not (_41192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_41193_, _41187_, _41192_);
  or (_43452_, _41193_, _41191_);
  and (_41194_, _41187_, _41144_);
  not (_41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_41196_, _41187_, _41195_);
  or (_43456_, _41196_, _41194_);
  and (_41197_, _41187_, _41147_);
  not (_41198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_41199_, _41187_, _41198_);
  or (_43460_, _41199_, _41197_);
  and (_41200_, _41187_, _41150_);
  not (_41201_, _41187_);
  and (_41202_, _41201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_43464_, _41202_, _41200_);
  and (_41203_, _41187_, _41154_);
  and (_41204_, _41201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_43468_, _41204_, _41203_);
  and (_41205_, _41187_, _41158_);
  and (_41206_, _41201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_43472_, _41206_, _41205_);
  and (_41207_, _41187_, _41050_);
  nor (_41208_, _41187_, _40889_);
  or (_43475_, _41208_, _41207_);
  and (_41209_, _41038_, _40851_);
  and (_41210_, _41209_, _41055_);
  and (_41211_, _41210_, _41135_);
  not (_41212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41213_, _41210_, _41212_);
  or (_43483_, _41213_, _41211_);
  and (_41214_, _41210_, _41141_);
  not (_41215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41216_, _41210_, _41215_);
  or (_43487_, _41216_, _41214_);
  and (_41217_, _41210_, _41144_);
  not (_41218_, _41210_);
  and (_41219_, _41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_43491_, _41219_, _41217_);
  and (_41220_, _41210_, _41147_);
  and (_41221_, _41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_43495_, _41221_, _41220_);
  and (_41222_, _41210_, _41150_);
  and (_41223_, _41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_43499_, _41223_, _41222_);
  and (_41224_, _41210_, _41154_);
  and (_41225_, _41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_43503_, _41225_, _41224_);
  and (_41226_, _41210_, _41158_);
  not (_41227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41228_, _41210_, _41227_);
  or (_43506_, _41228_, _41226_);
  and (_41229_, _41210_, _41050_);
  and (_41230_, _41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_43509_, _41230_, _41229_);
  and (_41231_, _41209_, _41136_);
  and (_41232_, _41231_, _41135_);
  not (_41233_, _41231_);
  and (_41234_, _41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_43514_, _41234_, _41232_);
  and (_41235_, _41231_, _41141_);
  and (_41236_, _41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_43518_, _41236_, _41235_);
  and (_41237_, _41231_, _41144_);
  and (_41238_, _41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_43522_, _41238_, _41237_);
  and (_41239_, _41231_, _41147_);
  and (_41240_, _41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_43526_, _41240_, _41239_);
  and (_41241_, _41231_, _41150_);
  not (_41242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_41243_, _41231_, _41242_);
  or (_43530_, _41243_, _41241_);
  and (_41244_, _41231_, _41154_);
  not (_41245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_41246_, _41231_, _41245_);
  or (_43534_, _41246_, _41244_);
  and (_41247_, _41231_, _41158_);
  not (_41248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_41249_, _41231_, _41248_);
  or (_43538_, _41249_, _41247_);
  and (_41250_, _41231_, _41050_);
  and (_41251_, _41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_43541_, _41251_, _41250_);
  and (_41252_, _41209_, _41163_);
  and (_41253_, _41252_, _41135_);
  not (_41254_, _41252_);
  and (_41255_, _41254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43546_, _41255_, _41253_);
  and (_41256_, _41252_, _41141_);
  and (_41257_, _41254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43550_, _41257_, _41256_);
  and (_41258_, _41252_, _41144_);
  not (_41259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_41260_, _41252_, _41259_);
  or (_43554_, _41260_, _41258_);
  and (_41261_, _41252_, _41147_);
  not (_41262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_41263_, _41252_, _41262_);
  or (_43558_, _41263_, _41261_);
  and (_41264_, _41252_, _41150_);
  not (_41265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_41266_, _41252_, _41265_);
  or (_43562_, _41266_, _41264_);
  and (_41267_, _41252_, _41154_);
  not (_41268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_41269_, _41252_, _41268_);
  or (_43566_, _41269_, _41267_);
  and (_41270_, _41252_, _41158_);
  not (_41271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_41272_, _41252_, _41271_);
  or (_43570_, _41272_, _41270_);
  and (_41273_, _41252_, _41050_);
  not (_41274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_41275_, _41252_, _41274_);
  or (_43573_, _41275_, _41273_);
  and (_41276_, _41209_, _41036_);
  and (_41277_, _41276_, _41135_);
  not (_41278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_41279_, _41276_, _41278_);
  or (_43578_, _41279_, _41277_);
  and (_41280_, _41276_, _41141_);
  not (_41281_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_41282_, _41276_, _41281_);
  or (_43582_, _41282_, _41280_);
  and (_41283_, _41276_, _41144_);
  not (_41284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_41285_, _41276_, _41284_);
  or (_43586_, _41285_, _41283_);
  and (_41286_, _41276_, _41147_);
  not (_41287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_41288_, _41276_, _41287_);
  or (_43590_, _41288_, _41286_);
  and (_41289_, _41276_, _41150_);
  not (_41290_, _41276_);
  and (_41291_, _41290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_43594_, _41291_, _41289_);
  and (_41292_, _41276_, _41154_);
  and (_41293_, _41290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_43598_, _41293_, _41292_);
  and (_41294_, _41276_, _41158_);
  not (_41295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_41296_, _41276_, _41295_);
  or (_43602_, _41296_, _41294_);
  and (_41297_, _41276_, _41050_);
  nor (_41298_, _41276_, _40925_);
  or (_43605_, _41298_, _41297_);
  and (_41299_, _41037_, _40681_);
  and (_41300_, _41299_, _41055_);
  and (_41301_, _41300_, _41135_);
  not (_41302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_41303_, _41300_, _41302_);
  or (_43613_, _41303_, _41301_);
  and (_41304_, _41300_, _41141_);
  not (_41305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_41306_, _41300_, _41305_);
  or (_43617_, _41306_, _41304_);
  and (_41307_, _41300_, _41144_);
  not (_41308_, _41300_);
  and (_41309_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_43621_, _41309_, _41307_);
  and (_41310_, _41300_, _41147_);
  and (_41311_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_43625_, _41311_, _41310_);
  and (_41312_, _41300_, _41150_);
  and (_41313_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_43629_, _41313_, _41312_);
  and (_41314_, _41300_, _41154_);
  and (_41315_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_43633_, _41315_, _41314_);
  and (_41316_, _41300_, _41158_);
  and (_41317_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_43637_, _41317_, _41316_);
  and (_41318_, _41300_, _41050_);
  and (_41319_, _41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_43640_, _41319_, _41318_);
  and (_41320_, _41299_, _41136_);
  and (_41321_, _41320_, _41135_);
  not (_41322_, _41320_);
  and (_41323_, _41322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_43645_, _41323_, _41321_);
  and (_41324_, _41320_, _41141_);
  and (_41325_, _41322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_43649_, _41325_, _41324_);
  and (_41326_, _41320_, _41144_);
  and (_41327_, _41322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_43653_, _41327_, _41326_);
  and (_41328_, _41320_, _41147_);
  not (_41329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_41330_, _41320_, _41329_);
  or (_43657_, _41330_, _41328_);
  and (_41331_, _41320_, _41150_);
  not (_41332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_41333_, _41320_, _41332_);
  or (_43661_, _41333_, _41331_);
  and (_41334_, _41320_, _41154_);
  not (_41335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_41336_, _41320_, _41335_);
  or (_43665_, _41336_, _41334_);
  and (_41337_, _41320_, _41158_);
  not (_41338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_41339_, _41320_, _41338_);
  or (_43669_, _41339_, _41337_);
  and (_41340_, _41320_, _41050_);
  and (_41341_, _41322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_43672_, _41341_, _41340_);
  and (_41342_, _41299_, _41163_);
  and (_41343_, _41342_, _41135_);
  not (_41344_, _41342_);
  and (_41345_, _41344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_43677_, _41345_, _41343_);
  and (_41346_, _41342_, _41141_);
  and (_41347_, _41344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_43681_, _41347_, _41346_);
  and (_41348_, _41342_, _41144_);
  not (_41349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_41350_, _41342_, _41349_);
  or (_43685_, _41350_, _41348_);
  and (_41351_, _41342_, _41147_);
  not (_41352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_41353_, _41342_, _41352_);
  or (_43689_, _41353_, _41351_);
  and (_41354_, _41342_, _41150_);
  not (_41355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_41356_, _41342_, _41355_);
  or (_43693_, _41356_, _41354_);
  and (_41357_, _41342_, _41154_);
  not (_41358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_41359_, _41342_, _41358_);
  or (_43697_, _41359_, _41357_);
  and (_41360_, _41342_, _41158_);
  not (_41361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_41362_, _41342_, _41361_);
  or (_43701_, _41362_, _41360_);
  and (_41363_, _41342_, _41050_);
  nor (_41364_, _41342_, _40964_);
  or (_43704_, _41364_, _41363_);
  and (_41365_, _41299_, _41036_);
  and (_41366_, _41365_, _41135_);
  not (_41367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_41368_, _41365_, _41367_);
  or (_43709_, _41368_, _41366_);
  and (_41369_, _41365_, _41141_);
  not (_41370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_41371_, _41365_, _41370_);
  or (_43713_, _41371_, _41369_);
  and (_41372_, _41365_, _41144_);
  not (_41373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_41374_, _41365_, _41373_);
  or (_43717_, _41374_, _41372_);
  and (_41375_, _41365_, _41147_);
  not (_41376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_41377_, _41365_, _41376_);
  or (_43721_, _41377_, _41375_);
  and (_41378_, _41365_, _41150_);
  not (_41379_, _41365_);
  and (_41380_, _41379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_43725_, _41380_, _41378_);
  and (_41381_, _41365_, _41154_);
  and (_41382_, _41379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_43729_, _41382_, _41381_);
  and (_41383_, _41365_, _41158_);
  and (_41384_, _41379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_43735_, _41384_, _41383_);
  and (_41385_, _41365_, _41050_);
  not (_41386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_41387_, _41365_, _41386_);
  or (_43750_, _41387_, _41385_);
  and (_41388_, _41055_, _41039_);
  and (_41389_, _41388_, _41135_);
  not (_41390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_41391_, _41388_, _41390_);
  or (_43779_, _41391_, _41389_);
  and (_41392_, _41388_, _41141_);
  not (_41393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_41394_, _41388_, _41393_);
  or (_43799_, _41394_, _41392_);
  and (_41395_, _41388_, _41144_);
  not (_41396_, _41388_);
  and (_41397_, _41396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_43819_, _41397_, _41395_);
  and (_41398_, _41388_, _41147_);
  not (_41399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_41400_, _41388_, _41399_);
  or (_43838_, _41400_, _41398_);
  and (_41401_, _41388_, _41150_);
  and (_41402_, _41396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_43856_, _41402_, _41401_);
  and (_41405_, _41388_, _41154_);
  and (_41407_, _41396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_43874_, _41407_, _41405_);
  and (_41410_, _41388_, _41158_);
  not (_41412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_41414_, _41388_, _41412_);
  or (_43892_, _41414_, _41410_);
  and (_41417_, _41388_, _41050_);
  and (_41419_, _41396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_43908_, _41419_, _41417_);
  and (_41422_, _41136_, _41039_);
  and (_41424_, _41422_, _41135_);
  not (_41426_, _41422_);
  and (_41428_, _41426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_43931_, _41428_, _41424_);
  and (_41431_, _41422_, _41141_);
  and (_41433_, _41426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_43951_, _41433_, _41431_);
  and (_41436_, _41422_, _41144_);
  and (_41438_, _41426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_43971_, _41438_, _41436_);
  and (_41441_, _41422_, _41147_);
  and (_41443_, _41426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_43976_, _41443_, _41441_);
  and (_41446_, _41422_, _41150_);
  not (_41448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_41450_, _41422_, _41448_);
  or (_43980_, _41450_, _41446_);
  and (_41451_, _41422_, _41154_);
  not (_41452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_41453_, _41422_, _41452_);
  or (_43984_, _41453_, _41451_);
  and (_41454_, _41422_, _41158_);
  not (_41455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_41456_, _41422_, _41455_);
  or (_43988_, _41456_, _41454_);
  and (_41457_, _41422_, _41050_);
  and (_41458_, _41426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_43991_, _41458_, _41457_);
  and (_41459_, _41163_, _41039_);
  and (_41460_, _41459_, _41135_);
  not (_41461_, _41459_);
  and (_41462_, _41461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_43996_, _41462_, _41460_);
  and (_41463_, _41459_, _41141_);
  and (_41464_, _41461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_44000_, _41464_, _41463_);
  and (_41465_, _41459_, _41144_);
  not (_41466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_41467_, _41459_, _41466_);
  or (_44002_, _41467_, _41465_);
  and (_41468_, _41459_, _41147_);
  and (_41469_, _41461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_44005_, _41469_, _41468_);
  and (_41470_, _41459_, _41150_);
  not (_41471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_41472_, _41459_, _41471_);
  or (_44009_, _41472_, _41470_);
  and (_41473_, _41459_, _41154_);
  not (_41474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_41475_, _41459_, _41474_);
  or (_44013_, _41475_, _41473_);
  and (_41476_, _41459_, _41158_);
  not (_41477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_41478_, _41459_, _41477_);
  or (_44017_, _41478_, _41476_);
  and (_41479_, _41459_, _41050_);
  nor (_41480_, _41459_, _40998_);
  or (_44020_, _41480_, _41479_);
  and (_41481_, _41135_, _41040_);
  not (_41482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_41483_, _41040_, _41482_);
  or (_44023_, _41483_, _41481_);
  and (_41484_, _41141_, _41040_);
  not (_41485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_41486_, _41040_, _41485_);
  or (_44027_, _41486_, _41484_);
  and (_41487_, _41144_, _41040_);
  not (_41488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_41489_, _41040_, _41488_);
  or (_44031_, _41489_, _41487_);
  and (_41490_, _41147_, _41040_);
  not (_41491_, _41040_);
  and (_41492_, _41491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_44035_, _41492_, _41490_);
  and (_41493_, _41150_, _41040_);
  and (_41494_, _41491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_44039_, _41494_, _41493_);
  and (_41495_, _41154_, _41040_);
  and (_41496_, _41491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_44043_, _41496_, _41495_);
  and (_41497_, _41158_, _41040_);
  not (_41498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_41499_, _41040_, _41498_);
  or (_44046_, _41499_, _41497_);
  or (_41500_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_41501_, _40593_, _41068_);
  and (_41502_, _41501_, _40765_);
  and (_41503_, _41502_, _41500_);
  nor (_41504_, _40593_, _41189_);
  and (_41505_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41506_, _41505_, _41504_);
  and (_41507_, _41506_, _40888_);
  or (_41508_, _41507_, _41503_);
  or (_41509_, _41508_, _40873_);
  or (_41510_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_41511_, _40593_, _41212_);
  and (_41512_, _41511_, _40765_);
  and (_41513_, _41512_, _41510_);
  nor (_41514_, _40593_, _41278_);
  and (_41515_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41516_, _41515_, _41514_);
  and (_41517_, _41516_, _40888_);
  or (_41518_, _41517_, _41513_);
  or (_41519_, _41518_, _40678_);
  and (_41520_, _41519_, _40912_);
  and (_41521_, _41520_, _41509_);
  nand (_41522_, _40593_, _41302_);
  or (_41523_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_41524_, _41523_, _41522_);
  and (_41525_, _41524_, _40765_);
  and (_41526_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_41527_, _40593_, _41367_);
  or (_41528_, _41527_, _41526_);
  and (_41529_, _41528_, _40888_);
  or (_41530_, _41529_, _41525_);
  or (_41531_, _41530_, _40873_);
  nand (_41532_, _40593_, _41390_);
  or (_41533_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_41534_, _41533_, _41532_);
  and (_41535_, _41534_, _40765_);
  and (_41536_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_41537_, _40593_, _41482_);
  or (_41538_, _41537_, _41536_);
  and (_41539_, _41538_, _40888_);
  or (_41540_, _41539_, _41535_);
  or (_41541_, _41540_, _40678_);
  and (_41542_, _41541_, _40842_);
  and (_41543_, _41542_, _41531_);
  or (_41544_, _41543_, _41521_);
  or (_41545_, _41544_, _40867_);
  or (_41546_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_41547_, _41546_, _42003_);
  and (_01414_, _41547_, _41545_);
  or (_41548_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_41549_, _40593_, _41081_);
  and (_41550_, _41549_, _40765_);
  and (_41551_, _41550_, _41548_);
  nor (_41552_, _40593_, _41192_);
  and (_41553_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41554_, _41553_, _41552_);
  and (_41555_, _41554_, _40888_);
  or (_41556_, _41555_, _41551_);
  or (_41557_, _41556_, _40873_);
  or (_41558_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_41559_, _40593_, _41215_);
  and (_41560_, _41559_, _40765_);
  and (_41561_, _41560_, _41558_);
  nor (_41562_, _40593_, _41281_);
  and (_41563_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41564_, _41563_, _41562_);
  and (_41565_, _41564_, _40888_);
  or (_41566_, _41565_, _41561_);
  or (_41567_, _41566_, _40678_);
  and (_41568_, _41567_, _40912_);
  and (_41569_, _41568_, _41557_);
  nand (_41570_, _40593_, _41305_);
  or (_41571_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_41572_, _41571_, _41570_);
  and (_41573_, _41572_, _40765_);
  and (_41574_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_41575_, _40593_, _41370_);
  or (_41576_, _41575_, _41574_);
  and (_41577_, _41576_, _40888_);
  or (_41578_, _41577_, _41573_);
  or (_41579_, _41578_, _40873_);
  nand (_41580_, _40593_, _41393_);
  or (_41581_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_41582_, _41581_, _41580_);
  and (_41583_, _41582_, _40765_);
  and (_41584_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_41585_, _40593_, _41485_);
  or (_41586_, _41585_, _41584_);
  and (_41587_, _41586_, _40888_);
  or (_41588_, _41587_, _41583_);
  or (_41589_, _41588_, _40678_);
  and (_41590_, _41589_, _40842_);
  and (_41591_, _41590_, _41579_);
  or (_41592_, _41591_, _41569_);
  or (_41593_, _41592_, _40867_);
  or (_41594_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_41595_, _41594_, _42003_);
  and (_01416_, _41595_, _41593_);
  and (_41596_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_41597_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_41598_, _41597_, _41596_);
  and (_41599_, _41598_, _40765_);
  nor (_41600_, _40593_, _41195_);
  and (_41601_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_41602_, _41601_, _41600_);
  and (_41603_, _41602_, _40888_);
  or (_41604_, _41603_, _41599_);
  or (_41605_, _41604_, _40873_);
  and (_41606_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_41607_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_41608_, _41607_, _41606_);
  and (_41609_, _41608_, _40765_);
  nor (_41610_, _40593_, _41284_);
  and (_41611_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_41612_, _41611_, _41610_);
  and (_41613_, _41612_, _40888_);
  or (_41614_, _41613_, _41609_);
  or (_41615_, _41614_, _40678_);
  and (_41616_, _41615_, _40912_);
  and (_41617_, _41616_, _41605_);
  or (_41618_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_41619_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_41620_, _41619_, _41618_);
  and (_41621_, _41620_, _40765_);
  or (_41622_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_41623_, _40593_, _41349_);
  and (_41624_, _41623_, _41622_);
  and (_41625_, _41624_, _40888_);
  or (_41626_, _41625_, _41621_);
  or (_41627_, _41626_, _40873_);
  or (_41628_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_41629_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_41630_, _41629_, _41628_);
  and (_41631_, _41630_, _40765_);
  or (_41632_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_41633_, _40593_, _41466_);
  and (_41634_, _41633_, _41632_);
  and (_41635_, _41634_, _40888_);
  or (_41636_, _41635_, _41631_);
  or (_41637_, _41636_, _40678_);
  and (_41638_, _41637_, _40842_);
  and (_41639_, _41638_, _41627_);
  or (_41640_, _41639_, _41617_);
  or (_41641_, _41640_, _40867_);
  or (_41642_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41643_, _41642_, _42003_);
  and (_01418_, _41643_, _41641_);
  or (_41644_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_41645_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_41646_, _41645_, _41644_);
  or (_41647_, _41646_, _40765_);
  nand (_41648_, _40593_, _41399_);
  or (_41649_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41650_, _41649_, _41648_);
  or (_41651_, _41650_, _40888_);
  and (_41652_, _41651_, _40842_);
  and (_41653_, _41652_, _41647_);
  and (_41654_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_41655_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_41656_, _41655_, _40888_);
  or (_41657_, _41656_, _41654_);
  nor (_41658_, _40593_, _41287_);
  and (_41659_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41660_, _41659_, _40765_);
  or (_41661_, _41660_, _41658_);
  and (_41662_, _41661_, _40912_);
  and (_41663_, _41662_, _41657_);
  or (_41664_, _41663_, _41653_);
  and (_41665_, _41664_, _40873_);
  or (_41666_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41667_, _40593_, _41352_);
  and (_41668_, _41667_, _41666_);
  or (_41669_, _41668_, _40765_);
  and (_41670_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_41671_, _40593_, _41329_);
  or (_41672_, _41671_, _41670_);
  or (_41673_, _41672_, _40888_);
  and (_41674_, _41673_, _40842_);
  and (_41675_, _41674_, _41669_);
  and (_41676_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_41677_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_41678_, _41677_, _40888_);
  or (_41679_, _41678_, _41676_);
  nor (_41680_, _40593_, _41198_);
  and (_41681_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41682_, _41681_, _40765_);
  or (_41683_, _41682_, _41680_);
  and (_41684_, _41683_, _40912_);
  and (_41685_, _41684_, _41679_);
  or (_41686_, _41685_, _41675_);
  and (_41687_, _41686_, _40678_);
  or (_41688_, _41687_, _40867_);
  or (_41689_, _41688_, _41665_);
  or (_41690_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41691_, _41690_, _42003_);
  and (_01420_, _41691_, _41689_);
  and (_41692_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41693_, _40593_, _41152_);
  or (_41694_, _41693_, _41692_);
  and (_41695_, _41694_, _40765_);
  or (_41696_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_41697_, _40593_, _41177_);
  and (_41698_, _41697_, _41696_);
  and (_41699_, _41698_, _40888_);
  or (_41700_, _41699_, _41695_);
  or (_41701_, _41700_, _40873_);
  and (_41702_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41703_, _40593_, _41242_);
  or (_41704_, _41703_, _41702_);
  and (_41705_, _41704_, _40765_);
  or (_41706_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_41707_, _40593_, _41265_);
  and (_41708_, _41707_, _41706_);
  and (_41709_, _41708_, _40888_);
  or (_41710_, _41709_, _41705_);
  or (_41711_, _41710_, _40678_);
  and (_41712_, _41711_, _40912_);
  and (_41713_, _41712_, _41701_);
  and (_41714_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41715_, _40593_, _41332_);
  or (_41716_, _41715_, _41714_);
  and (_41717_, _41716_, _40765_);
  or (_41718_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41719_, _40593_, _41355_);
  and (_41720_, _41719_, _41718_);
  and (_41721_, _41720_, _40888_);
  or (_41722_, _41721_, _41717_);
  or (_41723_, _41722_, _40873_);
  and (_41724_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41725_, _40593_, _41448_);
  or (_41726_, _41725_, _41724_);
  and (_41727_, _41726_, _40765_);
  or (_41728_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41729_, _40593_, _41471_);
  and (_41730_, _41729_, _41728_);
  and (_41731_, _41730_, _40888_);
  or (_41732_, _41731_, _41727_);
  or (_41733_, _41732_, _40678_);
  and (_41734_, _41733_, _40842_);
  and (_41735_, _41734_, _41723_);
  or (_41736_, _41735_, _41713_);
  or (_41737_, _41736_, _40867_);
  or (_41738_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41739_, _41738_, _42003_);
  and (_01422_, _41739_, _41737_);
  and (_41740_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41741_, _40593_, _41156_);
  or (_41742_, _41741_, _41740_);
  and (_41743_, _41742_, _40765_);
  or (_41744_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_41745_, _40593_, _41180_);
  and (_41746_, _41745_, _41744_);
  and (_41747_, _41746_, _40888_);
  or (_41748_, _41747_, _41743_);
  or (_41749_, _41748_, _40873_);
  and (_41750_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41751_, _40593_, _41245_);
  or (_41752_, _41751_, _41750_);
  and (_41753_, _41752_, _40765_);
  or (_41754_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_41755_, _40593_, _41268_);
  and (_41756_, _41755_, _41754_);
  and (_41757_, _41756_, _40888_);
  or (_41758_, _41757_, _41753_);
  or (_41759_, _41758_, _40678_);
  and (_41760_, _41759_, _40912_);
  and (_41761_, _41760_, _41749_);
  and (_41762_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41763_, _40593_, _41335_);
  or (_41764_, _41763_, _41762_);
  and (_41765_, _41764_, _40765_);
  or (_41766_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41767_, _40593_, _41358_);
  and (_41768_, _41767_, _41766_);
  and (_41769_, _41768_, _40888_);
  or (_41770_, _41769_, _41765_);
  or (_41771_, _41770_, _40873_);
  and (_41772_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41773_, _40593_, _41452_);
  or (_41774_, _41773_, _41772_);
  and (_41775_, _41774_, _40765_);
  or (_41776_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41777_, _40593_, _41474_);
  and (_41778_, _41777_, _41776_);
  and (_41779_, _41778_, _40888_);
  or (_41780_, _41779_, _41775_);
  or (_41781_, _41780_, _40678_);
  and (_41782_, _41781_, _40842_);
  and (_41783_, _41782_, _41771_);
  or (_41784_, _41783_, _41761_);
  or (_41785_, _41784_, _40867_);
  or (_41786_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41787_, _41786_, _42003_);
  and (_01424_, _41787_, _41785_);
  and (_41788_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_41789_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_41790_, _41789_, _41788_);
  and (_41791_, _41790_, _40765_);
  and (_41792_, _40876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_41793_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_41794_, _41793_, _41792_);
  and (_41795_, _41794_, _40888_);
  or (_41796_, _41795_, _41791_);
  or (_41797_, _41796_, _40873_);
  and (_41798_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41799_, _40593_, _41248_);
  or (_41800_, _41799_, _41798_);
  and (_41801_, _41800_, _40765_);
  nor (_41802_, _40593_, _41295_);
  and (_41803_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41804_, _41803_, _41802_);
  and (_41805_, _41804_, _40888_);
  or (_41806_, _41805_, _41801_);
  or (_41807_, _41806_, _40678_);
  and (_41808_, _41807_, _40912_);
  and (_41809_, _41808_, _41797_);
  and (_41810_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_41811_, _40593_, _41338_);
  or (_41812_, _41811_, _41810_);
  and (_41813_, _41812_, _40765_);
  or (_41814_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_41815_, _40593_, _41361_);
  and (_41816_, _41815_, _41814_);
  and (_41817_, _41816_, _40888_);
  or (_41818_, _41817_, _41813_);
  or (_41819_, _41818_, _40873_);
  nand (_41820_, _40593_, _41412_);
  or (_41821_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41822_, _41821_, _41820_);
  and (_41823_, _41822_, _40765_);
  or (_41824_, _40593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41825_, _40593_, _41477_);
  and (_41826_, _41825_, _41824_);
  and (_41827_, _41826_, _40888_);
  or (_41828_, _41827_, _41823_);
  or (_41829_, _41828_, _40678_);
  and (_41830_, _41829_, _40842_);
  and (_41831_, _41830_, _41819_);
  or (_41832_, _41831_, _41809_);
  or (_41833_, _41832_, _40867_);
  or (_41834_, _41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41835_, _41834_, _42003_);
  and (_01425_, _41835_, _41833_);
  or (_41836_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41837_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41838_, _41837_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41839_, _41838_, _41836_);
  nand (_41840_, _41839_, _42003_);
  or (_41841_, \oc8051_gm_cxrom_1.cell0.data [7], _42003_);
  and (_01433_, _41841_, _41840_);
  or (_41842_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41843_, \oc8051_gm_cxrom_1.cell0.data [0], _41837_);
  nand (_41844_, _41843_, _41842_);
  nand (_41845_, _41844_, _42003_);
  or (_41846_, \oc8051_gm_cxrom_1.cell0.data [0], _42003_);
  and (_01440_, _41846_, _41845_);
  or (_41847_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41848_, \oc8051_gm_cxrom_1.cell0.data [1], _41837_);
  nand (_41849_, _41848_, _41847_);
  nand (_41850_, _41849_, _42003_);
  or (_41851_, \oc8051_gm_cxrom_1.cell0.data [1], _42003_);
  and (_01444_, _41851_, _41850_);
  or (_41852_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41853_, \oc8051_gm_cxrom_1.cell0.data [2], _41837_);
  nand (_41854_, _41853_, _41852_);
  nand (_41855_, _41854_, _42003_);
  or (_41856_, \oc8051_gm_cxrom_1.cell0.data [2], _42003_);
  and (_01448_, _41856_, _41855_);
  or (_41857_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41858_, \oc8051_gm_cxrom_1.cell0.data [3], _41837_);
  nand (_41859_, _41858_, _41857_);
  nand (_41860_, _41859_, _42003_);
  or (_41861_, \oc8051_gm_cxrom_1.cell0.data [3], _42003_);
  and (_01452_, _41861_, _41860_);
  or (_41862_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41863_, \oc8051_gm_cxrom_1.cell0.data [4], _41837_);
  nand (_41864_, _41863_, _41862_);
  nand (_41865_, _41864_, _42003_);
  or (_41866_, \oc8051_gm_cxrom_1.cell0.data [4], _42003_);
  and (_01456_, _41866_, _41865_);
  or (_41867_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41868_, \oc8051_gm_cxrom_1.cell0.data [5], _41837_);
  nand (_41869_, _41868_, _41867_);
  nand (_41870_, _41869_, _42003_);
  or (_41871_, \oc8051_gm_cxrom_1.cell0.data [5], _42003_);
  and (_01460_, _41871_, _41870_);
  or (_41872_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41873_, \oc8051_gm_cxrom_1.cell0.data [6], _41837_);
  nand (_41874_, _41873_, _41872_);
  nand (_41875_, _41874_, _42003_);
  or (_41876_, \oc8051_gm_cxrom_1.cell0.data [6], _42003_);
  and (_01464_, _41876_, _41875_);
  or (_41877_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41878_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41879_, _41878_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41880_, _41879_, _41877_);
  nand (_41881_, _41880_, _42003_);
  or (_41882_, \oc8051_gm_cxrom_1.cell1.data [7], _42003_);
  and (_01485_, _41882_, _41881_);
  or (_41883_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41884_, \oc8051_gm_cxrom_1.cell1.data [0], _41878_);
  nand (_41885_, _41884_, _41883_);
  nand (_41886_, _41885_, _42003_);
  or (_41887_, \oc8051_gm_cxrom_1.cell1.data [0], _42003_);
  and (_01492_, _41887_, _41886_);
  or (_41888_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41889_, \oc8051_gm_cxrom_1.cell1.data [1], _41878_);
  nand (_41890_, _41889_, _41888_);
  nand (_41891_, _41890_, _42003_);
  or (_41892_, \oc8051_gm_cxrom_1.cell1.data [1], _42003_);
  and (_01496_, _41892_, _41891_);
  or (_41893_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41894_, \oc8051_gm_cxrom_1.cell1.data [2], _41878_);
  nand (_41895_, _41894_, _41893_);
  nand (_41896_, _41895_, _42003_);
  or (_41897_, \oc8051_gm_cxrom_1.cell1.data [2], _42003_);
  and (_01500_, _41897_, _41896_);
  or (_41898_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41899_, \oc8051_gm_cxrom_1.cell1.data [3], _41878_);
  nand (_41900_, _41899_, _41898_);
  nand (_41901_, _41900_, _42003_);
  or (_41902_, \oc8051_gm_cxrom_1.cell1.data [3], _42003_);
  and (_01503_, _41902_, _41901_);
  or (_41903_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41904_, \oc8051_gm_cxrom_1.cell1.data [4], _41878_);
  nand (_41905_, _41904_, _41903_);
  nand (_41906_, _41905_, _42003_);
  or (_41907_, \oc8051_gm_cxrom_1.cell1.data [4], _42003_);
  and (_01507_, _41907_, _41906_);
  or (_41908_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41909_, \oc8051_gm_cxrom_1.cell1.data [5], _41878_);
  nand (_41910_, _41909_, _41908_);
  nand (_41911_, _41910_, _42003_);
  or (_41912_, \oc8051_gm_cxrom_1.cell1.data [5], _42003_);
  and (_01511_, _41912_, _41911_);
  or (_41913_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41914_, \oc8051_gm_cxrom_1.cell1.data [6], _41878_);
  nand (_41915_, _41914_, _41913_);
  nand (_41916_, _41915_, _42003_);
  or (_41917_, \oc8051_gm_cxrom_1.cell1.data [6], _42003_);
  and (_01515_, _41917_, _41916_);
  or (_41918_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41919_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41920_, _41919_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41921_, _41920_, _41918_);
  nand (_41922_, _41921_, _42003_);
  or (_41923_, \oc8051_gm_cxrom_1.cell2.data [7], _42003_);
  and (_01537_, _41923_, _41922_);
  or (_41924_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41925_, \oc8051_gm_cxrom_1.cell2.data [0], _41919_);
  nand (_41926_, _41925_, _41924_);
  nand (_41927_, _41926_, _42003_);
  or (_41928_, \oc8051_gm_cxrom_1.cell2.data [0], _42003_);
  and (_01543_, _41928_, _41927_);
  or (_41929_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41930_, \oc8051_gm_cxrom_1.cell2.data [1], _41919_);
  nand (_41931_, _41930_, _41929_);
  nand (_41932_, _41931_, _42003_);
  or (_41933_, \oc8051_gm_cxrom_1.cell2.data [1], _42003_);
  and (_01547_, _41933_, _41932_);
  or (_41934_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41935_, \oc8051_gm_cxrom_1.cell2.data [2], _41919_);
  nand (_41936_, _41935_, _41934_);
  nand (_41937_, _41936_, _42003_);
  or (_41938_, \oc8051_gm_cxrom_1.cell2.data [2], _42003_);
  and (_01551_, _41938_, _41937_);
  or (_41939_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41940_, \oc8051_gm_cxrom_1.cell2.data [3], _41919_);
  nand (_41941_, _41940_, _41939_);
  nand (_41942_, _41941_, _42003_);
  or (_41943_, \oc8051_gm_cxrom_1.cell2.data [3], _42003_);
  and (_01555_, _41943_, _41942_);
  or (_41944_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41946_, \oc8051_gm_cxrom_1.cell2.data [4], _41919_);
  nand (_41947_, _41946_, _41944_);
  nand (_41949_, _41947_, _42003_);
  or (_41951_, \oc8051_gm_cxrom_1.cell2.data [4], _42003_);
  and (_01559_, _41951_, _41949_);
  or (_41953_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41955_, \oc8051_gm_cxrom_1.cell2.data [5], _41919_);
  nand (_41957_, _41955_, _41953_);
  nand (_41959_, _41957_, _42003_);
  or (_41960_, \oc8051_gm_cxrom_1.cell2.data [5], _42003_);
  and (_01563_, _41960_, _41959_);
  or (_41961_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41962_, \oc8051_gm_cxrom_1.cell2.data [6], _41919_);
  nand (_41963_, _41962_, _41961_);
  nand (_41964_, _41963_, _42003_);
  or (_41965_, \oc8051_gm_cxrom_1.cell2.data [6], _42003_);
  and (_01567_, _41965_, _41964_);
  or (_41966_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_41967_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_41968_, _41967_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_41969_, _41968_, _41966_);
  nand (_41970_, _41969_, _42003_);
  or (_41971_, \oc8051_gm_cxrom_1.cell3.data [7], _42003_);
  and (_01588_, _41971_, _41970_);
  or (_41972_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41973_, \oc8051_gm_cxrom_1.cell3.data [0], _41967_);
  nand (_41974_, _41973_, _41972_);
  nand (_41975_, _41974_, _42003_);
  or (_41976_, \oc8051_gm_cxrom_1.cell3.data [0], _42003_);
  and (_01595_, _41976_, _41975_);
  or (_41977_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41978_, \oc8051_gm_cxrom_1.cell3.data [1], _41967_);
  nand (_41979_, _41978_, _41977_);
  nand (_41980_, _41979_, _42003_);
  or (_41981_, \oc8051_gm_cxrom_1.cell3.data [1], _42003_);
  and (_01599_, _41981_, _41980_);
  or (_41982_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41983_, \oc8051_gm_cxrom_1.cell3.data [2], _41967_);
  nand (_41984_, _41983_, _41982_);
  nand (_41985_, _41984_, _42003_);
  or (_41986_, \oc8051_gm_cxrom_1.cell3.data [2], _42003_);
  and (_01603_, _41986_, _41985_);
  or (_41987_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41988_, \oc8051_gm_cxrom_1.cell3.data [3], _41967_);
  nand (_41989_, _41988_, _41987_);
  nand (_41991_, _41989_, _42003_);
  or (_41993_, \oc8051_gm_cxrom_1.cell3.data [3], _42003_);
  and (_01607_, _41993_, _41991_);
  or (_41996_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41998_, \oc8051_gm_cxrom_1.cell3.data [4], _41967_);
  nand (_42000_, _41998_, _41996_);
  nand (_42002_, _42000_, _42003_);
  or (_42004_, \oc8051_gm_cxrom_1.cell3.data [4], _42003_);
  and (_01611_, _42004_, _42002_);
  or (_42005_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42006_, \oc8051_gm_cxrom_1.cell3.data [5], _41967_);
  nand (_42007_, _42006_, _42005_);
  nand (_42008_, _42007_, _42003_);
  or (_42009_, \oc8051_gm_cxrom_1.cell3.data [5], _42003_);
  and (_01615_, _42009_, _42008_);
  or (_42010_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42011_, \oc8051_gm_cxrom_1.cell3.data [6], _41967_);
  nand (_42012_, _42011_, _42010_);
  nand (_42013_, _42012_, _42003_);
  or (_42014_, \oc8051_gm_cxrom_1.cell3.data [6], _42003_);
  and (_01616_, _42014_, _42013_);
  or (_42015_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_42016_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_42017_, _42016_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_42018_, _42017_, _42015_);
  nand (_42019_, _42018_, _42003_);
  or (_42020_, \oc8051_gm_cxrom_1.cell4.data [7], _42003_);
  and (_01627_, _42020_, _42019_);
  or (_42021_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42022_, \oc8051_gm_cxrom_1.cell4.data [0], _42016_);
  nand (_42023_, _42022_, _42021_);
  nand (_42024_, _42023_, _42003_);
  or (_42025_, \oc8051_gm_cxrom_1.cell4.data [0], _42003_);
  and (_01634_, _42025_, _42024_);
  or (_42026_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42027_, \oc8051_gm_cxrom_1.cell4.data [1], _42016_);
  nand (_42028_, _42027_, _42026_);
  nand (_42029_, _42028_, _42003_);
  or (_42030_, \oc8051_gm_cxrom_1.cell4.data [1], _42003_);
  and (_01638_, _42030_, _42029_);
  or (_42031_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42032_, \oc8051_gm_cxrom_1.cell4.data [2], _42016_);
  nand (_42033_, _42032_, _42031_);
  nand (_42034_, _42033_, _42003_);
  or (_42035_, \oc8051_gm_cxrom_1.cell4.data [2], _42003_);
  and (_01642_, _42035_, _42034_);
  or (_42036_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42037_, \oc8051_gm_cxrom_1.cell4.data [3], _42016_);
  nand (_42038_, _42037_, _42036_);
  nand (_42039_, _42038_, _42003_);
  or (_42040_, \oc8051_gm_cxrom_1.cell4.data [3], _42003_);
  and (_01646_, _42040_, _42039_);
  or (_42041_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42042_, \oc8051_gm_cxrom_1.cell4.data [4], _42016_);
  nand (_42043_, _42042_, _42041_);
  nand (_42044_, _42043_, _42003_);
  or (_42045_, \oc8051_gm_cxrom_1.cell4.data [4], _42003_);
  and (_01650_, _42045_, _42044_);
  or (_42046_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42047_, \oc8051_gm_cxrom_1.cell4.data [5], _42016_);
  nand (_42048_, _42047_, _42046_);
  nand (_42049_, _42048_, _42003_);
  or (_42050_, \oc8051_gm_cxrom_1.cell4.data [5], _42003_);
  and (_01654_, _42050_, _42049_);
  or (_42051_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42052_, \oc8051_gm_cxrom_1.cell4.data [6], _42016_);
  nand (_42053_, _42052_, _42051_);
  nand (_42054_, _42053_, _42003_);
  or (_42055_, \oc8051_gm_cxrom_1.cell4.data [6], _42003_);
  and (_01658_, _42055_, _42054_);
  or (_42056_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_42057_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_42058_, _42057_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_42059_, _42058_, _42056_);
  nand (_42060_, _42059_, _42003_);
  or (_42061_, \oc8051_gm_cxrom_1.cell5.data [7], _42003_);
  and (_01680_, _42061_, _42060_);
  or (_42062_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42063_, \oc8051_gm_cxrom_1.cell5.data [0], _42057_);
  nand (_42064_, _42063_, _42062_);
  nand (_42065_, _42064_, _42003_);
  or (_42066_, \oc8051_gm_cxrom_1.cell5.data [0], _42003_);
  and (_01687_, _42066_, _42065_);
  or (_42067_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42068_, \oc8051_gm_cxrom_1.cell5.data [1], _42057_);
  nand (_42069_, _42068_, _42067_);
  nand (_42070_, _42069_, _42003_);
  or (_42071_, \oc8051_gm_cxrom_1.cell5.data [1], _42003_);
  and (_01691_, _42071_, _42070_);
  or (_42072_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42073_, \oc8051_gm_cxrom_1.cell5.data [2], _42057_);
  nand (_42074_, _42073_, _42072_);
  nand (_42075_, _42074_, _42003_);
  or (_42076_, \oc8051_gm_cxrom_1.cell5.data [2], _42003_);
  and (_01695_, _42076_, _42075_);
  or (_42077_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42078_, \oc8051_gm_cxrom_1.cell5.data [3], _42057_);
  nand (_42079_, _42078_, _42077_);
  nand (_42080_, _42079_, _42003_);
  or (_42081_, \oc8051_gm_cxrom_1.cell5.data [3], _42003_);
  and (_01699_, _42081_, _42080_);
  or (_42082_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42083_, \oc8051_gm_cxrom_1.cell5.data [4], _42057_);
  nand (_42084_, _42083_, _42082_);
  nand (_42085_, _42084_, _42003_);
  or (_42086_, \oc8051_gm_cxrom_1.cell5.data [4], _42003_);
  and (_01703_, _42086_, _42085_);
  or (_42087_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42088_, \oc8051_gm_cxrom_1.cell5.data [5], _42057_);
  nand (_42089_, _42088_, _42087_);
  nand (_42090_, _42089_, _42003_);
  or (_42091_, \oc8051_gm_cxrom_1.cell5.data [5], _42003_);
  and (_01707_, _42091_, _42090_);
  or (_42092_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42093_, \oc8051_gm_cxrom_1.cell5.data [6], _42057_);
  nand (_42094_, _42093_, _42092_);
  nand (_42095_, _42094_, _42003_);
  or (_42096_, \oc8051_gm_cxrom_1.cell5.data [6], _42003_);
  and (_01711_, _42096_, _42095_);
  or (_42097_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_42098_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_42099_, _42098_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_42100_, _42099_, _42097_);
  nand (_42101_, _42100_, _42003_);
  or (_42102_, \oc8051_gm_cxrom_1.cell6.data [7], _42003_);
  and (_01732_, _42102_, _42101_);
  or (_42103_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42104_, \oc8051_gm_cxrom_1.cell6.data [0], _42098_);
  nand (_42105_, _42104_, _42103_);
  nand (_42106_, _42105_, _42003_);
  or (_42107_, \oc8051_gm_cxrom_1.cell6.data [0], _42003_);
  and (_01739_, _42107_, _42106_);
  or (_42108_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42109_, \oc8051_gm_cxrom_1.cell6.data [1], _42098_);
  nand (_42110_, _42109_, _42108_);
  nand (_42111_, _42110_, _42003_);
  or (_42112_, \oc8051_gm_cxrom_1.cell6.data [1], _42003_);
  and (_01743_, _42112_, _42111_);
  or (_42113_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42114_, \oc8051_gm_cxrom_1.cell6.data [2], _42098_);
  nand (_42115_, _42114_, _42113_);
  nand (_42116_, _42115_, _42003_);
  or (_42117_, \oc8051_gm_cxrom_1.cell6.data [2], _42003_);
  and (_01747_, _42117_, _42116_);
  or (_42118_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42119_, \oc8051_gm_cxrom_1.cell6.data [3], _42098_);
  nand (_42120_, _42119_, _42118_);
  nand (_42121_, _42120_, _42003_);
  or (_42122_, \oc8051_gm_cxrom_1.cell6.data [3], _42003_);
  and (_01751_, _42122_, _42121_);
  or (_42123_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42124_, \oc8051_gm_cxrom_1.cell6.data [4], _42098_);
  nand (_42125_, _42124_, _42123_);
  nand (_42126_, _42125_, _42003_);
  or (_42127_, \oc8051_gm_cxrom_1.cell6.data [4], _42003_);
  and (_01755_, _42127_, _42126_);
  or (_42128_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42129_, \oc8051_gm_cxrom_1.cell6.data [5], _42098_);
  nand (_42130_, _42129_, _42128_);
  nand (_42131_, _42130_, _42003_);
  or (_42132_, \oc8051_gm_cxrom_1.cell6.data [5], _42003_);
  and (_01759_, _42132_, _42131_);
  or (_42133_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42134_, \oc8051_gm_cxrom_1.cell6.data [6], _42098_);
  nand (_42135_, _42134_, _42133_);
  nand (_42136_, _42135_, _42003_);
  or (_42137_, \oc8051_gm_cxrom_1.cell6.data [6], _42003_);
  and (_01763_, _42137_, _42136_);
  or (_42138_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_42139_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_42140_, _42139_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_42141_, _42140_, _42138_);
  nand (_42142_, _42141_, _42003_);
  or (_42143_, \oc8051_gm_cxrom_1.cell7.data [7], _42003_);
  and (_01784_, _42143_, _42142_);
  or (_42144_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42145_, \oc8051_gm_cxrom_1.cell7.data [0], _42139_);
  nand (_42146_, _42145_, _42144_);
  nand (_42147_, _42146_, _42003_);
  or (_42148_, \oc8051_gm_cxrom_1.cell7.data [0], _42003_);
  and (_01791_, _42148_, _42147_);
  or (_42149_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42150_, \oc8051_gm_cxrom_1.cell7.data [1], _42139_);
  nand (_42151_, _42150_, _42149_);
  nand (_42152_, _42151_, _42003_);
  or (_42153_, \oc8051_gm_cxrom_1.cell7.data [1], _42003_);
  and (_01795_, _42153_, _42152_);
  or (_42154_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42155_, \oc8051_gm_cxrom_1.cell7.data [2], _42139_);
  nand (_42156_, _42155_, _42154_);
  nand (_42157_, _42156_, _42003_);
  or (_42158_, \oc8051_gm_cxrom_1.cell7.data [2], _42003_);
  and (_01799_, _42158_, _42157_);
  or (_42159_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42160_, \oc8051_gm_cxrom_1.cell7.data [3], _42139_);
  nand (_42161_, _42160_, _42159_);
  nand (_42162_, _42161_, _42003_);
  or (_42163_, \oc8051_gm_cxrom_1.cell7.data [3], _42003_);
  and (_01802_, _42163_, _42162_);
  or (_42164_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42165_, \oc8051_gm_cxrom_1.cell7.data [4], _42139_);
  nand (_42166_, _42165_, _42164_);
  nand (_42167_, _42166_, _42003_);
  or (_42168_, \oc8051_gm_cxrom_1.cell7.data [4], _42003_);
  and (_01806_, _42168_, _42167_);
  or (_42169_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42170_, \oc8051_gm_cxrom_1.cell7.data [5], _42139_);
  nand (_42171_, _42170_, _42169_);
  nand (_42172_, _42171_, _42003_);
  or (_42173_, \oc8051_gm_cxrom_1.cell7.data [5], _42003_);
  and (_01810_, _42173_, _42172_);
  or (_42174_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42175_, \oc8051_gm_cxrom_1.cell7.data [6], _42139_);
  nand (_42176_, _42175_, _42174_);
  nand (_42177_, _42176_, _42003_);
  or (_42178_, \oc8051_gm_cxrom_1.cell7.data [6], _42003_);
  and (_01814_, _42178_, _42177_);
  or (_42179_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_42180_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_42181_, _42180_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_42182_, _42181_, _42179_);
  nand (_42183_, _42182_, _42003_);
  or (_42184_, \oc8051_gm_cxrom_1.cell8.data [7], _42003_);
  and (_01835_, _42184_, _42183_);
  or (_42185_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42186_, \oc8051_gm_cxrom_1.cell8.data [0], _42180_);
  nand (_42187_, _42186_, _42185_);
  nand (_42188_, _42187_, _42003_);
  or (_42189_, \oc8051_gm_cxrom_1.cell8.data [0], _42003_);
  and (_01842_, _42189_, _42188_);
  or (_42190_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42191_, \oc8051_gm_cxrom_1.cell8.data [1], _42180_);
  nand (_42192_, _42191_, _42190_);
  nand (_42193_, _42192_, _42003_);
  or (_42194_, \oc8051_gm_cxrom_1.cell8.data [1], _42003_);
  and (_01846_, _42194_, _42193_);
  or (_42195_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42196_, \oc8051_gm_cxrom_1.cell8.data [2], _42180_);
  nand (_42197_, _42196_, _42195_);
  nand (_42198_, _42197_, _42003_);
  or (_42199_, \oc8051_gm_cxrom_1.cell8.data [2], _42003_);
  and (_01850_, _42199_, _42198_);
  or (_42200_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42201_, \oc8051_gm_cxrom_1.cell8.data [3], _42180_);
  nand (_42202_, _42201_, _42200_);
  nand (_42203_, _42202_, _42003_);
  or (_42204_, \oc8051_gm_cxrom_1.cell8.data [3], _42003_);
  and (_01854_, _42204_, _42203_);
  or (_42205_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42206_, \oc8051_gm_cxrom_1.cell8.data [4], _42180_);
  nand (_42207_, _42206_, _42205_);
  nand (_42208_, _42207_, _42003_);
  or (_42209_, \oc8051_gm_cxrom_1.cell8.data [4], _42003_);
  and (_01858_, _42209_, _42208_);
  or (_42210_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42211_, \oc8051_gm_cxrom_1.cell8.data [5], _42180_);
  nand (_42212_, _42211_, _42210_);
  nand (_42213_, _42212_, _42003_);
  or (_42214_, \oc8051_gm_cxrom_1.cell8.data [5], _42003_);
  and (_01862_, _42214_, _42213_);
  or (_42215_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42216_, \oc8051_gm_cxrom_1.cell8.data [6], _42180_);
  nand (_42217_, _42216_, _42215_);
  nand (_42218_, _42217_, _42003_);
  or (_42219_, \oc8051_gm_cxrom_1.cell8.data [6], _42003_);
  and (_01866_, _42219_, _42218_);
  or (_42220_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_42221_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_42222_, _42221_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_42223_, _42222_, _42220_);
  nand (_42224_, _42223_, _42003_);
  or (_42225_, \oc8051_gm_cxrom_1.cell9.data [7], _42003_);
  and (_01888_, _42225_, _42224_);
  or (_42226_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42227_, \oc8051_gm_cxrom_1.cell9.data [0], _42221_);
  nand (_42228_, _42227_, _42226_);
  nand (_42229_, _42228_, _42003_);
  or (_42230_, \oc8051_gm_cxrom_1.cell9.data [0], _42003_);
  and (_01894_, _42230_, _42229_);
  or (_42231_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42232_, \oc8051_gm_cxrom_1.cell9.data [1], _42221_);
  nand (_42233_, _42232_, _42231_);
  nand (_42234_, _42233_, _42003_);
  or (_42235_, \oc8051_gm_cxrom_1.cell9.data [1], _42003_);
  and (_01898_, _42235_, _42234_);
  or (_42236_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42237_, \oc8051_gm_cxrom_1.cell9.data [2], _42221_);
  nand (_42238_, _42237_, _42236_);
  nand (_42239_, _42238_, _42003_);
  or (_42240_, \oc8051_gm_cxrom_1.cell9.data [2], _42003_);
  and (_01902_, _42240_, _42239_);
  or (_42241_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42242_, \oc8051_gm_cxrom_1.cell9.data [3], _42221_);
  nand (_42243_, _42242_, _42241_);
  nand (_42244_, _42243_, _42003_);
  or (_42245_, \oc8051_gm_cxrom_1.cell9.data [3], _42003_);
  and (_01906_, _42245_, _42244_);
  or (_42246_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42247_, \oc8051_gm_cxrom_1.cell9.data [4], _42221_);
  nand (_42248_, _42247_, _42246_);
  nand (_42249_, _42248_, _42003_);
  or (_42250_, \oc8051_gm_cxrom_1.cell9.data [4], _42003_);
  and (_01910_, _42250_, _42249_);
  or (_42251_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42252_, \oc8051_gm_cxrom_1.cell9.data [5], _42221_);
  nand (_42253_, _42252_, _42251_);
  nand (_42254_, _42253_, _42003_);
  or (_42255_, \oc8051_gm_cxrom_1.cell9.data [5], _42003_);
  and (_01914_, _42255_, _42254_);
  or (_42256_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42257_, \oc8051_gm_cxrom_1.cell9.data [6], _42221_);
  nand (_42258_, _42257_, _42256_);
  nand (_42259_, _42258_, _42003_);
  or (_42260_, \oc8051_gm_cxrom_1.cell9.data [6], _42003_);
  and (_01918_, _42260_, _42259_);
  or (_42261_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_42262_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_42263_, _42262_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_42264_, _42263_, _42261_);
  nand (_42265_, _42264_, _42003_);
  or (_42266_, \oc8051_gm_cxrom_1.cell10.data [7], _42003_);
  and (_01940_, _42266_, _42265_);
  or (_42267_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42268_, \oc8051_gm_cxrom_1.cell10.data [0], _42262_);
  nand (_42269_, _42268_, _42267_);
  nand (_42270_, _42269_, _42003_);
  or (_42271_, \oc8051_gm_cxrom_1.cell10.data [0], _42003_);
  and (_01946_, _42271_, _42270_);
  or (_42272_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42273_, \oc8051_gm_cxrom_1.cell10.data [1], _42262_);
  nand (_42274_, _42273_, _42272_);
  nand (_42275_, _42274_, _42003_);
  or (_42276_, \oc8051_gm_cxrom_1.cell10.data [1], _42003_);
  and (_01950_, _42276_, _42275_);
  or (_42277_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42278_, \oc8051_gm_cxrom_1.cell10.data [2], _42262_);
  nand (_42279_, _42278_, _42277_);
  nand (_42280_, _42279_, _42003_);
  or (_42281_, \oc8051_gm_cxrom_1.cell10.data [2], _42003_);
  and (_01954_, _42281_, _42280_);
  or (_42282_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42283_, \oc8051_gm_cxrom_1.cell10.data [3], _42262_);
  nand (_42284_, _42283_, _42282_);
  nand (_42285_, _42284_, _42003_);
  or (_42286_, \oc8051_gm_cxrom_1.cell10.data [3], _42003_);
  and (_01958_, _42286_, _42285_);
  or (_42287_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42288_, \oc8051_gm_cxrom_1.cell10.data [4], _42262_);
  nand (_42289_, _42288_, _42287_);
  nand (_42290_, _42289_, _42003_);
  or (_42291_, \oc8051_gm_cxrom_1.cell10.data [4], _42003_);
  and (_01962_, _42291_, _42290_);
  or (_42292_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42293_, \oc8051_gm_cxrom_1.cell10.data [5], _42262_);
  nand (_42294_, _42293_, _42292_);
  nand (_42295_, _42294_, _42003_);
  or (_42296_, \oc8051_gm_cxrom_1.cell10.data [5], _42003_);
  and (_01966_, _42296_, _42295_);
  or (_42297_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42298_, \oc8051_gm_cxrom_1.cell10.data [6], _42262_);
  nand (_42299_, _42298_, _42297_);
  nand (_42300_, _42299_, _42003_);
  or (_42301_, \oc8051_gm_cxrom_1.cell10.data [6], _42003_);
  and (_01970_, _42301_, _42300_);
  or (_42302_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_42303_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_42304_, _42303_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_42305_, _42304_, _42302_);
  nand (_42306_, _42305_, _42003_);
  or (_42307_, \oc8051_gm_cxrom_1.cell11.data [7], _42003_);
  and (_01992_, _42307_, _42306_);
  or (_42308_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42309_, \oc8051_gm_cxrom_1.cell11.data [0], _42303_);
  nand (_42310_, _42309_, _42308_);
  nand (_42311_, _42310_, _42003_);
  or (_42312_, \oc8051_gm_cxrom_1.cell11.data [0], _42003_);
  and (_01999_, _42312_, _42311_);
  or (_42313_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42314_, \oc8051_gm_cxrom_1.cell11.data [1], _42303_);
  nand (_42315_, _42314_, _42313_);
  nand (_42316_, _42315_, _42003_);
  or (_42317_, \oc8051_gm_cxrom_1.cell11.data [1], _42003_);
  and (_02002_, _42317_, _42316_);
  or (_42318_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42319_, \oc8051_gm_cxrom_1.cell11.data [2], _42303_);
  nand (_42320_, _42319_, _42318_);
  nand (_42321_, _42320_, _42003_);
  or (_42322_, \oc8051_gm_cxrom_1.cell11.data [2], _42003_);
  and (_02006_, _42322_, _42321_);
  or (_42323_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42324_, \oc8051_gm_cxrom_1.cell11.data [3], _42303_);
  nand (_42325_, _42324_, _42323_);
  nand (_42326_, _42325_, _42003_);
  or (_42327_, \oc8051_gm_cxrom_1.cell11.data [3], _42003_);
  and (_02010_, _42327_, _42326_);
  or (_42328_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42329_, \oc8051_gm_cxrom_1.cell11.data [4], _42303_);
  nand (_42330_, _42329_, _42328_);
  nand (_42331_, _42330_, _42003_);
  or (_42332_, \oc8051_gm_cxrom_1.cell11.data [4], _42003_);
  and (_02014_, _42332_, _42331_);
  or (_42333_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42334_, \oc8051_gm_cxrom_1.cell11.data [5], _42303_);
  nand (_42335_, _42334_, _42333_);
  nand (_42336_, _42335_, _42003_);
  or (_42337_, \oc8051_gm_cxrom_1.cell11.data [5], _42003_);
  and (_02018_, _42337_, _42336_);
  or (_42338_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42339_, \oc8051_gm_cxrom_1.cell11.data [6], _42303_);
  nand (_42340_, _42339_, _42338_);
  nand (_42341_, _42340_, _42003_);
  or (_42342_, \oc8051_gm_cxrom_1.cell11.data [6], _42003_);
  and (_02022_, _42342_, _42341_);
  or (_42343_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_42344_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_42345_, _42344_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_42346_, _42345_, _42343_);
  nand (_42347_, _42346_, _42003_);
  or (_42348_, \oc8051_gm_cxrom_1.cell12.data [7], _42003_);
  and (_02044_, _42348_, _42347_);
  or (_42349_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42350_, \oc8051_gm_cxrom_1.cell12.data [0], _42344_);
  nand (_42351_, _42350_, _42349_);
  nand (_42352_, _42351_, _42003_);
  or (_42353_, \oc8051_gm_cxrom_1.cell12.data [0], _42003_);
  and (_02051_, _42353_, _42352_);
  or (_42354_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42355_, \oc8051_gm_cxrom_1.cell12.data [1], _42344_);
  nand (_42356_, _42355_, _42354_);
  nand (_42357_, _42356_, _42003_);
  or (_42358_, \oc8051_gm_cxrom_1.cell12.data [1], _42003_);
  and (_02055_, _42358_, _42357_);
  or (_42359_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42360_, \oc8051_gm_cxrom_1.cell12.data [2], _42344_);
  nand (_42361_, _42360_, _42359_);
  nand (_42362_, _42361_, _42003_);
  or (_42363_, \oc8051_gm_cxrom_1.cell12.data [2], _42003_);
  and (_02058_, _42363_, _42362_);
  or (_42364_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42365_, \oc8051_gm_cxrom_1.cell12.data [3], _42344_);
  nand (_42366_, _42365_, _42364_);
  nand (_42367_, _42366_, _42003_);
  or (_42368_, \oc8051_gm_cxrom_1.cell12.data [3], _42003_);
  and (_02062_, _42368_, _42367_);
  or (_42369_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42370_, \oc8051_gm_cxrom_1.cell12.data [4], _42344_);
  nand (_42371_, _42370_, _42369_);
  nand (_42372_, _42371_, _42003_);
  or (_42373_, \oc8051_gm_cxrom_1.cell12.data [4], _42003_);
  and (_02066_, _42373_, _42372_);
  or (_42374_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42375_, \oc8051_gm_cxrom_1.cell12.data [5], _42344_);
  nand (_42376_, _42375_, _42374_);
  nand (_42377_, _42376_, _42003_);
  or (_42378_, \oc8051_gm_cxrom_1.cell12.data [5], _42003_);
  and (_02070_, _42378_, _42377_);
  or (_42379_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42380_, \oc8051_gm_cxrom_1.cell12.data [6], _42344_);
  nand (_42381_, _42380_, _42379_);
  nand (_42382_, _42381_, _42003_);
  or (_42383_, \oc8051_gm_cxrom_1.cell12.data [6], _42003_);
  and (_02074_, _42383_, _42382_);
  or (_42384_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_42385_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_42386_, _42385_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_42387_, _42386_, _42384_);
  nand (_42388_, _42387_, _42003_);
  or (_42389_, \oc8051_gm_cxrom_1.cell13.data [7], _42003_);
  and (_02096_, _42389_, _42388_);
  or (_42390_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42391_, \oc8051_gm_cxrom_1.cell13.data [0], _42385_);
  nand (_42392_, _42391_, _42390_);
  nand (_42393_, _42392_, _42003_);
  or (_42394_, \oc8051_gm_cxrom_1.cell13.data [0], _42003_);
  and (_02103_, _42394_, _42393_);
  or (_42395_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42396_, \oc8051_gm_cxrom_1.cell13.data [1], _42385_);
  nand (_42397_, _42396_, _42395_);
  nand (_42398_, _42397_, _42003_);
  or (_42399_, \oc8051_gm_cxrom_1.cell13.data [1], _42003_);
  and (_02107_, _42399_, _42398_);
  or (_42400_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42401_, \oc8051_gm_cxrom_1.cell13.data [2], _42385_);
  nand (_42402_, _42401_, _42400_);
  nand (_42403_, _42402_, _42003_);
  or (_42404_, \oc8051_gm_cxrom_1.cell13.data [2], _42003_);
  and (_02111_, _42404_, _42403_);
  or (_42405_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42406_, \oc8051_gm_cxrom_1.cell13.data [3], _42385_);
  nand (_42407_, _42406_, _42405_);
  nand (_42408_, _42407_, _42003_);
  or (_42409_, \oc8051_gm_cxrom_1.cell13.data [3], _42003_);
  and (_02114_, _42409_, _42408_);
  or (_42410_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42411_, \oc8051_gm_cxrom_1.cell13.data [4], _42385_);
  nand (_42412_, _42411_, _42410_);
  nand (_42413_, _42412_, _42003_);
  or (_42414_, \oc8051_gm_cxrom_1.cell13.data [4], _42003_);
  and (_02118_, _42414_, _42413_);
  or (_42415_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42416_, \oc8051_gm_cxrom_1.cell13.data [5], _42385_);
  nand (_42417_, _42416_, _42415_);
  nand (_42418_, _42417_, _42003_);
  or (_42419_, \oc8051_gm_cxrom_1.cell13.data [5], _42003_);
  and (_02122_, _42419_, _42418_);
  or (_42420_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42421_, \oc8051_gm_cxrom_1.cell13.data [6], _42385_);
  nand (_42422_, _42421_, _42420_);
  nand (_42423_, _42422_, _42003_);
  or (_42424_, \oc8051_gm_cxrom_1.cell13.data [6], _42003_);
  and (_02126_, _42424_, _42423_);
  or (_42425_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_42426_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_42427_, _42426_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_42428_, _42427_, _42425_);
  nand (_42429_, _42428_, _42003_);
  or (_42430_, \oc8051_gm_cxrom_1.cell14.data [7], _42003_);
  and (_02148_, _42430_, _42429_);
  or (_42431_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42432_, \oc8051_gm_cxrom_1.cell14.data [0], _42426_);
  nand (_42433_, _42432_, _42431_);
  nand (_42434_, _42433_, _42003_);
  or (_42435_, \oc8051_gm_cxrom_1.cell14.data [0], _42003_);
  and (_02155_, _42435_, _42434_);
  or (_42436_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42437_, \oc8051_gm_cxrom_1.cell14.data [1], _42426_);
  nand (_42438_, _42437_, _42436_);
  nand (_42439_, _42438_, _42003_);
  or (_42440_, \oc8051_gm_cxrom_1.cell14.data [1], _42003_);
  and (_02159_, _42440_, _42439_);
  or (_42441_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42442_, \oc8051_gm_cxrom_1.cell14.data [2], _42426_);
  nand (_42443_, _42442_, _42441_);
  nand (_42444_, _42443_, _42003_);
  or (_42445_, \oc8051_gm_cxrom_1.cell14.data [2], _42003_);
  and (_02163_, _42445_, _42444_);
  or (_42446_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42447_, \oc8051_gm_cxrom_1.cell14.data [3], _42426_);
  nand (_42448_, _42447_, _42446_);
  nand (_42449_, _42448_, _42003_);
  or (_42450_, \oc8051_gm_cxrom_1.cell14.data [3], _42003_);
  and (_02167_, _42450_, _42449_);
  or (_42451_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42452_, \oc8051_gm_cxrom_1.cell14.data [4], _42426_);
  nand (_42453_, _42452_, _42451_);
  nand (_42454_, _42453_, _42003_);
  or (_42455_, \oc8051_gm_cxrom_1.cell14.data [4], _42003_);
  and (_02170_, _42455_, _42454_);
  or (_42456_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42457_, \oc8051_gm_cxrom_1.cell14.data [5], _42426_);
  nand (_42458_, _42457_, _42456_);
  nand (_42459_, _42458_, _42003_);
  or (_42460_, \oc8051_gm_cxrom_1.cell14.data [5], _42003_);
  and (_02174_, _42460_, _42459_);
  or (_42461_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42462_, \oc8051_gm_cxrom_1.cell14.data [6], _42426_);
  nand (_42463_, _42462_, _42461_);
  nand (_42464_, _42463_, _42003_);
  or (_42465_, \oc8051_gm_cxrom_1.cell14.data [6], _42003_);
  and (_02178_, _42465_, _42464_);
  or (_42466_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_42467_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_42468_, _42467_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_42469_, _42468_, _42466_);
  nand (_42470_, _42469_, _42003_);
  or (_42471_, \oc8051_gm_cxrom_1.cell15.data [7], _42003_);
  and (_02200_, _42471_, _42470_);
  or (_42472_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42473_, \oc8051_gm_cxrom_1.cell15.data [0], _42467_);
  nand (_42474_, _42473_, _42472_);
  nand (_42475_, _42474_, _42003_);
  or (_42476_, \oc8051_gm_cxrom_1.cell15.data [0], _42003_);
  and (_02207_, _42476_, _42475_);
  or (_42477_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42478_, \oc8051_gm_cxrom_1.cell15.data [1], _42467_);
  nand (_42479_, _42478_, _42477_);
  nand (_42480_, _42479_, _42003_);
  or (_42481_, \oc8051_gm_cxrom_1.cell15.data [1], _42003_);
  and (_02211_, _42481_, _42480_);
  or (_42482_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42483_, \oc8051_gm_cxrom_1.cell15.data [2], _42467_);
  nand (_42484_, _42483_, _42482_);
  nand (_42485_, _42484_, _42003_);
  or (_42486_, \oc8051_gm_cxrom_1.cell15.data [2], _42003_);
  and (_02215_, _42486_, _42485_);
  or (_42487_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42488_, \oc8051_gm_cxrom_1.cell15.data [3], _42467_);
  nand (_42489_, _42488_, _42487_);
  nand (_42490_, _42489_, _42003_);
  or (_42491_, \oc8051_gm_cxrom_1.cell15.data [3], _42003_);
  and (_02219_, _42491_, _42490_);
  or (_42492_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42493_, \oc8051_gm_cxrom_1.cell15.data [4], _42467_);
  nand (_42494_, _42493_, _42492_);
  nand (_42495_, _42494_, _42003_);
  or (_42496_, \oc8051_gm_cxrom_1.cell15.data [4], _42003_);
  and (_02223_, _42496_, _42495_);
  or (_42497_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42498_, \oc8051_gm_cxrom_1.cell15.data [5], _42467_);
  nand (_42499_, _42498_, _42497_);
  nand (_42500_, _42499_, _42003_);
  or (_42501_, \oc8051_gm_cxrom_1.cell15.data [5], _42003_);
  and (_02226_, _42501_, _42500_);
  or (_42502_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42503_, \oc8051_gm_cxrom_1.cell15.data [6], _42467_);
  nand (_42504_, _42503_, _42502_);
  nand (_42505_, _42504_, _42003_);
  or (_42506_, \oc8051_gm_cxrom_1.cell15.data [6], _42003_);
  and (_02230_, _42506_, _42505_);
  nor (_06004_, _38068_, rst);
  and (_42507_, _33939_, _42003_);
  nand (_42508_, _42507_, _36707_);
  nor (_42509_, _36652_, _36389_);
  or (_06007_, _42509_, _42508_);
  not (_42510_, _34312_);
  and (_42511_, _34806_, _42510_);
  and (_42512_, _42511_, _34565_);
  not (_42513_, _36313_);
  and (_42514_, _35322_, _35091_);
  and (_42515_, _42514_, _35578_);
  and (_42516_, _42515_, _42513_);
  and (_42517_, _42516_, _42512_);
  not (_42518_, _34565_);
  and (_42519_, _34806_, _34312_);
  and (_42520_, _42519_, _42518_);
  and (_42521_, _42515_, _36313_);
  and (_42522_, _42521_, _42520_);
  or (_42523_, _42522_, _42517_);
  not (_42524_, _35830_);
  and (_42525_, _42524_, _34565_);
  nor (_42526_, _42524_, _34565_);
  nor (_42527_, _42526_, _42525_);
  and (_42528_, _35578_, _35322_);
  not (_42529_, _35091_);
  and (_42530_, _36313_, _42529_);
  and (_42531_, _42530_, _42528_);
  and (_42532_, _42531_, _42519_);
  and (_42533_, _42532_, _42527_);
  not (_42534_, _34806_);
  and (_42535_, _42534_, _34312_);
  and (_42536_, _42531_, _35830_);
  and (_42537_, _42536_, _42535_);
  or (_42538_, _42537_, _42533_);
  or (_42539_, _42538_, _42523_);
  and (_42540_, _42535_, _42526_);
  and (_42541_, _42540_, _42516_);
  and (_42542_, _35830_, _34565_);
  nor (_42543_, _34806_, _34312_);
  and (_42544_, _42543_, _42542_);
  not (_42545_, _35578_);
  nor (_42546_, _42545_, _35322_);
  and (_42547_, _42546_, _42529_);
  and (_42548_, _42547_, _42513_);
  and (_42549_, _42548_, _42544_);
  or (_42550_, _42549_, _42541_);
  and (_42551_, _42544_, _42545_);
  and (_42552_, _35830_, _35578_);
  and (_42553_, _42543_, _42518_);
  and (_42554_, _42553_, _42514_);
  and (_42555_, _42554_, _42552_);
  or (_42556_, _42555_, _42551_);
  or (_42557_, _42556_, _42550_);
  and (_42558_, _42546_, _42530_);
  and (_42559_, _42511_, _42524_);
  and (_42560_, _42559_, _42558_);
  and (_42561_, _42553_, _42531_);
  or (_42562_, _42561_, _42560_);
  and (_42563_, _42525_, _42511_);
  and (_42564_, _42531_, _42563_);
  and (_42565_, _42519_, _34565_);
  and (_42566_, _42565_, _42521_);
  or (_42567_, _42566_, _42564_);
  or (_42568_, _42567_, _42562_);
  or (_42569_, _42568_, _42557_);
  nor (_42570_, _35830_, _34565_);
  and (_42571_, _42535_, _42570_);
  nor (_42572_, _42571_, _42513_);
  and (_42573_, _42528_, _42529_);
  not (_42574_, _42573_);
  nor (_42575_, _42574_, _42572_);
  not (_42576_, _42575_);
  and (_42577_, _42526_, _42519_);
  and (_42578_, _42531_, _42577_);
  and (_42579_, _42535_, _42525_);
  and (_42580_, _42579_, _42531_);
  nor (_42581_, _42580_, _42578_);
  and (_42582_, _42581_, _42576_);
  and (_42583_, _42526_, _42511_);
  and (_42584_, _42583_, _42547_);
  nor (_42585_, _35322_, _42529_);
  nor (_42586_, _42585_, _42545_);
  not (_42587_, _42586_);
  and (_42588_, _42587_, _42583_);
  and (_42589_, _42543_, _42570_);
  and (_42590_, _42589_, _42515_);
  or (_42591_, _42590_, _42588_);
  nor (_42592_, _42591_, _42584_);
  nand (_42593_, _42592_, _42582_);
  or (_42594_, _42593_, _42569_);
  or (_42595_, _42594_, _42539_);
  and (_42596_, _42595_, _33950_);
  not (_42597_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42598_, _33929_, _15704_);
  and (_42599_, _42598_, _36817_);
  nor (_42600_, _42599_, _42597_);
  or (_42601_, _42600_, rst);
  or (_06010_, _42601_, _42596_);
  nand (_42602_, _34312_, _33885_);
  or (_42603_, _33885_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42604_, _42603_, _42003_);
  and (_06013_, _42604_, _42602_);
  and (_42605_, \oc8051_top_1.oc8051_sfr1.wait_data , _42003_);
  and (_42606_, _42605_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42607_, _36532_, _36093_);
  and (_42608_, _37936_, _37025_);
  or (_42609_, _42608_, _42607_);
  and (_42610_, _36652_, _36093_);
  or (_42611_, _42610_, _37760_);
  or (_42612_, _42611_, _37430_);
  and (_42613_, _37201_, _36532_);
  and (_42614_, _36663_, _36389_);
  or (_42615_, _42614_, _42613_);
  or (_42616_, _42615_, _42612_);
  or (_42617_, _42616_, _37650_);
  or (_42618_, _42617_, _42609_);
  and (_42619_, _42618_, _42507_);
  or (_06016_, _42619_, _42606_);
  and (_42620_, _36652_, _36455_);
  or (_42621_, _42620_, _36554_);
  and (_42622_, _37113_, _36433_);
  or (_42623_, _42622_, _36444_);
  and (_42624_, _36970_, _35135_);
  and (_42625_, _42624_, _37201_);
  or (_42626_, _42625_, _42623_);
  or (_42627_, _42626_, _42621_);
  and (_42628_, _42627_, _33939_);
  and (_42629_, \oc8051_top_1.oc8051_decoder1.state [0], _15704_);
  and (_42630_, _42629_, _42597_);
  not (_42631_, _37969_);
  and (_42632_, _42631_, _42630_);
  and (_42633_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42634_, _42633_, _42632_);
  or (_42635_, _42634_, _42628_);
  and (_06019_, _42635_, _42003_);
  and (_42636_, _42605_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_42637_, _37936_, _37135_);
  not (_42638_, _36992_);
  nor (_42639_, _37135_, _36663_);
  nor (_42640_, _42639_, _42638_);
  or (_42641_, _42640_, _42637_);
  and (_42642_, _42624_, _37310_);
  or (_42643_, _42642_, _42641_);
  nor (_42644_, _42639_, _35622_);
  not (_42645_, _35622_);
  and (_42646_, _37310_, _42645_);
  or (_42647_, _42646_, _42644_);
  or (_42648_, _42647_, _36071_);
  nor (_42649_, _35874_, _35622_);
  and (_42650_, _42649_, _36038_);
  and (_42651_, _37936_, _37003_);
  or (_42652_, _42651_, _42650_);
  or (_42653_, _42652_, _42621_);
  or (_42654_, _42653_, _42648_);
  or (_42655_, _42654_, _42643_);
  and (_42656_, _42655_, _42507_);
  or (_06022_, _42656_, _42636_);
  and (_42657_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42658_, _37485_, _33939_);
  or (_42659_, _42658_, _42657_);
  or (_42660_, _42659_, _42632_);
  and (_06025_, _42660_, _42003_);
  and (_42661_, _36532_, _36082_);
  not (_42662_, _37025_);
  nor (_42663_, _42509_, _42662_);
  nor (_42664_, _42663_, _42661_);
  not (_42665_, _42664_);
  and (_42666_, _42665_, _42630_);
  or (_42667_, _42666_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42668_, _37310_, _36400_);
  and (_42669_, _36981_, _36378_);
  and (_42670_, _42669_, _35885_);
  or (_42671_, _42670_, _42668_);
  or (_42672_, _42671_, _42607_);
  and (_42673_, _42671_, _36839_);
  or (_42674_, _42673_, _36949_);
  and (_42675_, _42674_, _42672_);
  or (_42676_, _42675_, _42667_);
  or (_42677_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15704_);
  and (_42678_, _42677_, _42003_);
  and (_06028_, _42678_, _42676_);
  and (_42679_, _42605_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_42680_, _36663_, _42645_);
  nor (_42681_, _42680_, _37353_);
  nor (_42682_, _42646_, _36554_);
  nand (_42683_, _42682_, _42681_);
  and (_42684_, _36400_, _36038_);
  or (_42685_, _42642_, _42614_);
  or (_42686_, _42685_, _42684_);
  or (_42687_, _42622_, _37212_);
  or (_42688_, _37310_, _37201_);
  and (_42689_, _42688_, _35929_);
  or (_42690_, _42689_, _42687_);
  or (_42691_, _42690_, _42686_);
  or (_42692_, _42691_, _42683_);
  and (_42693_, _42692_, _42507_);
  or (_06031_, _42693_, _42679_);
  and (_42694_, _42605_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_42695_, _42625_, _37323_);
  and (_42696_, _36532_, _35940_);
  and (_42697_, _42624_, _36740_);
  or (_42698_, _42697_, _42696_);
  or (_42699_, _42698_, _42695_);
  or (_42700_, _42699_, _42647_);
  and (_42701_, _37936_, _37294_);
  or (_42702_, _37342_, _37302_);
  or (_42703_, _42702_, _42701_);
  and (_42704_, _36696_, _34861_);
  or (_42705_, _42704_, _36751_);
  and (_42706_, _36663_, _35929_);
  or (_42707_, _42706_, _42705_);
  or (_42708_, _42707_, _42703_);
  or (_42709_, _42708_, _42700_);
  nor (_42710_, _37518_, _36006_);
  not (_42711_, _42710_);
  not (_42712_, _37408_);
  and (_42713_, _37113_, _34861_);
  and (_42714_, _37113_, _36587_);
  or (_42715_, _42714_, _42713_);
  or (_42716_, _42715_, _42712_);
  or (_42717_, _42716_, _42711_);
  or (_42718_, _42717_, _42643_);
  or (_42719_, _42718_, _42709_);
  and (_42720_, _42719_, _42507_);
  or (_06034_, _42720_, _42694_);
  and (_42721_, _36082_, _35907_);
  and (_42722_, _42624_, _35951_);
  or (_42723_, _42722_, _42721_);
  and (_42724_, _42649_, _36082_);
  or (_42725_, _42724_, _35962_);
  and (_42726_, _35951_, _42645_);
  or (_42727_, _42726_, _42725_);
  or (_42728_, _42727_, _42723_);
  and (_42729_, _36992_, _36455_);
  and (_42730_, _37936_, _36455_);
  or (_42731_, _42730_, _42729_);
  or (_42732_, _42731_, _42728_);
  and (_42733_, _42732_, _33939_);
  and (_42734_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42735_, _42734_, _38035_);
  or (_42736_, _42735_, _42733_);
  and (_06037_, _42736_, _42003_);
  or (_42737_, _37245_, _37212_);
  not (_42738_, _37441_);
  or (_42739_, _42640_, _42738_);
  or (_42740_, _42739_, _42737_);
  and (_42741_, _36576_, _35885_);
  and (_42742_, _42741_, _36992_);
  or (_42743_, _42742_, _37317_);
  or (_42744_, _42743_, _37302_);
  or (_42745_, _42744_, _42668_);
  or (_42746_, _42745_, _37540_);
  or (_42747_, _42746_, _42740_);
  and (_42748_, _37113_, _36082_);
  or (_42749_, _42748_, _42670_);
  and (_42750_, _42649_, _36576_);
  or (_42751_, _42750_, _37124_);
  or (_42752_, _42751_, _42623_);
  or (_42753_, _42752_, _42749_);
  and (_42754_, _42741_, _35929_);
  or (_42755_, _42754_, _36006_);
  or (_42756_, _42755_, _37047_);
  or (_42757_, _37562_, _36104_);
  or (_42758_, _42757_, _42756_);
  or (_42759_, _42758_, _42753_);
  or (_42760_, _42759_, _42647_);
  or (_42761_, _42760_, _42747_);
  and (_42762_, _42761_, _33939_);
  or (_42763_, _42673_, _42632_);
  and (_42764_, _37815_, _36839_);
  or (_42765_, _42764_, _42763_);
  and (_42766_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42767_, _42766_, _42765_);
  or (_42768_, _42767_, _42762_);
  and (_06040_, _42768_, _42003_);
  nor (_06099_, _36905_, rst);
  nor (_06101_, _37881_, rst);
  not (_42769_, _42507_);
  or (_06104_, _42664_, _42769_);
  and (_42770_, _36707_, _36652_);
  nor (_42771_, _42770_, _42661_);
  or (_06107_, _42771_, _42769_);
  or (_42772_, _42560_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42773_, _42772_, _42523_);
  and (_42774_, _42773_, _42599_);
  nor (_42775_, _42598_, _36817_);
  or (_42776_, _42775_, rst);
  or (_06110_, _42776_, _42774_);
  nand (_42777_, _36313_, _33885_);
  or (_42778_, _33885_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42779_, _42778_, _42003_);
  and (_06113_, _42779_, _42777_);
  or (_42780_, _35091_, _38002_);
  or (_42781_, _33885_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42782_, _42781_, _42003_);
  and (_06116_, _42782_, _42780_);
  nand (_42783_, _35322_, _33885_);
  or (_42784_, _33885_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42785_, _42784_, _42003_);
  and (_06119_, _42785_, _42783_);
  nand (_42786_, _35578_, _33885_);
  or (_42787_, _33885_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42788_, _42787_, _42003_);
  and (_06122_, _42788_, _42786_);
  or (_42789_, _35830_, _38002_);
  or (_42790_, _33885_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42791_, _42790_, _42003_);
  and (_06125_, _42791_, _42789_);
  nand (_42792_, _34565_, _33885_);
  or (_42793_, _33885_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42794_, _42793_, _42003_);
  and (_06128_, _42794_, _42792_);
  nand (_42795_, _34806_, _33885_);
  or (_42796_, _33885_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42797_, _42796_, _42003_);
  and (_06131_, _42797_, _42795_);
  or (_42798_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _15704_);
  and (_42799_, _42798_, _42667_);
  and (_42800_, _42715_, _34356_);
  and (_42801_, _36707_, _35885_);
  and (_42802_, _42801_, _37936_);
  and (_42803_, _37113_, _36707_);
  and (_42804_, _42624_, _37080_);
  or (_42805_, _42804_, _42803_);
  or (_42806_, _42805_, _42802_);
  or (_42807_, _42725_, _42697_);
  and (_42808_, _37936_, _36598_);
  or (_42809_, _42808_, _35918_);
  or (_42810_, _42809_, _42807_);
  or (_42811_, _42810_, _42806_);
  or (_42812_, _42811_, _42800_);
  and (_42813_, _42624_, _37294_);
  or (_42814_, _42813_, _42620_);
  and (_42815_, _37091_, _42645_);
  or (_42816_, _42815_, _42814_);
  and (_42817_, _37936_, _37310_);
  and (_42818_, _37936_, _36663_);
  or (_42819_, _42818_, _42817_);
  or (_42820_, _42819_, _42637_);
  or (_42821_, _42820_, _42816_);
  or (_42822_, _37036_, _36751_);
  or (_42823_, _42696_, _42608_);
  or (_42824_, _42823_, _42822_);
  and (_42825_, _42624_, _36455_);
  or (_42826_, _42722_, _36466_);
  or (_42827_, _42826_, _42825_);
  or (_42828_, _36729_, _36554_);
  or (_42829_, _42828_, _42827_);
  or (_42830_, _42829_, _42824_);
  or (_42831_, _42830_, _42821_);
  or (_42832_, _42831_, _42812_);
  and (_42833_, _42832_, _33939_);
  or (_42834_, _42833_, _42799_);
  and (_30470_, _42834_, _42003_);
  and (_42835_, _42605_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_42836_, _37294_, _36740_);
  and (_42837_, _42836_, _36400_);
  or (_42838_, _42814_, _42715_);
  or (_42839_, _42838_, _42837_);
  nor (_42840_, _42650_, _36049_);
  not (_42841_, _42840_);
  or (_42842_, _42841_, _42651_);
  or (_42843_, _42842_, _37223_);
  or (_42844_, _42843_, _42609_);
  or (_42845_, _36740_, _37091_);
  and (_42846_, _42845_, _37936_);
  or (_42847_, _42846_, _42707_);
  or (_42848_, _42847_, _42844_);
  or (_42849_, _42848_, _42839_);
  and (_42850_, _42849_, _42507_);
  or (_30473_, _42850_, _42835_);
  or (_42851_, _42757_, _42749_);
  or (_42852_, _42851_, _42747_);
  and (_42853_, _42852_, _33939_);
  and (_42854_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42855_, _42854_, _42765_);
  or (_42856_, _42855_, _42853_);
  and (_30475_, _42856_, _42003_);
  and (_42857_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42858_, _37507_, _35874_);
  or (_42859_, _42858_, _36444_);
  or (_42860_, _42859_, _42756_);
  or (_42861_, _42860_, _42671_);
  and (_42862_, _42861_, _33939_);
  or (_42863_, _42862_, _42857_);
  or (_42864_, _42863_, _42763_);
  and (_30477_, _42864_, _42003_);
  or (_42865_, _42666_, _38046_);
  or (_42866_, _42836_, _36598_);
  and (_42867_, _42866_, _37936_);
  or (_42868_, _42724_, _35973_);
  or (_42869_, _42815_, _42696_);
  or (_42870_, _42869_, _42868_);
  or (_42871_, _42870_, _42867_);
  and (_42872_, _37936_, _37201_);
  or (_42873_, _42731_, _42872_);
  or (_42874_, _42802_, _37947_);
  and (_42875_, _42624_, _37322_);
  or (_42876_, _42875_, _42608_);
  or (_42877_, _42876_, _42874_);
  or (_42878_, _42877_, _42820_);
  or (_42879_, _42878_, _42873_);
  and (_42880_, _42722_, _35874_);
  or (_42881_, _42880_, _36609_);
  or (_42882_, _42750_, _36466_);
  or (_42883_, _42882_, _42754_);
  and (_42884_, _36400_, _37080_);
  and (_42885_, _42801_, _36992_);
  or (_42886_, _42885_, _42884_);
  or (_42887_, _42886_, _42883_);
  or (_42888_, _42887_, _42881_);
  or (_42889_, _42661_, _37958_);
  and (_42890_, _42722_, _35885_);
  or (_42891_, _42890_, _42804_);
  or (_42892_, _42891_, _42889_);
  or (_42893_, _42892_, _42671_);
  or (_42894_, _42893_, _42888_);
  or (_42895_, _42894_, _42879_);
  or (_42896_, _42895_, _42871_);
  and (_42897_, _42896_, _33939_);
  or (_42898_, _42897_, _42865_);
  and (_42899_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42900_, _42899_, _42898_);
  and (_30479_, _42900_, _42003_);
  and (_42901_, _42801_, _35929_);
  or (_42902_, _37958_, _36466_);
  or (_42903_, _42902_, _37562_);
  or (_42904_, _42903_, _42901_);
  and (_42905_, _42649_, _36707_);
  or (_42906_, _42742_, _42620_);
  or (_42907_, _42906_, _42905_);
  or (_42908_, _42907_, _36620_);
  or (_42909_, _42908_, _42904_);
  or (_42910_, _42909_, _42870_);
  and (_42911_, _37518_, _36521_);
  and (_42912_, _37302_, _36521_);
  or (_42913_, _42912_, _37102_);
  or (_42914_, _42913_, _42911_);
  or (_42915_, _42914_, _42879_);
  or (_42916_, _42915_, _42910_);
  and (_42917_, _42916_, _33939_);
  or (_42918_, _42917_, _42865_);
  and (_42919_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42920_, _42919_, _42918_);
  and (_30481_, _42920_, _42003_);
  and (_42921_, _42605_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_42922_, _40504_);
  or (_42923_, _42825_, _42922_);
  and (_42924_, _36532_, _35995_);
  and (_42925_, _42924_, _35885_);
  and (_42926_, _42614_, _36521_);
  or (_42927_, _42926_, _42925_);
  or (_42929_, _42927_, _42683_);
  or (_42931_, _42929_, _42923_);
  not (_42933_, _40503_);
  or (_42935_, _42689_, _42933_);
  or (_42937_, _42818_, _42642_);
  or (_42939_, _42937_, _42737_);
  or (_42941_, _42939_, _42935_);
  and (_42943_, _36532_, _37322_);
  or (_42945_, _42724_, _42622_);
  and (_42947_, _35962_, _35885_);
  or (_42949_, _42947_, _42945_);
  or (_42951_, _42949_, _42943_);
  and (_42953_, _37606_, _42645_);
  or (_42955_, _42953_, _36466_);
  or (_42957_, _42955_, _37474_);
  and (_42959_, _37606_, _36532_);
  or (_42961_, _42890_, _42959_);
  or (_42963_, _42961_, _42957_);
  or (_42965_, _42963_, _42951_);
  or (_42967_, _42965_, _42941_);
  or (_42969_, _42967_, _42931_);
  and (_42971_, _42969_, _42507_);
  or (_30483_, _42971_, _42921_);
  or (_42974_, _42625_, _37397_);
  or (_42976_, _42706_, _42704_);
  or (_42978_, _42976_, _42974_);
  or (_42980_, _42978_, _42703_);
  or (_42982_, _42980_, _42892_);
  or (_42984_, _42818_, _42959_);
  or (_42986_, _42925_, _42881_);
  or (_42988_, _42986_, _42984_);
  or (_42989_, _42713_, _36554_);
  or (_42990_, _42989_, _35973_);
  or (_42991_, _42815_, _37573_);
  or (_42992_, _42991_, _42990_);
  or (_42993_, _42992_, _42988_);
  or (_42994_, _42993_, _42982_);
  and (_42995_, _42994_, _42507_);
  and (_42996_, _33896_, _42003_);
  and (_42997_, _42996_, _37958_);
  and (_42998_, _42605_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_42999_, _42998_, _42997_);
  or (_30485_, _42999_, _42995_);
  or (_43000_, _42875_, _42825_);
  or (_43001_, _43000_, _42608_);
  nor (_43002_, _42650_, _37386_);
  nand (_43003_, _43002_, _36477_);
  or (_43004_, _43003_, _43001_);
  and (_43005_, _36389_, _37322_);
  or (_43006_, _43005_, _42802_);
  and (_43007_, _42649_, _34872_);
  or (_43008_, _43007_, _35918_);
  or (_43009_, _43008_, _43006_);
  or (_43010_, _43009_, _43004_);
  nor (_43011_, _42804_, _37562_);
  not (_43012_, _43011_);
  nor (_43013_, _43012_, _37551_);
  and (_43014_, _36532_, _35951_);
  or (_43015_, _42945_, _42625_);
  nor (_43016_, _43015_, _43014_);
  nand (_43017_, _43016_, _43013_);
  or (_43018_, _43017_, _43010_);
  or (_43019_, _42648_, _42643_);
  or (_43020_, _43019_, _43018_);
  and (_43021_, _43020_, _33939_);
  and (_43022_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_43023_, _43022_, _38013_);
  or (_43024_, _43023_, _43021_);
  and (_30487_, _43024_, _42003_);
  or (_43025_, _43012_, _43006_);
  or (_43026_, _43025_, _43008_);
  or (_43027_, _36444_, _36006_);
  nor (_43028_, _43027_, _42924_);
  nand (_43029_, _43028_, _40504_);
  or (_43030_, _42937_, _42687_);
  or (_43031_, _43030_, _43029_);
  or (_43032_, _42647_, _42641_);
  or (_43033_, _43032_, _43031_);
  or (_43034_, _43033_, _43026_);
  and (_43035_, _43034_, _33939_);
  and (_43036_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_43037_, _43036_, _38024_);
  or (_43038_, _43037_, _43035_);
  and (_30489_, _43038_, _42003_);
  and (_43039_, _42605_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_43040_, _36378_);
  and (_43041_, _43040_, _37322_);
  or (_43042_, _43041_, _37234_);
  or (_43043_, _42943_, _42613_);
  or (_43044_, _43043_, _43042_);
  or (_43045_, _42984_, _42933_);
  or (_43046_, _43045_, _43044_);
  or (_43047_, _42927_, _42728_);
  or (_43048_, _43047_, _42923_);
  or (_43049_, _43048_, _43046_);
  and (_43050_, _43049_, _42507_);
  or (_30491_, _43050_, _43039_);
  nor (_39013_, _34312_, rst);
  nor (_39015_, _40496_, rst);
  and (_43051_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_43052_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_43053_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43054_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_43055_, _43054_, _43053_);
  and (_43056_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_43057_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_43058_, _43057_, _43056_);
  and (_43059_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_43060_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_43061_, _43060_, _43059_);
  and (_43062_, _43061_, _43058_);
  and (_43064_, _43062_, _43055_);
  nor (_43065_, _43064_, _33994_);
  nor (_43066_, _43065_, _43052_);
  nor (_43067_, _43066_, _40480_);
  nor (_43068_, _43067_, _43051_);
  nor (_39016_, _43068_, rst);
  nor (_39025_, _36313_, rst);
  and (_39026_, _35091_, _42003_);
  nor (_39027_, _35322_, rst);
  nor (_39028_, _35578_, rst);
  and (_39029_, _35830_, _42003_);
  nor (_39030_, _34565_, rst);
  nor (_39031_, _34806_, rst);
  nor (_39032_, _40583_, rst);
  nor (_39034_, _40739_, rst);
  nor (_39035_, _40656_, rst);
  nor (_39036_, _40534_, rst);
  nor (_39037_, _40717_, rst);
  nor (_39038_, _40635_, rst);
  nor (_39040_, _40832_, rst);
  and (_43070_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_43071_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_43072_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_43073_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_43074_, _43073_, _43072_);
  and (_43075_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_43076_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_43077_, _43076_, _43075_);
  and (_43078_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_43079_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_43080_, _43079_, _43078_);
  and (_43081_, _43080_, _43077_);
  and (_43082_, _43081_, _43074_);
  nor (_43083_, _43082_, _33994_);
  nor (_43084_, _43083_, _43071_);
  nor (_43085_, _43084_, _40480_);
  nor (_43086_, _43085_, _43070_);
  nor (_39041_, _43086_, rst);
  and (_43087_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_43088_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_43089_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_43090_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_43091_, _43090_, _43089_);
  and (_43092_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_43093_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_43094_, _43093_, _43092_);
  and (_43095_, _43094_, _43091_);
  and (_43096_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_43097_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_43098_, _43097_, _43096_);
  and (_43099_, _43098_, _43095_);
  nor (_43100_, _43099_, _33994_);
  nor (_43101_, _43100_, _43088_);
  nor (_43102_, _43101_, _40480_);
  nor (_43103_, _43102_, _43087_);
  nor (_39042_, _43103_, rst);
  and (_43104_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_43105_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_43106_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_43107_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_43108_, _43107_, _43106_);
  and (_43109_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_43110_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_43111_, _43110_, _43109_);
  and (_43112_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_43113_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_43114_, _43113_, _43112_);
  and (_43115_, _43114_, _43111_);
  and (_43116_, _43115_, _43108_);
  nor (_43117_, _43116_, _33994_);
  nor (_43118_, _43117_, _43105_);
  nor (_43119_, _43118_, _40480_);
  nor (_43120_, _43119_, _43104_);
  nor (_39043_, _43120_, rst);
  and (_43121_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_43122_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_43123_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_43124_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_43125_, _43124_, _43123_);
  and (_43126_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_43127_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_43128_, _43127_, _43126_);
  and (_43129_, _43128_, _43125_);
  and (_43130_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_43131_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_43132_, _43131_, _43130_);
  and (_43133_, _43132_, _43129_);
  nor (_43134_, _43133_, _33994_);
  nor (_43135_, _43134_, _43122_);
  nor (_43136_, _43135_, _40480_);
  nor (_43137_, _43136_, _43121_);
  nor (_39044_, _43137_, rst);
  and (_43138_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_43139_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_43140_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_43141_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_43142_, _43141_, _43140_);
  and (_43143_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_43144_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_43145_, _43144_, _43143_);
  and (_43146_, _43145_, _43142_);
  and (_43147_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_43148_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_43149_, _43148_, _43147_);
  and (_43150_, _43149_, _43146_);
  nor (_43151_, _43150_, _33994_);
  nor (_43152_, _43151_, _43139_);
  nor (_43153_, _43152_, _40480_);
  nor (_43154_, _43153_, _43138_);
  nor (_39046_, _43154_, rst);
  and (_43155_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_43156_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_43157_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_43158_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_43159_, _43158_, _43157_);
  and (_43160_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_43161_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_43162_, _43161_, _43160_);
  and (_43163_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_43164_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_43165_, _43164_, _43163_);
  and (_43166_, _43165_, _43162_);
  and (_43167_, _43166_, _43159_);
  nor (_43168_, _43167_, _33994_);
  nor (_43169_, _43168_, _43156_);
  nor (_43170_, _43169_, _40480_);
  nor (_43171_, _43170_, _43155_);
  nor (_39047_, _43171_, rst);
  and (_43172_, _40480_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_43173_, _33994_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_43174_, _34038_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_43175_, _34082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_43176_, _43175_, _43174_);
  and (_43177_, _34126_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_43178_, _34203_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_43179_, _43178_, _43177_);
  and (_43180_, _34225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_43181_, _34170_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_43182_, _43181_, _43180_);
  and (_43183_, _43182_, _43179_);
  and (_43184_, _43183_, _43176_);
  nor (_43185_, _43184_, _33994_);
  nor (_43186_, _43185_, _43173_);
  nor (_43187_, _43186_, _40480_);
  nor (_43188_, _43187_, _43172_);
  nor (_39048_, _43188_, rst);
  and (_43189_, _33950_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_43190_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_43191_, _43189_, _38780_);
  and (_43192_, _43191_, _42003_);
  and (_39073_, _43192_, _43190_);
  not (_43193_, _43189_);
  or (_43194_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00001_, _43189_, _42003_);
  and (_43195_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42003_);
  or (_43196_, _43195_, _00001_);
  and (_39075_, _43196_, _43194_);
  nor (_39112_, _40501_, rst);
  and (_39114_, _39161_, _42003_);
  nor (_39115_, _40474_, rst);
  nor (_43197_, _40723_, _25344_);
  and (_43198_, _40723_, _25344_);
  nor (_43199_, _43198_, _43197_);
  nor (_43200_, _40639_, _24886_);
  and (_43201_, _40639_, _24886_);
  nor (_43202_, _43201_, _43200_);
  nor (_43203_, _43202_, _43199_);
  nor (_43204_, _40501_, _25061_);
  and (_43205_, _40501_, _25061_);
  nor (_43206_, _43205_, _43204_);
  nor (_43207_, _40836_, _24754_);
  and (_43208_, _40836_, _24754_);
  nor (_43209_, _43208_, _43207_);
  nor (_43210_, _43209_, _43206_);
  nor (_43211_, _40555_, _25213_);
  and (_43212_, _40555_, _25213_);
  nor (_43213_, _43212_, _43211_);
  not (_43214_, _43213_);
  and (_43215_, _43214_, _43210_);
  and (_43216_, _43215_, _43203_);
  nor (_43217_, _37639_, _42629_);
  and (_43218_, _39050_, _28199_);
  and (_43219_, _43218_, _43217_);
  and (_43220_, _43219_, _43216_);
  nor (_43221_, _26977_, _26943_);
  nor (_43222_, _28939_, _26705_);
  and (_43223_, _43222_, _43221_);
  nand (_43224_, _43223_, _30960_);
  nor (_43225_, _43224_, _31698_);
  and (_43226_, _43225_, _32482_);
  nor (_43227_, _43217_, _37771_);
  and (_43228_, _43227_, _43226_);
  and (_43229_, _43228_, _27162_);
  and (_43230_, _43217_, _26128_);
  nor (_43231_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_43232_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_43233_, _43232_, _43231_);
  nor (_43234_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_43235_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_43236_, _43235_, _43234_);
  and (_43237_, _43236_, _43233_);
  and (_43238_, _43237_, _36861_);
  not (_43239_, _37771_);
  nor (_43240_, _43217_, _34609_);
  nor (_43241_, _43240_, _43239_);
  and (_43242_, _43241_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_43243_, _43242_, _43238_);
  or (_43244_, _43243_, _43230_);
  nor (_43245_, _43244_, _43229_);
  not (_43246_, _42875_);
  and (_43247_, _43246_, _42681_);
  or (_43248_, _37606_, _36598_);
  or (_43249_, _43248_, _37080_);
  and (_43250_, _43249_, _36652_);
  nor (_43251_, _43250_, _42841_);
  and (_43252_, _43251_, _43247_);
  not (_43253_, _43252_);
  and (_43254_, _43253_, _43245_);
  and (_43255_, _37760_, _35874_);
  not (_43256_, _43255_);
  and (_43257_, _43256_, _37826_);
  nor (_43258_, _43257_, _43245_);
  nor (_43259_, _42610_, _36609_);
  not (_43260_, _43259_);
  or (_43261_, _43260_, _43258_);
  nor (_43262_, _43261_, _43254_);
  nor (_43263_, _43262_, _37782_);
  and (_43264_, _36400_, _35995_);
  nor (_43265_, _43264_, _42669_);
  nor (_43266_, _43265_, _33896_);
  nor (_43267_, _43266_, _36872_);
  not (_43268_, _43267_);
  nor (_43269_, _43268_, _43263_);
  nor (_43270_, _39049_, _39061_);
  and (_43271_, _43270_, _39070_);
  not (_43272_, _43271_);
  and (_43273_, _43272_, _43241_);
  not (_43274_, _39290_);
  and (_43275_, _43274_, _36861_);
  nor (_43276_, _43275_, _43273_);
  not (_43277_, _43276_);
  nor (_43278_, _43277_, _43269_);
  not (_43279_, _43278_);
  nor (_43280_, _43279_, _43220_);
  nand (_43281_, _43203_, _43210_);
  or (_43282_, _43213_, _39619_);
  or (_43283_, _40591_, _24535_);
  nand (_43284_, _40591_, _24535_);
  and (_43285_, _43284_, _43283_);
  and (_43286_, _40763_, _30776_);
  nor (_43287_, _40763_, _30776_);
  or (_43288_, _43287_, _43286_);
  or (_43289_, _43288_, _43285_);
  or (_43290_, _40676_, _24293_);
  nand (_43291_, _40676_, _24293_);
  and (_43292_, _43291_, _43290_);
  or (_43293_, _43292_, _43289_);
  or (_43294_, _43293_, _43282_);
  nor (_43295_, _43294_, _43281_);
  nor (_43296_, _25061_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_43297_, _43296_, _43295_);
  not (_43298_, _43297_);
  and (_43299_, _43298_, _43280_);
  nor (_43300_, _36883_, rst);
  and (_39119_, _43300_, _43299_);
  and (_39120_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42003_);
  and (_39121_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42003_);
  and (_43301_, _36883_, _28133_);
  and (_43302_, _36839_, _36609_);
  not (_43303_, _43302_);
  nor (_43304_, _43303_, _38791_);
  nor (_43305_, _42875_, _37353_);
  and (_43306_, _42840_, _37639_);
  and (_43307_, _43306_, _43305_);
  nor (_43308_, _43307_, _37782_);
  and (_43309_, _43264_, _36949_);
  nor (_43310_, _43309_, _37727_);
  not (_43311_, _43310_);
  nor (_43312_, _43311_, _43308_);
  and (_43313_, _43312_, _43266_);
  and (_43314_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43315_, _43314_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43316_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43317_, _43316_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43318_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43319_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43320_, _43319_, _43318_);
  and (_43321_, _43320_, _43317_);
  and (_43322_, _43321_, _43315_);
  and (_43323_, _43322_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43324_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43325_, _43324_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_43326_, _43325_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43327_, _43326_, _38780_);
  or (_43328_, _43326_, _38780_);
  and (_43329_, _43328_, _43327_);
  and (_43330_, _43329_, _43313_);
  and (_43331_, _43309_, _40497_);
  nor (_43332_, _43302_, _43266_);
  nand (_43334_, _43332_, _43312_);
  nor (_43335_, _43260_, _37760_);
  and (_43336_, _43335_, _43247_);
  and (_43337_, _43336_, _43306_);
  nor (_43338_, _43337_, _37782_);
  and (_43340_, _37584_, _36949_);
  or (_43341_, _43340_, _43338_);
  nor (_43342_, _43341_, _43334_);
  and (_43343_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_43344_, _43343_, _43331_);
  or (_43346_, _43344_, _43330_);
  nor (_43347_, _43346_, _43304_);
  nand (_43348_, _43347_, _43299_);
  or (_43349_, _43348_, _43301_);
  not (_43350_, _43068_);
  not (_43352_, _43340_);
  and (_43353_, _43352_, _43312_);
  nor (_43354_, _43353_, _43350_);
  and (_43355_, _43353_, _40496_);
  nor (_43356_, _43355_, _43354_);
  and (_43358_, _43356_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_43359_, _43356_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_43360_, _43188_);
  nor (_43361_, _43353_, _43360_);
  and (_43362_, _43353_, _40832_);
  nor (_43364_, _43362_, _43361_);
  and (_43365_, _43364_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43366_, _43364_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43367_, _43366_, _43365_);
  not (_43368_, _43171_);
  nor (_43370_, _43353_, _43368_);
  and (_43371_, _43353_, _40635_);
  nor (_43373_, _43371_, _43370_);
  and (_43374_, _43373_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_43375_, _43373_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_43376_, _43154_);
  nor (_43377_, _43353_, _43376_);
  and (_43378_, _43353_, _40717_);
  nor (_43379_, _43378_, _43377_);
  nand (_43381_, _43379_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_43382_, _43137_);
  nor (_43383_, _43353_, _43382_);
  and (_43385_, _43353_, _40534_);
  nor (_43386_, _43385_, _43383_);
  and (_43387_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_43389_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_43390_, _43120_);
  nor (_43391_, _43353_, _43390_);
  and (_43393_, _43353_, _40656_);
  nor (_43394_, _43393_, _43391_);
  and (_43395_, _43394_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_43397_, _43103_);
  nor (_43398_, _43353_, _43397_);
  and (_43399_, _43353_, _40739_);
  nor (_43401_, _43399_, _43398_);
  and (_43402_, _43401_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_43403_, _43086_);
  nor (_43405_, _43353_, _43403_);
  and (_43406_, _43353_, _40583_);
  nor (_43408_, _43406_, _43405_);
  and (_43409_, _43408_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_43410_, _43401_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_43411_, _43410_, _43402_);
  and (_43412_, _43411_, _43409_);
  nor (_43413_, _43412_, _43402_);
  not (_43414_, _43413_);
  nor (_43416_, _43394_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_43417_, _43416_, _43395_);
  and (_43418_, _43417_, _43414_);
  nor (_43420_, _43418_, _43395_);
  nor (_43421_, _43420_, _43389_);
  or (_43422_, _43421_, _43387_);
  or (_43424_, _43379_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43425_, _43424_, _43381_);
  nand (_43426_, _43425_, _43422_);
  and (_43428_, _43426_, _43381_);
  nor (_43429_, _43428_, _43375_);
  or (_43430_, _43429_, _43374_);
  and (_43432_, _43430_, _43367_);
  nor (_43433_, _43432_, _43365_);
  nor (_43434_, _43433_, _43359_);
  or (_43436_, _43434_, _43358_);
  and (_43437_, _43436_, _43315_);
  and (_43438_, _43437_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43440_, _43438_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43441_, _43440_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43443_, _43441_, _43356_);
  not (_43444_, _43356_);
  nor (_43445_, _43436_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43446_, _43445_, _38758_);
  and (_43447_, _43446_, _38763_);
  and (_43449_, _43447_, _38748_);
  nor (_43450_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43451_, _43450_, _43449_);
  nor (_43453_, _43451_, _43444_);
  nor (_43454_, _43453_, _43443_);
  or (_43455_, _43356_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43457_, _43356_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43458_, _43457_, _43455_);
  and (_43459_, _43458_, _43454_);
  or (_43461_, _43459_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_43462_, _43459_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_43463_, _43462_, _43461_);
  not (_43465_, _43332_);
  and (_43466_, _43465_, _43353_);
  and (_43467_, _36652_, _36949_);
  and (_43469_, _43467_, _35951_);
  nor (_43470_, _43469_, _43338_);
  nor (_43471_, _43470_, _43466_);
  and (_43473_, _43471_, _43463_);
  or (_43474_, _43473_, _43349_);
  not (_43476_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43478_, _43477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43479_, _43478_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43480_, _43479_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43481_, _43480_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43482_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43484_, _43482_, _43481_);
  and (_43485_, _43484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43486_, _43485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43488_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43489_, _34115_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43490_, _43489_, _40480_);
  nor (_43492_, _43490_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_43493_, _43492_);
  and (_43494_, _43493_, _43488_);
  and (_43496_, _43494_, _43486_);
  nand (_43497_, _43496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_43498_, _43497_, _43476_);
  or (_43500_, _43497_, _43476_);
  and (_43501_, _43500_, _43498_);
  or (_43502_, _43501_, _43299_);
  and (_43504_, _43502_, _42003_);
  and (_39123_, _43504_, _43474_);
  and (_43505_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42003_);
  and (_43507_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_43508_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_43510_, _33939_, _43508_);
  not (_43511_, _43510_);
  not (_43512_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_43513_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43515_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_43516_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_43517_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43519_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43520_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43521_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43523_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43524_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43525_, _43524_, _43523_);
  and (_43527_, _43525_, _43521_);
  and (_43528_, _43527_, _43520_);
  and (_43529_, _43528_, _43519_);
  and (_43531_, _43529_, _43517_);
  and (_43532_, _43531_, _43516_);
  and (_43533_, _43532_, _43515_);
  and (_43535_, _43533_, _43513_);
  and (_43536_, _43535_, _43512_);
  nor (_43537_, _43536_, _43476_);
  and (_43539_, _43536_, _43476_);
  nor (_43540_, _43539_, _43537_);
  nor (_43542_, _43535_, _43512_);
  nor (_43543_, _43542_, _43536_);
  not (_43544_, _43543_);
  not (_43545_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_43548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_43551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43552_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_43553_, _43552_, _43549_);
  and (_43555_, _43553_, _43551_);
  nor (_43556_, _43555_, _43549_);
  nor (_43557_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43559_, _43557_, _43548_);
  not (_43560_, _43559_);
  nor (_43561_, _43560_, _43556_);
  nor (_43563_, _43561_, _43548_);
  not (_43564_, _43563_);
  and (_43565_, _43564_, _43533_);
  and (_43567_, _43565_, _43547_);
  and (_43568_, _43567_, _43545_);
  and (_43569_, _43568_, _43544_);
  nor (_43571_, _43568_, _43544_);
  or (_43572_, _43571_, _43569_);
  not (_43574_, _43572_);
  and (_43575_, _43563_, _43535_);
  and (_43576_, _43563_, _43533_);
  and (_43577_, _43576_, _43547_);
  nor (_43579_, _43577_, _43545_);
  or (_43580_, _43579_, _43575_);
  nor (_43581_, _43576_, _43547_);
  nor (_43583_, _43581_, _43577_);
  not (_43584_, _43583_);
  and (_43585_, _43563_, _43532_);
  nor (_43587_, _43585_, _43515_);
  nor (_43588_, _43587_, _43576_);
  not (_43589_, _43588_);
  and (_43591_, _43563_, _43529_);
  and (_43592_, _43591_, _43517_);
  nor (_43593_, _43592_, _43516_);
  nor (_43595_, _43593_, _43585_);
  not (_43596_, _43595_);
  nor (_43597_, _43591_, _43517_);
  nor (_43599_, _43597_, _43592_);
  and (_43600_, _43563_, _43527_);
  and (_43601_, _43600_, _43520_);
  nor (_43603_, _43600_, _43520_);
  nor (_43604_, _43603_, _43601_);
  not (_43606_, _43604_);
  and (_43607_, _43563_, _43525_);
  nor (_43608_, _43607_, _43521_);
  nor (_43609_, _43608_, _43600_);
  not (_43610_, _43609_);
  and (_43611_, _43563_, _43524_);
  nor (_43612_, _43611_, _43523_);
  nor (_43614_, _43612_, _43607_);
  not (_43615_, _43614_);
  not (_43616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43618_, _43563_, _43616_);
  nor (_43619_, _43563_, _43616_);
  nor (_43620_, _43619_, _43618_);
  not (_43622_, _43620_);
  and (_43623_, _42583_, _42558_);
  not (_43624_, _43623_);
  nor (_43626_, _42549_, _42533_);
  and (_43627_, _43626_, _43624_);
  not (_43628_, _42547_);
  and (_43630_, _42542_, _42511_);
  nor (_43631_, _42571_, _43630_);
  nor (_43632_, _42589_, _42520_);
  nor (_43634_, _43632_, _36313_);
  not (_43635_, _43634_);
  and (_43636_, _43635_, _43631_);
  nor (_43638_, _43636_, _43628_);
  not (_43639_, _43638_);
  and (_43641_, _43639_, _43627_);
  and (_43642_, _42579_, _42558_);
  nor (_43643_, _43642_, _42521_);
  nor (_43644_, _42579_, _42540_);
  and (_43646_, _42543_, _42525_);
  not (_43647_, _43646_);
  nor (_43648_, _42583_, _42544_);
  and (_43650_, _43648_, _43647_);
  and (_43651_, _43650_, _43644_);
  nor (_43652_, _43651_, _43643_);
  not (_43654_, _42548_);
  and (_43655_, _42579_, _42516_);
  nor (_43656_, _43655_, _42566_);
  and (_43658_, _43656_, _43654_);
  nor (_43659_, _42579_, _42565_);
  and (_43660_, _42543_, _42526_);
  nor (_43662_, _43646_, _43660_);
  and (_43663_, _43662_, _43659_);
  nor (_43664_, _43663_, _43658_);
  nor (_43666_, _43664_, _43652_);
  and (_43667_, _43666_, _43641_);
  nor (_43668_, _42588_, _42551_);
  and (_43670_, _42558_, _42540_);
  and (_43671_, _42563_, _42545_);
  nor (_43673_, _43671_, _43670_);
  and (_43674_, _43673_, _43668_);
  and (_43675_, _42585_, _35578_);
  and (_43676_, _43675_, _42559_);
  or (_43678_, _43676_, _42564_);
  nor (_43679_, _43678_, _42537_);
  and (_43680_, _43679_, _43674_);
  and (_43682_, _42570_, _42519_);
  and (_43683_, _42558_, _43682_);
  and (_43684_, _42535_, _42518_);
  and (_43686_, _42585_, _43684_);
  and (_43687_, _43686_, _42552_);
  nor (_43688_, _43687_, _43683_);
  and (_43690_, _42571_, _42515_);
  and (_43691_, _42558_, _42577_);
  nor (_43692_, _43691_, _43690_);
  and (_43694_, _43692_, _43688_);
  and (_43695_, _43694_, _42582_);
  and (_43696_, _43695_, _43680_);
  and (_43698_, _42570_, _42511_);
  nor (_43699_, _43698_, _42540_);
  nor (_43700_, _43699_, _35578_);
  and (_43702_, _42535_, _42542_);
  not (_43703_, _43702_);
  nor (_43705_, _42547_, _42521_);
  nor (_43706_, _43705_, _43703_);
  nor (_43707_, _43706_, _43700_);
  nor (_43708_, _42540_, _42563_);
  nor (_43710_, _43708_, _43654_);
  not (_43711_, _43710_);
  and (_43712_, _42583_, _42548_);
  and (_43714_, _43702_, _42516_);
  nor (_43715_, _43714_, _43712_);
  and (_43716_, _43715_, _43711_);
  and (_43718_, _43716_, _43707_);
  and (_43719_, _42536_, _42511_);
  and (_43720_, _42521_, _42511_);
  and (_43722_, _43720_, _42525_);
  nor (_43723_, _43722_, _43719_);
  not (_43724_, _42531_);
  and (_43726_, _42543_, _34565_);
  nor (_43727_, _43698_, _43726_);
  nor (_43728_, _43727_, _43724_);
  and (_43730_, _43720_, _42527_);
  nor (_43731_, _43730_, _43728_);
  and (_43734_, _43731_, _43723_);
  and (_43741_, _43734_, _43718_);
  and (_43742_, _43741_, _43696_);
  and (_43755_, _43742_, _43667_);
  nor (_43756_, _43553_, _43551_);
  nor (_43760_, _43756_, _43555_);
  not (_43768_, _43760_);
  nor (_43778_, _43768_, _43755_);
  and (_43785_, _43715_, _43627_);
  nor (_43786_, _42588_, _42566_);
  and (_43798_, _43786_, _43711_);
  nor (_43803_, _43655_, _42578_);
  and (_43804_, _42531_, _43630_);
  and (_43818_, _42571_, _42516_);
  nor (_43823_, _43818_, _43804_);
  and (_43824_, _43823_, _43803_);
  and (_43837_, _43824_, _43798_);
  and (_43843_, _43837_, _43785_);
  not (_43844_, _43843_);
  nor (_43855_, _43844_, _43755_);
  not (_43863_, _43855_);
  nor (_43864_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43873_, _43864_, _43551_);
  and (_43882_, _43873_, _43863_);
  and (_43883_, _43768_, _43755_);
  nor (_43891_, _43883_, _43778_);
  and (_43900_, _43891_, _43882_);
  nor (_43901_, _43900_, _43778_);
  not (_43912_, _43901_);
  and (_43913_, _43560_, _43556_);
  nor (_43919_, _43913_, _43561_);
  and (_43930_, _43919_, _43912_);
  and (_43937_, _43930_, _43622_);
  not (_43938_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43950_, _43618_, _43938_);
  or (_43955_, _43950_, _43611_);
  and (_43956_, _43955_, _43937_);
  and (_43970_, _43956_, _43615_);
  and (_43973_, _43970_, _43610_);
  and (_43974_, _43973_, _43606_);
  nor (_43975_, _43601_, _43519_);
  or (_43977_, _43975_, _43591_);
  nand (_43978_, _43977_, _43974_);
  nor (_43979_, _43978_, _43599_);
  and (_43981_, _43979_, _43596_);
  and (_43982_, _43981_, _43589_);
  and (_43983_, _43982_, _43584_);
  and (_43985_, _43983_, _43580_);
  and (_43986_, _43985_, _43574_);
  nor (_43987_, _43986_, _43569_);
  not (_43989_, _43987_);
  nor (_43990_, _43989_, _43540_);
  and (_43992_, _43989_, _43540_);
  or (_43993_, _43992_, _43990_);
  or (_43994_, _43993_, _43511_);
  or (_43995_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_43997_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_43998_, _43997_, _43995_);
  and (_43999_, _43998_, _43994_);
  or (_39124_, _43999_, _43507_);
  nor (_44001_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_39125_, _44001_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_39126_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42003_);
  not (_44003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_44004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_44006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_44007_, _44006_, _44004_);
  not (_44008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_44010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_44011_, _44010_, _44008_);
  and (_44012_, _44011_, _44007_);
  and (_44014_, _44012_, _44003_);
  and (_44015_, \oc8051_top_1.oc8051_rom1.ea_int , _33907_);
  nand (_44016_, _44015_, _33939_);
  nand (_44018_, _44016_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_44019_, _44018_, _44014_);
  and (_39128_, _44019_, _42003_);
  and (_44021_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_44022_, _44021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_39129_, _44022_, _42003_);
  nor (_44024_, _43492_, _40480_);
  nor (_44025_, _43755_, _34060_);
  nor (_44026_, _43855_, _34158_);
  and (_44028_, _43755_, _34060_);
  nor (_44029_, _44028_, _44025_);
  and (_44030_, _44029_, _44026_);
  nor (_44032_, _44030_, _44025_);
  nor (_44033_, _44032_, _40480_);
  and (_44034_, _44033_, _34016_);
  nor (_44036_, _44033_, _34016_);
  nor (_44037_, _44036_, _44034_);
  nor (_44038_, _44037_, _44024_);
  and (_44040_, _34071_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_44041_, _44040_, _44024_);
  nor (_44042_, _44041_, _43843_);
  or (_44044_, _44042_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_44045_, _44044_, _44038_);
  and (_39130_, _44045_, _42003_);
  not (_44047_, _35015_);
  and (_44048_, _34269_, _44047_);
  not (_44049_, _35764_);
  and (_44050_, _44049_, _34762_);
  and (_44051_, _44050_, _44048_);
  and (_44052_, _33950_, _42003_);
  nand (_44053_, _44052_, _35278_);
  nor (_44054_, _44053_, _35543_);
  not (_44055_, _34521_);
  nor (_44056_, _36269_, _44055_);
  and (_44057_, _44056_, _44054_);
  and (_39133_, _44057_, _44051_);
  nor (_44058_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_44059_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_44060_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_39136_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42003_);
  and (_44061_, _39136_, _44060_);
  or (_39135_, _44061_, _44059_);
  not (_44062_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_44063_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44064_, _44063_, _44062_);
  and (_44065_, _44063_, _44062_);
  nor (_44066_, _44065_, _44064_);
  not (_44067_, _44066_);
  and (_44068_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44069_, _44068_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44070_, _44068_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44071_, _44070_, _44069_);
  or (_44072_, _44071_, _44063_);
  and (_44073_, _44072_, _44067_);
  nor (_44074_, _44064_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44075_, _44064_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_44076_, _44075_, _44074_);
  or (_44077_, _44069_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_39138_, _44077_, _42003_);
  and (_44078_, _39138_, _44076_);
  and (_39137_, _44078_, _44073_);
  not (_44079_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_44080_, _43492_, _44079_);
  and (_44081_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_44082_, _44080_);
  and (_44083_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_44084_, _44083_, _44081_);
  and (_39139_, _44084_, _42003_);
  and (_44085_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_44086_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_44087_, _44086_, _44085_);
  and (_39140_, _44087_, _42003_);
  and (_44088_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_44089_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44090_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _44089_);
  and (_44091_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_44092_, _44091_, _44088_);
  and (_39142_, _44092_, _42003_);
  and (_44093_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44094_, _44093_, _44090_);
  and (_39143_, _44094_, _42003_);
  or (_44095_, _44089_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_39144_, _44095_, _42003_);
  not (_44096_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_44097_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_44098_, _44097_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44099_, _44089_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_44100_, _44099_, _42003_);
  and (_39145_, _44100_, _44098_);
  or (_44101_, _44089_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_39146_, _44101_, _42003_);
  nor (_44102_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_44103_, _44102_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44104_, _44103_, _42003_);
  and (_44105_, _39136_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39147_, _44105_, _44104_);
  and (_44106_, _44079_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_44107_, _44106_, _44103_);
  and (_39148_, _44107_, _42003_);
  nand (_44108_, _44103_, _38791_);
  or (_44109_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_44110_, _44109_, _42003_);
  and (_39149_, _44110_, _44108_);
  and (_39150_, _38101_, _40443_);
  or (_44111_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_44112_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_44113_, _43189_, _44112_);
  and (_44114_, _44113_, _42003_);
  and (_39185_, _44114_, _44111_);
  or (_44115_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_44116_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_44117_, _43189_, _44116_);
  and (_44118_, _44117_, _42003_);
  and (_39186_, _44118_, _44115_);
  or (_44119_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_44120_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_44121_, _43189_, _44120_);
  and (_44122_, _44121_, _42003_);
  and (_39187_, _44122_, _44119_);
  or (_44123_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_44124_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _42003_);
  or (_44125_, _44124_, _00001_);
  and (_39189_, _44125_, _44123_);
  or (_44126_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_44127_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_44128_, _43189_, _44127_);
  and (_44129_, _44128_, _42003_);
  and (_39190_, _44129_, _44126_);
  or (_44130_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_44131_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_44132_, _43189_, _44131_);
  and (_44133_, _44132_, _42003_);
  and (_39191_, _44133_, _44130_);
  or (_44134_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_44135_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_44136_, _43189_, _44135_);
  and (_44137_, _44136_, _42003_);
  and (_39192_, _44137_, _44134_);
  or (_44138_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_44139_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_44140_, _43189_, _44139_);
  and (_44141_, _44140_, _42003_);
  and (_39193_, _44141_, _44138_);
  or (_44142_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_44143_, _43189_, _38752_);
  and (_44144_, _44143_, _42003_);
  and (_39194_, _44144_, _44142_);
  or (_44145_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_44146_, _43189_, _38758_);
  and (_44147_, _44146_, _42003_);
  and (_39195_, _44147_, _44145_);
  or (_44148_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_44149_, _43189_, _38763_);
  and (_44150_, _44149_, _42003_);
  and (_39196_, _44150_, _44148_);
  or (_44151_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_44152_, _43189_, _38748_);
  and (_44153_, _44152_, _42003_);
  and (_39197_, _44153_, _44151_);
  or (_44154_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_44155_, _43189_, _38769_);
  and (_44156_, _44155_, _42003_);
  and (_39198_, _44156_, _44154_);
  or (_44157_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_44158_, _43189_, _38744_);
  and (_44159_, _44158_, _42003_);
  and (_39200_, _44159_, _44157_);
  or (_44160_, _43189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_44161_, _43189_, _38775_);
  and (_44162_, _44161_, _42003_);
  and (_39201_, _44162_, _44160_);
  or (_44163_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_44164_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _42003_);
  or (_44165_, _44164_, _00001_);
  and (_39205_, _44165_, _44163_);
  or (_44166_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_44167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _42003_);
  or (_44168_, _44167_, _00001_);
  and (_39206_, _44168_, _44166_);
  or (_44169_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_44170_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _42003_);
  or (_44171_, _44170_, _00001_);
  and (_39207_, _44171_, _44169_);
  or (_44172_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_44173_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _42003_);
  or (_44174_, _44173_, _00001_);
  and (_39208_, _44174_, _44172_);
  or (_44175_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_44176_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _42003_);
  or (_44177_, _44176_, _00001_);
  and (_39209_, _44177_, _44175_);
  or (_44178_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_44179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _42003_);
  or (_44180_, _44179_, _00001_);
  and (_39210_, _44180_, _44178_);
  or (_44181_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_44182_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _42003_);
  or (_44183_, _44182_, _00001_);
  and (_39211_, _44183_, _44181_);
  or (_44184_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_44185_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _42003_);
  or (_44186_, _44185_, _00001_);
  and (_39212_, _44186_, _44184_);
  or (_44187_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_44188_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _42003_);
  or (_44189_, _44188_, _00001_);
  and (_39214_, _44189_, _44187_);
  or (_44190_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_44191_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _42003_);
  or (_44192_, _44191_, _00001_);
  and (_39215_, _44192_, _44190_);
  or (_44193_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_44194_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _42003_);
  or (_44195_, _44194_, _00001_);
  and (_39216_, _44195_, _44193_);
  or (_44196_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_44197_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _42003_);
  or (_44198_, _44197_, _00001_);
  and (_39217_, _44198_, _44196_);
  or (_44199_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_44200_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _42003_);
  or (_44201_, _44200_, _00001_);
  and (_39218_, _44201_, _44199_);
  or (_44202_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_44203_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _42003_);
  or (_44204_, _44203_, _00001_);
  and (_39219_, _44204_, _44202_);
  or (_44205_, _43193_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_44206_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _42003_);
  or (_44207_, _44206_, _00001_);
  and (_39220_, _44207_, _44205_);
  and (_44208_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_44209_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_44210_, _44209_, _44208_);
  and (_39397_, _44210_, _42003_);
  and (_44211_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_44212_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_44213_, _44212_, _44211_);
  and (_39398_, _44213_, _42003_);
  and (_44214_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_44215_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_44216_, _44215_, _44214_);
  and (_39399_, _44216_, _42003_);
  and (_44217_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_44218_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_44219_, _44218_, _44217_);
  and (_39400_, _44219_, _42003_);
  and (_44220_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_44221_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_44222_, _44221_, _44220_);
  and (_39401_, _44222_, _42003_);
  and (_44223_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_44224_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_44225_, _44224_, _44223_);
  and (_39402_, _44225_, _42003_);
  and (_44226_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_44227_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_44228_, _44227_, _44226_);
  and (_39404_, _44228_, _42003_);
  and (_44229_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_44230_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_44231_, _44230_, _44229_);
  and (_39405_, _44231_, _42003_);
  and (_44232_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_44233_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_44234_, _44233_, _44232_);
  and (_39406_, _44234_, _42003_);
  and (_44235_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_44236_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_44237_, _44236_, _44235_);
  and (_39407_, _44237_, _42003_);
  and (_44238_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_44239_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_44240_, _44239_, _44238_);
  and (_39408_, _44240_, _42003_);
  and (_44241_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_44242_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_44243_, _44242_, _44241_);
  and (_39409_, _44243_, _42003_);
  and (_44244_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_44245_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_44246_, _44245_, _44244_);
  and (_39410_, _44246_, _42003_);
  and (_44247_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_44248_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_44249_, _44248_, _44247_);
  and (_39411_, _44249_, _42003_);
  and (_44250_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_44251_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_44252_, _44251_, _44250_);
  and (_39412_, _44252_, _42003_);
  and (_44253_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_44254_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_44255_, _44254_, _44253_);
  and (_39413_, _44255_, _42003_);
  and (_00011_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_00012_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_00013_, _00012_, _00011_);
  and (_39415_, _00013_, _42003_);
  and (_00014_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_00015_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_00016_, _00015_, _00014_);
  and (_39416_, _00016_, _42003_);
  and (_00017_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_00018_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_00019_, _00018_, _00017_);
  and (_39417_, _00019_, _42003_);
  and (_00020_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_00021_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_00022_, _00021_, _00020_);
  and (_39418_, _00022_, _42003_);
  and (_00023_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_00024_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_00025_, _00024_, _00023_);
  and (_39419_, _00025_, _42003_);
  and (_00026_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_00027_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_00028_, _00027_, _00026_);
  and (_39420_, _00028_, _42003_);
  and (_00029_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_00030_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00031_, _00030_, _00029_);
  and (_39421_, _00031_, _42003_);
  and (_00032_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_00033_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_00034_, _00033_, _00032_);
  and (_39422_, _00034_, _42003_);
  and (_00035_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_00036_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_00037_, _00036_, _00035_);
  and (_39423_, _00037_, _42003_);
  and (_00038_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_00039_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_00040_, _00039_, _00038_);
  and (_39424_, _00040_, _42003_);
  and (_00041_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_00042_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_00043_, _00042_, _00041_);
  and (_39426_, _00043_, _42003_);
  and (_00044_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_00045_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_00046_, _00045_, _00044_);
  and (_39427_, _00046_, _42003_);
  and (_00047_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_00048_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_00049_, _00048_, _00047_);
  and (_39428_, _00049_, _42003_);
  and (_00050_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_00051_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_00052_, _00051_, _00050_);
  and (_39429_, _00052_, _42003_);
  and (_00053_, _44080_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_00054_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_00055_, _00054_, _00053_);
  and (_39430_, _00055_, _42003_);
  nor (_39431_, _36356_, rst);
  nor (_39432_, _35135_, rst);
  nor (_39433_, _35366_, rst);
  nor (_39434_, _40447_, rst);
  nor (_39436_, _40567_, rst);
  nor (_39437_, _40752_, rst);
  nor (_39438_, _40672_, rst);
  nor (_39439_, _40551_, rst);
  nor (_39440_, _40697_, rst);
  nor (_39442_, _40611_, rst);
  nor (_39443_, _40814_, rst);
  and (_39459_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42003_);
  and (_39460_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42003_);
  and (_39461_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42003_);
  and (_39463_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42003_);
  and (_39464_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42003_);
  and (_39465_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42003_);
  and (_39466_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42003_);
  or (_00056_, _43342_, _43302_);
  and (_00057_, _00056_, _29299_);
  and (_00058_, _43313_, _40584_);
  and (_00059_, _43309_, _43403_);
  or (_00060_, _00059_, _00058_);
  and (_00061_, _37727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00062_, _00061_, _00060_);
  nor (_00063_, _43408_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00064_, _00063_, _43409_);
  and (_00065_, _00064_, _43471_);
  nor (_00066_, _00065_, _00062_);
  nand (_00067_, _00066_, _43299_);
  or (_00068_, _00067_, _00057_);
  or (_00069_, _43299_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00070_, _00069_, _42003_);
  and (_39467_, _00070_, _00068_);
  and (_00071_, _00056_, _29972_);
  and (_00072_, _43313_, _40740_);
  and (_00073_, _43309_, _43397_);
  and (_00074_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00075_, _00074_, _00073_);
  or (_00076_, _00075_, _00072_);
  or (_00077_, _00076_, _00071_);
  nor (_00078_, _43411_, _43409_);
  nor (_00079_, _00078_, _43412_);
  nand (_00080_, _00079_, _43471_);
  nand (_00081_, _00080_, _43299_);
  or (_00082_, _00081_, _00077_);
  or (_00083_, _43299_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00084_, _00083_, _42003_);
  and (_39468_, _00084_, _00082_);
  and (_00085_, _00056_, _30667_);
  and (_00086_, _43313_, _40657_);
  and (_00087_, _43309_, _43390_);
  or (_00088_, _00087_, _00086_);
  or (_00089_, _43417_, _43414_);
  not (_00090_, _43471_);
  nor (_00091_, _00090_, _43418_);
  and (_00092_, _00091_, _00089_);
  or (_00093_, _00092_, _00088_);
  or (_00094_, _00093_, _00085_);
  nand (_00095_, _37727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand (_00096_, _00095_, _43299_);
  or (_00097_, _00096_, _00094_);
  not (_00098_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00099_, _43492_, _00098_);
  and (_00100_, _43492_, _00098_);
  nor (_00101_, _00100_, _00099_);
  or (_00102_, _00101_, _43299_);
  and (_00103_, _00102_, _42003_);
  and (_39469_, _00103_, _00097_);
  and (_00104_, _00056_, _31427_);
  or (_00105_, _43389_, _43387_);
  and (_00106_, _00105_, _43420_);
  not (_00107_, _43466_);
  and (_00108_, _43341_, _00107_);
  or (_00109_, _00105_, _43420_);
  nand (_00110_, _00109_, _00108_);
  or (_00111_, _00110_, _00106_);
  and (_00112_, _43313_, _40535_);
  and (_00113_, _43309_, _43382_);
  and (_00114_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00115_, _00114_, _00113_);
  nor (_00116_, _00115_, _00112_);
  and (_00117_, _00116_, _00111_);
  nand (_00118_, _00117_, _43299_);
  or (_00119_, _00118_, _00104_);
  and (_00120_, _00099_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00121_, _00099_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00122_, _00121_, _00120_);
  or (_00123_, _00122_, _43299_);
  and (_00124_, _00123_, _42003_);
  and (_39470_, _00124_, _00119_);
  and (_00125_, _00056_, _32144_);
  and (_00126_, _43313_, _40718_);
  and (_00127_, _43309_, _43376_);
  and (_00128_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00129_, _00128_, _00127_);
  or (_00130_, _00129_, _00126_);
  or (_00131_, _43425_, _43422_);
  and (_00132_, _00108_, _43426_);
  and (_00133_, _00132_, _00131_);
  nor (_00134_, _00133_, _00130_);
  nand (_00135_, _00134_, _43299_);
  or (_00136_, _00135_, _00125_);
  and (_00137_, _43478_, _43493_);
  nor (_00138_, _00120_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00139_, _00138_, _00137_);
  or (_00140_, _00139_, _43299_);
  and (_00141_, _00140_, _42003_);
  and (_39471_, _00141_, _00136_);
  and (_00142_, _00056_, _32954_);
  or (_00143_, _43375_, _43374_);
  nand (_00144_, _00143_, _43428_);
  or (_00145_, _00143_, _43428_);
  and (_00146_, _00145_, _00108_);
  and (_00147_, _00146_, _00144_);
  and (_00148_, _43313_, _40636_);
  and (_00149_, _43309_, _43368_);
  and (_00150_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00151_, _00150_, _00149_);
  or (_00152_, _00151_, _00148_);
  nor (_00153_, _00152_, _00147_);
  nand (_00154_, _00153_, _43299_);
  or (_00155_, _00154_, _00142_);
  and (_00156_, _43479_, _43493_);
  nor (_00157_, _00137_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00158_, _00157_, _00156_);
  or (_00159_, _00158_, _43299_);
  and (_00160_, _00159_, _42003_);
  and (_39472_, _00160_, _00155_);
  not (_00161_, _43299_);
  nor (_00162_, _43430_, _43367_);
  nor (_00163_, _00162_, _43432_);
  and (_00164_, _00163_, _43471_);
  and (_00165_, _00056_, _33688_);
  and (_00166_, _43313_, _40833_);
  and (_00167_, _43309_, _43360_);
  and (_00168_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00169_, _00168_, _00167_);
  or (_00170_, _00169_, _00166_);
  or (_00171_, _00170_, _00165_);
  or (_00172_, _00171_, _00164_);
  or (_00173_, _00172_, _00161_);
  and (_00174_, _00156_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00175_, _00156_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00176_, _00175_, _00174_);
  or (_00177_, _00176_, _43299_);
  and (_00178_, _00177_, _42003_);
  and (_39474_, _00178_, _00173_);
  or (_00179_, _43358_, _43359_);
  and (_00180_, _00179_, _43433_);
  nor (_00181_, _00179_, _43433_);
  or (_00182_, _00181_, _00180_);
  or (_00183_, _00182_, _00090_);
  and (_00184_, _00056_, _28133_);
  and (_00185_, _43313_, _40497_);
  and (_00186_, _43309_, _43350_);
  and (_00187_, _36883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00188_, _00187_, _00186_);
  or (_00189_, _00188_, _00185_);
  nor (_00190_, _00189_, _00184_);
  and (_00191_, _00190_, _00183_);
  nand (_00192_, _00191_, _43299_);
  and (_00193_, _00174_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00194_, _00174_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00195_, _00194_, _00193_);
  or (_00196_, _00195_, _43299_);
  and (_00197_, _00196_, _42003_);
  and (_39475_, _00197_, _00192_);
  nor (_00198_, _37738_, _29288_);
  and (_00199_, _43436_, _38752_);
  nor (_00200_, _43436_, _38752_);
  nor (_00201_, _00200_, _00199_);
  nor (_00202_, _00201_, _43356_);
  and (_00203_, _00201_, _43356_);
  or (_00204_, _00203_, _00202_);
  and (_00205_, _00204_, _43471_);
  nor (_00206_, _43303_, _38828_);
  and (_00207_, _43313_, _42518_);
  and (_00208_, _43309_, _40584_);
  and (_00209_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00210_, _00209_, _00208_);
  or (_00211_, _00210_, _00207_);
  or (_00212_, _00211_, _00206_);
  or (_00213_, _00212_, _00205_);
  or (_00214_, _00213_, _00198_);
  or (_00215_, _00214_, _00161_);
  and (_00216_, _00193_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00217_, _00193_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00218_, _00217_, _00216_);
  or (_00219_, _00218_, _43299_);
  and (_00220_, _00219_, _42003_);
  and (_39476_, _00220_, _00215_);
  and (_00221_, _43436_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00222_, _00221_, _43444_);
  and (_00223_, _43445_, _43356_);
  nor (_00224_, _00223_, _00222_);
  nand (_00225_, _00224_, _38758_);
  or (_00226_, _00224_, _38758_);
  and (_00227_, _00226_, _00108_);
  and (_00228_, _00227_, _00225_);
  nor (_00229_, _43303_, _38856_);
  and (_00230_, _43313_, _42534_);
  and (_00231_, _43309_, _40740_);
  and (_00232_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00233_, _00232_, _00231_);
  or (_00234_, _00233_, _00230_);
  nor (_00235_, _00234_, _00229_);
  nand (_00236_, _00235_, _43299_);
  or (_00237_, _00236_, _00228_);
  nor (_00238_, _37738_, _29961_);
  or (_00239_, _00238_, _00237_);
  and (_00240_, _43484_, _43493_);
  nor (_00241_, _00216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00242_, _00241_, _00240_);
  or (_00243_, _00242_, _43299_);
  and (_00244_, _00243_, _42003_);
  and (_39477_, _00244_, _00239_);
  and (_00245_, _36883_, _30667_);
  and (_00246_, _43446_, _43356_);
  and (_00247_, _00222_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_00248_, _00247_, _00246_);
  nand (_00249_, _00248_, _38763_);
  or (_00250_, _00248_, _38763_);
  and (_00251_, _00250_, _00108_);
  and (_00252_, _00251_, _00249_);
  nor (_00253_, _43303_, _38884_);
  and (_00254_, _43313_, _42510_);
  and (_00255_, _43309_, _40657_);
  and (_00256_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_00257_, _00256_, _00255_);
  or (_00258_, _00257_, _00254_);
  nor (_00259_, _00258_, _00253_);
  nand (_00260_, _00259_, _43299_);
  or (_00261_, _00260_, _00252_);
  or (_00262_, _00261_, _00245_);
  and (_00263_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00264_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00265_, _00264_, _00263_);
  or (_00266_, _00265_, _43299_);
  and (_00267_, _00266_, _42003_);
  and (_39478_, _00267_, _00262_);
  or (_00268_, _37738_, _31416_);
  or (_00269_, _43303_, _38913_);
  nor (_00270_, _43322_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00271_, _00270_, _43323_);
  nand (_00272_, _00271_, _43313_);
  nand (_00273_, _43309_, _40535_);
  nand (_00274_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00275_, _00274_, _00273_);
  and (_00276_, _00275_, _00272_);
  and (_00277_, _00276_, _00269_);
  and (_00278_, _43437_, _43444_);
  and (_00279_, _43447_, _43356_);
  nor (_00280_, _00279_, _00278_);
  and (_00281_, _00280_, _38748_);
  nor (_00282_, _00280_, _38748_);
  or (_00283_, _00282_, _00090_);
  or (_00284_, _00283_, _00281_);
  and (_00285_, _00284_, _00277_);
  and (_00286_, _00285_, _00268_);
  nand (_00287_, _00286_, _43299_);
  and (_00288_, _00263_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00289_, _00263_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00290_, _00289_, _00288_);
  or (_00291_, _00290_, _43299_);
  and (_00292_, _00291_, _42003_);
  and (_39479_, _00292_, _00287_);
  and (_00293_, _36883_, _32144_);
  and (_00294_, _43438_, _43444_);
  and (_00295_, _43449_, _43356_);
  nor (_00296_, _00295_, _00294_);
  nor (_00297_, _00296_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00298_, _00296_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_00299_, _00298_, _00297_);
  and (_00300_, _00299_, _00108_);
  nor (_00301_, _43303_, _38941_);
  nor (_00302_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00303_, _00302_, _43324_);
  and (_00304_, _00303_, _43313_);
  and (_00305_, _43309_, _40718_);
  and (_00306_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_00307_, _00306_, _00305_);
  or (_00308_, _00307_, _00304_);
  nor (_00309_, _00308_, _00301_);
  nand (_00310_, _00309_, _43299_);
  or (_00311_, _00310_, _00300_);
  or (_00312_, _00311_, _00293_);
  and (_00313_, _00288_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00314_, _00288_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00315_, _00314_, _00313_);
  or (_00316_, _00315_, _43299_);
  and (_00317_, _00316_, _42003_);
  and (_39480_, _00317_, _00312_);
  and (_00318_, _43440_, _43444_);
  and (_00319_, _00295_, _38769_);
  nor (_00320_, _00319_, _00318_);
  nand (_00321_, _00320_, _38744_);
  or (_00322_, _00320_, _38744_);
  and (_00323_, _00322_, _00108_);
  and (_00324_, _00323_, _00321_);
  and (_00325_, _36883_, _32954_);
  nor (_00326_, _43303_, _38970_);
  nor (_00327_, _43324_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00328_, _00327_, _43325_);
  and (_00329_, _00328_, _43313_);
  and (_00330_, _43309_, _40636_);
  and (_00331_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00332_, _00331_, _00330_);
  or (_00333_, _00332_, _00329_);
  nor (_00334_, _00333_, _00326_);
  nand (_00335_, _00334_, _43299_);
  or (_00336_, _00335_, _00325_);
  or (_00337_, _00336_, _00324_);
  or (_00338_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_00339_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00340_, _00339_, _00338_);
  or (_00341_, _00340_, _43299_);
  and (_00342_, _00341_, _42003_);
  and (_39481_, _00342_, _00337_);
  or (_00343_, _43454_, _38775_);
  nand (_00344_, _43454_, _38775_);
  nand (_00345_, _00344_, _00343_);
  and (_00346_, _00345_, _00108_);
  and (_00347_, _36883_, _33688_);
  or (_00348_, _43303_, _38996_);
  or (_00349_, _43325_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00350_, _00349_, _43326_);
  nand (_00351_, _00350_, _43313_);
  nand (_00352_, _43309_, _40833_);
  nand (_00353_, _43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00354_, _00353_, _00352_);
  and (_00355_, _00354_, _00351_);
  and (_00356_, _00355_, _00348_);
  nand (_00357_, _00356_, _43299_);
  or (_00358_, _00357_, _00347_);
  or (_00359_, _00358_, _00346_);
  or (_00360_, _43496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00361_, _00360_, _43497_);
  or (_00362_, _00361_, _43299_);
  and (_00363_, _00362_, _42003_);
  and (_39482_, _00363_, _00359_);
  or (_00364_, _43873_, _43863_);
  nor (_00365_, _43511_, _43882_);
  and (_00366_, _00365_, _00364_);
  nor (_00367_, _43510_, _44112_);
  or (_00368_, _00367_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00369_, _00368_, _00366_);
  or (_00370_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _33907_);
  and (_00371_, _00370_, _42003_);
  and (_39483_, _00371_, _00369_);
  nor (_00372_, _43891_, _43882_);
  nor (_00373_, _00372_, _43900_);
  or (_00374_, _00373_, _43511_);
  or (_00375_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00376_, _00375_, _43997_);
  and (_00377_, _00376_, _00374_);
  and (_00378_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39484_, _00378_, _00377_);
  and (_00379_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00380_, _43919_, _43912_);
  nor (_00381_, _00380_, _43930_);
  or (_00382_, _00381_, _43511_);
  or (_00383_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00384_, _00383_, _43997_);
  and (_00385_, _00384_, _00382_);
  or (_39485_, _00385_, _00379_);
  and (_00386_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00387_, _43930_, _43622_);
  nor (_00388_, _00387_, _43937_);
  or (_00389_, _00388_, _43511_);
  or (_00390_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00391_, _00390_, _43997_);
  and (_00392_, _00391_, _00389_);
  or (_39486_, _00392_, _00386_);
  and (_00393_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00394_, _43955_, _43937_);
  nor (_00395_, _00394_, _43956_);
  or (_00396_, _00395_, _43511_);
  or (_00397_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00398_, _00397_, _43997_);
  and (_00399_, _00398_, _00396_);
  or (_39487_, _00399_, _00393_);
  and (_00400_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00401_, _43956_, _43615_);
  nor (_00402_, _00401_, _43970_);
  or (_00403_, _00402_, _43511_);
  or (_00404_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00405_, _00404_, _43997_);
  and (_00406_, _00405_, _00403_);
  or (_39488_, _00406_, _00400_);
  and (_00407_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00408_, _43970_, _43610_);
  nor (_00409_, _00408_, _43973_);
  or (_00410_, _00409_, _43511_);
  or (_00411_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00412_, _00411_, _43997_);
  and (_00413_, _00412_, _00410_);
  or (_39489_, _00413_, _00407_);
  nor (_00414_, _43973_, _43606_);
  nor (_00415_, _00414_, _43974_);
  or (_00416_, _00415_, _43511_);
  or (_00417_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00418_, _00417_, _43997_);
  and (_00419_, _00418_, _00416_);
  and (_00420_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_39490_, _00420_, _00419_);
  or (_00421_, _43977_, _43974_);
  and (_00422_, _00421_, _43978_);
  or (_00423_, _00422_, _43511_);
  or (_00424_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00425_, _00424_, _43997_);
  and (_00426_, _00425_, _00423_);
  and (_00427_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_39491_, _00427_, _00426_);
  and (_00428_, _43978_, _43599_);
  nor (_00429_, _00428_, _43979_);
  or (_00430_, _00429_, _43511_);
  or (_00431_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00432_, _00431_, _43997_);
  and (_00433_, _00432_, _00430_);
  and (_00434_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39492_, _00434_, _00433_);
  nor (_00435_, _43979_, _43596_);
  nor (_00436_, _00435_, _43981_);
  or (_00437_, _00436_, _43511_);
  or (_00438_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00439_, _00438_, _43997_);
  and (_00440_, _00439_, _00437_);
  and (_00441_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39493_, _00441_, _00440_);
  nor (_00442_, _43981_, _43589_);
  nor (_00443_, _00442_, _43982_);
  or (_00444_, _00443_, _43511_);
  or (_00445_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00446_, _00445_, _43997_);
  and (_00447_, _00446_, _00444_);
  and (_00448_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39495_, _00448_, _00447_);
  nor (_00449_, _43982_, _43584_);
  nor (_00450_, _00449_, _43983_);
  or (_00451_, _00450_, _43511_);
  or (_00452_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00453_, _00452_, _43997_);
  and (_00454_, _00453_, _00451_);
  and (_00455_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39496_, _00455_, _00454_);
  nor (_00456_, _43983_, _43580_);
  nor (_00457_, _00456_, _43985_);
  or (_00458_, _00457_, _43511_);
  or (_00459_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00460_, _00459_, _43997_);
  and (_00461_, _00460_, _00458_);
  and (_00462_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39497_, _00462_, _00461_);
  and (_00463_, _43505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00464_, _43985_, _43574_);
  nor (_00465_, _00464_, _43986_);
  or (_00466_, _00465_, _43511_);
  or (_00467_, _43510_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00468_, _00467_, _43997_);
  and (_00469_, _00468_, _00466_);
  or (_39498_, _00469_, _00463_);
  and (_00470_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00471_, _00470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39499_, _00471_, _42003_);
  and (_00472_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_00473_, _00472_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39500_, _00473_, _42003_);
  and (_00474_, _44012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_00475_, _00474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39501_, _00475_, _42003_);
  and (_00476_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00477_, _00476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39502_, _00477_, _42003_);
  and (_00478_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00479_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39503_, _00479_, _42003_);
  and (_00480_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00481_, _00480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39504_, _00481_, _42003_);
  and (_00482_, _44014_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39506_, _00483_, _42003_);
  nor (_00484_, _43855_, _40480_);
  nand (_00485_, _00484_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00486_, _00484_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00487_, _00486_, _43997_);
  and (_39507_, _00487_, _00485_);
  nor (_00488_, _44029_, _44026_);
  nor (_00489_, _00488_, _44030_);
  or (_00490_, _00489_, _40480_);
  or (_00491_, _33939_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00492_, _00491_, _43997_);
  and (_39508_, _00492_, _00490_);
  and (_00493_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00494_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00495_, _00494_, _39136_);
  or (_39524_, _00495_, _00493_);
  and (_00496_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00497_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00498_, _00497_, _39136_);
  or (_39525_, _00498_, _00496_);
  and (_00499_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00500_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00501_, _00500_, _39136_);
  or (_39526_, _00501_, _00499_);
  and (_00502_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00503_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00504_, _00503_, _39136_);
  or (_39528_, _00504_, _00502_);
  and (_00505_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00506_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00507_, _00506_, _39136_);
  or (_39529_, _00507_, _00505_);
  and (_00508_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00509_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00510_, _00509_, _39136_);
  or (_39530_, _00510_, _00508_);
  and (_00511_, _44058_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00512_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00513_, _00512_, _39136_);
  or (_39531_, _00513_, _00511_);
  and (_39532_, _44066_, _42003_);
  nor (_39533_, _44076_, rst);
  and (_39534_, _44072_, _42003_);
  and (_00514_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00515_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00516_, _00515_, _00514_);
  and (_39535_, _00516_, _42003_);
  and (_00517_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00518_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00519_, _00518_, _00517_);
  and (_39536_, _00519_, _42003_);
  and (_00520_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00521_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00522_, _00521_, _00520_);
  and (_39537_, _00522_, _42003_);
  and (_00523_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00524_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00525_, _00524_, _00523_);
  and (_39539_, _00525_, _42003_);
  and (_00526_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00527_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00528_, _00527_, _00526_);
  and (_39540_, _00528_, _42003_);
  and (_00529_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00530_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00531_, _00530_, _00529_);
  and (_39541_, _00531_, _42003_);
  and (_00532_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00533_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00534_, _00533_, _00532_);
  and (_39542_, _00534_, _42003_);
  and (_00535_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00536_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00537_, _00536_, _00535_);
  and (_39543_, _00537_, _42003_);
  and (_00538_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00539_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00540_, _00539_, _00538_);
  and (_39544_, _00540_, _42003_);
  and (_00541_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00542_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00543_, _00542_, _00541_);
  and (_39545_, _00543_, _42003_);
  and (_00544_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00545_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00546_, _00545_, _00544_);
  and (_39546_, _00546_, _42003_);
  and (_00547_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00548_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00549_, _00548_, _00547_);
  and (_39547_, _00549_, _42003_);
  and (_00550_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00551_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00552_, _00551_, _00550_);
  and (_39548_, _00552_, _42003_);
  and (_00553_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00554_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00555_, _00554_, _00553_);
  and (_39550_, _00555_, _42003_);
  and (_00556_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00557_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00558_, _00557_, _00556_);
  and (_39551_, _00558_, _42003_);
  and (_00559_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00560_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00561_, _00560_, _00559_);
  and (_39552_, _00561_, _42003_);
  and (_00562_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00563_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00564_, _00563_, _00562_);
  and (_39553_, _00564_, _42003_);
  and (_00565_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00566_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00567_, _00566_, _00565_);
  and (_39554_, _00567_, _42003_);
  and (_00568_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00569_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00570_, _00569_, _00568_);
  and (_39555_, _00570_, _42003_);
  and (_00571_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00572_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00573_, _00572_, _00571_);
  and (_39556_, _00573_, _42003_);
  and (_00574_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00575_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00576_, _00575_, _00574_);
  and (_39557_, _00576_, _42003_);
  and (_00577_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00578_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00579_, _00578_, _00577_);
  and (_39558_, _00579_, _42003_);
  and (_00580_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00581_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00582_, _00581_, _00580_);
  and (_39559_, _00582_, _42003_);
  and (_00583_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00584_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00585_, _00584_, _00583_);
  and (_39561_, _00585_, _42003_);
  and (_00586_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00587_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00588_, _00587_, _00586_);
  and (_39562_, _00588_, _42003_);
  and (_00589_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00590_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00591_, _00590_, _00589_);
  and (_39563_, _00591_, _42003_);
  and (_00592_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00593_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00594_, _00593_, _00592_);
  and (_39564_, _00594_, _42003_);
  and (_00595_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00596_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00597_, _00596_, _00595_);
  and (_39565_, _00597_, _42003_);
  and (_00598_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00599_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00600_, _00599_, _00598_);
  and (_39566_, _00600_, _42003_);
  and (_00601_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00602_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00603_, _00602_, _00601_);
  and (_39567_, _00603_, _42003_);
  and (_00604_, _44080_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00605_, _44082_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00606_, _00605_, _00604_);
  and (_39568_, _00606_, _42003_);
  and (_00607_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00608_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00609_, _00608_, _00607_);
  and (_39569_, _00609_, _42003_);
  and (_00610_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00611_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00612_, _00611_, _00610_);
  and (_39570_, _00612_, _42003_);
  and (_00613_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00614_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00615_, _00614_, _00613_);
  and (_39572_, _00615_, _42003_);
  and (_00616_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00617_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00618_, _00617_, _00616_);
  and (_39573_, _00618_, _42003_);
  and (_00619_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00620_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00621_, _00620_, _00619_);
  and (_39574_, _00621_, _42003_);
  and (_00622_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00623_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00624_, _00623_, _00622_);
  and (_39575_, _00624_, _42003_);
  and (_00625_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00626_, _44090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00627_, _00626_, _00625_);
  and (_39576_, _00627_, _42003_);
  and (_00628_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00629_, _40567_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00630_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00631_, _00630_, _44089_);
  and (_00632_, _00631_, _00629_);
  or (_00633_, _00632_, _00628_);
  and (_39577_, _00633_, _42003_);
  and (_00634_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00635_, _40752_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00636_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00637_, _00636_, _44089_);
  and (_00638_, _00637_, _00635_);
  or (_00639_, _00638_, _00634_);
  and (_39578_, _00639_, _42003_);
  and (_00640_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00641_, _40672_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00642_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00643_, _00642_, _44089_);
  and (_00644_, _00643_, _00641_);
  or (_00645_, _00644_, _00640_);
  and (_39579_, _00645_, _42003_);
  and (_00646_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00647_, _40551_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00648_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00649_, _00648_, _44089_);
  and (_00650_, _00649_, _00647_);
  or (_00651_, _00650_, _00646_);
  and (_39580_, _00651_, _42003_);
  and (_00652_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00653_, _40697_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00654_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00655_, _00654_, _44089_);
  and (_00656_, _00655_, _00653_);
  or (_00657_, _00656_, _00652_);
  and (_39581_, _00657_, _42003_);
  and (_00658_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00659_, _40611_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00660_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00661_, _00660_, _44089_);
  and (_00662_, _00661_, _00659_);
  or (_00663_, _00662_, _00658_);
  and (_39583_, _00663_, _42003_);
  and (_00664_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00665_, _40814_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00666_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00667_, _00666_, _44089_);
  and (_00668_, _00667_, _00665_);
  or (_00669_, _00668_, _00664_);
  and (_39584_, _00669_, _42003_);
  and (_00670_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00671_, _40474_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00672_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00673_, _00672_, _44089_);
  and (_00674_, _00673_, _00671_);
  or (_00675_, _00674_, _00670_);
  and (_39585_, _00675_, _42003_);
  and (_00676_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00677_, _00676_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00678_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _44089_);
  and (_00679_, _00678_, _42003_);
  and (_39586_, _00679_, _00677_);
  and (_00680_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00681_, _00680_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00682_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _44089_);
  and (_00683_, _00682_, _42003_);
  and (_39587_, _00683_, _00681_);
  and (_00684_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00685_, _00684_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00686_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _44089_);
  and (_00687_, _00686_, _42003_);
  and (_39588_, _00687_, _00685_);
  and (_00688_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00689_, _00688_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00690_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _44089_);
  and (_00691_, _00690_, _42003_);
  and (_39589_, _00691_, _00689_);
  and (_00692_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00693_, _00692_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00694_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _44089_);
  and (_00695_, _00694_, _42003_);
  and (_39590_, _00695_, _00693_);
  and (_00696_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00697_, _00696_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00698_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _44089_);
  and (_00699_, _00698_, _42003_);
  and (_39591_, _00699_, _00697_);
  and (_00700_, _44096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00701_, _00700_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00702_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _44089_);
  and (_00703_, _00702_, _42003_);
  and (_39592_, _00703_, _00701_);
  nand (_00704_, _44103_, _29288_);
  or (_00705_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00706_, _00705_, _42003_);
  and (_39594_, _00706_, _00704_);
  nand (_00707_, _44103_, _29961_);
  or (_00708_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00709_, _00708_, _42003_);
  and (_39595_, _00709_, _00707_);
  nand (_00710_, _44103_, _30656_);
  or (_00711_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00712_, _00711_, _42003_);
  and (_39596_, _00712_, _00710_);
  nand (_00713_, _44103_, _31416_);
  or (_00714_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00715_, _00714_, _42003_);
  and (_39597_, _00715_, _00713_);
  nand (_00716_, _44103_, _32133_);
  or (_00717_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00718_, _00717_, _42003_);
  and (_39598_, _00718_, _00716_);
  nand (_00719_, _44103_, _32943_);
  or (_00720_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00721_, _00720_, _42003_);
  and (_39599_, _00721_, _00719_);
  nand (_00722_, _44103_, _33677_);
  or (_00723_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00724_, _00723_, _42003_);
  and (_39600_, _00724_, _00722_);
  nand (_00725_, _44103_, _28122_);
  or (_00726_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00727_, _00726_, _42003_);
  and (_39601_, _00727_, _00725_);
  nand (_00728_, _44103_, _38828_);
  or (_00729_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00730_, _00729_, _42003_);
  and (_39602_, _00730_, _00728_);
  nand (_00731_, _44103_, _38856_);
  or (_00732_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00733_, _00732_, _42003_);
  and (_39603_, _00733_, _00731_);
  nand (_00734_, _44103_, _38884_);
  or (_00735_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00736_, _00735_, _42003_);
  and (_39605_, _00736_, _00734_);
  nand (_00737_, _44103_, _38913_);
  or (_00738_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00739_, _00738_, _42003_);
  and (_39606_, _00739_, _00737_);
  nand (_00740_, _44103_, _38941_);
  or (_00741_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00742_, _00741_, _42003_);
  and (_39607_, _00742_, _00740_);
  nand (_00743_, _44103_, _38970_);
  or (_00744_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00745_, _00744_, _42003_);
  and (_39608_, _00745_, _00743_);
  nand (_00746_, _44103_, _38996_);
  or (_00747_, _44103_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00748_, _00747_, _42003_);
  and (_39609_, _00748_, _00746_);
  nor (_39816_, _40513_, rst);
  nor (_00749_, _40556_, _40723_);
  and (_00750_, _00749_, _40639_);
  nor (_00751_, _40836_, _40501_);
  and (_00752_, _00751_, _00750_);
  not (_00753_, _40676_);
  nor (_00754_, _39303_, _39287_);
  and (_00755_, _39303_, _39287_);
  nor (_00756_, _00755_, _00754_);
  and (_00757_, _39276_, _39264_);
  nor (_00758_, _39276_, _39264_);
  or (_00759_, _00758_, _00757_);
  nor (_00760_, _00759_, _00756_);
  and (_00761_, _00759_, _00756_);
  nor (_00762_, _00761_, _00760_);
  nor (_00763_, _39325_, _39314_);
  and (_00764_, _39325_, _39314_);
  nor (_00765_, _00764_, _00763_);
  not (_00766_, _39252_);
  nor (_00767_, _39336_, _00766_);
  and (_00768_, _39336_, _00766_);
  nor (_00769_, _00768_, _00767_);
  nor (_00770_, _00769_, _00765_);
  and (_00771_, _00769_, _00765_);
  or (_00772_, _00771_, _00770_);
  or (_00773_, _00772_, _00762_);
  nand (_00774_, _00772_, _00762_);
  and (_00775_, _00774_, _00773_);
  or (_00776_, _00775_, _00753_);
  and (_00777_, _40591_, _40763_);
  or (_00778_, _40676_, _39168_);
  and (_00779_, _00778_, _00777_);
  and (_00780_, _00779_, _00776_);
  or (_00781_, _00753_, _39081_);
  not (_00782_, _40591_);
  and (_00783_, _00782_, _40763_);
  or (_00784_, _40676_, _39176_);
  and (_00785_, _00784_, _00783_);
  and (_00786_, _00785_, _00781_);
  nor (_00787_, _40591_, _40763_);
  and (_00788_, _00787_, _40676_);
  and (_00789_, _00788_, _39157_);
  and (_00790_, _00787_, _00753_);
  and (_00791_, _00790_, _39069_);
  or (_00792_, _00791_, _00789_);
  or (_00793_, _00792_, _00786_);
  or (_00794_, _00753_, _39141_);
  nor (_00795_, _00782_, _40763_);
  or (_00796_, _40676_, _39223_);
  and (_00797_, _00796_, _00795_);
  and (_00798_, _00797_, _00794_);
  or (_00799_, _00798_, _00793_);
  or (_00800_, _00799_, _00780_);
  and (_00801_, _00800_, _00752_);
  and (_00802_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_00803_, _00802_, _00753_);
  and (_00804_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00805_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_00806_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_00807_, _00806_, _00805_);
  or (_00808_, _00807_, _00804_);
  or (_00809_, _00808_, _00803_);
  and (_00810_, _40836_, _40640_);
  not (_00811_, _40501_);
  and (_00812_, _40723_, _00811_);
  and (_00813_, _00812_, _40556_);
  and (_00814_, _00813_, _00810_);
  and (_00815_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_00816_, _00815_, _40676_);
  and (_00817_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_00818_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00819_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_00820_, _00819_, _00818_);
  or (_00821_, _00820_, _00817_);
  or (_00822_, _00821_, _00816_);
  and (_00823_, _00822_, _00814_);
  and (_00824_, _00823_, _00809_);
  and (_00825_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_00826_, _00825_, _40676_);
  and (_00827_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_00828_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_00829_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_00830_, _00829_, _00828_);
  or (_00831_, _00830_, _00827_);
  or (_00832_, _00831_, _00826_);
  and (_00833_, _40836_, _40639_);
  and (_00834_, _00833_, _00812_);
  and (_00835_, _00834_, _40556_);
  and (_00836_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_00837_, _00836_, _00753_);
  and (_00838_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_00839_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_00840_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_00841_, _00840_, _00839_);
  or (_00842_, _00841_, _00838_);
  or (_00843_, _00842_, _00837_);
  and (_00844_, _00843_, _00835_);
  and (_00845_, _00844_, _00832_);
  and (_00846_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00847_, _00846_, _00753_);
  and (_00848_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00849_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00850_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00851_, _00850_, _00849_);
  or (_00852_, _00851_, _00848_);
  or (_00853_, _00852_, _00847_);
  nor (_00854_, _40836_, _40639_);
  and (_00855_, _00812_, _40555_);
  and (_00856_, _00855_, _00854_);
  and (_00857_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00858_, _00857_, _40676_);
  and (_00859_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00860_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00861_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00862_, _00861_, _00860_);
  or (_00863_, _00862_, _00859_);
  or (_00864_, _00863_, _00858_);
  and (_00865_, _00864_, _00856_);
  and (_00866_, _00865_, _00853_);
  or (_00867_, _00866_, _00845_);
  or (_00868_, _00867_, _00824_);
  and (_00869_, _00749_, _00811_);
  and (_00871_, _00869_, _00854_);
  and (_00872_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00873_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00874_, _00873_, _00872_);
  and (_00875_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00876_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00877_, _00876_, _00875_);
  or (_00878_, _00877_, _00874_);
  and (_00879_, _00878_, _40676_);
  and (_00880_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00881_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_00882_, _00881_, _00880_);
  and (_00883_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_00884_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00885_, _00884_, _00883_);
  or (_00886_, _00885_, _00882_);
  and (_00887_, _00886_, _00753_);
  or (_00888_, _00887_, _00879_);
  and (_00889_, _00888_, _00871_);
  and (_00890_, _34872_, _42645_);
  not (_00891_, _00890_);
  nor (_00892_, _42646_, _37146_);
  and (_00893_, _00892_, _00891_);
  nor (_00894_, _37245_, _37190_);
  and (_00895_, _00894_, _00893_);
  nor (_00896_, _42711_, _42644_);
  and (_00897_, _00896_, _00895_);
  nor (_00898_, _42714_, _35918_);
  and (_00899_, _36696_, _37749_);
  not (_00900_, _00899_);
  and (_00902_, _00900_, _00898_);
  and (_00903_, _00902_, _43013_);
  and (_00904_, _00903_, _00897_);
  and (_00905_, _00904_, _37463_);
  nor (_00906_, _00905_, _33896_);
  and (_00907_, _43193_, p2in_reg[6]);
  and (_00908_, _43189_, p2_in[6]);
  or (_00909_, _00908_, _00907_);
  or (_00910_, _00909_, _00906_);
  not (_00911_, _00906_);
  or (_00912_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_00913_, _00912_, _00910_);
  and (_00914_, _00913_, _00795_);
  or (_00915_, _00914_, _40676_);
  and (_00916_, _43193_, p2in_reg[7]);
  and (_00917_, _43189_, p2_in[7]);
  or (_00918_, _00917_, _00916_);
  or (_00919_, _00918_, _00906_);
  nand (_00920_, _00906_, _39380_);
  and (_00921_, _00920_, _00919_);
  and (_00923_, _00921_, _00787_);
  and (_00924_, _43193_, p2in_reg[4]);
  and (_00925_, _43189_, p2_in[4]);
  or (_00926_, _00925_, _00924_);
  or (_00927_, _00926_, _00906_);
  or (_00928_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00929_, _00928_, _00927_);
  and (_00930_, _00929_, _00777_);
  and (_00931_, _43193_, p2in_reg[5]);
  and (_00932_, _43189_, p2_in[5]);
  or (_00933_, _00932_, _00931_);
  or (_00934_, _00933_, _00906_);
  or (_00935_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00936_, _00935_, _00934_);
  and (_00937_, _00936_, _00783_);
  or (_00938_, _00937_, _00930_);
  or (_00939_, _00938_, _00923_);
  or (_00940_, _00939_, _00915_);
  and (_00941_, _00855_, _00810_);
  and (_00942_, _43193_, p2in_reg[2]);
  and (_00943_, _43189_, p2_in[2]);
  or (_00944_, _00943_, _00942_);
  or (_00945_, _00944_, _00906_);
  nand (_00946_, _00906_, _39805_);
  and (_00947_, _00946_, _00945_);
  and (_00948_, _00947_, _00795_);
  or (_00949_, _00948_, _00753_);
  and (_00950_, _43193_, p2in_reg[3]);
  and (_00951_, _43189_, p2_in[3]);
  or (_00952_, _00951_, _00950_);
  or (_00953_, _00952_, _00906_);
  or (_00954_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00955_, _00954_, _00953_);
  and (_00956_, _00955_, _00787_);
  and (_00957_, _43193_, p2in_reg[0]);
  and (_00958_, _43189_, p2_in[0]);
  or (_00959_, _00958_, _00957_);
  or (_00960_, _00959_, _00906_);
  or (_00961_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_00962_, _00961_, _00960_);
  and (_00963_, _00962_, _00777_);
  and (_00964_, _43193_, p2in_reg[1]);
  and (_00965_, _43189_, p2_in[1]);
  or (_00966_, _00965_, _00964_);
  or (_00967_, _00966_, _00906_);
  or (_00968_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_00969_, _00968_, _00967_);
  and (_00970_, _00969_, _00783_);
  or (_00971_, _00970_, _00963_);
  or (_00972_, _00971_, _00956_);
  or (_00973_, _00972_, _00949_);
  and (_00974_, _00973_, _00941_);
  and (_00975_, _00974_, _00940_);
  or (_00976_, _00975_, _00889_);
  nor (_00977_, _40555_, _40501_);
  and (_00978_, _40836_, _40724_);
  and (_00979_, _00978_, _00977_);
  and (_00980_, _00979_, _40640_);
  and (_00981_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_00982_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_00983_, _00982_, _00981_);
  and (_00984_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00985_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_00986_, _00985_, _00984_);
  or (_00987_, _00986_, _00983_);
  and (_00988_, _00987_, _40676_);
  and (_00989_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_00990_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_00991_, _00990_, _00989_);
  and (_00992_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00993_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _00991_);
  and (_00996_, _00995_, _00753_);
  or (_00997_, _00996_, _00988_);
  and (_00998_, _00997_, _00980_);
  and (_00999_, _43193_, p1in_reg[5]);
  and (_01000_, _43189_, p1_in[5]);
  or (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00906_);
  or (_01003_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01004_, _01003_, _01002_);
  and (_01005_, _01004_, _00783_);
  or (_01006_, _01005_, _40676_);
  and (_01007_, _43193_, p1in_reg[7]);
  and (_01008_, _43189_, p1_in[7]);
  or (_01009_, _01008_, _01007_);
  or (_01010_, _01009_, _00906_);
  nand (_01011_, _00906_, _39361_);
  and (_01012_, _01011_, _01010_);
  and (_01013_, _01012_, _00787_);
  and (_01014_, _43193_, p1in_reg[4]);
  and (_01015_, _43189_, p1_in[4]);
  or (_01016_, _01015_, _01014_);
  or (_01017_, _01016_, _00906_);
  or (_01018_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01019_, _01018_, _01017_);
  and (_01020_, _01019_, _00777_);
  and (_01021_, _43193_, p1in_reg[6]);
  and (_01022_, _43189_, p1_in[6]);
  or (_01023_, _01022_, _01021_);
  or (_01024_, _01023_, _00906_);
  or (_01025_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01026_, _01025_, _01024_);
  and (_01027_, _01026_, _00795_);
  or (_01028_, _01027_, _01020_);
  or (_01029_, _01028_, _01013_);
  or (_01030_, _01029_, _01006_);
  and (_01031_, _00869_, _00833_);
  and (_01032_, _43193_, p1in_reg[1]);
  and (_01033_, _43189_, p1_in[1]);
  or (_01034_, _01033_, _01032_);
  or (_01035_, _01034_, _00906_);
  or (_01036_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_01037_, _01036_, _01035_);
  and (_01038_, _01037_, _00783_);
  or (_01039_, _01038_, _00753_);
  and (_01040_, _43193_, p1in_reg[3]);
  and (_01041_, _43189_, p1_in[3]);
  or (_01042_, _01041_, _01040_);
  or (_01043_, _01042_, _00906_);
  or (_01044_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_01045_, _01044_, _01043_);
  and (_01046_, _01045_, _00787_);
  and (_01047_, _43193_, p1in_reg[0]);
  and (_01048_, _43189_, p1_in[0]);
  or (_01049_, _01048_, _01047_);
  or (_01050_, _01049_, _00906_);
  or (_01051_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01052_, _01051_, _01050_);
  and (_01053_, _01052_, _00777_);
  and (_01054_, _43193_, p1in_reg[2]);
  and (_01055_, _43189_, p1_in[2]);
  or (_01056_, _01055_, _01054_);
  or (_01057_, _01056_, _00906_);
  nand (_01058_, _00906_, _39721_);
  and (_01059_, _01058_, _01057_);
  and (_01060_, _01059_, _00795_);
  or (_01061_, _01060_, _01053_);
  or (_01062_, _01061_, _01046_);
  or (_01063_, _01062_, _01039_);
  and (_01064_, _01063_, _01031_);
  and (_01065_, _01064_, _01030_);
  or (_01066_, _01065_, _00998_);
  or (_01067_, _01066_, _00976_);
  and (_01068_, _00813_, _40836_);
  nor (_01069_, _01068_, _00752_);
  nor (_01070_, _00979_, _00871_);
  and (_01071_, _01070_, _01069_);
  nor (_01072_, _40556_, _40501_);
  and (_01073_, _01072_, _40836_);
  nor (_01074_, _01073_, _00856_);
  and (_01075_, _01074_, _01071_);
  nand (_01076_, _43295_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_01077_, _01076_, _01075_);
  and (_01078_, _43193_, p0in_reg[6]);
  and (_01079_, _43189_, p0_in[6]);
  or (_01080_, _01079_, _01078_);
  or (_01081_, _01080_, _00906_);
  or (_01082_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01083_, _01082_, _01081_);
  and (_01084_, _01083_, _00795_);
  or (_01085_, _01084_, _40676_);
  and (_01086_, _43193_, p0in_reg[7]);
  and (_01087_, _43189_, p0_in[7]);
  or (_01088_, _01087_, _01086_);
  or (_01089_, _01088_, _00906_);
  nand (_01090_, _00906_, _39347_);
  and (_01091_, _01090_, _01089_);
  and (_01092_, _01091_, _00787_);
  and (_01093_, _43193_, p0in_reg[5]);
  and (_01094_, _43189_, p0_in[5]);
  or (_01095_, _01094_, _01093_);
  or (_01096_, _01095_, _00906_);
  or (_01097_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01098_, _01097_, _01096_);
  and (_01099_, _01098_, _00783_);
  and (_01100_, _43193_, p0in_reg[4]);
  and (_01101_, _43189_, p0_in[4]);
  or (_01102_, _01101_, _01100_);
  or (_01103_, _01102_, _00906_);
  or (_01104_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01105_, _01104_, _01103_);
  and (_01106_, _01105_, _00777_);
  or (_01107_, _01106_, _01099_);
  or (_01108_, _01107_, _01092_);
  or (_01109_, _01108_, _01085_);
  and (_01110_, _00834_, _40555_);
  and (_01111_, _43193_, p0in_reg[2]);
  and (_01112_, _43189_, p0_in[2]);
  or (_01113_, _01112_, _01111_);
  or (_01114_, _01113_, _00906_);
  nand (_01115_, _00906_, _39635_);
  and (_01116_, _01115_, _01114_);
  and (_01117_, _01116_, _00795_);
  or (_01118_, _01117_, _00753_);
  and (_01119_, _43193_, p0in_reg[3]);
  and (_01120_, _43189_, p0_in[3]);
  or (_01121_, _01120_, _01119_);
  or (_01122_, _01121_, _00906_);
  nand (_01123_, _00906_, _39639_);
  and (_01124_, _01123_, _01122_);
  and (_01125_, _01124_, _00787_);
  and (_01126_, _43193_, p0in_reg[1]);
  and (_01127_, _43189_, p0_in[1]);
  or (_01128_, _01127_, _01126_);
  or (_01129_, _01128_, _00906_);
  or (_01130_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01131_, _01130_, _01129_);
  and (_01132_, _01131_, _00783_);
  and (_01133_, _43193_, p0in_reg[0]);
  and (_01134_, _43189_, p0_in[0]);
  or (_01135_, _01134_, _01133_);
  or (_01136_, _01135_, _00906_);
  nand (_01137_, _00906_, _39494_);
  and (_01138_, _01137_, _01136_);
  and (_01139_, _01138_, _00777_);
  or (_01140_, _01139_, _01132_);
  or (_01141_, _01140_, _01125_);
  or (_01142_, _01141_, _01118_);
  and (_01143_, _01142_, _01110_);
  and (_01144_, _01143_, _01109_);
  and (_01145_, _43193_, p3in_reg[1]);
  and (_01146_, _43189_, p3_in[1]);
  or (_01147_, _01146_, _01145_);
  or (_01148_, _01147_, _00906_);
  or (_01149_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01150_, _01149_, _01148_);
  and (_01151_, _01150_, _00783_);
  or (_01152_, _01151_, _00753_);
  and (_01153_, _43193_, p3in_reg[3]);
  and (_01154_, _43189_, p3_in[3]);
  or (_01155_, _01154_, _01153_);
  or (_01156_, _01155_, _00906_);
  or (_01157_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_01158_, _01157_, _01156_);
  and (_01159_, _01158_, _00787_);
  and (_01160_, _43193_, p3in_reg[2]);
  and (_01161_, _43189_, p3_in[2]);
  or (_01162_, _01161_, _01160_);
  or (_01163_, _01162_, _00906_);
  nand (_01164_, _00906_, _39895_);
  and (_01165_, _01164_, _01163_);
  and (_01166_, _01165_, _00795_);
  and (_01167_, _43193_, p3in_reg[0]);
  and (_01168_, _43189_, p3_in[0]);
  or (_01169_, _01168_, _01167_);
  or (_01170_, _01169_, _00906_);
  or (_01171_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01172_, _01171_, _01170_);
  and (_01173_, _01172_, _00777_);
  or (_01174_, _01173_, _01166_);
  or (_01175_, _01174_, _01159_);
  or (_01176_, _01175_, _01152_);
  and (_01177_, _00869_, _00810_);
  and (_01178_, _43193_, p3in_reg[5]);
  and (_01179_, _43189_, p3_in[5]);
  or (_01180_, _01179_, _01178_);
  or (_01181_, _01180_, _00906_);
  or (_01182_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01183_, _01182_, _01181_);
  and (_01184_, _01183_, _00783_);
  or (_01185_, _01184_, _40676_);
  and (_01186_, _43193_, p3in_reg[7]);
  and (_01187_, _43189_, p3_in[7]);
  or (_01188_, _01187_, _01186_);
  or (_01189_, _01188_, _00906_);
  nand (_01190_, _00906_, _39414_);
  and (_01191_, _01190_, _01189_);
  and (_01192_, _01191_, _00787_);
  and (_01193_, _43193_, p3in_reg[6]);
  and (_01194_, _43189_, p3_in[6]);
  or (_01195_, _01194_, _01193_);
  or (_01196_, _01195_, _00906_);
  or (_01197_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_01198_, _01197_, _01196_);
  and (_01199_, _01198_, _00795_);
  and (_01200_, _43193_, p3in_reg[4]);
  and (_01201_, _43189_, p3_in[4]);
  or (_01202_, _01201_, _01200_);
  or (_01203_, _01202_, _00906_);
  or (_01204_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01205_, _01204_, _01203_);
  and (_01206_, _01205_, _00777_);
  or (_01207_, _01206_, _01199_);
  or (_01208_, _01207_, _01192_);
  or (_01209_, _01208_, _01185_);
  and (_01210_, _01209_, _01177_);
  and (_01211_, _01210_, _01176_);
  nor (_01212_, _01211_, _01144_);
  nand (_01213_, _01212_, _01077_);
  or (_01214_, _01213_, _01067_);
  or (_01215_, _01214_, _00868_);
  or (_01216_, _01215_, _00801_);
  and (_01217_, _00856_, _39228_);
  nor (_01218_, _01077_, _29375_);
  nor (_01219_, _01218_, _01217_);
  and (_01220_, _01219_, _01216_);
  and (_01221_, _00790_, _39252_);
  and (_01222_, _00783_, _39325_);
  or (_01223_, _01222_, _40676_);
  and (_01224_, _00777_, _39314_);
  and (_01225_, _00795_, _39336_);
  or (_01226_, _01225_, _01224_);
  or (_01227_, _01226_, _01223_);
  and (_01228_, _00795_, _39287_);
  and (_01229_, _00783_, _39276_);
  or (_01230_, _01229_, _00753_);
  or (_01231_, _01230_, _01228_);
  and (_01232_, _00777_, _39264_);
  not (_01233_, _00787_);
  nor (_01234_, _01233_, _39303_);
  or (_01235_, _01234_, _01232_);
  or (_01236_, _01235_, _01231_);
  and (_01237_, _01236_, _01227_);
  or (_01238_, _01237_, _01221_);
  and (_01239_, _01238_, _01217_);
  not (_01240_, _01075_);
  not (_01241_, _39056_);
  and (_01242_, _01073_, _00911_);
  nor (_01243_, _01242_, _01241_);
  and (_01244_, _01243_, _43216_);
  and (_01245_, _01244_, _01240_);
  or (_01246_, _01245_, _01239_);
  or (_01247_, _01246_, _01220_);
  and (_01248_, _00783_, _40750_);
  or (_01249_, _01248_, _00753_);
  and (_01250_, _00795_, _40670_);
  and (_01251_, _00787_, _40549_);
  and (_01252_, _00777_, _38629_);
  or (_01253_, _01252_, _01251_);
  or (_01254_, _01253_, _01250_);
  or (_01255_, _01254_, _01249_);
  and (_01256_, _00783_, _40601_);
  or (_01257_, _01256_, _40676_);
  and (_01258_, _00795_, _40812_);
  and (_01259_, _00787_, _40472_);
  and (_01260_, _00777_, _40695_);
  or (_01261_, _01260_, _01259_);
  or (_01262_, _01261_, _01258_);
  or (_01263_, _01262_, _01257_);
  nand (_01264_, _01263_, _01255_);
  nand (_01265_, _01264_, _01245_);
  and (_01266_, _01265_, _42003_);
  and (_39847_, _01266_, _01247_);
  and (_01267_, _00777_, _40676_);
  and (_01268_, _01267_, _00752_);
  and (_01269_, _01268_, _39061_);
  and (_01270_, _01110_, _00788_);
  and (_01271_, _01270_, _38702_);
  nor (_01272_, _01271_, _01269_);
  nor (_01273_, _01272_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01274_, _00790_);
  and (_01275_, _01274_, _39045_);
  and (_01276_, _01275_, _43216_);
  and (_01277_, _01267_, _00856_);
  and (_01278_, _01277_, _39243_);
  or (_01279_, _01278_, _43297_);
  or (_01280_, _01279_, _01276_);
  or (_01281_, _01280_, _01273_);
  and (_01282_, _40555_, _40676_);
  and (_01283_, _01282_, _00795_);
  and (_01284_, _01283_, _00834_);
  and (_01285_, _01284_, _38702_);
  nor (_01286_, _01285_, rst);
  and (_39848_, _01286_, _01281_);
  not (_01287_, _01285_);
  and (_01288_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01289_, _40836_, _00811_);
  nor (_01290_, _40723_, _40639_);
  and (_01291_, _01290_, _01289_);
  and (_01292_, _01267_, _40556_);
  and (_01293_, _01292_, _01291_);
  and (_01294_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01295_, _01294_, _01288_);
  and (_01296_, _01292_, _00834_);
  and (_01297_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01298_, _00810_, _00812_);
  and (_01299_, _01292_, _01298_);
  and (_01300_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01301_, _01300_, _01297_);
  or (_01302_, _01301_, _01295_);
  and (_01303_, _01282_, _00777_);
  and (_01304_, _01290_, _00751_);
  and (_01305_, _01304_, _01303_);
  and (_01306_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01307_, _01282_, _00787_);
  and (_01308_, _01307_, _00834_);
  and (_01309_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01310_, _01309_, _01306_);
  and (_01311_, _01282_, _00783_);
  and (_01312_, _01311_, _00834_);
  and (_01313_, _01312_, _38653_);
  and (_01314_, _01291_, _01303_);
  and (_01315_, _01314_, _01191_);
  or (_01316_, _01315_, _01313_);
  or (_01317_, _01316_, _01310_);
  or (_01318_, _01317_, _01302_);
  and (_01319_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01320_, _01303_, _01298_);
  and (_01321_, _01320_, _00921_);
  and (_01322_, _40724_, _40639_);
  and (_01323_, _01289_, _01322_);
  and (_01324_, _01323_, _01303_);
  and (_01325_, _01324_, _01012_);
  or (_01326_, _01325_, _01321_);
  and (_01327_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01328_, _01303_, _00834_);
  and (_01329_, _01328_, _01091_);
  or (_01330_, _01329_, _01327_);
  or (_01331_, _01330_, _01326_);
  or (_01332_, _01331_, _01319_);
  nor (_01333_, _01332_, _01318_);
  nor (_01334_, _01333_, _01281_);
  and (_01335_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_01336_, _01335_, _01334_);
  and (_01337_, _01336_, _01287_);
  nor (_01338_, _01287_, _28122_);
  or (_01339_, _01338_, _01337_);
  and (_39849_, _01339_, _42003_);
  and (_01340_, _01268_, _00775_);
  and (_01341_, _01267_, _00835_);
  and (_01342_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01343_, _01267_, _00814_);
  and (_01344_, _01343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01345_, _01267_, _01110_);
  and (_01346_, _01345_, _01138_);
  or (_01347_, _01346_, _01344_);
  or (_01348_, _01347_, _01342_);
  and (_01349_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01350_, _01320_, _00962_);
  and (_01351_, _01303_, _01322_);
  and (_01352_, _01351_, _01289_);
  and (_01353_, _01352_, _01052_);
  or (_01354_, _01353_, _01350_);
  or (_01355_, _01354_, _01349_);
  and (_01356_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01357_, _01314_, _01172_);
  or (_01358_, _01357_, _01356_);
  and (_01359_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01360_, _01312_, _40587_);
  or (_01361_, _01360_, _01359_);
  or (_01362_, _01361_, _01358_);
  and (_01363_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01364_, _01270_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_01365_, _01364_, _01363_);
  or (_01366_, _01365_, _01362_);
  or (_01367_, _01366_, _01355_);
  or (_01368_, _01367_, _01348_);
  or (_01369_, _01368_, _01281_);
  or (_01370_, _01369_, _01340_);
  and (_01371_, _43295_, _25072_);
  and (_01372_, _01371_, _28155_);
  and (_01373_, _01274_, _43216_);
  and (_01374_, _01373_, _39045_);
  nor (_01375_, _01374_, _01372_);
  and (_01376_, _01277_, _39228_);
  and (_01377_, _01277_, _39225_);
  not (_01378_, _01377_);
  and (_01379_, _01378_, _01272_);
  nor (_01380_, _01379_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_01381_, _01380_, _01376_);
  and (_01382_, _01381_, _01375_);
  or (_01383_, _01382_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01384_, _01383_, _01370_);
  or (_01385_, _01384_, _01285_);
  nand (_01386_, _01285_, _29288_);
  and (_01387_, _01386_, _42003_);
  and (_39912_, _01387_, _01385_);
  and (_01388_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_01389_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_01390_, _01389_, _01388_);
  and (_01391_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01392_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01393_, _01392_, _01391_);
  or (_01394_, _01393_, _01390_);
  and (_01395_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01396_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_01397_, _01396_, _01395_);
  and (_01398_, _01312_, _40756_);
  and (_01399_, _01314_, _01150_);
  or (_01400_, _01399_, _01398_);
  or (_01401_, _01400_, _01397_);
  or (_01402_, _01401_, _01394_);
  and (_01403_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01404_, _01320_, _00969_);
  and (_01405_, _01324_, _01037_);
  or (_01406_, _01405_, _01404_);
  and (_01407_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01408_, _01328_, _01131_);
  or (_01409_, _01408_, _01407_);
  or (_01410_, _01409_, _01406_);
  or (_01411_, _01410_, _01403_);
  nor (_01412_, _01411_, _01402_);
  nor (_01413_, _01412_, _01281_);
  and (_01415_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_01417_, _01415_, _01413_);
  and (_01419_, _01417_, _01287_);
  nor (_01421_, _01287_, _29961_);
  or (_01423_, _01421_, _01419_);
  and (_39913_, _01423_, _42003_);
  and (_01426_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01427_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01428_, _01427_, _01426_);
  and (_01429_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01430_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01431_, _01430_, _01429_);
  or (_01432_, _01431_, _01428_);
  and (_01434_, _01314_, _01165_);
  and (_01435_, _01312_, _40660_);
  or (_01437_, _01435_, _01434_);
  and (_01438_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01439_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_01441_, _01439_, _01438_);
  or (_01442_, _01441_, _01437_);
  or (_01443_, _01442_, _01432_);
  and (_01445_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01446_, _01320_, _00947_);
  and (_01447_, _01324_, _01059_);
  or (_01449_, _01447_, _01446_);
  and (_01450_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01451_, _01328_, _01116_);
  or (_01453_, _01451_, _01450_);
  or (_01454_, _01453_, _01449_);
  or (_01455_, _01454_, _01445_);
  nor (_01457_, _01455_, _01443_);
  nor (_01458_, _01457_, _01281_);
  and (_01459_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_01461_, _01459_, _01458_);
  and (_01462_, _01461_, _01287_);
  nor (_01463_, _01287_, _30656_);
  or (_01465_, _01463_, _01462_);
  and (_39914_, _01465_, _42003_);
  and (_01466_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_01467_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01468_, _01467_, _01466_);
  and (_01469_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01470_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01471_, _01470_, _01469_);
  or (_01472_, _01471_, _01468_);
  and (_01473_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01474_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_01475_, _01474_, _01473_);
  and (_01476_, _01314_, _01158_);
  and (_01477_, _01312_, _40538_);
  or (_01478_, _01477_, _01476_);
  or (_01479_, _01478_, _01475_);
  or (_01480_, _01479_, _01472_);
  and (_01481_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01482_, _01320_, _00955_);
  and (_01483_, _01324_, _01045_);
  or (_01484_, _01483_, _01482_);
  and (_01486_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01487_, _01328_, _01124_);
  or (_01489_, _01487_, _01486_);
  or (_01490_, _01489_, _01484_);
  or (_01491_, _01490_, _01481_);
  nor (_01493_, _01491_, _01480_);
  nor (_01494_, _01493_, _01281_);
  and (_01495_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_01497_, _01495_, _01494_);
  and (_01498_, _01497_, _01287_);
  nor (_01499_, _01287_, _31416_);
  or (_01501_, _01499_, _01498_);
  and (_39915_, _01501_, _42003_);
  and (_01502_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_01504_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_01505_, _01504_, _01502_);
  and (_01506_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01508_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01509_, _01508_, _01506_);
  or (_01510_, _01509_, _01505_);
  and (_01512_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01513_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01514_, _01513_, _01512_);
  and (_01516_, _01312_, _40701_);
  and (_01517_, _01314_, _01205_);
  or (_01518_, _01517_, _01516_);
  or (_01519_, _01518_, _01514_);
  or (_01520_, _01519_, _01510_);
  and (_01521_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01522_, _01320_, _00929_);
  and (_01523_, _01324_, _01019_);
  or (_01524_, _01523_, _01522_);
  and (_01525_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01526_, _01328_, _01105_);
  or (_01527_, _01526_, _01525_);
  or (_01528_, _01527_, _01524_);
  or (_01529_, _01528_, _01521_);
  nor (_01530_, _01529_, _01520_);
  nor (_01531_, _01530_, _01281_);
  and (_01532_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_01533_, _01532_, _01531_);
  and (_01534_, _01533_, _01287_);
  nor (_01535_, _01287_, _32133_);
  or (_01536_, _01535_, _01534_);
  and (_39916_, _01536_, _42003_);
  and (_01538_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01540_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_01541_, _01540_, _01538_);
  and (_01542_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01544_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01545_, _01544_, _01542_);
  or (_01546_, _01545_, _01541_);
  and (_01548_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01549_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01550_, _01549_, _01548_);
  and (_01552_, _01312_, _40617_);
  and (_01553_, _01314_, _01183_);
  or (_01554_, _01553_, _01552_);
  or (_01556_, _01554_, _01550_);
  or (_01557_, _01556_, _01546_);
  and (_01558_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01560_, _01320_, _00936_);
  and (_01561_, _01324_, _01004_);
  or (_01562_, _01561_, _01560_);
  and (_01564_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01565_, _01328_, _01098_);
  or (_01566_, _01565_, _01564_);
  or (_01568_, _01566_, _01562_);
  or (_01569_, _01568_, _01558_);
  nor (_01570_, _01569_, _01557_);
  nor (_01571_, _01570_, _01281_);
  and (_01572_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_01573_, _01572_, _01571_);
  and (_01574_, _01573_, _01287_);
  nor (_01575_, _01287_, _32943_);
  or (_01576_, _01575_, _01574_);
  and (_39917_, _01576_, _42003_);
  and (_01577_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01578_, _01284_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_01579_, _01578_, _01577_);
  and (_01580_, _01296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01581_, _01299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01582_, _01581_, _01580_);
  or (_01583_, _01582_, _01579_);
  and (_01584_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01585_, _01308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01586_, _01585_, _01584_);
  and (_01587_, _01312_, _40802_);
  and (_01589_, _01314_, _01198_);
  or (_01590_, _01589_, _01587_);
  or (_01592_, _01590_, _01586_);
  or (_01593_, _01592_, _01583_);
  and (_01594_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01596_, _01320_, _00913_);
  and (_01597_, _01324_, _01026_);
  or (_01598_, _01597_, _01596_);
  and (_01600_, _01268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01601_, _01328_, _01083_);
  or (_01602_, _01601_, _01600_);
  or (_01604_, _01602_, _01598_);
  or (_01605_, _01604_, _01594_);
  nor (_01606_, _01605_, _01593_);
  nor (_01608_, _01606_, _01281_);
  and (_01609_, _01281_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_01610_, _01609_, _01608_);
  and (_01612_, _01610_, _01287_);
  nor (_01613_, _01287_, _33677_);
  or (_01614_, _01613_, _01612_);
  and (_39918_, _01614_, _42003_);
  and (_39962_, _40867_, _42003_);
  and (_39963_, _41049_, _42003_);
  nor (_39965_, _40676_, rst);
  and (_39981_, _41066_, _42003_);
  and (_39982_, _41079_, _42003_);
  and (_39983_, _41092_, _42003_);
  and (_39984_, _41100_, _42003_);
  and (_39985_, _41110_, _42003_);
  and (_39986_, _41121_, _42003_);
  and (_39987_, _41130_, _42003_);
  nor (_39988_, _40591_, rst);
  nor (_39989_, _40763_, rst);
  not (_01617_, _42059_);
  nor (_01618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01619_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01620_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01619_);
  nor (_01621_, _01620_, _01618_);
  nor (_01622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01623_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01619_);
  nor (_01624_, _01623_, _01622_);
  not (_01625_, _01624_);
  nor (_01626_, _01625_, _01621_);
  nor (_01628_, _01624_, _01621_);
  not (_01629_, _01628_);
  nor (_01631_, _00101_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01632_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01619_);
  nor (_01633_, _01632_, _01631_);
  and (_01635_, _01633_, _01629_);
  nor (_01636_, _00122_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01637_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01619_);
  nor (_01639_, _01637_, _01636_);
  nor (_01640_, _01633_, _01629_);
  or (_01641_, _01640_, _01639_);
  nor (_01643_, _01641_, _01635_);
  and (_01644_, _01643_, _01626_);
  and (_01645_, _01644_, _01617_);
  not (_01647_, _42100_);
  and (_01648_, _01624_, _01621_);
  and (_01649_, _01643_, _01648_);
  and (_01651_, _01649_, _01647_);
  or (_01652_, _01651_, _01645_);
  not (_01653_, _42018_);
  and (_01655_, _01625_, _01621_);
  and (_01656_, _01655_, _01643_);
  and (_01657_, _01656_, _01653_);
  not (_01659_, _41969_);
  not (_01660_, _01639_);
  and (_01661_, _01640_, _01660_);
  and (_01662_, _01661_, _01659_);
  or (_01663_, _01662_, _01657_);
  or (_01664_, _01663_, _01652_);
  not (_01665_, _41839_);
  nor (_01666_, _01660_, _01635_);
  not (_01667_, _01666_);
  and (_01668_, _01667_, _01641_);
  and (_01669_, _01655_, _01668_);
  and (_01670_, _01669_, _01665_);
  not (_01671_, _41880_);
  and (_01672_, _01668_, _01626_);
  and (_01673_, _01672_, _01671_);
  not (_01674_, _41921_);
  and (_01675_, _01668_, _01648_);
  and (_01676_, _01675_, _01674_);
  or (_01677_, _01676_, _01673_);
  or (_01678_, _01677_, _01670_);
  or (_01679_, _01678_, _01664_);
  not (_01681_, _42305_);
  and (_01682_, _01640_, _01639_);
  and (_01684_, _01682_, _01681_);
  not (_01685_, _42264_);
  and (_01686_, _01660_, _01633_);
  and (_01688_, _01686_, _01648_);
  and (_01689_, _01688_, _01685_);
  not (_01690_, _42223_);
  and (_01692_, _01686_, _01626_);
  and (_01693_, _01692_, _01690_);
  or (_01694_, _01693_, _01689_);
  not (_01696_, _42141_);
  and (_01697_, _01633_, _01628_);
  and (_01698_, _01697_, _01660_);
  and (_01700_, _01698_, _01696_);
  not (_01701_, _42182_);
  and (_01702_, _01686_, _01655_);
  and (_01704_, _01702_, _01701_);
  or (_01705_, _01704_, _01700_);
  or (_01706_, _01705_, _01694_);
  or (_01708_, _01706_, _01684_);
  not (_01709_, _42469_);
  and (_01710_, _01697_, _01639_);
  and (_01712_, _01710_, _01709_);
  not (_01713_, _42346_);
  and (_01714_, _01655_, _01666_);
  and (_01715_, _01714_, _01713_);
  not (_01716_, _42428_);
  and (_01717_, _01666_, _01648_);
  and (_01718_, _01717_, _01716_);
  not (_01719_, _42387_);
  and (_01720_, _01666_, _01626_);
  and (_01721_, _01720_, _01719_);
  or (_01722_, _01721_, _01718_);
  or (_01723_, _01722_, _01715_);
  or (_01724_, _01723_, _01712_);
  or (_01725_, _01724_, _01708_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01725_, _01679_);
  and (_01726_, _01669_, _01716_);
  and (_01727_, _01644_, _01659_);
  or (_01728_, _01727_, _01726_);
  and (_01729_, _01656_, _01674_);
  and (_01730_, _01649_, _01653_);
  or (_01731_, _01730_, _01729_);
  or (_01733_, _01731_, _01728_);
  and (_01734_, _01692_, _01696_);
  and (_01736_, _01714_, _01685_);
  or (_01737_, _01736_, _01734_);
  and (_01738_, _01720_, _01681_);
  and (_01740_, _01702_, _01647_);
  or (_01741_, _01740_, _01738_);
  or (_01742_, _01741_, _01737_);
  and (_01744_, _01710_, _01719_);
  and (_01745_, _01698_, _01617_);
  or (_01746_, _01745_, _01744_);
  and (_01748_, _01682_, _01690_);
  and (_01749_, _01661_, _01671_);
  or (_01750_, _01749_, _01748_);
  or (_01752_, _01750_, _01746_);
  and (_01753_, _01717_, _01713_);
  and (_01754_, _01688_, _01701_);
  or (_01756_, _01754_, _01753_);
  or (_01757_, _01756_, _01752_);
  and (_01758_, _01672_, _01709_);
  and (_01760_, _01675_, _01665_);
  or (_01761_, _01760_, _01758_);
  or (_01762_, _01761_, _01757_);
  or (_01764_, _01762_, _01742_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01764_, _01733_);
  and (_01765_, _01672_, _01665_);
  and (_01766_, _01656_, _01659_);
  or (_01767_, _01766_, _01765_);
  and (_01768_, _01649_, _01617_);
  and (_01769_, _01644_, _01653_);
  or (_01770_, _01769_, _01768_);
  or (_01771_, _01770_, _01767_);
  and (_01772_, _01692_, _01701_);
  and (_01773_, _01702_, _01696_);
  or (_01774_, _01773_, _01772_);
  and (_01775_, _01714_, _01681_);
  and (_01776_, _01688_, _01690_);
  or (_01777_, _01776_, _01775_);
  or (_01778_, _01777_, _01774_);
  and (_01779_, _01661_, _01674_);
  and (_01780_, _01698_, _01647_);
  or (_01781_, _01780_, _01779_);
  and (_01782_, _01710_, _01716_);
  and (_01783_, _01682_, _01685_);
  or (_01785_, _01783_, _01782_);
  or (_01786_, _01785_, _01781_);
  and (_01788_, _01717_, _01719_);
  and (_01789_, _01720_, _01713_);
  or (_01790_, _01789_, _01788_);
  or (_01792_, _01790_, _01786_);
  and (_01793_, _01669_, _01709_);
  and (_01794_, _01675_, _01671_);
  or (_01796_, _01794_, _01793_);
  or (_01797_, _01796_, _01792_);
  or (_01798_, _01797_, _01778_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01798_, _01771_);
  and (_01800_, _01672_, _01716_);
  and (_01801_, _01669_, _01719_);
  or (_01803_, _01801_, _01800_);
  and (_01804_, _01649_, _01659_);
  and (_01805_, _01656_, _01671_);
  or (_01807_, _01805_, _01804_);
  or (_01808_, _01807_, _01803_);
  and (_01809_, _01688_, _01696_);
  and (_01811_, _01720_, _01685_);
  or (_01812_, _01811_, _01809_);
  and (_01813_, _01714_, _01690_);
  and (_01815_, _01692_, _01647_);
  or (_01816_, _01815_, _01813_);
  or (_01817_, _01816_, _01812_);
  and (_01818_, _01710_, _01713_);
  and (_01819_, _01661_, _01665_);
  or (_01820_, _01819_, _01818_);
  and (_01821_, _01682_, _01701_);
  and (_01822_, _01698_, _01653_);
  or (_01823_, _01822_, _01821_);
  or (_01824_, _01823_, _01820_);
  and (_01825_, _01717_, _01681_);
  and (_01826_, _01702_, _01617_);
  or (_01827_, _01826_, _01825_);
  or (_01828_, _01827_, _01824_);
  and (_01829_, _01675_, _01709_);
  and (_01830_, _01644_, _01674_);
  or (_01831_, _01830_, _01829_);
  or (_01832_, _01831_, _01828_);
  or (_01833_, _01832_, _01817_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01833_, _01808_);
  not (_01834_, _42023_);
  and (_01836_, _01656_, _01834_);
  not (_01837_, _41885_);
  and (_01839_, _01672_, _01837_);
  or (_01840_, _01839_, _01836_);
  not (_01841_, _42064_);
  and (_01843_, _01644_, _01841_);
  not (_01844_, _41926_);
  and (_01845_, _01675_, _01844_);
  or (_01847_, _01845_, _01843_);
  or (_01848_, _01847_, _01840_);
  not (_01849_, _42433_);
  and (_01851_, _01717_, _01849_);
  not (_01852_, _42228_);
  and (_01853_, _01692_, _01852_);
  or (_01855_, _01853_, _01851_);
  not (_01856_, _42392_);
  and (_01857_, _01720_, _01856_);
  not (_01859_, _42187_);
  and (_01860_, _01702_, _01859_);
  or (_01861_, _01860_, _01857_);
  or (_01863_, _01861_, _01855_);
  not (_01864_, _42146_);
  and (_01865_, _01698_, _01864_);
  not (_01867_, _41974_);
  and (_01868_, _01661_, _01867_);
  or (_01869_, _01868_, _01865_);
  not (_01870_, _42474_);
  and (_01871_, _01710_, _01870_);
  not (_01872_, _42310_);
  and (_01873_, _01682_, _01872_);
  or (_01874_, _01873_, _01871_);
  or (_01875_, _01874_, _01869_);
  not (_01876_, _42351_);
  and (_01877_, _01714_, _01876_);
  not (_01878_, _42269_);
  and (_01879_, _01688_, _01878_);
  or (_01880_, _01879_, _01877_);
  or (_01881_, _01880_, _01875_);
  not (_01882_, _42105_);
  and (_01883_, _01649_, _01882_);
  not (_01884_, _41844_);
  and (_01885_, _01669_, _01884_);
  or (_01886_, _01885_, _01883_);
  or (_01887_, _01886_, _01881_);
  or (_01889_, _01887_, _01863_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01889_, _01848_);
  not (_01891_, _42069_);
  and (_01892_, _01644_, _01891_);
  not (_01893_, _42110_);
  and (_01895_, _01649_, _01893_);
  or (_01896_, _01895_, _01892_);
  not (_01897_, _41849_);
  and (_01899_, _01669_, _01897_);
  not (_01900_, _42028_);
  and (_01901_, _01656_, _01900_);
  or (_01903_, _01901_, _01899_);
  or (_01904_, _01903_, _01896_);
  not (_01905_, _42274_);
  and (_01907_, _01688_, _01905_);
  not (_01908_, _42233_);
  and (_01909_, _01692_, _01908_);
  or (_01911_, _01909_, _01907_);
  not (_01912_, _42397_);
  and (_01913_, _01720_, _01912_);
  not (_01915_, _42192_);
  and (_01916_, _01702_, _01915_);
  or (_01917_, _01916_, _01913_);
  or (_01919_, _01917_, _01911_);
  not (_01920_, _41890_);
  and (_01921_, _01672_, _01920_);
  not (_01922_, _41931_);
  and (_01923_, _01675_, _01922_);
  or (_01924_, _01923_, _01921_);
  not (_01925_, _42479_);
  and (_01926_, _01710_, _01925_);
  not (_01927_, _42315_);
  and (_01928_, _01682_, _01927_);
  or (_01929_, _01928_, _01926_);
  not (_01930_, _42151_);
  and (_01931_, _01698_, _01930_);
  not (_01932_, _41979_);
  and (_01933_, _01661_, _01932_);
  or (_01934_, _01933_, _01931_);
  or (_01935_, _01934_, _01929_);
  not (_01936_, _42438_);
  and (_01937_, _01717_, _01936_);
  not (_01938_, _42356_);
  and (_01939_, _01714_, _01938_);
  or (_01941_, _01939_, _01937_);
  or (_01942_, _01941_, _01935_);
  or (_01944_, _01942_, _01924_);
  or (_01945_, _01944_, _01919_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01945_, _01904_);
  not (_01947_, _42074_);
  and (_01948_, _01644_, _01947_);
  not (_01949_, _42033_);
  and (_01951_, _01656_, _01949_);
  or (_01952_, _01951_, _01948_);
  not (_01953_, _42115_);
  and (_01955_, _01649_, _01953_);
  not (_01956_, _41854_);
  and (_01957_, _01669_, _01956_);
  or (_01959_, _01957_, _01955_);
  or (_01960_, _01959_, _01952_);
  not (_01961_, _42279_);
  and (_01963_, _01688_, _01961_);
  not (_01964_, _42443_);
  and (_01965_, _01717_, _01964_);
  or (_01967_, _01965_, _01963_);
  not (_01968_, _42238_);
  and (_01969_, _01692_, _01968_);
  not (_01971_, _42402_);
  and (_01972_, _01720_, _01971_);
  or (_01973_, _01972_, _01969_);
  or (_01974_, _01973_, _01967_);
  not (_01975_, _41895_);
  and (_01976_, _01672_, _01975_);
  not (_01977_, _41936_);
  and (_01978_, _01675_, _01977_);
  or (_01979_, _01978_, _01976_);
  not (_01980_, _42484_);
  and (_01981_, _01710_, _01980_);
  not (_01982_, _41984_);
  and (_01983_, _01661_, _01982_);
  or (_01984_, _01983_, _01981_);
  not (_01985_, _42156_);
  and (_01986_, _01698_, _01985_);
  not (_01987_, _42320_);
  and (_01988_, _01682_, _01987_);
  or (_01989_, _01988_, _01986_);
  or (_01990_, _01989_, _01984_);
  not (_01991_, _42197_);
  and (_01993_, _01702_, _01991_);
  not (_01994_, _42361_);
  and (_01996_, _01714_, _01994_);
  or (_01997_, _01996_, _01993_);
  or (_01998_, _01997_, _01990_);
  or (_02000_, _01998_, _01979_);
  or (_02001_, _02000_, _01974_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02001_, _01960_);
  not (_02003_, _42038_);
  and (_02004_, _01656_, _02003_);
  not (_02005_, _41941_);
  and (_02007_, _01675_, _02005_);
  or (_02008_, _02007_, _02004_);
  not (_02009_, _41859_);
  and (_02011_, _01669_, _02009_);
  not (_02012_, _41900_);
  and (_02013_, _01672_, _02012_);
  or (_02015_, _02013_, _02011_);
  or (_02016_, _02015_, _02008_);
  not (_02017_, _42284_);
  and (_02019_, _01688_, _02017_);
  not (_02020_, _42243_);
  and (_02021_, _01692_, _02020_);
  or (_02023_, _02021_, _02019_);
  not (_02024_, _42407_);
  and (_02025_, _01720_, _02024_);
  not (_02026_, _42202_);
  and (_02027_, _01702_, _02026_);
  or (_02028_, _02027_, _02025_);
  or (_02029_, _02028_, _02023_);
  not (_02030_, _42120_);
  and (_02031_, _01649_, _02030_);
  not (_02032_, _42079_);
  and (_02033_, _01644_, _02032_);
  or (_02034_, _02033_, _02031_);
  not (_02035_, _42489_);
  and (_02036_, _01710_, _02035_);
  not (_02037_, _42325_);
  and (_02038_, _01682_, _02037_);
  or (_02039_, _02038_, _02036_);
  not (_02040_, _42161_);
  and (_02041_, _01698_, _02040_);
  not (_02042_, _41989_);
  and (_02043_, _01661_, _02042_);
  or (_02045_, _02043_, _02041_);
  or (_02046_, _02045_, _02039_);
  not (_02048_, _42448_);
  and (_02049_, _01717_, _02048_);
  not (_02050_, _42366_);
  and (_02052_, _01714_, _02050_);
  or (_02053_, _02052_, _02049_);
  or (_02054_, _02053_, _02046_);
  or (_02056_, _02054_, _02034_);
  or (_02057_, _02056_, _02029_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02057_, _02016_);
  not (_02059_, _42125_);
  and (_02060_, _01649_, _02059_);
  not (_02061_, _41947_);
  and (_02063_, _01675_, _02061_);
  or (_02064_, _02063_, _02060_);
  not (_02065_, _41864_);
  and (_02067_, _01669_, _02065_);
  not (_02068_, _41905_);
  and (_02069_, _01672_, _02068_);
  or (_02071_, _02069_, _02067_);
  or (_02072_, _02071_, _02064_);
  not (_02073_, _42412_);
  and (_02075_, _01720_, _02073_);
  not (_02076_, _42453_);
  and (_02077_, _01717_, _02076_);
  or (_02078_, _02077_, _02075_);
  not (_02079_, _42248_);
  and (_02080_, _01692_, _02079_);
  not (_02081_, _42207_);
  and (_02082_, _01702_, _02081_);
  or (_02083_, _02082_, _02080_);
  or (_02084_, _02083_, _02078_);
  not (_02085_, _42000_);
  and (_02086_, _01661_, _02085_);
  not (_02087_, _42330_);
  and (_02088_, _01682_, _02087_);
  or (_02089_, _02088_, _02086_);
  not (_02090_, _42494_);
  and (_02091_, _01710_, _02090_);
  not (_02092_, _42166_);
  and (_02093_, _01698_, _02092_);
  or (_02094_, _02093_, _02091_);
  or (_02095_, _02094_, _02089_);
  not (_02097_, _42289_);
  and (_02098_, _01688_, _02097_);
  not (_02100_, _42371_);
  and (_02101_, _01714_, _02100_);
  or (_02102_, _02101_, _02098_);
  or (_02104_, _02102_, _02095_);
  not (_02105_, _42084_);
  and (_02106_, _01644_, _02105_);
  not (_02108_, _42043_);
  and (_02109_, _01656_, _02108_);
  or (_02110_, _02109_, _02106_);
  or (_02112_, _02110_, _02104_);
  or (_02113_, _02112_, _02084_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02113_, _02072_);
  not (_02115_, _42048_);
  and (_02116_, _01656_, _02115_);
  not (_02117_, _41957_);
  and (_02119_, _01675_, _02117_);
  or (_02120_, _02119_, _02116_);
  not (_02121_, _42089_);
  and (_02123_, _01644_, _02121_);
  not (_02124_, _41910_);
  and (_02125_, _01672_, _02124_);
  or (_02127_, _02125_, _02123_);
  or (_02128_, _02127_, _02120_);
  not (_02129_, _42458_);
  and (_02130_, _01717_, _02129_);
  not (_02131_, _42253_);
  and (_02132_, _01692_, _02131_);
  or (_02133_, _02132_, _02130_);
  not (_02134_, _42417_);
  and (_02135_, _01720_, _02134_);
  not (_02136_, _42376_);
  and (_02137_, _01714_, _02136_);
  or (_02138_, _02137_, _02135_);
  or (_02139_, _02138_, _02133_);
  not (_02140_, _42335_);
  and (_02141_, _01682_, _02140_);
  not (_02142_, _42171_);
  and (_02143_, _01698_, _02142_);
  or (_02144_, _02143_, _02141_);
  not (_02145_, _42499_);
  and (_02146_, _01710_, _02145_);
  not (_02147_, _42007_);
  and (_02149_, _01661_, _02147_);
  or (_02150_, _02149_, _02146_);
  or (_02152_, _02150_, _02144_);
  not (_02153_, _42294_);
  and (_02154_, _01688_, _02153_);
  not (_02156_, _42212_);
  and (_02157_, _01702_, _02156_);
  or (_02158_, _02157_, _02154_);
  or (_02160_, _02158_, _02152_);
  not (_02161_, _42130_);
  and (_02162_, _01649_, _02161_);
  not (_02164_, _41869_);
  and (_02165_, _01669_, _02164_);
  or (_02166_, _02165_, _02162_);
  or (_02168_, _02166_, _02160_);
  or (_02169_, _02168_, _02139_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02169_, _02128_);
  not (_02171_, _41915_);
  and (_02172_, _01672_, _02171_);
  not (_02173_, _41963_);
  and (_02175_, _01675_, _02173_);
  or (_02176_, _02175_, _02172_);
  not (_02177_, _42094_);
  and (_02179_, _01644_, _02177_);
  not (_02180_, _41874_);
  and (_02181_, _01669_, _02180_);
  or (_02182_, _02181_, _02179_);
  or (_02183_, _02182_, _02176_);
  not (_02184_, _42299_);
  and (_02185_, _01688_, _02184_);
  not (_02186_, _42258_);
  and (_02187_, _01692_, _02186_);
  or (_02188_, _02187_, _02185_);
  not (_02189_, _42422_);
  and (_02190_, _01720_, _02189_);
  not (_02191_, _42217_);
  and (_02192_, _01702_, _02191_);
  or (_02193_, _02192_, _02190_);
  or (_02194_, _02193_, _02188_);
  not (_02195_, _42340_);
  and (_02196_, _01682_, _02195_);
  not (_02197_, _42176_);
  and (_02198_, _01698_, _02197_);
  or (_02199_, _02198_, _02196_);
  not (_02201_, _42504_);
  and (_02202_, _01710_, _02201_);
  not (_02204_, _42012_);
  and (_02205_, _01661_, _02204_);
  or (_02206_, _02205_, _02202_);
  or (_02208_, _02206_, _02199_);
  not (_02209_, _42463_);
  and (_02210_, _01717_, _02209_);
  not (_02212_, _42381_);
  and (_02213_, _01714_, _02212_);
  or (_02214_, _02213_, _02210_);
  or (_02216_, _02214_, _02208_);
  not (_02217_, _42135_);
  and (_02218_, _01649_, _02217_);
  not (_02220_, _42053_);
  and (_02221_, _01656_, _02220_);
  or (_02222_, _02221_, _02218_);
  or (_02224_, _02222_, _02216_);
  or (_02225_, _02224_, _02194_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02225_, _02183_);
  and (_02227_, _01656_, _01867_);
  and (_02228_, _01675_, _01837_);
  or (_02229_, _02228_, _02227_);
  and (_02231_, _01644_, _01834_);
  and (_02232_, _01672_, _01884_);
  or (_02233_, _02232_, _02231_);
  or (_02234_, _02233_, _02229_);
  and (_02235_, _01720_, _01876_);
  and (_02236_, _01688_, _01852_);
  or (_02237_, _02236_, _02235_);
  and (_02238_, _01717_, _01856_);
  and (_02239_, _01692_, _01859_);
  or (_02240_, _02239_, _02238_);
  or (_02241_, _02240_, _02237_);
  and (_02242_, _01714_, _01872_);
  and (_02243_, _01702_, _01864_);
  or (_02244_, _02243_, _02242_);
  and (_02245_, _01698_, _01882_);
  and (_02246_, _01661_, _01844_);
  or (_02247_, _02246_, _02245_);
  and (_02248_, _01710_, _01849_);
  and (_02249_, _01682_, _01878_);
  or (_02250_, _02249_, _02248_);
  or (_02251_, _02250_, _02247_);
  or (_02252_, _02251_, _02244_);
  and (_02253_, _01669_, _01870_);
  and (_02254_, _01649_, _01841_);
  or (_02255_, _02254_, _02253_);
  or (_02256_, _02255_, _02252_);
  or (_02257_, _02256_, _02241_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02257_, _02234_);
  and (_02258_, _01656_, _01932_);
  and (_02259_, _01675_, _01920_);
  or (_02260_, _02259_, _02258_);
  and (_02261_, _01644_, _01900_);
  and (_02262_, _01672_, _01897_);
  or (_02263_, _02262_, _02261_);
  or (_02264_, _02263_, _02260_);
  and (_02265_, _01720_, _01938_);
  and (_02266_, _01688_, _01908_);
  or (_02267_, _02266_, _02265_);
  and (_02268_, _01717_, _01912_);
  and (_02269_, _01692_, _01915_);
  or (_02270_, _02269_, _02268_);
  or (_02271_, _02270_, _02267_);
  and (_02272_, _01714_, _01927_);
  and (_02273_, _01702_, _01930_);
  or (_02274_, _02273_, _02272_);
  and (_02275_, _01698_, _01893_);
  and (_02276_, _01661_, _01922_);
  or (_02277_, _02276_, _02275_);
  and (_02278_, _01710_, _01936_);
  and (_02279_, _01682_, _01905_);
  or (_02280_, _02279_, _02278_);
  or (_02281_, _02280_, _02277_);
  or (_02282_, _02281_, _02274_);
  and (_02283_, _01669_, _01925_);
  and (_02284_, _01649_, _01891_);
  or (_02285_, _02284_, _02283_);
  or (_02286_, _02285_, _02282_);
  or (_02287_, _02286_, _02271_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02287_, _02264_);
  and (_02288_, _01669_, _01980_);
  and (_02289_, _01644_, _01949_);
  or (_02290_, _02289_, _02288_);
  and (_02291_, _01672_, _01956_);
  and (_02292_, _01675_, _01975_);
  or (_02293_, _02292_, _02291_);
  or (_02294_, _02293_, _02290_);
  and (_02295_, _01692_, _01991_);
  and (_02296_, _01720_, _01994_);
  or (_02297_, _02296_, _02295_);
  and (_02298_, _01717_, _01971_);
  and (_02299_, _01714_, _01987_);
  or (_02300_, _02299_, _02298_);
  or (_02301_, _02300_, _02297_);
  and (_02302_, _01698_, _01953_);
  and (_02303_, _01710_, _01964_);
  or (_02304_, _02303_, _02302_);
  and (_02305_, _01661_, _01977_);
  and (_02306_, _01682_, _01961_);
  or (_02307_, _02306_, _02305_);
  or (_02308_, _02307_, _02304_);
  and (_02309_, _01688_, _01968_);
  and (_02310_, _01702_, _01985_);
  or (_02311_, _02310_, _02309_);
  or (_02312_, _02311_, _02308_);
  and (_02313_, _01649_, _01947_);
  and (_02314_, _01656_, _01982_);
  or (_02315_, _02314_, _02313_);
  or (_02316_, _02315_, _02312_);
  or (_02317_, _02316_, _02301_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02317_, _02294_);
  and (_02318_, _01669_, _02035_);
  and (_02319_, _01644_, _02003_);
  or (_02320_, _02319_, _02318_);
  and (_02321_, _01672_, _02009_);
  and (_02322_, _01675_, _02012_);
  or (_02323_, _02322_, _02321_);
  or (_02324_, _02323_, _02320_);
  and (_02325_, _01702_, _02040_);
  and (_02326_, _01692_, _02026_);
  or (_02327_, _02326_, _02325_);
  and (_02328_, _01688_, _02020_);
  and (_02329_, _01720_, _02050_);
  or (_02330_, _02329_, _02328_);
  or (_02331_, _02330_, _02327_);
  and (_02332_, _01682_, _02017_);
  and (_02333_, _01710_, _02048_);
  or (_02334_, _02333_, _02332_);
  and (_02335_, _01698_, _02030_);
  and (_02336_, _01661_, _02005_);
  or (_02337_, _02336_, _02335_);
  or (_02338_, _02337_, _02334_);
  and (_02339_, _01717_, _02024_);
  and (_02340_, _01714_, _02037_);
  or (_02341_, _02340_, _02339_);
  or (_02342_, _02341_, _02338_);
  and (_02343_, _01649_, _02032_);
  and (_02344_, _01656_, _02042_);
  or (_02345_, _02344_, _02343_);
  or (_02346_, _02345_, _02342_);
  or (_02347_, _02346_, _02331_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02347_, _02324_);
  and (_02348_, _01669_, _02090_);
  and (_02349_, _01672_, _02065_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _01644_, _02108_);
  and (_02352_, _01675_, _02068_);
  or (_02353_, _02352_, _02351_);
  or (_02354_, _02353_, _02350_);
  and (_02355_, _01692_, _02081_);
  and (_02356_, _01702_, _02092_);
  or (_02357_, _02356_, _02355_);
  and (_02358_, _01717_, _02073_);
  and (_02359_, _01714_, _02087_);
  or (_02360_, _02359_, _02358_);
  or (_02361_, _02360_, _02357_);
  and (_02362_, _01698_, _02059_);
  and (_02363_, _01710_, _02076_);
  or (_02364_, _02363_, _02362_);
  and (_02365_, _01661_, _02061_);
  and (_02366_, _01682_, _02097_);
  or (_02367_, _02366_, _02365_);
  or (_02368_, _02367_, _02364_);
  and (_02369_, _01688_, _02079_);
  and (_02370_, _01720_, _02100_);
  or (_02371_, _02370_, _02369_);
  or (_02372_, _02371_, _02368_);
  and (_02373_, _01649_, _02105_);
  and (_02374_, _01656_, _02085_);
  or (_02375_, _02374_, _02373_);
  or (_02376_, _02375_, _02372_);
  or (_02377_, _02376_, _02361_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02377_, _02354_);
  and (_02378_, _01656_, _02147_);
  and (_02379_, _01644_, _02115_);
  or (_02380_, _02379_, _02378_);
  and (_02381_, _01675_, _02124_);
  and (_02382_, _01649_, _02121_);
  or (_02383_, _02382_, _02381_);
  or (_02384_, _02383_, _02380_);
  and (_02385_, _01720_, _02136_);
  and (_02386_, _01702_, _02142_);
  or (_02387_, _02386_, _02385_);
  and (_02388_, _01717_, _02134_);
  and (_02389_, _01688_, _02131_);
  or (_02390_, _02389_, _02388_);
  or (_02391_, _02390_, _02387_);
  and (_02392_, _01682_, _02153_);
  and (_02393_, _01698_, _02161_);
  or (_02394_, _02393_, _02392_);
  and (_02395_, _01710_, _02129_);
  and (_02396_, _01661_, _02117_);
  or (_02397_, _02396_, _02395_);
  or (_02398_, _02397_, _02394_);
  and (_02399_, _01714_, _02140_);
  and (_02400_, _01692_, _02156_);
  or (_02401_, _02400_, _02399_);
  or (_02402_, _02401_, _02398_);
  and (_02403_, _01669_, _02145_);
  and (_02404_, _01672_, _02164_);
  or (_02405_, _02404_, _02403_);
  or (_02406_, _02405_, _02402_);
  or (_02407_, _02406_, _02391_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02407_, _02384_);
  and (_02408_, _01669_, _02201_);
  and (_02409_, _01644_, _02220_);
  or (_02410_, _02409_, _02408_);
  and (_02411_, _01672_, _02180_);
  and (_02412_, _01675_, _02171_);
  or (_02413_, _02412_, _02411_);
  or (_02414_, _02413_, _02410_);
  and (_02415_, _01692_, _02191_);
  and (_02416_, _01720_, _02212_);
  or (_02417_, _02416_, _02415_);
  and (_02418_, _01717_, _02189_);
  and (_02419_, _01714_, _02195_);
  or (_02420_, _02419_, _02418_);
  or (_02421_, _02420_, _02417_);
  and (_02422_, _01698_, _02217_);
  and (_02423_, _01710_, _02209_);
  or (_02424_, _02423_, _02422_);
  and (_02425_, _01661_, _02173_);
  and (_02426_, _01682_, _02184_);
  or (_02427_, _02426_, _02425_);
  or (_02428_, _02427_, _02424_);
  and (_02429_, _01688_, _02186_);
  and (_02430_, _01702_, _02197_);
  or (_02431_, _02430_, _02429_);
  or (_02432_, _02431_, _02428_);
  and (_02433_, _01649_, _02177_);
  and (_02434_, _01656_, _02204_);
  or (_02435_, _02434_, _02433_);
  or (_02436_, _02435_, _02432_);
  or (_02437_, _02436_, _02421_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02437_, _02414_);
  and (_02438_, _01644_, _01867_);
  and (_02439_, _01669_, _01849_);
  or (_02440_, _02439_, _02438_);
  and (_02441_, _01672_, _01870_);
  and (_02442_, _01656_, _01844_);
  or (_02443_, _02442_, _02441_);
  or (_02444_, _02443_, _02440_);
  and (_02445_, _01688_, _01859_);
  and (_02446_, _01692_, _01864_);
  or (_02447_, _02446_, _02445_);
  and (_02448_, _01714_, _01878_);
  and (_02449_, _01717_, _01876_);
  or (_02450_, _02449_, _02448_);
  or (_02451_, _02450_, _02447_);
  and (_02452_, _01661_, _01837_);
  and (_02453_, _01710_, _01856_);
  or (_02454_, _02453_, _02452_);
  and (_02455_, _01698_, _01841_);
  and (_02456_, _01682_, _01852_);
  or (_02457_, _02456_, _02455_);
  or (_02458_, _02457_, _02454_);
  and (_02459_, _01702_, _01882_);
  and (_02460_, _01720_, _01872_);
  or (_02461_, _02460_, _02459_);
  or (_02462_, _02461_, _02458_);
  and (_02463_, _01649_, _01834_);
  and (_02464_, _01675_, _01884_);
  or (_02465_, _02464_, _02463_);
  or (_02466_, _02465_, _02462_);
  or (_02467_, _02466_, _02451_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02467_, _02444_);
  and (_02468_, _01644_, _01932_);
  and (_02469_, _01649_, _01900_);
  or (_02470_, _02469_, _02468_);
  and (_02471_, _01669_, _01936_);
  and (_02473_, _01656_, _01922_);
  or (_02474_, _02473_, _02471_);
  or (_02475_, _02474_, _02470_);
  and (_02476_, _01692_, _01930_);
  and (_02477_, _01702_, _01893_);
  or (_02478_, _02477_, _02476_);
  and (_02479_, _01720_, _01927_);
  and (_02480_, _01714_, _01905_);
  or (_02481_, _02480_, _02479_);
  or (_02482_, _02481_, _02478_);
  and (_02483_, _01682_, _01908_);
  and (_02484_, _01698_, _01891_);
  or (_02485_, _02484_, _02483_);
  and (_02486_, _01710_, _01912_);
  and (_02487_, _01661_, _01920_);
  or (_02488_, _02487_, _02486_);
  or (_02489_, _02488_, _02485_);
  and (_02490_, _01717_, _01938_);
  and (_02491_, _01688_, _01915_);
  or (_02492_, _02491_, _02490_);
  or (_02493_, _02492_, _02489_);
  and (_02494_, _01672_, _01925_);
  and (_02495_, _01675_, _01897_);
  or (_02496_, _02495_, _02494_);
  or (_02497_, _02496_, _02493_);
  or (_02498_, _02497_, _02482_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02498_, _02475_);
  and (_02499_, _01644_, _01982_);
  and (_02500_, _01669_, _01964_);
  or (_02501_, _02500_, _02499_);
  and (_02502_, _01672_, _01980_);
  and (_02503_, _01675_, _01956_);
  or (_02504_, _02503_, _02502_);
  or (_02505_, _02504_, _02501_);
  and (_02506_, _01688_, _01991_);
  and (_02507_, _01692_, _01985_);
  or (_02508_, _02507_, _02506_);
  and (_02509_, _01717_, _01994_);
  and (_02510_, _01720_, _01987_);
  or (_02511_, _02510_, _02509_);
  or (_02512_, _02511_, _02508_);
  and (_02513_, _01698_, _01947_);
  and (_02514_, _01710_, _01971_);
  or (_02515_, _02514_, _02513_);
  and (_02516_, _01661_, _01975_);
  and (_02517_, _01682_, _01968_);
  or (_02518_, _02517_, _02516_);
  or (_02519_, _02518_, _02515_);
  and (_02520_, _01702_, _01953_);
  and (_02521_, _01714_, _01961_);
  or (_02522_, _02521_, _02520_);
  or (_02523_, _02522_, _02519_);
  and (_02524_, _01649_, _01949_);
  and (_02525_, _01656_, _01977_);
  or (_02526_, _02525_, _02524_);
  or (_02527_, _02526_, _02523_);
  or (_02528_, _02527_, _02512_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02528_, _02505_);
  and (_02529_, _01672_, _02035_);
  and (_02530_, _01644_, _02042_);
  or (_02531_, _02530_, _02529_);
  and (_02532_, _01669_, _02048_);
  and (_02533_, _01649_, _02003_);
  or (_02534_, _02533_, _02532_);
  or (_02535_, _02534_, _02531_);
  and (_02536_, _01717_, _02050_);
  and (_02537_, _01688_, _02026_);
  or (_02538_, _02537_, _02536_);
  and (_02539_, _01720_, _02037_);
  and (_02540_, _01702_, _02030_);
  or (_02541_, _02540_, _02539_);
  or (_02542_, _02541_, _02538_);
  and (_02543_, _01675_, _02009_);
  and (_02544_, _01656_, _02005_);
  or (_02545_, _02544_, _02543_);
  and (_02546_, _01682_, _02020_);
  and (_02547_, _01698_, _02032_);
  or (_02548_, _02547_, _02546_);
  and (_02549_, _01710_, _02024_);
  and (_02550_, _01661_, _02012_);
  or (_02551_, _02550_, _02549_);
  or (_02552_, _02551_, _02548_);
  and (_02553_, _01692_, _02040_);
  and (_02554_, _01714_, _02017_);
  or (_02555_, _02554_, _02553_);
  or (_02556_, _02555_, _02552_);
  or (_02557_, _02556_, _02545_);
  or (_02558_, _02557_, _02542_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02558_, _02535_);
  and (_02559_, _01644_, _02085_);
  and (_02560_, _01649_, _02108_);
  or (_02561_, _02560_, _02559_);
  and (_02562_, _01672_, _02090_);
  and (_02563_, _01656_, _02061_);
  or (_02564_, _02563_, _02562_);
  or (_02565_, _02564_, _02561_);
  and (_02566_, _01692_, _02092_);
  and (_02567_, _01702_, _02059_);
  or (_02568_, _02567_, _02566_);
  and (_02569_, _01714_, _02097_);
  and (_02570_, _01720_, _02087_);
  or (_02571_, _02570_, _02569_);
  or (_02572_, _02571_, _02568_);
  and (_02573_, _01710_, _02073_);
  and (_02574_, _01698_, _02105_);
  or (_02575_, _02574_, _02573_);
  and (_02576_, _01682_, _02079_);
  and (_02577_, _01661_, _02068_);
  or (_02578_, _02577_, _02576_);
  or (_02579_, _02578_, _02575_);
  and (_02580_, _01688_, _02081_);
  and (_02581_, _01717_, _02100_);
  or (_02582_, _02581_, _02580_);
  or (_02583_, _02582_, _02579_);
  and (_02584_, _01669_, _02076_);
  and (_02585_, _01675_, _02065_);
  or (_02586_, _02585_, _02584_);
  or (_02587_, _02586_, _02583_);
  or (_02588_, _02587_, _02572_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02588_, _02565_);
  and (_02589_, _01644_, _02147_);
  and (_02590_, _01649_, _02115_);
  or (_02591_, _02590_, _02589_);
  and (_02592_, _01672_, _02145_);
  and (_02593_, _01656_, _02117_);
  or (_02594_, _02593_, _02592_);
  or (_02595_, _02594_, _02591_);
  and (_02596_, _01692_, _02142_);
  and (_02597_, _01702_, _02161_);
  or (_02598_, _02597_, _02596_);
  and (_02599_, _01720_, _02140_);
  and (_02600_, _01714_, _02153_);
  or (_02601_, _02600_, _02599_);
  or (_02602_, _02601_, _02598_);
  and (_02603_, _01682_, _02131_);
  and (_02604_, _01698_, _02121_);
  or (_02605_, _02604_, _02603_);
  and (_02606_, _01710_, _02134_);
  and (_02607_, _01661_, _02124_);
  or (_02608_, _02607_, _02606_);
  or (_02609_, _02608_, _02605_);
  and (_02610_, _01717_, _02136_);
  and (_02611_, _01688_, _02156_);
  or (_02612_, _02611_, _02610_);
  or (_02613_, _02612_, _02609_);
  and (_02614_, _01669_, _02129_);
  and (_02615_, _01675_, _02164_);
  or (_02616_, _02615_, _02614_);
  or (_02617_, _02616_, _02613_);
  or (_02618_, _02617_, _02602_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02618_, _02595_);
  and (_02619_, _01672_, _02201_);
  and (_02620_, _01656_, _02173_);
  or (_02621_, _02620_, _02619_);
  and (_02622_, _01669_, _02209_);
  and (_02623_, _01675_, _02180_);
  or (_02624_, _02623_, _02622_);
  or (_02625_, _02624_, _02621_);
  and (_02626_, _01717_, _02212_);
  and (_02627_, _01714_, _02184_);
  or (_02628_, _02627_, _02626_);
  and (_02629_, _01720_, _02195_);
  and (_02630_, _01702_, _02217_);
  or (_02631_, _02630_, _02629_);
  or (_02632_, _02631_, _02628_);
  and (_02633_, _01644_, _02204_);
  and (_02634_, _01649_, _02220_);
  or (_02635_, _02634_, _02633_);
  and (_02636_, _01688_, _02191_);
  and (_02637_, _01692_, _02197_);
  or (_02638_, _02637_, _02636_);
  and (_02639_, _01710_, _02189_);
  and (_02640_, _01661_, _02171_);
  or (_02641_, _02640_, _02639_);
  and (_02642_, _01682_, _02186_);
  and (_02643_, _01698_, _02177_);
  or (_02644_, _02643_, _02642_);
  or (_02645_, _02644_, _02641_);
  or (_02646_, _02645_, _02638_);
  or (_02647_, _02646_, _02635_);
  or (_02648_, _02647_, _02632_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02648_, _02625_);
  and (_02649_, _01675_, _01870_);
  and (_02650_, _01672_, _01849_);
  or (_02651_, _02650_, _02649_);
  and (_02652_, _01669_, _01856_);
  and (_02653_, _01656_, _01837_);
  or (_02654_, _02653_, _02652_);
  or (_02655_, _02654_, _02651_);
  and (_02656_, _01720_, _01878_);
  and (_02657_, _01692_, _01882_);
  or (_02658_, _02657_, _02656_);
  and (_02659_, _01717_, _01872_);
  and (_02660_, _01714_, _01852_);
  or (_02661_, _02660_, _02659_);
  or (_02662_, _02661_, _02658_);
  and (_02663_, _01698_, _01834_);
  and (_02664_, _01661_, _01884_);
  or (_02665_, _02664_, _02663_);
  and (_02666_, _01710_, _01876_);
  and (_02668_, _01682_, _01859_);
  or (_02669_, _02668_, _02666_);
  or (_02670_, _02669_, _02665_);
  and (_02671_, _01688_, _01864_);
  and (_02672_, _01702_, _01841_);
  or (_02673_, _02672_, _02671_);
  or (_02674_, _02673_, _02670_);
  and (_02675_, _01649_, _01867_);
  and (_02676_, _01644_, _01844_);
  or (_02677_, _02676_, _02675_);
  or (_02678_, _02677_, _02674_);
  or (_02679_, _02678_, _02662_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02679_, _02655_);
  and (_02680_, _01675_, _01925_);
  and (_02681_, _01644_, _01922_);
  or (_02682_, _02681_, _02680_);
  and (_02683_, _01669_, _01912_);
  and (_02684_, _01649_, _01932_);
  or (_02685_, _02684_, _02683_);
  or (_02686_, _02685_, _02682_);
  and (_02687_, _01714_, _01908_);
  and (_02688_, _01720_, _01905_);
  or (_02689_, _02688_, _02687_);
  and (_02690_, _01702_, _01891_);
  and (_02691_, _01692_, _01893_);
  or (_02692_, _02691_, _02690_);
  or (_02693_, _02692_, _02689_);
  and (_02694_, _01698_, _01900_);
  and (_02695_, _01661_, _01897_);
  or (_02696_, _02695_, _02694_);
  and (_02697_, _01710_, _01938_);
  and (_02698_, _01682_, _01915_);
  or (_02699_, _02698_, _02697_);
  or (_02700_, _02699_, _02696_);
  and (_02701_, _01717_, _01927_);
  and (_02702_, _01688_, _01930_);
  or (_02703_, _02702_, _02701_);
  or (_02704_, _02703_, _02700_);
  and (_02705_, _01672_, _01936_);
  and (_02706_, _01656_, _01920_);
  or (_02707_, _02706_, _02705_);
  or (_02708_, _02707_, _02704_);
  or (_02709_, _02708_, _02693_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02709_, _02686_);
  and (_02710_, _01672_, _01964_);
  and (_02711_, _01675_, _01980_);
  or (_02712_, _02711_, _02710_);
  and (_02713_, _01717_, _01987_);
  and (_02714_, _01714_, _01968_);
  and (_02715_, _01720_, _01961_);
  or (_02716_, _02715_, _02714_);
  and (_02717_, _01688_, _01985_);
  and (_02718_, _01682_, _01991_);
  or (_02719_, _02718_, _02717_);
  or (_02720_, _02719_, _02716_);
  or (_02721_, _02720_, _02713_);
  or (_02722_, _02721_, _02712_);
  and (_02723_, _01692_, _01953_);
  and (_02724_, _01702_, _01947_);
  or (_02725_, _02724_, _02723_);
  and (_02726_, _01698_, _01949_);
  and (_02727_, _01649_, _01982_);
  or (_02728_, _02727_, _02726_);
  or (_02729_, _02728_, _02725_);
  and (_02730_, _01661_, _01956_);
  and (_02731_, _01656_, _01975_);
  and (_02732_, _01644_, _01977_);
  or (_02733_, _02732_, _02731_);
  or (_02734_, _02733_, _02730_);
  or (_02735_, _02734_, _02729_);
  and (_02736_, _01669_, _01971_);
  and (_02737_, _01710_, _01994_);
  or (_02738_, _02737_, _02736_);
  or (_02739_, _02738_, _02735_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02739_, _02722_);
  and (_02740_, _01675_, _02035_);
  and (_02741_, _01644_, _02005_);
  or (_02742_, _02741_, _02740_);
  and (_02743_, _01669_, _02024_);
  and (_02744_, _01656_, _02012_);
  or (_02745_, _02744_, _02743_);
  or (_02746_, _02745_, _02742_);
  and (_02747_, _01688_, _02040_);
  and (_02748_, _01714_, _02020_);
  or (_02749_, _02748_, _02747_);
  and (_02750_, _01720_, _02017_);
  and (_02751_, _01692_, _02030_);
  or (_02752_, _02751_, _02750_);
  or (_02753_, _02752_, _02749_);
  and (_02754_, _01682_, _02026_);
  and (_02755_, _01698_, _02003_);
  or (_02756_, _02755_, _02754_);
  and (_02757_, _01710_, _02050_);
  and (_02758_, _01661_, _02009_);
  or (_02759_, _02758_, _02757_);
  or (_02760_, _02759_, _02756_);
  and (_02761_, _01717_, _02037_);
  and (_02762_, _01702_, _02032_);
  or (_02763_, _02762_, _02761_);
  or (_02764_, _02763_, _02760_);
  and (_02765_, _01672_, _02048_);
  and (_02766_, _01649_, _02042_);
  or (_02767_, _02766_, _02765_);
  or (_02768_, _02767_, _02764_);
  or (_02769_, _02768_, _02753_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02769_, _02746_);
  and (_02770_, _01675_, _02090_);
  and (_02771_, _01672_, _02076_);
  or (_02772_, _02771_, _02770_);
  and (_02773_, _01669_, _02073_);
  and (_02774_, _01720_, _02097_);
  and (_02775_, _01714_, _02079_);
  or (_02776_, _02775_, _02774_);
  and (_02777_, _01688_, _02092_);
  and (_02778_, _01682_, _02081_);
  or (_02779_, _02778_, _02777_);
  or (_02780_, _02779_, _02776_);
  or (_02781_, _02780_, _02773_);
  or (_02782_, _02781_, _02772_);
  and (_02783_, _01692_, _02059_);
  and (_02784_, _01702_, _02105_);
  or (_02785_, _02784_, _02783_);
  and (_02786_, _01649_, _02085_);
  and (_02787_, _01698_, _02108_);
  or (_02788_, _02787_, _02786_);
  or (_02789_, _02788_, _02785_);
  and (_02790_, _01661_, _02065_);
  and (_02791_, _01656_, _02068_);
  and (_02792_, _01644_, _02061_);
  or (_02793_, _02792_, _02791_);
  or (_02794_, _02793_, _02790_);
  or (_02795_, _02794_, _02789_);
  and (_02796_, _01717_, _02087_);
  and (_02797_, _01710_, _02100_);
  or (_02798_, _02797_, _02796_);
  or (_02799_, _02798_, _02795_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02799_, _02782_);
  and (_02800_, _01669_, _02134_);
  and (_02801_, _01649_, _02147_);
  or (_02802_, _02801_, _02800_);
  and (_02803_, _01672_, _02129_);
  and (_02804_, _01656_, _02124_);
  or (_02805_, _02804_, _02803_);
  or (_02806_, _02805_, _02802_);
  and (_02807_, _01714_, _02131_);
  and (_02808_, _01720_, _02153_);
  or (_02809_, _02808_, _02807_);
  and (_02810_, _01702_, _02121_);
  and (_02811_, _01692_, _02161_);
  or (_02812_, _02811_, _02810_);
  or (_02813_, _02812_, _02809_);
  and (_02814_, _01682_, _02156_);
  and (_02815_, _01698_, _02115_);
  or (_02816_, _02815_, _02814_);
  and (_02817_, _01710_, _02136_);
  and (_02818_, _01661_, _02164_);
  or (_02819_, _02818_, _02817_);
  or (_02820_, _02819_, _02816_);
  and (_02821_, _01717_, _02140_);
  and (_02822_, _01688_, _02142_);
  or (_02823_, _02822_, _02821_);
  or (_02824_, _02823_, _02820_);
  and (_02825_, _01675_, _02145_);
  and (_02826_, _01644_, _02117_);
  or (_02827_, _02826_, _02825_);
  or (_02828_, _02827_, _02824_);
  or (_02829_, _02828_, _02813_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02829_, _02806_);
  and (_02830_, _01656_, _02171_);
  and (_02831_, _01644_, _02173_);
  or (_02832_, _02831_, _02830_);
  and (_02833_, _01675_, _02201_);
  and (_02834_, _01649_, _02204_);
  or (_02835_, _02834_, _02833_);
  or (_02836_, _02835_, _02832_);
  and (_02837_, _01714_, _02186_);
  and (_02838_, _01720_, _02184_);
  or (_02839_, _02838_, _02837_);
  and (_02840_, _01692_, _02217_);
  and (_02841_, _01702_, _02177_);
  or (_02842_, _02841_, _02840_);
  or (_02843_, _02842_, _02839_);
  and (_02844_, _01669_, _02189_);
  and (_02845_, _01672_, _02209_);
  or (_02846_, _02845_, _02844_);
  and (_02847_, _01682_, _02191_);
  and (_02848_, _01698_, _02220_);
  or (_02849_, _02848_, _02847_);
  and (_02850_, _01710_, _02212_);
  and (_02851_, _01661_, _02180_);
  or (_02852_, _02851_, _02850_);
  or (_02853_, _02852_, _02849_);
  and (_02854_, _01717_, _02195_);
  and (_02855_, _01688_, _02197_);
  or (_02856_, _02855_, _02854_);
  or (_02857_, _02856_, _02853_);
  or (_02858_, _02857_, _02846_);
  or (_02859_, _02858_, _02843_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02859_, _02836_);
  not (_02860_, \oc8051_golden_model_1.PC [1]);
  nand (_02862_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  nor (_02863_, _02862_, _02860_);
  and (_02864_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02865_, _02864_, \oc8051_golden_model_1.PC [3]);
  nor (_02866_, _02865_, _02863_);
  nand (_02867_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02868_, \oc8051_golden_model_1.PC [3]);
  or (_02869_, \oc8051_golden_model_1.PC [2], _02868_);
  or (_02870_, _02869_, _02867_);
  or (_02871_, _02870_, _42320_);
  or (_02872_, _02860_, \oc8051_golden_model_1.PC [0]);
  or (_02873_, _02872_, _02869_);
  or (_02874_, _02873_, _42279_);
  and (_02875_, _02874_, _02871_);
  not (_02876_, \oc8051_golden_model_1.PC [2]);
  or (_02877_, _02876_, \oc8051_golden_model_1.PC [3]);
  or (_02878_, _02877_, _02867_);
  or (_02879_, _02878_, _42156_);
  or (_02880_, _02877_, _02872_);
  or (_02881_, _02880_, _42115_);
  and (_02882_, _02881_, _02879_);
  and (_02883_, _02882_, _02875_);
  or (_02884_, _02862_, _02867_);
  or (_02885_, _02884_, _42484_);
  or (_02886_, _02862_, _02872_);
  or (_02887_, _02886_, _42443_);
  and (_02888_, _02887_, _02885_);
  or (_02889_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02890_, _02889_, _02867_);
  or (_02891_, _02890_, _41984_);
  or (_02892_, _02889_, _02872_);
  or (_02893_, _02892_, _41936_);
  and (_02894_, _02893_, _02891_);
  and (_02895_, _02894_, _02888_);
  and (_02896_, _02895_, _02883_);
  not (_02897_, \oc8051_golden_model_1.PC [0]);
  or (_02898_, \oc8051_golden_model_1.PC [1], _02897_);
  or (_02899_, _02898_, _02862_);
  or (_02900_, _02899_, _42402_);
  or (_02901_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02902_, _02901_, _02862_);
  or (_02903_, _02902_, _42361_);
  and (_02904_, _02903_, _02900_);
  or (_02905_, _02889_, _02901_);
  or (_02906_, _02905_, _41854_);
  or (_02907_, _02889_, _02898_);
  or (_02908_, _02907_, _41895_);
  and (_02909_, _02908_, _02906_);
  and (_02910_, _02909_, _02904_);
  or (_02911_, _02898_, _02869_);
  or (_02912_, _02911_, _42238_);
  or (_02913_, _02901_, _02869_);
  or (_02914_, _02913_, _42197_);
  and (_02915_, _02914_, _02912_);
  or (_02916_, _02898_, _02877_);
  or (_02917_, _02916_, _42074_);
  or (_02918_, _02901_, _02877_);
  or (_02919_, _02918_, _42033_);
  and (_02920_, _02919_, _02917_);
  and (_02921_, _02920_, _02915_);
  and (_02922_, _02921_, _02910_);
  nand (_02923_, _02922_, _02896_);
  or (_02924_, _02870_, _42325_);
  or (_02925_, _02873_, _42284_);
  and (_02926_, _02925_, _02924_);
  or (_02927_, _02878_, _42161_);
  or (_02928_, _02880_, _42120_);
  and (_02929_, _02928_, _02927_);
  and (_02930_, _02929_, _02926_);
  or (_02931_, _02884_, _42489_);
  or (_02932_, _02886_, _42448_);
  and (_02933_, _02932_, _02931_);
  or (_02934_, _02890_, _41989_);
  or (_02935_, _02892_, _41941_);
  and (_02936_, _02935_, _02934_);
  and (_02937_, _02936_, _02933_);
  and (_02938_, _02937_, _02930_);
  or (_02939_, _02899_, _42407_);
  or (_02940_, _02902_, _42366_);
  and (_02941_, _02940_, _02939_);
  or (_02942_, _02905_, _41859_);
  or (_02943_, _02907_, _41900_);
  and (_02944_, _02943_, _02942_);
  and (_02945_, _02944_, _02941_);
  or (_02946_, _02911_, _42243_);
  or (_02947_, _02913_, _42202_);
  and (_02948_, _02947_, _02946_);
  or (_02949_, _02916_, _42079_);
  or (_02950_, _02918_, _42038_);
  and (_02951_, _02950_, _02949_);
  and (_02952_, _02951_, _02948_);
  and (_02953_, _02952_, _02945_);
  nand (_02954_, _02953_, _02938_);
  or (_02955_, _02954_, _02923_);
  or (_02956_, _02870_, _42310_);
  or (_02957_, _02873_, _42269_);
  and (_02958_, _02957_, _02956_);
  or (_02959_, _02878_, _42146_);
  or (_02960_, _02880_, _42105_);
  and (_02961_, _02960_, _02959_);
  and (_02962_, _02961_, _02958_);
  or (_02963_, _02884_, _42474_);
  or (_02964_, _02886_, _42433_);
  and (_02965_, _02964_, _02963_);
  or (_02966_, _02890_, _41974_);
  or (_02967_, _02892_, _41926_);
  and (_02968_, _02967_, _02966_);
  and (_02969_, _02968_, _02965_);
  and (_02970_, _02969_, _02962_);
  or (_02971_, _02899_, _42392_);
  or (_02972_, _02902_, _42351_);
  and (_02973_, _02972_, _02971_);
  or (_02974_, _02905_, _41844_);
  or (_02975_, _02907_, _41885_);
  and (_02976_, _02975_, _02974_);
  and (_02977_, _02976_, _02973_);
  or (_02978_, _02911_, _42228_);
  or (_02979_, _02913_, _42187_);
  and (_02980_, _02979_, _02978_);
  or (_02981_, _02916_, _42064_);
  or (_02982_, _02918_, _42023_);
  and (_02983_, _02982_, _02981_);
  and (_02984_, _02983_, _02980_);
  and (_02985_, _02984_, _02977_);
  and (_02986_, _02985_, _02970_);
  or (_02987_, _02870_, _42315_);
  or (_02988_, _02873_, _42274_);
  and (_02989_, _02988_, _02987_);
  or (_02990_, _02878_, _42151_);
  or (_02991_, _02880_, _42110_);
  and (_02992_, _02991_, _02990_);
  and (_02993_, _02992_, _02989_);
  or (_02994_, _02884_, _42479_);
  or (_02995_, _02886_, _42438_);
  and (_02996_, _02995_, _02994_);
  or (_02997_, _02890_, _41979_);
  or (_02998_, _02892_, _41931_);
  and (_02999_, _02998_, _02997_);
  and (_03000_, _02999_, _02996_);
  and (_03001_, _03000_, _02993_);
  or (_03002_, _02899_, _42397_);
  or (_03003_, _02902_, _42356_);
  and (_03004_, _03003_, _03002_);
  or (_03005_, _02905_, _41849_);
  or (_03006_, _02907_, _41890_);
  and (_03007_, _03006_, _03005_);
  and (_03008_, _03007_, _03004_);
  or (_03009_, _02911_, _42233_);
  or (_03010_, _02913_, _42192_);
  and (_03011_, _03010_, _03009_);
  or (_03012_, _02916_, _42069_);
  or (_03013_, _02918_, _42028_);
  and (_03014_, _03013_, _03012_);
  and (_03015_, _03014_, _03011_);
  and (_03016_, _03015_, _03008_);
  nand (_03017_, _03016_, _03001_);
  or (_03018_, _03017_, _02986_);
  or (_03019_, _03018_, _02955_);
  not (_03020_, _03019_);
  or (_03021_, _02870_, _42340_);
  or (_03023_, _02873_, _42299_);
  and (_03024_, _03023_, _03021_);
  or (_03025_, _02878_, _42176_);
  or (_03026_, _02880_, _42135_);
  and (_03027_, _03026_, _03025_);
  and (_03028_, _03027_, _03024_);
  or (_03029_, _02884_, _42504_);
  or (_03030_, _02886_, _42463_);
  and (_03031_, _03030_, _03029_);
  or (_03032_, _02890_, _42012_);
  or (_03034_, _02892_, _41963_);
  and (_03035_, _03034_, _03032_);
  and (_03036_, _03035_, _03031_);
  and (_03037_, _03036_, _03028_);
  or (_03038_, _02899_, _42422_);
  or (_03039_, _02902_, _42381_);
  and (_03040_, _03039_, _03038_);
  or (_03041_, _02905_, _41874_);
  or (_03042_, _02907_, _41915_);
  and (_03043_, _03042_, _03041_);
  and (_03044_, _03043_, _03040_);
  or (_03045_, _02911_, _42258_);
  or (_03046_, _02913_, _42217_);
  and (_03047_, _03046_, _03045_);
  or (_03048_, _02916_, _42094_);
  or (_03049_, _02918_, _42053_);
  and (_03050_, _03049_, _03048_);
  and (_03051_, _03050_, _03047_);
  and (_03052_, _03051_, _03044_);
  nand (_03053_, _03052_, _03037_);
  or (_03055_, _02870_, _42305_);
  or (_03056_, _02873_, _42264_);
  and (_03057_, _03056_, _03055_);
  or (_03058_, _02878_, _42141_);
  or (_03059_, _02880_, _42100_);
  and (_03060_, _03059_, _03058_);
  and (_03061_, _03060_, _03057_);
  or (_03062_, _02884_, _42469_);
  or (_03063_, _02886_, _42428_);
  and (_03064_, _03063_, _03062_);
  or (_03066_, _02890_, _41969_);
  or (_03067_, _02892_, _41921_);
  and (_03068_, _03067_, _03066_);
  and (_03069_, _03068_, _03064_);
  and (_03070_, _03069_, _03061_);
  or (_03071_, _02899_, _42387_);
  or (_03072_, _02902_, _42346_);
  and (_03073_, _03072_, _03071_);
  or (_03074_, _02905_, _41839_);
  or (_03075_, _02907_, _41880_);
  and (_03077_, _03075_, _03074_);
  and (_03078_, _03077_, _03073_);
  or (_03079_, _02911_, _42223_);
  or (_03080_, _02913_, _42182_);
  and (_03081_, _03080_, _03079_);
  or (_03082_, _02916_, _42059_);
  or (_03083_, _02918_, _42018_);
  and (_03084_, _03083_, _03082_);
  and (_03085_, _03084_, _03081_);
  and (_03086_, _03085_, _03078_);
  and (_03087_, _03086_, _03070_);
  or (_03088_, _03087_, _03053_);
  or (_03089_, _02870_, _42330_);
  or (_03090_, _02873_, _42289_);
  and (_03091_, _03090_, _03089_);
  or (_03092_, _02878_, _42166_);
  or (_03093_, _02880_, _42125_);
  and (_03094_, _03093_, _03092_);
  and (_03095_, _03094_, _03091_);
  or (_03096_, _02884_, _42494_);
  or (_03098_, _02886_, _42453_);
  and (_03099_, _03098_, _03096_);
  or (_03100_, _02890_, _42000_);
  or (_03101_, _02892_, _41947_);
  and (_03102_, _03101_, _03100_);
  and (_03103_, _03102_, _03099_);
  and (_03104_, _03103_, _03095_);
  or (_03105_, _02899_, _42412_);
  or (_03106_, _02902_, _42371_);
  and (_03107_, _03106_, _03105_);
  or (_03109_, _02905_, _41864_);
  or (_03110_, _02907_, _41905_);
  and (_03111_, _03110_, _03109_);
  and (_03112_, _03111_, _03107_);
  or (_03113_, _02911_, _42248_);
  or (_03114_, _02913_, _42207_);
  and (_03115_, _03114_, _03113_);
  or (_03116_, _02916_, _42084_);
  or (_03117_, _02918_, _42043_);
  and (_03118_, _03117_, _03116_);
  and (_03120_, _03118_, _03115_);
  and (_03121_, _03120_, _03112_);
  nand (_03122_, _03121_, _03104_);
  or (_03123_, _02870_, _42335_);
  or (_03124_, _02873_, _42294_);
  and (_03125_, _03124_, _03123_);
  or (_03126_, _02878_, _42171_);
  or (_03127_, _02880_, _42130_);
  and (_03128_, _03127_, _03126_);
  and (_03129_, _03128_, _03125_);
  or (_03131_, _02884_, _42499_);
  or (_03132_, _02886_, _42458_);
  and (_03133_, _03132_, _03131_);
  or (_03134_, _02890_, _42007_);
  or (_03135_, _02892_, _41957_);
  and (_03136_, _03135_, _03134_);
  and (_03137_, _03136_, _03133_);
  and (_03138_, _03137_, _03129_);
  or (_03139_, _02899_, _42417_);
  or (_03140_, _02902_, _42376_);
  and (_03142_, _03140_, _03139_);
  or (_03143_, _02905_, _41869_);
  or (_03144_, _02907_, _41910_);
  and (_03145_, _03144_, _03143_);
  and (_03146_, _03145_, _03142_);
  or (_03147_, _02911_, _42253_);
  or (_03148_, _02913_, _42212_);
  and (_03149_, _03148_, _03147_);
  or (_03150_, _02916_, _42089_);
  or (_03151_, _02918_, _42048_);
  and (_03153_, _03151_, _03150_);
  and (_03154_, _03153_, _03149_);
  and (_03155_, _03154_, _03146_);
  nand (_03156_, _03155_, _03138_);
  or (_03157_, _03156_, _03122_);
  nor (_03158_, _03157_, _03088_);
  and (_03159_, _03158_, _03020_);
  not (_03160_, _03159_);
  and (_03161_, _03121_, _03104_);
  and (_03162_, _03155_, _03138_);
  or (_03164_, _03162_, _03161_);
  not (_03165_, _03164_);
  and (_03166_, _03087_, _03053_);
  and (_03167_, _03166_, _03165_);
  and (_03168_, _03167_, _03020_);
  or (_03169_, _03162_, _03122_);
  not (_03170_, _03169_);
  and (_03171_, _03170_, _03166_);
  and (_03172_, _03171_, _03020_);
  nor (_03173_, _03172_, _03168_);
  and (_03175_, _03173_, _03160_);
  not (_03176_, _03157_);
  and (_03177_, _03176_, _03166_);
  and (_03178_, _03177_, _03020_);
  or (_03179_, _03156_, _03161_);
  not (_03180_, _03179_);
  and (_03181_, _03180_, _03166_);
  and (_03182_, _03181_, _03020_);
  nor (_03183_, _03182_, _03178_);
  and (_03184_, _03183_, _03175_);
  and (_03186_, _03052_, _03037_);
  and (_03187_, _03087_, _03186_);
  and (_03188_, _03170_, _03187_);
  and (_03189_, _03188_, _03020_);
  and (_03190_, _03187_, _03165_);
  and (_03191_, _03190_, _03020_);
  nor (_03192_, _03191_, _03189_);
  and (_03193_, _03176_, _03187_);
  and (_03194_, _03193_, _03020_);
  and (_03195_, _03187_, _03180_);
  and (_03196_, _03195_, _03020_);
  nor (_03197_, _03196_, _03194_);
  and (_03198_, _03197_, _03192_);
  and (_03199_, _03198_, _03184_);
  or (_03200_, _03087_, _03186_);
  or (_03201_, _03200_, _03179_);
  or (_03202_, _03201_, _03019_);
  or (_03203_, _03200_, _03164_);
  or (_03204_, _03203_, _03019_);
  and (_03205_, _03204_, _03202_);
  or (_03206_, _03088_, _03164_);
  or (_03207_, _03206_, _03019_);
  or (_03208_, _03200_, _03169_);
  or (_03209_, _03208_, _03019_);
  and (_03210_, _03209_, _03207_);
  or (_03211_, _03200_, _03157_);
  or (_03212_, _03211_, _03019_);
  or (_03213_, _03169_, _03088_);
  or (_03214_, _03213_, _03019_);
  and (_03215_, _03214_, _03212_);
  and (_03216_, _03215_, _03210_);
  and (_03217_, _03216_, _03205_);
  nor (_03218_, _03088_, _03179_);
  and (_03219_, _03218_, _03020_);
  not (_03220_, _03018_);
  not (_03221_, _02954_);
  and (_03222_, _03221_, _02923_);
  and (_03223_, _03222_, _03220_);
  and (_03224_, _03223_, _03158_);
  nor (_03225_, _03224_, _03219_);
  and (_03226_, _03225_, _03217_);
  and (_03227_, _03226_, _03199_);
  or (_03228_, _03227_, _02866_);
  not (_03229_, _03218_);
  not (_03230_, _03017_);
  or (_03231_, _03230_, _02986_);
  or (_03232_, _03231_, _02955_);
  or (_03233_, _03232_, _03229_);
  and (_03234_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  and (_03235_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_03236_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03237_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03238_, _03237_, _03235_);
  and (_03239_, _03238_, _03236_);
  nor (_03240_, _03239_, _03235_);
  nor (_03241_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03242_, _03241_, _03234_);
  not (_03243_, _03242_);
  nor (_03244_, _03243_, _03240_);
  nor (_03245_, _03244_, _03234_);
  and (_03246_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03247_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03248_, _03247_, _03246_);
  not (_03249_, _03248_);
  nor (_03250_, _03249_, _03245_);
  and (_03251_, _03249_, _03245_);
  nor (_03252_, _03251_, _03250_);
  or (_03253_, _03252_, _03233_);
  not (_03254_, _02878_);
  nor (_03255_, _02867_, _02876_);
  nor (_03256_, _03255_, _02868_);
  nor (_03257_, _03256_, _03254_);
  and (_03258_, _03233_, _03257_);
  nand (_03259_, _03258_, _03217_);
  nand (_03260_, _03259_, _03253_);
  not (_03261_, _03158_);
  nor (_03262_, _03232_, _03261_);
  not (_03263_, _03262_);
  and (_03264_, _03263_, _03225_);
  and (_03265_, _03264_, _03260_);
  and (_03266_, _02867_, _02876_);
  nor (_03267_, _03266_, _03255_);
  and (_03268_, _03267_, \oc8051_golden_model_1.ACC [2]);
  not (_03269_, \oc8051_golden_model_1.ACC [1]);
  and (_03270_, _02898_, _02872_);
  nor (_03271_, _03270_, _03269_);
  and (_03272_, \oc8051_golden_model_1.ACC [0], _02897_);
  and (_03273_, _03270_, _03269_);
  nor (_03274_, _03273_, _03271_);
  and (_03275_, _03274_, _03272_);
  nor (_03277_, _03275_, _03271_);
  nor (_03278_, _03267_, \oc8051_golden_model_1.ACC [2]);
  nor (_03279_, _03278_, _03268_);
  not (_03280_, _03279_);
  nor (_03281_, _03280_, _03277_);
  nor (_03282_, _03281_, _03268_);
  nor (_03283_, _03257_, \oc8051_golden_model_1.ACC [3]);
  and (_03284_, _03257_, \oc8051_golden_model_1.ACC [3]);
  nor (_03285_, _03284_, _03283_);
  and (_03286_, _03285_, _03282_);
  nor (_03287_, _03285_, _03282_);
  nor (_03288_, _03287_, _03286_);
  nor (_03289_, _03288_, _03263_);
  or (_03290_, _03289_, _03265_);
  nand (_03291_, _03290_, _03199_);
  nand (_03292_, _03291_, _03228_);
  nor (_03293_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03294_, _03293_, _02864_);
  or (_03295_, _03294_, _03227_);
  and (_03296_, _03243_, _03240_);
  nor (_03297_, _03296_, _03244_);
  or (_03298_, _03297_, _03233_);
  not (_03299_, _03267_);
  and (_03300_, _03299_, _03233_);
  nand (_03301_, _03300_, _03217_);
  nand (_03302_, _03301_, _03298_);
  and (_03303_, _03302_, _03264_);
  and (_03304_, _03280_, _03277_);
  nor (_03305_, _03304_, _03281_);
  nor (_03306_, _03305_, _03263_);
  or (_03307_, _03306_, _03303_);
  nand (_03308_, _03307_, _03199_);
  nand (_03309_, _03308_, _03295_);
  or (_03310_, _03309_, _03292_);
  or (_03311_, _03199_, _02860_);
  or (_03312_, _03217_, \oc8051_golden_model_1.PC [1]);
  not (_03313_, _03270_);
  nand (_03314_, _03313_, _03217_);
  nand (_03315_, _03314_, _03312_);
  nand (_03316_, _03315_, _03233_);
  nor (_03317_, _03238_, _03236_);
  nor (_03318_, _03317_, _03239_);
  not (_03319_, _03318_);
  or (_03320_, _03319_, _03233_);
  and (_03321_, _03320_, _03225_);
  nand (_03322_, _03321_, _03316_);
  or (_03323_, _03225_, _02860_);
  and (_03324_, _03323_, _03263_);
  nand (_03325_, _03324_, _03322_);
  not (_03326_, _03199_);
  nor (_03327_, _03274_, _03272_);
  nor (_03328_, _03327_, _03275_);
  and (_03329_, _03328_, _03262_);
  nor (_03330_, _03329_, _03326_);
  nand (_03331_, _03330_, _03325_);
  and (_03332_, _03331_, _03311_);
  or (_03333_, _03226_, _02897_);
  not (_03334_, _03233_);
  nor (_03335_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03336_, _03335_, _03236_);
  nand (_03337_, _03336_, _03334_);
  and (_03338_, _03233_, _02897_);
  nand (_03339_, _03338_, _03217_);
  nand (_03340_, _03339_, _03337_);
  nand (_03341_, _03340_, _03225_);
  nand (_03342_, _03341_, _03333_);
  nand (_03343_, _03342_, _03263_);
  not (_03344_, \oc8051_golden_model_1.ACC [0]);
  and (_03345_, _03344_, \oc8051_golden_model_1.PC [0]);
  nor (_03346_, _03345_, _03272_);
  and (_03347_, _03346_, _03262_);
  nor (_03348_, _03347_, _03326_);
  nand (_03349_, _03348_, _03343_);
  or (_03350_, _03199_, \oc8051_golden_model_1.PC [0]);
  and (_03351_, _03350_, _03349_);
  or (_03352_, _03351_, _03332_);
  or (_03353_, _03352_, _03310_);
  or (_03354_, _03353_, _42346_);
  and (_03355_, _03291_, _03228_);
  and (_03356_, _03308_, _03295_);
  or (_03357_, _03356_, _03355_);
  or (_03358_, _03357_, _03352_);
  or (_03359_, _03358_, _41839_);
  and (_03360_, _03359_, _03354_);
  nand (_03361_, _03350_, _03349_);
  or (_03362_, _03361_, _03332_);
  or (_03363_, _03362_, _03310_);
  or (_03364_, _03363_, _42387_);
  nand (_03365_, _03331_, _03311_);
  or (_03366_, _03361_, _03365_);
  or (_03367_, _03309_, _03355_);
  or (_03368_, _03367_, _03366_);
  or (_03369_, _03368_, _42141_);
  and (_03370_, _03369_, _03364_);
  and (_03371_, _03370_, _03360_);
  or (_03372_, _03351_, _03365_);
  or (_03373_, _03372_, _03357_);
  or (_03374_, _03373_, _41921_);
  or (_03375_, _03362_, _03357_);
  or (_03376_, _03375_, _41880_);
  and (_03377_, _03376_, _03374_);
  or (_03378_, _03372_, _03310_);
  or (_03379_, _03378_, _42428_);
  or (_03380_, _03356_, _03292_);
  or (_03381_, _03380_, _03372_);
  or (_03382_, _03381_, _42264_);
  and (_03383_, _03382_, _03379_);
  and (_03384_, _03383_, _03377_);
  and (_03385_, _03384_, _03371_);
  or (_03386_, _03380_, _03362_);
  or (_03387_, _03386_, _42223_);
  or (_03388_, _03367_, _03352_);
  or (_03389_, _03388_, _42018_);
  and (_03390_, _03389_, _03387_);
  or (_03391_, _03366_, _03310_);
  or (_03392_, _03391_, _42469_);
  or (_03393_, _03380_, _03366_);
  or (_03394_, _03393_, _42305_);
  and (_03395_, _03394_, _03392_);
  and (_03396_, _03395_, _03390_);
  or (_03397_, _03380_, _03352_);
  or (_03398_, _03397_, _42182_);
  or (_03399_, _03367_, _03362_);
  or (_03400_, _03399_, _42059_);
  and (_03401_, _03400_, _03398_);
  or (_03402_, _03372_, _03367_);
  or (_03403_, _03402_, _42100_);
  or (_03404_, _03366_, _03357_);
  or (_03405_, _03404_, _41969_);
  and (_03406_, _03405_, _03403_);
  and (_03407_, _03406_, _03401_);
  and (_03408_, _03407_, _03396_);
  nand (_03409_, _03408_, _03385_);
  or (_03410_, _03391_, _42489_);
  or (_03411_, _03375_, _41900_);
  and (_03412_, _03411_, _03410_);
  or (_03413_, _03393_, _42325_);
  or (_03414_, _03358_, _41859_);
  and (_03415_, _03414_, _03413_);
  and (_03416_, _03415_, _03412_);
  or (_03417_, _03397_, _42202_);
  or (_03418_, _03373_, _41941_);
  and (_03419_, _03418_, _03417_);
  or (_03420_, _03368_, _42161_);
  or (_03421_, _03388_, _42038_);
  and (_03422_, _03421_, _03420_);
  and (_03423_, _03422_, _03419_);
  and (_03424_, _03423_, _03416_);
  or (_03425_, _03399_, _42079_);
  or (_03426_, _03404_, _41989_);
  and (_03427_, _03426_, _03425_);
  or (_03428_, _03378_, _42448_);
  or (_03429_, _03381_, _42284_);
  and (_03430_, _03429_, _03428_);
  and (_03431_, _03430_, _03427_);
  or (_03432_, _03353_, _42366_);
  or (_03433_, _03386_, _42243_);
  and (_03434_, _03433_, _03432_);
  or (_03435_, _03363_, _42407_);
  or (_03436_, _03402_, _42120_);
  and (_03437_, _03436_, _03435_);
  and (_03438_, _03437_, _03434_);
  and (_03439_, _03438_, _03431_);
  and (_03440_, _03439_, _03424_);
  or (_03441_, _03440_, _03409_);
  not (_03442_, _02955_);
  and (_03443_, _03230_, _02986_);
  and (_03444_, _03443_, _03442_);
  and (_03445_, _03444_, _03195_);
  not (_03446_, _03445_);
  nor (_03447_, _03446_, _03441_);
  nor (_03448_, _03446_, _03409_);
  not (_03449_, _03448_);
  and (_03450_, _03017_, _02986_);
  and (_03451_, _03450_, _03442_);
  and (_03452_, _03451_, _03218_);
  not (_03453_, _03452_);
  nor (_03454_, _03441_, _03453_);
  not (_03455_, \oc8051_golden_model_1.SP [0]);
  nor (_03456_, _03207_, _03455_);
  not (_03457_, _03206_);
  and (_03458_, _03457_, _03451_);
  not (_03459_, _03458_);
  nor (_03460_, _03459_, _03441_);
  nor (_03461_, _03459_, _03409_);
  not (_03462_, _03461_);
  not (_03463_, _03211_);
  and (_03464_, _03444_, _03463_);
  and (_03465_, _03463_, _03451_);
  not (_03466_, _03465_);
  nor (_03467_, _03466_, _03441_);
  not (_03468_, _03201_);
  and (_03469_, _03468_, _03451_);
  not (_03470_, _03469_);
  or (_03471_, _03470_, _03441_);
  nor (_03472_, _03470_, _03409_);
  and (_03473_, _03223_, _03193_);
  not (_03474_, _03473_);
  and (_03475_, _03188_, _03451_);
  not (_03476_, _03475_);
  and (_03478_, _03223_, _03188_);
  and (_03479_, _03478_, _03440_);
  not (_03480_, _03478_);
  nor (_03481_, _03368_, _42176_);
  nor (_03482_, _03404_, _42012_);
  nor (_03483_, _03482_, _03481_);
  nor (_03484_, _03378_, _42463_);
  nor (_03485_, _03386_, _42258_);
  nor (_03486_, _03485_, _03484_);
  and (_03487_, _03486_, _03483_);
  nor (_03488_, _03402_, _42135_);
  nor (_03489_, _03399_, _42094_);
  nor (_03490_, _03489_, _03488_);
  nor (_03491_, _03373_, _41963_);
  nor (_03492_, _03375_, _41915_);
  nor (_03493_, _03492_, _03491_);
  and (_03494_, _03493_, _03490_);
  and (_03495_, _03494_, _03487_);
  nor (_03496_, _03363_, _42422_);
  nor (_03497_, _03393_, _42340_);
  nor (_03498_, _03497_, _03496_);
  nor (_03499_, _03391_, _42504_);
  nor (_03500_, _03353_, _42381_);
  nor (_03501_, _03500_, _03499_);
  and (_03502_, _03501_, _03498_);
  nor (_03503_, _03388_, _42053_);
  nor (_03504_, _03358_, _41874_);
  nor (_03505_, _03504_, _03503_);
  nor (_03506_, _03381_, _42299_);
  nor (_03507_, _03397_, _42217_);
  nor (_03508_, _03507_, _03506_);
  and (_03509_, _03508_, _03505_);
  and (_03510_, _03509_, _03502_);
  and (_03511_, _03510_, _03495_);
  nor (_03512_, _03511_, _03409_);
  not (_03513_, _03440_);
  and (_03514_, _03513_, _03409_);
  nor (_03515_, _03514_, _03512_);
  and (_03516_, _03451_, _03167_);
  and (_03517_, _03158_, _03451_);
  nor (_03518_, _03517_, _03516_);
  not (_03519_, _03518_);
  and (_03520_, _03519_, _03515_);
  not (_03521_, _03224_);
  and (_03522_, _03444_, _03457_);
  nor (_03523_, _03458_, _03522_);
  nor (_03524_, _03523_, _03515_);
  and (_03525_, _03515_, _03469_);
  not (_03526_, \oc8051_golden_model_1.SP [3]);
  and (_03527_, _03444_, _03468_);
  and (_03528_, _03527_, _03526_);
  nor (_03529_, _03528_, _03525_);
  and (_03530_, _03223_, _03463_);
  not (_03531_, _03530_);
  nor (_03532_, _03527_, _03469_);
  not (_03533_, _03532_);
  and (_03534_, _03223_, _03468_);
  not (_03535_, _03208_);
  and (_03536_, _03223_, _03535_);
  nor (_03537_, _03536_, _03534_);
  and (_03538_, _03537_, \oc8051_golden_model_1.PSW [3]);
  or (_03539_, _03538_, _03533_);
  and (_03540_, _03539_, _03531_);
  and (_03541_, _03537_, _03531_);
  nor (_03542_, _03541_, _03440_);
  or (_03543_, _03542_, _03540_);
  and (_03544_, _03543_, _03466_);
  and (_03545_, _03544_, _03529_);
  nor (_03546_, _03515_, _03466_);
  and (_03547_, _03223_, _03457_);
  nor (_03548_, _03547_, _03464_);
  not (_03549_, _03548_);
  nor (_03550_, _03549_, _03546_);
  not (_03551_, _03550_);
  nor (_03552_, _03551_, _03545_);
  not (_03553_, _03523_);
  and (_03554_, _03549_, _03440_);
  or (_03555_, _03554_, _03553_);
  nor (_03556_, _03555_, _03552_);
  nor (_03557_, _03556_, _03524_);
  not (_03558_, _03213_);
  not (_03559_, _02923_);
  and (_03560_, _02954_, _03559_);
  and (_03561_, _03560_, _03443_);
  and (_03562_, _03561_, _03558_);
  not (_03563_, _03562_);
  and (_03564_, _03560_, _03450_);
  and (_03565_, _02954_, _02923_);
  and (_03566_, _03565_, _03443_);
  or (_03567_, _03566_, _03564_);
  and (_03568_, _03567_, _03558_);
  not (_03569_, _03568_);
  and (_03570_, _03565_, _03220_);
  and (_03571_, _03565_, _03017_);
  or (_03572_, _03571_, _03570_);
  and (_03573_, _03572_, _03558_);
  not (_03574_, _03573_);
  and (_03575_, _03560_, _03220_);
  and (_03576_, _03575_, _03558_);
  not (_03577_, _03231_);
  and (_03578_, _03560_, _03577_);
  and (_03579_, _03578_, _03558_);
  nor (_03580_, _03579_, _03576_);
  and (_03581_, _03580_, _03574_);
  and (_03582_, _03581_, _03569_);
  and (_03583_, _03582_, _03563_);
  not (_03584_, _03583_);
  nor (_03585_, _03584_, _03557_);
  and (_03586_, _03444_, _03558_);
  and (_03587_, _03558_, _03451_);
  nor (_03588_, _03587_, _03586_);
  not (_03589_, _03588_);
  nor (_03590_, _03583_, _03440_);
  nor (_03591_, _03590_, _03589_);
  not (_03592_, _03591_);
  nor (_03593_, _03592_, _03585_);
  and (_03594_, _03223_, _03218_);
  and (_03595_, _03589_, _03515_);
  nor (_03596_, _03595_, _03594_);
  not (_03597_, _03596_);
  nor (_03598_, _03597_, _03593_);
  not (_03599_, _03594_);
  nor (_03600_, _03599_, _03440_);
  or (_03601_, _03600_, _03598_);
  and (_03602_, _03601_, _03453_);
  nor (_03603_, _03515_, _03453_);
  or (_03604_, _03603_, _03602_);
  and (_03605_, _03604_, _03521_);
  and (_03606_, _03570_, _03457_);
  and (_03607_, _03443_, _03222_);
  and (_03608_, _03607_, _03457_);
  nor (_03609_, _03608_, _03606_);
  not (_03610_, _03232_);
  and (_03611_, _03610_, _03181_);
  and (_03612_, _03565_, _03450_);
  and (_03613_, _03612_, _03457_);
  nor (_03614_, _03613_, _03611_);
  and (_03615_, _03193_, _03451_);
  nor (_03616_, _03615_, _03445_);
  and (_03617_, _03444_, _03190_);
  and (_03618_, _03610_, _03177_);
  nor (_03619_, _03618_, _03617_);
  and (_03620_, _03619_, _03616_);
  and (_03621_, _03444_, _03218_);
  not (_03622_, _03621_);
  and (_03623_, _03610_, _03171_);
  and (_03624_, _03223_, _03167_);
  nor (_03625_, _03624_, _03623_);
  and (_03626_, _03625_, _03622_);
  and (_03627_, _03626_, _03620_);
  and (_03628_, _03627_, _03614_);
  and (_03629_, _03577_, _03222_);
  and (_03630_, _03629_, _03457_);
  not (_03631_, _03630_);
  and (_03632_, _03565_, _03577_);
  and (_03633_, _03632_, _03457_);
  nor (_03634_, _03633_, _03534_);
  and (_03635_, _03634_, _03631_);
  and (_03636_, _03635_, _03628_);
  and (_03637_, _03578_, _03457_);
  and (_03638_, _03567_, _03457_);
  nor (_03639_, _03638_, _03637_);
  and (_03640_, _03560_, _03230_);
  and (_03641_, _03640_, _03457_);
  not (_03642_, _03641_);
  and (_03643_, _03642_, _03639_);
  and (_03644_, _03444_, _03188_);
  and (_03645_, _03195_, _03451_);
  nor (_03646_, _03645_, _03644_);
  and (_03647_, _03222_, _03450_);
  and (_03648_, _03647_, _03457_);
  nor (_03649_, _03648_, _03547_);
  and (_03650_, _03649_, _03646_);
  and (_03651_, _03650_, _03643_);
  and (_03652_, _03651_, _03636_);
  and (_03653_, _03652_, _03609_);
  nor (_03654_, _03653_, _02897_);
  and (_03655_, _03653_, _02897_);
  nor (_03656_, _03655_, _03654_);
  nor (_03657_, _03655_, _02860_);
  and (_03658_, _03655_, _02860_);
  nor (_03659_, _03658_, _03657_);
  and (_03660_, _03659_, _03656_);
  nor (_03661_, _03653_, _03294_);
  and (_03662_, _03653_, _03299_);
  nor (_03663_, _03662_, _03661_);
  not (_03664_, _03663_);
  not (_03665_, _02866_);
  nor (_03666_, _03653_, _03665_);
  not (_03667_, _03257_);
  and (_03668_, _03653_, _03667_);
  nor (_03669_, _03668_, _03666_);
  nor (_03670_, _03669_, _03664_);
  and (_03671_, _03670_, _03660_);
  and (_03672_, _03671_, _02048_);
  nor (_03673_, _03659_, _03656_);
  and (_03674_, _03673_, _03670_);
  and (_03675_, _03674_, _02024_);
  nor (_03676_, _03675_, _03672_);
  not (_03677_, _03659_);
  nor (_03679_, _03677_, _03656_);
  and (_03680_, _03669_, _03663_);
  and (_03681_, _03680_, _03679_);
  and (_03682_, _03681_, _02040_);
  and (_03683_, _03669_, _03664_);
  and (_03684_, _03683_, _03679_);
  and (_03685_, _03684_, _02042_);
  nor (_03686_, _03685_, _03682_);
  and (_03687_, _03686_, _03676_);
  and (_03688_, _03680_, _03660_);
  and (_03689_, _03688_, _02030_);
  and (_03690_, _03680_, _03673_);
  and (_03691_, _03690_, _02032_);
  nor (_03692_, _03691_, _03689_);
  and (_03693_, _03677_, _03656_);
  and (_03694_, _03693_, _03683_);
  and (_03695_, _03694_, _02009_);
  and (_03696_, _03683_, _03660_);
  and (_03697_, _03696_, _02005_);
  nor (_03698_, _03697_, _03695_);
  and (_03699_, _03698_, _03692_);
  and (_03700_, _03699_, _03687_);
  nor (_03701_, _03669_, _03663_);
  and (_03702_, _03701_, _03660_);
  and (_03703_, _03702_, _02017_);
  and (_03704_, _03701_, _03693_);
  and (_03705_, _03704_, _02026_);
  nor (_03706_, _03705_, _03703_);
  and (_03707_, _03679_, _03670_);
  and (_03708_, _03707_, _02035_);
  and (_03709_, _03693_, _03670_);
  and (_03710_, _03709_, _02050_);
  nor (_03711_, _03710_, _03708_);
  and (_03712_, _03711_, _03706_);
  and (_03713_, _03693_, _03680_);
  and (_03714_, _03713_, _02003_);
  and (_03715_, _03683_, _03673_);
  and (_03716_, _03715_, _02012_);
  nor (_03717_, _03716_, _03714_);
  and (_03718_, _03701_, _03679_);
  and (_03719_, _03718_, _02037_);
  and (_03720_, _03701_, _03673_);
  and (_03721_, _03720_, _02020_);
  nor (_03722_, _03721_, _03719_);
  and (_03723_, _03722_, _03717_);
  and (_03724_, _03723_, _03712_);
  and (_03725_, _03724_, _03700_);
  nor (_03726_, _03725_, _03521_);
  nor (_03727_, _03726_, _03519_);
  not (_03728_, _03727_);
  nor (_03729_, _03728_, _03605_);
  or (_03730_, _03729_, _03520_);
  and (_03731_, _03223_, _03190_);
  not (_03732_, _03731_);
  and (_03733_, _03181_, _03451_);
  not (_03734_, _03733_);
  and (_03735_, _03223_, _03181_);
  nor (_03736_, _03735_, _03611_);
  and (_03737_, _03736_, _03734_);
  and (_03738_, _03737_, _03732_);
  and (_03739_, _03223_, _03177_);
  not (_03740_, _03739_);
  and (_03741_, _03177_, _03451_);
  nor (_03742_, _03741_, _03618_);
  and (_03743_, _03742_, _03740_);
  and (_03744_, _03171_, _03451_);
  not (_03745_, _03744_);
  and (_03746_, _03223_, _03171_);
  nor (_03747_, _03746_, _03623_);
  and (_03748_, _03747_, _03745_);
  and (_03749_, _03748_, _03743_);
  and (_03750_, _03749_, _03738_);
  nand (_03751_, _03750_, _03730_);
  and (_03752_, _03190_, _03451_);
  nor (_03753_, _03750_, _03513_);
  nor (_03754_, _03753_, _03752_);
  and (_03755_, _03754_, _03751_);
  and (_03756_, _03752_, \oc8051_golden_model_1.SP [3]);
  or (_03757_, _03756_, _03617_);
  nor (_03758_, _03757_, _03755_);
  and (_03759_, _03515_, _03617_);
  or (_03760_, _03759_, _03758_);
  and (_03761_, _03760_, _03480_);
  or (_03762_, _03761_, _03479_);
  nand (_03763_, _03762_, _03476_);
  and (_03764_, _03475_, _03526_);
  nor (_03765_, _03764_, _03644_);
  nand (_03766_, _03765_, _03763_);
  and (_03767_, _03223_, _03195_);
  not (_03768_, _03644_);
  nor (_03769_, _03768_, _03515_);
  nor (_03770_, _03769_, _03767_);
  nand (_03771_, _03770_, _03766_);
  and (_03772_, _03767_, _03440_);
  nor (_03773_, _03772_, _03445_);
  and (_03774_, _03773_, _03771_);
  nor (_03775_, _03446_, _03515_);
  or (_03776_, _03775_, _03774_);
  nand (_03777_, _03776_, _03474_);
  nor (_03778_, _03474_, _03440_);
  not (_03779_, _03778_);
  and (_03780_, _03779_, _03777_);
  nor (_03781_, _03391_, _42499_);
  nor (_03782_, _03404_, _42007_);
  nor (_03783_, _03782_, _03781_);
  nor (_03784_, _03378_, _42458_);
  nor (_03785_, _03397_, _42212_);
  nor (_03786_, _03785_, _03784_);
  and (_03787_, _03786_, _03783_);
  nor (_03788_, _03399_, _42089_);
  nor (_03789_, _03402_, _42130_);
  nor (_03790_, _03789_, _03788_);
  nor (_03791_, _03393_, _42335_);
  nor (_03792_, _03368_, _42171_);
  nor (_03793_, _03792_, _03791_);
  and (_03794_, _03793_, _03790_);
  and (_03795_, _03794_, _03787_);
  nor (_03796_, _03363_, _42417_);
  nor (_03797_, _03353_, _42376_);
  nor (_03798_, _03797_, _03796_);
  nor (_03799_, _03386_, _42253_);
  nor (_03800_, _03373_, _41957_);
  nor (_03801_, _03800_, _03799_);
  and (_03802_, _03801_, _03798_);
  nor (_03803_, _03381_, _42294_);
  nor (_03804_, _03388_, _42048_);
  nor (_03805_, _03804_, _03803_);
  nor (_03806_, _03358_, _41869_);
  nor (_03807_, _03375_, _41910_);
  nor (_03808_, _03807_, _03806_);
  and (_03809_, _03808_, _03805_);
  and (_03810_, _03809_, _03802_);
  and (_03811_, _03810_, _03795_);
  nor (_03812_, _03811_, _03409_);
  and (_03813_, _03588_, _03523_);
  not (_03814_, _03617_);
  nor (_03815_, _03465_, _03452_);
  and (_03816_, _03815_, _03814_);
  and (_03817_, _03816_, _03813_);
  nor (_03818_, _03644_, _03445_);
  and (_03819_, _03518_, _03470_);
  and (_03820_, _03819_, _03818_);
  and (_03821_, _03820_, _03817_);
  not (_03822_, _03821_);
  and (_03823_, _03822_, _03812_);
  not (_03824_, _03823_);
  and (_03825_, _03681_, _01985_);
  and (_03826_, _03684_, _01982_);
  nor (_03827_, _03826_, _03825_);
  and (_03828_, _03671_, _01964_);
  and (_03829_, _03720_, _01968_);
  nor (_03830_, _03829_, _03828_);
  and (_03831_, _03830_, _03827_);
  and (_03832_, _03688_, _01953_);
  and (_03833_, _03690_, _01947_);
  nor (_03834_, _03833_, _03832_);
  and (_03835_, _03696_, _01977_);
  and (_03836_, _03715_, _01975_);
  nor (_03837_, _03836_, _03835_);
  and (_03838_, _03837_, _03834_);
  and (_03839_, _03838_, _03831_);
  and (_03840_, _03674_, _01971_);
  and (_03841_, _03718_, _01987_);
  nor (_03842_, _03841_, _03840_);
  and (_03843_, _03707_, _01980_);
  and (_03844_, _03709_, _01994_);
  nor (_03845_, _03844_, _03843_);
  and (_03846_, _03845_, _03842_);
  and (_03847_, _03713_, _01949_);
  and (_03848_, _03694_, _01956_);
  nor (_03849_, _03848_, _03847_);
  and (_03850_, _03702_, _01961_);
  and (_03851_, _03704_, _01991_);
  nor (_03852_, _03851_, _03850_);
  and (_03853_, _03852_, _03849_);
  and (_03854_, _03853_, _03846_);
  and (_03855_, _03854_, _03839_);
  nor (_03856_, _03855_, _03521_);
  not (_03857_, \oc8051_golden_model_1.SP [2]);
  nor (_03858_, _03752_, _03475_);
  nor (_03859_, _03858_, _03857_);
  not (_03860_, _03859_);
  and (_03861_, _03571_, _03195_);
  and (_03862_, _03571_, _03463_);
  nor (_03863_, _03862_, _03861_);
  and (_03864_, _03565_, _03230_);
  and (_03865_, _03864_, _03463_);
  and (_03866_, _03864_, _03468_);
  nor (_03867_, _03866_, _03865_);
  and (_03868_, _03867_, _03863_);
  not (_03869_, _03571_);
  and (_03870_, _03206_, _03229_);
  nor (_03871_, _03158_, _03171_);
  and (_03872_, _03871_, _03870_);
  nor (_03873_, _03872_, _03869_);
  not (_03874_, _03873_);
  and (_03875_, _03874_, _03868_);
  and (_03876_, _03875_, _03860_);
  not (_03877_, _03864_);
  nor (_03878_, _03053_, _03164_);
  not (_03880_, _03878_);
  nor (_03881_, _03181_, _03188_);
  and (_03882_, _03881_, _03880_);
  and (_03883_, _03882_, _03871_);
  nor (_03884_, _03883_, _03877_);
  not (_03885_, _03884_);
  and (_03886_, _03527_, \oc8051_golden_model_1.SP [2]);
  not (_03887_, _03886_);
  and (_03888_, _03565_, _03535_);
  not (_03889_, _03888_);
  and (_03890_, _03571_, _03193_);
  and (_03891_, _03571_, _03188_);
  nor (_03892_, _03891_, _03890_);
  and (_03893_, _03892_, _03889_);
  and (_03894_, _03893_, _03887_);
  and (_03895_, _03571_, _03190_);
  and (_03896_, _03864_, _03193_);
  nor (_03897_, _03896_, _03895_);
  and (_03898_, _03571_, _03468_);
  and (_03899_, _03864_, _03218_);
  nor (_03900_, _03899_, _03898_);
  and (_03901_, _03900_, _03897_);
  and (_03902_, _03565_, _03177_);
  not (_03903_, _03902_);
  and (_03904_, _03571_, _03181_);
  and (_03905_, _03864_, _03195_);
  nor (_03906_, _03905_, _03904_);
  and (_03907_, _03906_, _03903_);
  and (_03908_, _03907_, _03901_);
  and (_03909_, _03908_, _03894_);
  and (_03910_, _03909_, _03885_);
  and (_03911_, _03910_, _03876_);
  not (_03912_, _03911_);
  nor (_03913_, _03912_, _03856_);
  nor (_03914_, _03402_, _42115_);
  nor (_03915_, _03399_, _42074_);
  nor (_03916_, _03915_, _03914_);
  nor (_03917_, _03391_, _42484_);
  nor (_03918_, _03393_, _42320_);
  nor (_03919_, _03918_, _03917_);
  and (_03920_, _03919_, _03916_);
  nor (_03921_, _03378_, _42443_);
  nor (_03922_, _03363_, _42402_);
  nor (_03923_, _03922_, _03921_);
  nor (_03924_, _03381_, _42279_);
  nor (_03925_, _03386_, _42238_);
  nor (_03926_, _03925_, _03924_);
  and (_03927_, _03926_, _03923_);
  and (_03928_, _03927_, _03920_);
  nor (_03929_, _03358_, _41854_);
  nor (_03930_, _03373_, _41936_);
  nor (_03931_, _03930_, _03929_);
  nor (_03932_, _03368_, _42156_);
  nor (_03933_, _03388_, _42033_);
  nor (_03934_, _03933_, _03932_);
  and (_03935_, _03934_, _03931_);
  nor (_03936_, _03353_, _42361_);
  nor (_03937_, _03397_, _42197_);
  nor (_03938_, _03937_, _03936_);
  nor (_03939_, _03404_, _41984_);
  nor (_03940_, _03375_, _41895_);
  nor (_03941_, _03940_, _03939_);
  and (_03942_, _03941_, _03938_);
  and (_03943_, _03942_, _03935_);
  and (_03944_, _03943_, _03928_);
  and (_03945_, _03599_, _03548_);
  and (_03946_, _03945_, _03541_);
  and (_03947_, _03946_, _03583_);
  not (_03948_, _03767_);
  nor (_03949_, _03478_, _03473_);
  and (_03950_, _03949_, _03948_);
  and (_03951_, _03950_, _03738_);
  and (_03952_, _03951_, _03749_);
  and (_03953_, _03952_, _03947_);
  nor (_03954_, _03953_, _03944_);
  not (_03955_, _03954_);
  and (_03956_, _03955_, _03913_);
  and (_03957_, _03956_, _03824_);
  not (_03958_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_03959_, _03393_, _42310_);
  or (_03960_, _03381_, _42269_);
  and (_03961_, _03960_, _03959_);
  or (_03962_, _03378_, _42433_);
  or (_03963_, _03353_, _42351_);
  and (_03964_, _03963_, _03962_);
  and (_03965_, _03964_, _03961_);
  or (_03966_, _03358_, _41844_);
  or (_03967_, _03375_, _41885_);
  and (_03968_, _03967_, _03966_);
  or (_03969_, _03399_, _42064_);
  or (_03970_, _03388_, _42023_);
  and (_03971_, _03970_, _03969_);
  and (_03972_, _03971_, _03968_);
  and (_03973_, _03972_, _03965_);
  or (_03974_, _03386_, _42228_);
  or (_03975_, _03397_, _42187_);
  and (_03976_, _03975_, _03974_);
  or (_03977_, _03391_, _42474_);
  or (_03978_, _03363_, _42392_);
  and (_03979_, _03978_, _03977_);
  and (_03980_, _03979_, _03976_);
  or (_03981_, _03368_, _42146_);
  or (_03982_, _03402_, _42105_);
  and (_03983_, _03982_, _03981_);
  or (_03984_, _03404_, _41974_);
  or (_03985_, _03373_, _41926_);
  and (_03986_, _03985_, _03984_);
  and (_03987_, _03986_, _03983_);
  and (_03988_, _03987_, _03980_);
  and (_03989_, _03988_, _03973_);
  nor (_03990_, _03989_, _03474_);
  not (_03991_, _03990_);
  nor (_03992_, _03989_, _03599_);
  nor (_03993_, _03588_, _03441_);
  not (_03994_, _03547_);
  nor (_03995_, _03989_, _03994_);
  or (_03996_, _03989_, _03531_);
  nor (_03997_, _03989_, _03537_);
  nor (_03998_, _03561_, _03223_);
  and (_03999_, _03565_, _02986_);
  nor (_04000_, _03999_, _03564_);
  nand (_04001_, _04000_, _03998_);
  and (_04002_, _04001_, _03535_);
  not (_04003_, _03203_);
  and (_04004_, _04003_, _03451_);
  and (_04005_, _03222_, _03017_);
  and (_04006_, _04005_, _04003_);
  and (_04007_, _04005_, _03535_);
  or (_04008_, _04007_, _04006_);
  and (_04009_, _04008_, _02986_);
  or (_04010_, _04009_, _04004_);
  nor (_04011_, _04010_, _04002_);
  and (_04012_, _04005_, _03468_);
  or (_04013_, _04012_, _03898_);
  nand (_04014_, _04013_, _02986_);
  and (_04015_, _03566_, _03468_);
  nor (_04016_, _04015_, _03534_);
  and (_04017_, _03535_, _03451_);
  and (_04018_, _03560_, _02986_);
  and (_04019_, _04018_, _03468_);
  nor (_04020_, _04019_, _04017_);
  and (_04021_, _04020_, _04016_);
  and (_04022_, _04021_, _04014_);
  and (_04023_, _04022_, _04011_);
  or (_04024_, _04023_, _03997_);
  nand (_04025_, _04024_, _03470_);
  nand (_04026_, _03471_, _04025_);
  and (_04027_, _03527_, _03455_);
  nor (_04028_, _04027_, _03530_);
  and (_04029_, _04005_, _03463_);
  and (_04030_, _04029_, _02986_);
  and (_04031_, _02986_, _02954_);
  and (_04032_, _04031_, _03463_);
  nor (_04033_, _04032_, _04030_);
  and (_04034_, _04033_, _04028_);
  nand (_04035_, _04034_, _04026_);
  nand (_04036_, _04035_, _03996_);
  and (_04037_, _04036_, _03466_);
  or (_04038_, _03467_, _04037_);
  and (_04039_, _03989_, _03464_);
  and (_04040_, _03561_, _03457_);
  not (_04041_, _04040_);
  and (_04042_, _03649_, _04041_);
  nor (_04043_, _03638_, _03613_);
  and (_04044_, _04043_, _04042_);
  not (_04045_, _04044_);
  nor (_04046_, _04045_, _04039_);
  and (_04047_, _04046_, _04038_);
  or (_04048_, _04047_, _03995_);
  nand (_04049_, _04048_, _03523_);
  nor (_04050_, _03523_, _03441_);
  nor (_04051_, _04050_, _03584_);
  nand (_04052_, _04051_, _04049_);
  and (_04053_, _03989_, _03584_);
  and (_04054_, _03647_, _03558_);
  not (_04055_, _04054_);
  and (_04056_, _04055_, _03588_);
  not (_04057_, _04056_);
  nor (_04058_, _04057_, _04053_);
  and (_04059_, _04058_, _04052_);
  or (_04060_, _04059_, _03993_);
  and (_04061_, _03566_, _03218_);
  not (_04062_, _04061_);
  and (_04063_, _03564_, _03218_);
  nor (_04064_, _04063_, _03594_);
  and (_04065_, _04064_, _04062_);
  and (_04066_, _04005_, _03218_);
  and (_04067_, _04066_, _02986_);
  nor (_04068_, _03612_, _03561_);
  nor (_04069_, _04068_, _03229_);
  nor (_04070_, _04069_, _04067_);
  and (_04071_, _04070_, _04065_);
  and (_04072_, _04071_, _04060_);
  or (_04073_, _04072_, _03992_);
  and (_04074_, _04073_, _03453_);
  or (_04075_, _04074_, _03454_);
  and (_04076_, _03564_, _03158_);
  not (_04077_, _04076_);
  and (_04078_, _03566_, _03158_);
  nor (_04079_, _04078_, _03224_);
  and (_04081_, _04079_, _04077_);
  and (_04082_, _04005_, _03158_);
  nand (_04083_, _04082_, _02986_);
  or (_04084_, _04068_, _03261_);
  and (_04085_, _04084_, _04083_);
  and (_04086_, _04085_, _04081_);
  and (_04087_, _04086_, _04075_);
  and (_04088_, _03671_, _01849_);
  and (_04089_, _03674_, _01856_);
  nor (_04090_, _04089_, _04088_);
  and (_04091_, _03713_, _01834_);
  and (_04092_, _03684_, _01867_);
  nor (_04093_, _04092_, _04091_);
  and (_04094_, _04093_, _04090_);
  and (_04095_, _03696_, _01844_);
  and (_04096_, _03715_, _01837_);
  nor (_04097_, _04096_, _04095_);
  and (_04098_, _03681_, _01864_);
  and (_04099_, _03690_, _01841_);
  nor (_04100_, _04099_, _04098_);
  and (_04101_, _04100_, _04097_);
  and (_04102_, _04101_, _04094_);
  and (_04103_, _03702_, _01878_);
  and (_04104_, _03704_, _01859_);
  nor (_04105_, _04104_, _04103_);
  and (_04106_, _03707_, _01870_);
  and (_04107_, _03709_, _01876_);
  nor (_04108_, _04107_, _04106_);
  and (_04109_, _04108_, _04105_);
  and (_04110_, _03688_, _01882_);
  and (_04111_, _03694_, _01884_);
  nor (_04112_, _04111_, _04110_);
  and (_04113_, _03718_, _01872_);
  and (_04114_, _03720_, _01852_);
  nor (_04115_, _04114_, _04113_);
  and (_04116_, _04115_, _04112_);
  and (_04117_, _04116_, _04109_);
  and (_04118_, _04117_, _04102_);
  nor (_04119_, _04118_, _03521_);
  or (_04120_, _04119_, _04087_);
  not (_04121_, _03516_);
  and (_04122_, _03517_, _03441_);
  and (_04123_, _03647_, _03167_);
  nor (_04124_, _04123_, _04122_);
  and (_04125_, _04124_, _04121_);
  and (_04126_, _04125_, _04120_);
  nor (_04127_, _04121_, _03441_);
  or (_04128_, _04127_, _04126_);
  and (_04129_, _03647_, _03171_);
  not (_04130_, _04129_);
  and (_04131_, _03564_, _03171_);
  and (_04132_, _03561_, _03171_);
  nor (_04133_, _04132_, _04131_);
  and (_04134_, _03999_, _03171_);
  not (_04135_, _04134_);
  and (_04136_, _04135_, _04133_);
  and (_04137_, _04136_, _04130_);
  and (_04138_, _04137_, _04128_);
  not (_04139_, _03989_);
  nor (_04140_, _04139_, _03748_);
  and (_04141_, _04005_, _03181_);
  nand (_04142_, _04141_, _02986_);
  and (_04143_, _03561_, _03181_);
  not (_04144_, _04143_);
  and (_04145_, _03564_, _03181_);
  and (_04146_, _03999_, _03181_);
  nor (_04147_, _04146_, _04145_);
  and (_04148_, _04147_, _04144_);
  and (_04149_, _04148_, _04142_);
  not (_04150_, _04149_);
  nor (_04151_, _04150_, _04140_);
  and (_04152_, _04151_, _04138_);
  nor (_04153_, _04139_, _03737_);
  and (_04154_, _03999_, _03177_);
  and (_04155_, _03564_, _03177_);
  and (_04156_, _03647_, _03177_);
  and (_04157_, _03561_, _03177_);
  or (_04158_, _04157_, _04156_);
  or (_04159_, _04158_, _04155_);
  nor (_04160_, _04159_, _04154_);
  not (_04161_, _04160_);
  nor (_04162_, _04161_, _04153_);
  and (_04163_, _04162_, _04152_);
  nor (_04164_, _04139_, _03743_);
  and (_04165_, _03647_, _03190_);
  not (_04166_, _03190_);
  not (_04167_, _03612_);
  and (_04168_, _03998_, _04167_);
  nor (_04169_, _04168_, _04166_);
  and (_04170_, _03567_, _03190_);
  or (_04171_, _04170_, _04169_);
  nor (_04172_, _04171_, _04165_);
  not (_04173_, _04172_);
  nor (_04174_, _04173_, _04164_);
  and (_04175_, _04174_, _04163_);
  nor (_04176_, _03989_, _03732_);
  or (_04177_, _04176_, _04175_);
  and (_04178_, _03752_, _03455_);
  nor (_04179_, _04178_, _03617_);
  and (_04180_, _04179_, _04177_);
  nor (_04182_, _03814_, _03441_);
  or (_04183_, _04182_, _04180_);
  and (_04184_, _04005_, _03188_);
  or (_04185_, _04184_, _03891_);
  nand (_04186_, _04185_, _02986_);
  nand (_04187_, _03567_, _03188_);
  and (_04188_, _03561_, _03188_);
  nor (_04189_, _04188_, _03478_);
  and (_04190_, _04189_, _04187_);
  and (_04191_, _04190_, _04186_);
  and (_04192_, _04191_, _04183_);
  nor (_04193_, _03989_, _03480_);
  or (_04194_, _04193_, _04192_);
  and (_04195_, _03475_, _03455_);
  nor (_04196_, _04195_, _03644_);
  and (_04197_, _04196_, _04194_);
  nor (_04198_, _03768_, _03441_);
  or (_04199_, _04198_, _04197_);
  and (_04200_, _03612_, _03195_);
  and (_04201_, _03647_, _03195_);
  nor (_04202_, _04201_, _04200_);
  and (_04203_, _03566_, _03195_);
  not (_04204_, _04203_);
  and (_04205_, _04018_, _03195_);
  nor (_04206_, _04205_, _03767_);
  and (_04207_, _04206_, _04204_);
  and (_04208_, _04207_, _04202_);
  and (_04209_, _04208_, _04199_);
  nor (_04210_, _03989_, _03948_);
  or (_04211_, _04210_, _04209_);
  and (_04212_, _04211_, _03446_);
  or (_04213_, _03447_, _04212_);
  and (_04214_, _03612_, _03193_);
  and (_04215_, _04005_, _03193_);
  and (_04216_, _04215_, _02986_);
  nor (_04217_, _04216_, _04214_);
  and (_04218_, _03566_, _03193_);
  not (_04219_, _04218_);
  and (_04220_, _04018_, _03193_);
  nor (_04221_, _04220_, _03473_);
  and (_04222_, _04221_, _04219_);
  and (_04223_, _04222_, _04217_);
  nand (_04224_, _04223_, _04213_);
  nand (_04225_, _04224_, _03991_);
  or (_04226_, _04225_, _03958_);
  nor (_04227_, _03391_, _42494_);
  nor (_04228_, _03399_, _42084_);
  nor (_04229_, _04228_, _04227_);
  nor (_04230_, _03378_, _42453_);
  nor (_04231_, _03397_, _42207_);
  nor (_04232_, _04231_, _04230_);
  and (_04233_, _04232_, _04229_);
  nor (_04234_, _03375_, _41905_);
  nor (_04235_, _03373_, _41947_);
  nor (_04236_, _04235_, _04234_);
  nor (_04237_, _03393_, _42330_);
  nor (_04238_, _03404_, _42000_);
  nor (_04239_, _04238_, _04237_);
  and (_04240_, _04239_, _04236_);
  and (_04241_, _04240_, _04233_);
  nor (_04242_, _03363_, _42412_);
  nor (_04243_, _03353_, _42371_);
  nor (_04244_, _04243_, _04242_);
  nor (_04245_, _03386_, _42248_);
  nor (_04246_, _03368_, _42166_);
  nor (_04247_, _04246_, _04245_);
  and (_04248_, _04247_, _04244_);
  nor (_04249_, _03381_, _42289_);
  nor (_04250_, _03402_, _42125_);
  nor (_04251_, _04250_, _04249_);
  nor (_04252_, _03388_, _42043_);
  nor (_04253_, _03358_, _41864_);
  nor (_04254_, _04253_, _04252_);
  and (_04255_, _04254_, _04251_);
  and (_04256_, _04255_, _04248_);
  and (_04257_, _04256_, _04241_);
  nor (_04258_, _04257_, _03409_);
  and (_04259_, _04258_, _03822_);
  not (_04260_, _04259_);
  nor (_04261_, _03391_, _42479_);
  nor (_04262_, _03388_, _42028_);
  nor (_04263_, _04262_, _04261_);
  nor (_04264_, _03378_, _42438_);
  nor (_04265_, _03386_, _42233_);
  nor (_04266_, _04265_, _04264_);
  and (_04267_, _04266_, _04263_);
  nor (_04268_, _03375_, _41890_);
  nor (_04269_, _03373_, _41931_);
  nor (_04270_, _04269_, _04268_);
  nor (_04271_, _03393_, _42315_);
  nor (_04272_, _03404_, _41979_);
  nor (_04273_, _04272_, _04271_);
  and (_04274_, _04273_, _04270_);
  and (_04275_, _04274_, _04267_);
  nor (_04276_, _03368_, _42151_);
  nor (_04277_, _03397_, _42192_);
  nor (_04278_, _04277_, _04276_);
  nor (_04279_, _03363_, _42397_);
  nor (_04280_, _03353_, _42356_);
  nor (_04281_, _04280_, _04279_);
  and (_04283_, _04281_, _04278_);
  nor (_04284_, _03381_, _42274_);
  nor (_04285_, _03402_, _42110_);
  nor (_04286_, _04285_, _04284_);
  nor (_04287_, _03399_, _42069_);
  nor (_04288_, _03358_, _41849_);
  nor (_04289_, _04288_, _04287_);
  and (_04290_, _04289_, _04286_);
  and (_04291_, _04290_, _04283_);
  and (_04292_, _04291_, _04275_);
  nor (_04293_, _04292_, _03953_);
  not (_04294_, _04293_);
  and (_04295_, _03707_, _01925_);
  and (_04296_, _03718_, _01927_);
  nor (_04297_, _04296_, _04295_);
  and (_04298_, _03681_, _01930_);
  and (_04299_, _03713_, _01900_);
  nor (_04300_, _04299_, _04298_);
  and (_04301_, _04300_, _04297_);
  and (_04302_, _03702_, _01905_);
  and (_04303_, _03720_, _01908_);
  nor (_04304_, _04303_, _04302_);
  and (_04305_, _03674_, _01912_);
  and (_04306_, _03709_, _01938_);
  nor (_04307_, _04306_, _04305_);
  and (_04308_, _04307_, _04304_);
  and (_04309_, _04308_, _04301_);
  and (_04310_, _03688_, _01893_);
  and (_04311_, _03690_, _01891_);
  nor (_04312_, _04311_, _04310_);
  and (_04313_, _03694_, _01897_);
  and (_04314_, _03696_, _01922_);
  nor (_04315_, _04314_, _04313_);
  and (_04316_, _04315_, _04312_);
  and (_04317_, _03671_, _01936_);
  and (_04318_, _03704_, _01915_);
  nor (_04319_, _04318_, _04317_);
  and (_04320_, _03684_, _01932_);
  and (_04321_, _03715_, _01920_);
  nor (_04322_, _04321_, _04320_);
  and (_04323_, _04322_, _04319_);
  and (_04324_, _04323_, _04316_);
  and (_04325_, _04324_, _04309_);
  nor (_04326_, _04325_, _03521_);
  and (_04327_, _03560_, _03017_);
  and (_04328_, _04327_, _03195_);
  not (_04329_, _04328_);
  and (_04330_, _04327_, _03171_);
  and (_04331_, _04327_, _03468_);
  nor (_04332_, _04331_, _04330_);
  and (_04333_, _04332_, _04329_);
  and (_04334_, _03571_, _03177_);
  and (_04335_, _04327_, _03218_);
  nor (_04336_, _04335_, _04334_);
  and (_04337_, _04327_, _03158_);
  and (_04338_, _04327_, _03193_);
  nor (_04339_, _04338_, _04337_);
  and (_04340_, _04339_, _04336_);
  and (_04341_, _04340_, _04333_);
  not (_04342_, \oc8051_golden_model_1.SP [1]);
  nor (_04343_, _03858_, _04342_);
  nor (_04344_, _04343_, _03873_);
  and (_04345_, _04344_, _04341_);
  nor (_04346_, _04327_, _03571_);
  nor (_04347_, _04346_, _03208_);
  not (_04348_, _04327_);
  nor (_04349_, _03181_, _03177_);
  nor (_04350_, _04349_, _04348_);
  nor (_04351_, _04350_, _04347_);
  and (_04352_, _03527_, \oc8051_golden_model_1.SP [1]);
  and (_04353_, _03187_, _03156_);
  nor (_04354_, _04353_, _03457_);
  nor (_04355_, _04354_, _04348_);
  nor (_04356_, _04355_, _04352_);
  and (_04357_, _04356_, _04351_);
  nor (_04358_, _03904_, _03895_);
  and (_04359_, _04327_, _03463_);
  nor (_04360_, _04359_, _03898_);
  and (_04361_, _04360_, _04358_);
  and (_04362_, _03892_, _03863_);
  and (_04363_, _04362_, _04361_);
  and (_04364_, _04363_, _04357_);
  and (_04365_, _04364_, _04345_);
  not (_04366_, _04365_);
  nor (_04367_, _04366_, _04326_);
  and (_04368_, _04367_, _04294_);
  and (_04369_, _04368_, _04260_);
  not (_04370_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04371_, _04224_, _03991_);
  or (_04372_, _04371_, _04370_);
  and (_04373_, _04372_, _04369_);
  nand (_04374_, _04373_, _04226_);
  not (_04375_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_04376_, _04371_, _04375_);
  not (_04377_, _04369_);
  not (_04378_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_04379_, _04225_, _04378_);
  and (_04380_, _04379_, _04377_);
  nand (_04381_, _04380_, _04376_);
  nand (_04382_, _04381_, _04374_);
  nand (_04384_, _04382_, _03957_);
  not (_04385_, _03957_);
  not (_04386_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_04387_, _04371_, _04386_);
  not (_04388_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_04389_, _04225_, _04388_);
  and (_04390_, _04389_, _04377_);
  nand (_04391_, _04390_, _04387_);
  not (_04392_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_04393_, _04225_, _04392_);
  not (_04394_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_04395_, _04371_, _04394_);
  and (_04396_, _04395_, _04369_);
  nand (_04397_, _04396_, _04393_);
  nand (_04398_, _04397_, _04391_);
  nand (_04399_, _04398_, _04385_);
  nand (_04400_, _04399_, _04384_);
  nand (_04401_, _04400_, _03780_);
  not (_04402_, _03780_);
  not (_04403_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_04404_, _04371_, _04403_);
  nand (_04405_, _04371_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04406_, _04405_, _04377_);
  nand (_04407_, _04406_, _04404_);
  not (_04408_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_04409_, _04225_, _04408_);
  nand (_04410_, _04225_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04411_, _04410_, _04369_);
  nand (_04412_, _04411_, _04409_);
  nand (_04413_, _04412_, _04407_);
  nand (_04414_, _04413_, _03957_);
  not (_04415_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_04416_, _04371_, _04415_);
  nand (_04417_, _04371_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04418_, _04417_, _04377_);
  nand (_04419_, _04418_, _04416_);
  not (_04420_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_04421_, _04225_, _04420_);
  nand (_04422_, _04225_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04423_, _04422_, _04369_);
  nand (_04424_, _04423_, _04421_);
  nand (_04425_, _04424_, _04419_);
  nand (_04426_, _04425_, _04385_);
  nand (_04427_, _04426_, _04414_);
  nand (_04428_, _04427_, _04402_);
  and (_04429_, _04428_, _04401_);
  nor (_04430_, _04012_, _04006_);
  or (_04431_, _04430_, _04429_);
  not (_04432_, _03534_);
  nor (_04433_, _04432_, _03409_);
  not (_04434_, _04433_);
  not (_04435_, _03204_);
  and (_04436_, _03223_, _04003_);
  not (_04437_, _04436_);
  nor (_04438_, _04437_, _03409_);
  and (_04439_, _04438_, _04139_);
  or (_04440_, _04439_, _04435_);
  and (_04441_, _04031_, _04003_);
  nor (_04442_, _04441_, _04438_);
  or (_04443_, _04442_, _04440_);
  nor (_04444_, _03204_, _03455_);
  and (_04445_, _04031_, _03468_);
  nor (_04446_, _04445_, _04444_);
  and (_04447_, _04446_, _04443_);
  and (_04448_, _04447_, _04434_);
  and (_04449_, _04448_, _04431_);
  and (_04450_, _04433_, _04139_);
  nor (_04451_, _04450_, _04449_);
  nor (_04452_, _04451_, _03472_);
  not (_04453_, _04452_);
  and (_04454_, _04453_, _03471_);
  nor (_04455_, _03202_, _03455_);
  nor (_04456_, _04455_, _04454_);
  not (_04457_, _03527_);
  nor (_04458_, _04457_, _03409_);
  and (_04459_, _04458_, _03989_);
  nor (_04460_, _04459_, _04032_);
  and (_04461_, _04460_, _04456_);
  nand (_04462_, _04428_, _04401_);
  and (_04463_, _04462_, _04029_);
  not (_04464_, _04463_);
  and (_04465_, _04464_, _04461_);
  nor (_04466_, _03466_, _03409_);
  nor (_04467_, _03531_, _03409_);
  and (_04468_, _04467_, _03989_);
  nor (_04469_, _04468_, _04466_);
  and (_04470_, _04469_, _04465_);
  nor (_04471_, _04470_, _03467_);
  nor (_04472_, _04471_, _03464_);
  and (_04473_, _03464_, _03455_);
  or (_04474_, _04473_, _04472_);
  and (_04475_, _04474_, _03462_);
  nor (_04476_, _04475_, _03460_);
  and (_04477_, _04031_, _03558_);
  or (_04478_, _04477_, _04476_);
  nor (_04479_, _04478_, _03456_);
  nor (_04480_, _03409_, _03453_);
  and (_04481_, _04005_, _03558_);
  and (_04482_, _04462_, _04481_);
  nor (_04483_, _04482_, _04480_);
  and (_04485_, _04483_, _04479_);
  nor (_04486_, _04485_, _03454_);
  nor (_04487_, _04486_, _03219_);
  and (_04488_, _03219_, _03455_);
  nor (_04489_, _04488_, _04487_);
  nor (_04490_, _03409_, _03261_);
  and (_04491_, _04490_, _03572_);
  not (_04492_, _04491_);
  not (_04493_, _03409_);
  and (_04494_, _04337_, _04493_);
  and (_04495_, _03640_, _03158_);
  or (_04496_, _04495_, _04078_);
  and (_04497_, _04496_, _04493_);
  nor (_04498_, _04497_, _04494_);
  and (_04499_, _04498_, _04492_);
  not (_04500_, _04082_);
  nor (_04501_, _04500_, _03409_);
  and (_04502_, _04490_, _03223_);
  nor (_04503_, _04502_, _04501_);
  and (_04504_, _04503_, _04499_);
  nor (_04505_, _04504_, _04139_);
  nor (_04506_, _04505_, _04489_);
  and (_04507_, _04005_, _03167_);
  and (_04508_, _04462_, _04507_);
  not (_04509_, _03624_);
  nor (_04510_, _04509_, _03409_);
  and (_04511_, _04031_, _03167_);
  nor (_04512_, _04511_, _04510_);
  not (_04513_, _04512_);
  nor (_04514_, _04513_, _04508_);
  and (_04515_, _04514_, _04506_);
  and (_04516_, _04510_, _04139_);
  nor (_04517_, _04516_, _04515_);
  nor (_04518_, _04517_, _03168_);
  and (_04519_, _03168_, _03455_);
  nor (_04520_, _04519_, _04518_);
  nor (_04521_, _03734_, _03409_);
  not (_04522_, _04521_);
  not (_04523_, _03611_);
  nor (_04524_, _04523_, _03409_);
  not (_04525_, _04524_);
  nor (_04526_, _03745_, _03409_);
  not (_04527_, _03623_);
  nor (_04528_, _04527_, _03409_);
  nor (_04529_, _04528_, _04526_);
  and (_04530_, _04529_, _04525_);
  and (_04531_, _04530_, _04522_);
  nor (_04532_, _04531_, _04139_);
  nor (_04533_, _04532_, _03182_);
  not (_04534_, _04533_);
  nor (_04535_, _04534_, _04520_);
  and (_04536_, _03182_, _03455_);
  nor (_04537_, _04536_, _04535_);
  nor (_04538_, _03742_, _03409_);
  and (_04539_, _04538_, _03989_);
  or (_04540_, _04539_, _03191_);
  nor (_04541_, _04540_, _04537_);
  and (_04542_, _03191_, _03455_);
  nor (_04543_, _04542_, _04541_);
  and (_04544_, _04005_, _03195_);
  and (_04545_, _04462_, _04544_);
  nor (_04546_, _03948_, _03409_);
  and (_04547_, _04031_, _03195_);
  or (_04548_, _04547_, _04546_);
  or (_04549_, _04548_, _04545_);
  nor (_04550_, _04549_, _04543_);
  and (_04551_, _04546_, _04139_);
  nor (_04552_, _04551_, _04550_);
  nor (_04553_, _03645_, _03196_);
  nor (_04554_, _04553_, _03455_);
  nor (_04555_, _04554_, _04552_);
  and (_04556_, _04555_, _03449_);
  nor (_04557_, _04556_, _03447_);
  and (_04558_, _04462_, _04215_);
  nor (_04559_, _03474_, _03409_);
  and (_04560_, _04031_, _03193_);
  or (_04561_, _04560_, _04559_);
  or (_04562_, _04561_, _04558_);
  nor (_04563_, _04562_, _04557_);
  and (_04564_, _04559_, _04139_);
  nor (_04565_, _04564_, _04563_);
  not (_04566_, _04292_);
  and (_04567_, _04559_, _04566_);
  and (_04568_, _04258_, _03445_);
  and (_04569_, _04342_, \oc8051_golden_model_1.SP [0]);
  and (_04570_, \oc8051_golden_model_1.SP [1], _03455_);
  nor (_04571_, _04570_, _04569_);
  not (_04572_, _04571_);
  and (_04573_, _04572_, _03191_);
  and (_04574_, _04510_, _04566_);
  and (_04575_, _04258_, _03452_);
  and (_04576_, _04572_, _03464_);
  not (_04577_, _03464_);
  not (_04578_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_04579_, _04225_, _04578_);
  not (_04580_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_04581_, _04371_, _04580_);
  and (_04582_, _04581_, _04369_);
  nand (_04583_, _04582_, _04579_);
  not (_04584_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_04586_, _04371_, _04584_);
  not (_04587_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04588_, _04225_, _04587_);
  and (_04589_, _04588_, _04377_);
  nand (_04590_, _04589_, _04586_);
  nand (_04591_, _04590_, _04583_);
  nand (_04592_, _04591_, _03957_);
  not (_04593_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_04594_, _04371_, _04593_);
  not (_04595_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04596_, _04225_, _04595_);
  and (_04597_, _04596_, _04377_);
  nand (_04598_, _04597_, _04594_);
  not (_04599_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04600_, _04225_, _04599_);
  not (_04601_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_04602_, _04371_, _04601_);
  and (_04603_, _04602_, _04369_);
  nand (_04604_, _04603_, _04600_);
  nand (_04605_, _04604_, _04598_);
  nand (_04606_, _04605_, _04385_);
  nand (_04607_, _04606_, _04592_);
  nand (_04608_, _04607_, _03780_);
  not (_04609_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_04610_, _04371_, _04609_);
  nand (_04611_, _04371_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04612_, _04611_, _04377_);
  nand (_04613_, _04612_, _04610_);
  not (_04614_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_04615_, _04225_, _04614_);
  nand (_04616_, _04225_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04617_, _04616_, _04369_);
  nand (_04618_, _04617_, _04615_);
  nand (_04619_, _04618_, _04613_);
  nand (_04620_, _04619_, _03957_);
  not (_04621_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_04622_, _04371_, _04621_);
  nand (_04623_, _04371_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04624_, _04623_, _04377_);
  nand (_04625_, _04624_, _04622_);
  not (_04626_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_04627_, _04225_, _04626_);
  nand (_04628_, _04225_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04629_, _04628_, _04369_);
  nand (_04630_, _04629_, _04627_);
  nand (_04631_, _04630_, _04625_);
  nand (_04632_, _04631_, _04385_);
  nand (_04633_, _04632_, _04620_);
  nand (_04634_, _04633_, _04402_);
  nand (_04635_, _04634_, _04608_);
  not (_04636_, _04635_);
  or (_04637_, _04636_, _04430_);
  and (_04638_, _03230_, _02954_);
  and (_04639_, _04638_, _04003_);
  nor (_04640_, _04639_, _04438_);
  and (_04641_, _04438_, _04566_);
  or (_04642_, _04641_, _04435_);
  or (_04643_, _04642_, _04640_);
  and (_04644_, _03575_, _03468_);
  and (_04645_, _04019_, _03230_);
  nor (_04646_, _04645_, _04644_);
  nor (_04647_, _04572_, _03204_);
  nor (_04648_, _04647_, _03866_);
  and (_04649_, _04648_, _04646_);
  and (_04650_, _04649_, _04643_);
  and (_04651_, _04650_, _04434_);
  and (_04652_, _04651_, _04637_);
  and (_04653_, _04433_, _04566_);
  nor (_04654_, _04653_, _04652_);
  and (_04655_, _04257_, _03472_);
  nor (_04656_, _04655_, _04654_);
  or (_04657_, _04572_, _03202_);
  nand (_04658_, _04657_, _04656_);
  and (_04659_, _04458_, _04292_);
  and (_04660_, _03575_, _03463_);
  not (_04661_, _04660_);
  and (_04662_, _03561_, _03463_);
  nor (_04663_, _04662_, _03865_);
  and (_04664_, _04663_, _04661_);
  not (_04665_, _04664_);
  nor (_04666_, _04665_, _04659_);
  not (_04667_, _04666_);
  nor (_04668_, _04667_, _04658_);
  and (_04669_, _04635_, _04029_);
  nor (_04670_, _04669_, _04467_);
  and (_04671_, _04670_, _04668_);
  and (_04672_, _04467_, _04566_);
  nor (_04673_, _04672_, _04671_);
  and (_04674_, _04257_, _04466_);
  nor (_04675_, _04674_, _04673_);
  and (_04676_, _04675_, _04577_);
  nor (_04677_, _04676_, _04576_);
  and (_04678_, _03461_, _04257_);
  or (_04679_, _04678_, _04677_);
  nor (_04680_, _04572_, _03207_);
  not (_04681_, _04680_);
  and (_04682_, _03640_, _03558_);
  and (_04683_, _03864_, _03558_);
  nor (_04684_, _04683_, _04682_);
  and (_04685_, _04684_, _04681_);
  not (_04687_, _04685_);
  nor (_04688_, _04687_, _04679_);
  and (_04689_, _04635_, _04481_);
  nor (_04690_, _04689_, _04480_);
  and (_04691_, _04690_, _04688_);
  nor (_04692_, _04691_, _04575_);
  nor (_04693_, _04692_, _03219_);
  and (_04694_, _04572_, _03219_);
  nor (_04695_, _04694_, _04693_);
  nor (_04696_, _04504_, _04566_);
  and (_04697_, _04638_, _03167_);
  nor (_04698_, _04697_, _04696_);
  not (_04699_, _04698_);
  nor (_04700_, _04699_, _04695_);
  and (_04701_, _04635_, _04507_);
  nor (_04702_, _04701_, _04510_);
  and (_04703_, _04702_, _04700_);
  nor (_04704_, _04703_, _04574_);
  nor (_04705_, _04704_, _03168_);
  and (_04706_, _04572_, _03168_);
  nor (_04707_, _04706_, _04705_);
  nor (_04708_, _04531_, _04566_);
  nor (_04709_, _04708_, _03182_);
  not (_04710_, _04709_);
  nor (_04711_, _04710_, _04707_);
  and (_04712_, _04572_, _03182_);
  nor (_04713_, _04712_, _04711_);
  and (_04714_, _04538_, _04292_);
  or (_04715_, _04714_, _03191_);
  nor (_04716_, _04715_, _04713_);
  nor (_04717_, _04716_, _04573_);
  not (_04718_, _03905_);
  and (_04719_, _03561_, _03195_);
  and (_04720_, _03575_, _03195_);
  nor (_04721_, _04720_, _04719_);
  nand (_04722_, _04721_, _04718_);
  nor (_04723_, _04722_, _04717_);
  and (_04724_, _04635_, _04544_);
  nor (_04725_, _04724_, _04546_);
  and (_04726_, _04725_, _04723_);
  and (_04727_, _04546_, _04566_);
  nor (_04728_, _04727_, _04726_);
  nor (_04729_, _04572_, _04553_);
  nor (_04730_, _04729_, _03448_);
  not (_04731_, _04730_);
  nor (_04732_, _04731_, _04728_);
  nor (_04733_, _04732_, _04568_);
  and (_04734_, _03561_, _03193_);
  and (_04735_, _03575_, _03193_);
  nor (_04736_, _04735_, _04734_);
  not (_04737_, _04736_);
  nor (_04738_, _04737_, _03896_);
  not (_04739_, _04738_);
  nor (_04740_, _04739_, _04733_);
  and (_04741_, _04635_, _04215_);
  nor (_04742_, _04741_, _04559_);
  and (_04743_, _04742_, _04740_);
  nor (_04744_, _04743_, _04567_);
  not (_04745_, _00001_);
  not (_04746_, _04559_);
  nor (_04747_, _04546_, _03448_);
  and (_04748_, _04747_, _04746_);
  nor (_04749_, _03461_, _04480_);
  nor (_04750_, _04521_, _04510_);
  and (_04751_, _04750_, _04749_);
  and (_04752_, _04751_, _04748_);
  and (_04753_, _04752_, _04530_);
  not (_04754_, _04502_);
  not (_04755_, _03207_);
  or (_04756_, _04755_, _03219_);
  not (_04757_, _04756_);
  and (_04758_, _04757_, _04553_);
  nor (_04759_, _03182_, _03168_);
  and (_04760_, _03569_, _04759_);
  and (_04761_, _04760_, _04758_);
  nor (_04762_, _04029_, _03579_);
  nor (_04763_, _03905_, _03573_);
  and (_04764_, _04763_, _04762_);
  nor (_04765_, _04544_, _04507_);
  nor (_04766_, _04481_, _03464_);
  and (_04767_, _04766_, _04765_);
  and (_04768_, _04767_, _04764_);
  and (_04769_, _04768_, _04761_);
  nor (_04770_, _04331_, _03898_);
  and (_04771_, _03565_, _04003_);
  not (_04772_, _04771_);
  and (_04773_, _04772_, _04770_);
  nor (_04774_, _04660_, _04359_);
  not (_04775_, _04774_);
  not (_04776_, _03443_);
  and (_04777_, _03560_, _03167_);
  and (_04778_, _04777_, _04776_);
  nor (_04779_, _04778_, _04775_);
  and (_04780_, _04779_, _04773_);
  nor (_04781_, _04734_, _04216_);
  and (_04782_, _03561_, _03167_);
  and (_04783_, _03629_, _03193_);
  nor (_04784_, _04783_, _04782_);
  and (_04785_, _04784_, _04781_);
  and (_04786_, _04785_, _04780_);
  and (_04788_, _04786_, _04769_);
  nor (_04789_, _04735_, _04338_);
  and (_04790_, _04789_, _04219_);
  and (_04791_, _04790_, _04646_);
  and (_04792_, _04791_, _04721_);
  and (_04793_, _03565_, _03167_);
  nor (_04794_, _04793_, _04662_);
  and (_04795_, _03572_, _03193_);
  and (_04796_, _03560_, _04003_);
  nor (_04797_, _04796_, _04795_);
  and (_04798_, _04797_, _04794_);
  nor (_04799_, _04328_, _04012_);
  nor (_04800_, _04682_, _04006_);
  and (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04798_);
  not (_04803_, _03191_);
  and (_04804_, _03205_, _04803_);
  and (_04805_, _04804_, _03868_);
  and (_04806_, _04805_, _04802_);
  and (_04807_, _04806_, _04792_);
  and (_04808_, _04807_, _04788_);
  not (_04809_, _04808_);
  nor (_04810_, _04809_, _04538_);
  and (_04811_, _04810_, _04754_);
  nor (_04812_, _04494_, _04491_);
  and (_04813_, _04812_, _04811_);
  nor (_04814_, _04458_, _03472_);
  nor (_04815_, _04438_, _04433_);
  and (_04816_, _04815_, _04814_);
  nor (_04817_, _04501_, _04497_);
  nor (_04818_, _04467_, _04466_);
  and (_04819_, _04818_, _04817_);
  and (_04820_, _04819_, _04816_);
  and (_04821_, _04820_, _04813_);
  and (_04822_, _04821_, _04753_);
  nor (_04823_, _04822_, _04745_);
  not (_04824_, _04823_);
  nor (_04825_, _04824_, _04744_);
  not (_04826_, _04825_);
  nor (_04827_, _04826_, _04565_);
  and (_04828_, _04559_, _03513_);
  not (_04829_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04830_, _04225_, _04829_);
  not (_04831_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_04832_, _04371_, _04831_);
  and (_04833_, _04832_, _04369_);
  nand (_04834_, _04833_, _04830_);
  not (_04835_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_04836_, _04371_, _04835_);
  not (_04837_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04838_, _04225_, _04837_);
  and (_04839_, _04838_, _04377_);
  nand (_04840_, _04839_, _04836_);
  nand (_04841_, _04840_, _04834_);
  nand (_04842_, _04841_, _03957_);
  not (_04843_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04844_, _04371_, _04843_);
  not (_04845_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04846_, _04225_, _04845_);
  and (_04847_, _04846_, _04377_);
  nand (_04848_, _04847_, _04844_);
  not (_04849_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04850_, _04225_, _04849_);
  not (_04851_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04852_, _04371_, _04851_);
  and (_04853_, _04852_, _04369_);
  nand (_04854_, _04853_, _04850_);
  nand (_04855_, _04854_, _04848_);
  nand (_04856_, _04855_, _04385_);
  nand (_04857_, _04856_, _04842_);
  nand (_04858_, _04857_, _03780_);
  not (_04859_, \oc8051_golden_model_1.IRAM[11] [3]);
  or (_04860_, _04371_, _04859_);
  not (_04861_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_04862_, _04225_, _04861_);
  and (_04863_, _04862_, _04377_);
  nand (_04864_, _04863_, _04860_);
  nand (_04865_, _04371_, \oc8051_golden_model_1.IRAM[8] [3]);
  not (_04866_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_04867_, _04371_, _04866_);
  and (_04868_, _04867_, _04369_);
  nand (_04869_, _04868_, _04865_);
  nand (_04870_, _04869_, _04864_);
  nand (_04871_, _04870_, _03957_);
  nand (_04872_, _04225_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04873_, _04371_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04874_, _04873_, _04377_);
  nand (_04875_, _04874_, _04872_);
  not (_04876_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_04877_, _04225_, _04876_);
  nand (_04878_, _04225_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04879_, _04878_, _04369_);
  nand (_04880_, _04879_, _04877_);
  nand (_04881_, _04880_, _04875_);
  nand (_04882_, _04881_, _04385_);
  nand (_04883_, _04882_, _04871_);
  nand (_04884_, _04883_, _04402_);
  nand (_04885_, _04884_, _04858_);
  and (_04886_, _04885_, _04507_);
  and (_04887_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04888_, _04887_, \oc8051_golden_model_1.SP [2]);
  or (_04889_, _04888_, \oc8051_golden_model_1.SP [3]);
  and (_04890_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04891_, _04890_, \oc8051_golden_model_1.SP [3]);
  nand (_04892_, _04891_, \oc8051_golden_model_1.SP [0]);
  and (_04893_, _04892_, _04889_);
  not (_04894_, _04893_);
  nor (_04895_, _04894_, _03207_);
  not (_04896_, _04458_);
  and (_04897_, _03511_, _03472_);
  and (_04898_, _04885_, _04012_);
  nor (_04899_, _04894_, _03204_);
  nor (_04900_, _04006_, \oc8051_golden_model_1.PSW [3]);
  and (_04901_, _04885_, _04006_);
  nor (_04902_, _04901_, _04900_);
  nor (_04903_, _04902_, _04438_);
  and (_04904_, _04438_, _03440_);
  nor (_04905_, _04904_, _04435_);
  not (_04906_, _04905_);
  nor (_04907_, _04906_, _04903_);
  or (_04908_, _04907_, _04012_);
  nor (_04909_, _04908_, _04899_);
  or (_04910_, _04909_, _04433_);
  nor (_04911_, _04910_, _04898_);
  and (_04912_, _04433_, _03513_);
  or (_04913_, _04912_, _03472_);
  nor (_04914_, _04913_, _04911_);
  nor (_04915_, _04914_, _04897_);
  and (_04916_, _04915_, _03202_);
  nor (_04917_, _04894_, _03202_);
  or (_04918_, _04917_, _04916_);
  and (_04919_, _04918_, _04896_);
  and (_04920_, _04458_, _03513_);
  nor (_04921_, _04920_, _04029_);
  not (_04922_, _04921_);
  nor (_04923_, _04922_, _04919_);
  and (_04924_, _04885_, _04029_);
  nor (_04925_, _04924_, _04467_);
  not (_04926_, _04925_);
  nor (_04927_, _04926_, _04923_);
  and (_04928_, _04467_, _03513_);
  or (_04929_, _04928_, _04466_);
  nor (_04930_, _04929_, _04927_);
  and (_04931_, _03511_, _04466_);
  nor (_04932_, _04931_, _04930_);
  and (_04933_, _04932_, _04577_);
  and (_04934_, _04893_, _03464_);
  nor (_04935_, _04934_, _04933_);
  nor (_04936_, _04935_, _03461_);
  nor (_04937_, _03462_, _03515_);
  or (_04938_, _04937_, _04936_);
  and (_04939_, _04938_, _03207_);
  or (_04940_, _04939_, _04481_);
  nor (_04941_, _04940_, _04895_);
  and (_04942_, _04885_, _04481_);
  nor (_04943_, _04942_, _04480_);
  not (_04944_, _04943_);
  nor (_04945_, _04944_, _04941_);
  not (_04946_, _04480_);
  nor (_04947_, _04946_, _03515_);
  nor (_04948_, _04947_, _04945_);
  nor (_04949_, _04948_, _03219_);
  and (_04950_, _04893_, _03219_);
  not (_04951_, _04950_);
  and (_04952_, _04951_, _04504_);
  not (_04953_, _04952_);
  nor (_04954_, _04953_, _04949_);
  nor (_04955_, _04504_, _03513_);
  nor (_04956_, _04955_, _04954_);
  nor (_04957_, _04956_, _04507_);
  or (_04958_, _04957_, _04510_);
  nor (_04959_, _04958_, _04886_);
  and (_04960_, _04510_, _03513_);
  nor (_04961_, _04960_, _04959_);
  nor (_04962_, _04961_, _03168_);
  and (_04963_, _04893_, _03168_);
  not (_04964_, _04963_);
  and (_04965_, _04964_, _04531_);
  not (_04966_, _04965_);
  nor (_04967_, _04966_, _04962_);
  nor (_04968_, _04531_, _03513_);
  nor (_04969_, _04968_, _03182_);
  not (_04970_, _04969_);
  nor (_04971_, _04970_, _04967_);
  and (_04972_, _04893_, _03182_);
  or (_04973_, _04972_, _04538_);
  nor (_04974_, _04973_, _04971_);
  and (_04975_, _04538_, _03440_);
  or (_04976_, _04975_, _03191_);
  nor (_04977_, _04976_, _04974_);
  and (_04978_, _04893_, _03191_);
  nor (_04979_, _04978_, _04544_);
  not (_04980_, _04979_);
  nor (_04981_, _04980_, _04977_);
  and (_04982_, _04885_, _04544_);
  nor (_04983_, _04982_, _04546_);
  not (_04984_, _04983_);
  nor (_04985_, _04984_, _04981_);
  not (_04986_, _04553_);
  and (_04987_, _04546_, _03513_);
  nor (_04988_, _04987_, _04986_);
  not (_04989_, _04988_);
  nor (_04990_, _04989_, _04985_);
  nor (_04991_, _04893_, _04553_);
  nor (_04992_, _04991_, _03448_);
  not (_04993_, _04992_);
  nor (_04994_, _04993_, _04990_);
  not (_04995_, _03511_);
  and (_04996_, _03448_, _04995_);
  nor (_04997_, _04996_, _04215_);
  not (_04998_, _04997_);
  nor (_04999_, _04998_, _04994_);
  and (_05000_, _04885_, _04215_);
  nor (_05001_, _05000_, _04559_);
  not (_05002_, _05001_);
  nor (_05003_, _05002_, _04999_);
  nor (_05004_, _05003_, _04828_);
  not (_05005_, _03944_);
  and (_05006_, _04559_, _05005_);
  and (_05007_, _03812_, _03445_);
  nor (_05008_, _04887_, \oc8051_golden_model_1.SP [2]);
  nor (_05009_, _05008_, _04888_);
  and (_05010_, _05009_, _03191_);
  and (_05011_, _04510_, _05005_);
  nor (_05012_, _04504_, _05005_);
  and (_05013_, _03812_, _03452_);
  and (_05014_, _05009_, _03464_);
  and (_05015_, _03812_, _03469_);
  and (_05016_, _04433_, _05005_);
  not (_05017_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_05018_, _04225_, _05017_);
  not (_05019_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05020_, _04371_, _05019_);
  and (_05021_, _05020_, _04369_);
  nand (_05022_, _05021_, _05018_);
  not (_05023_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_05024_, _04371_, _05023_);
  not (_05025_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05026_, _04225_, _05025_);
  and (_05027_, _05026_, _04377_);
  nand (_05028_, _05027_, _05024_);
  nand (_05029_, _05028_, _05022_);
  nand (_05030_, _05029_, _03957_);
  not (_05031_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_05032_, _04371_, _05031_);
  not (_05033_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_05034_, _04225_, _05033_);
  and (_05035_, _05034_, _04377_);
  nand (_05036_, _05035_, _05032_);
  not (_05037_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_05038_, _04225_, _05037_);
  not (_05039_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_05040_, _04371_, _05039_);
  and (_05041_, _05040_, _04369_);
  nand (_05042_, _05041_, _05038_);
  nand (_05043_, _05042_, _05036_);
  nand (_05044_, _05043_, _04385_);
  nand (_05045_, _05044_, _05030_);
  nand (_05046_, _05045_, _03780_);
  not (_05047_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_05048_, _04371_, _05047_);
  not (_05049_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_05050_, _04225_, _05049_);
  and (_05051_, _05050_, _04377_);
  nand (_05052_, _05051_, _05048_);
  nand (_05053_, _04371_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_05054_, _04225_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_05055_, _05054_, _04369_);
  nand (_05056_, _05055_, _05053_);
  nand (_05057_, _05056_, _05052_);
  nand (_05058_, _05057_, _03957_);
  not (_05059_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_05060_, _04371_, _05059_);
  not (_05061_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_05062_, _04225_, _05061_);
  and (_05063_, _05062_, _04377_);
  nand (_05064_, _05063_, _05060_);
  nand (_05065_, _04371_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_05066_, _04225_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_05067_, _05066_, _04369_);
  nand (_05068_, _05067_, _05065_);
  nand (_05069_, _05068_, _05064_);
  nand (_05070_, _05069_, _04385_);
  nand (_05071_, _05070_, _05058_);
  nand (_05072_, _05071_, _04402_);
  nand (_05073_, _05072_, _05046_);
  not (_05074_, _05073_);
  or (_05075_, _05074_, _04430_);
  nor (_05076_, _04796_, _04438_);
  and (_05077_, _04438_, _05005_);
  or (_05078_, _05077_, _04435_);
  or (_05079_, _05078_, _05076_);
  nor (_05080_, _05009_, _03204_);
  nor (_05081_, _05080_, _04331_);
  and (_05082_, _05081_, _04646_);
  and (_05083_, _05082_, _05079_);
  and (_05084_, _05083_, _04434_);
  and (_05085_, _05084_, _05075_);
  nor (_05086_, _05085_, _05016_);
  nor (_05087_, _05086_, _03472_);
  nor (_05088_, _05087_, _05015_);
  nor (_05089_, _05009_, _03202_);
  nor (_05090_, _05089_, _05088_);
  and (_05091_, _04458_, _03944_);
  and (_05092_, _03560_, _03463_);
  nor (_05093_, _05092_, _05091_);
  and (_05094_, _05093_, _05090_);
  and (_05095_, _05073_, _04029_);
  nor (_05096_, _05095_, _04467_);
  and (_05097_, _05096_, _05094_);
  and (_05098_, _04467_, _05005_);
  nor (_05099_, _05098_, _05097_);
  and (_05100_, _03811_, _04466_);
  nor (_05101_, _05100_, _05099_);
  and (_05102_, _05101_, _04577_);
  nor (_05103_, _05102_, _05014_);
  and (_05104_, _03461_, _03811_);
  or (_05105_, _05104_, _05103_);
  nor (_05106_, _05009_, _03207_);
  and (_05107_, _03560_, _03558_);
  nor (_05108_, _05107_, _05106_);
  not (_05109_, _05108_);
  nor (_05110_, _05109_, _05105_);
  and (_05111_, _05073_, _04481_);
  nor (_05112_, _05111_, _04480_);
  and (_05113_, _05112_, _05110_);
  nor (_05114_, _05113_, _05013_);
  nor (_05115_, _05114_, _03219_);
  and (_05116_, _05009_, _03219_);
  nor (_05117_, _05116_, _05115_);
  or (_05118_, _05117_, _04777_);
  nor (_05119_, _05118_, _05012_);
  and (_05120_, _05073_, _04507_);
  nor (_05121_, _05120_, _04510_);
  and (_05122_, _05121_, _05119_);
  nor (_05123_, _05122_, _05011_);
  nor (_05124_, _05123_, _03168_);
  and (_05125_, _05009_, _03168_);
  nor (_05126_, _05125_, _05124_);
  nor (_05127_, _04531_, _05005_);
  nor (_05128_, _05127_, _03182_);
  not (_05129_, _05128_);
  nor (_05130_, _05129_, _05126_);
  and (_05131_, _05009_, _03182_);
  nor (_05132_, _05131_, _05130_);
  and (_05133_, _04538_, _03944_);
  or (_05134_, _05133_, _03191_);
  nor (_05135_, _05134_, _05132_);
  nor (_05136_, _05135_, _05010_);
  not (_05137_, _04719_);
  and (_05138_, _03578_, _03195_);
  not (_05139_, _03195_);
  nor (_05140_, _03575_, _03564_);
  nor (_05141_, _05140_, _05139_);
  nor (_05142_, _05141_, _05138_);
  and (_05143_, _05142_, _05137_);
  not (_05144_, _05143_);
  nor (_05145_, _05144_, _05136_);
  and (_05146_, _05073_, _04544_);
  nor (_05147_, _05146_, _04546_);
  and (_05148_, _05147_, _05145_);
  and (_05149_, _04546_, _05005_);
  nor (_05150_, _05149_, _05148_);
  nor (_05151_, _05009_, _04553_);
  nor (_05152_, _05151_, _03448_);
  not (_05153_, _05152_);
  nor (_05154_, _05153_, _05150_);
  nor (_05155_, _05154_, _05007_);
  and (_05156_, _03560_, _03193_);
  nor (_05157_, _05156_, _05155_);
  and (_05158_, _05073_, _04215_);
  nor (_05159_, _05158_, _04559_);
  and (_05160_, _05159_, _05157_);
  nor (_05161_, _05160_, _05006_);
  nor (_05162_, _05161_, _04824_);
  not (_05163_, _05162_);
  nor (_05164_, _05163_, _05004_);
  and (_05165_, _05164_, _04827_);
  or (_05166_, _05165_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05167_, _04890_, _03455_);
  nor (_05168_, _05009_, _04570_);
  nor (_05169_, _05168_, _05167_);
  and (_05170_, _04891_, _03455_);
  nor (_05171_, _05167_, _04893_);
  nor (_05172_, _05171_, _05170_);
  and (_05173_, _44052_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_05174_, _05173_);
  and (_05175_, _04758_, _04759_);
  and (_05176_, _05175_, _04804_);
  nor (_05177_, _05176_, _05174_);
  and (_05178_, _05177_, _05172_);
  and (_05179_, _05178_, _05169_);
  and (_05180_, _05179_, _04569_);
  not (_05181_, _05180_);
  and (_05182_, _05181_, _05166_);
  not (_05183_, _04744_);
  nor (_05184_, _05174_, _04822_);
  not (_05185_, _05184_);
  nor (_05186_, _05185_, _04565_);
  and (_05187_, _05186_, _05183_);
  not (_05188_, _05161_);
  nor (_05189_, _05185_, _05004_);
  and (_05190_, _05189_, _05188_);
  and (_05191_, _05190_, _05187_);
  not (_05192_, _05191_);
  not (_05193_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_05194_, _04225_, _05193_);
  not (_05195_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05196_, _04371_, _05195_);
  and (_05197_, _05196_, _04369_);
  nand (_05198_, _05197_, _05194_);
  not (_05199_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05200_, _04371_, _05199_);
  not (_05201_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_05202_, _04225_, _05201_);
  and (_05203_, _05202_, _04377_);
  nand (_05204_, _05203_, _05200_);
  nand (_05205_, _05204_, _05198_);
  nand (_05206_, _05205_, _03957_);
  not (_05207_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05208_, _04371_, _05207_);
  not (_05209_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_05210_, _04225_, _05209_);
  and (_05211_, _05210_, _04377_);
  nand (_05212_, _05211_, _05208_);
  not (_05213_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_05214_, _04225_, _05213_);
  not (_05215_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05216_, _04371_, _05215_);
  and (_05217_, _05216_, _04369_);
  nand (_05218_, _05217_, _05214_);
  nand (_05219_, _05218_, _05212_);
  nand (_05220_, _05219_, _04385_);
  nand (_05221_, _05220_, _05206_);
  nand (_05222_, _05221_, _03780_);
  not (_05223_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_05224_, _04371_, _05223_);
  not (_05225_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_05226_, _04225_, _05225_);
  and (_05227_, _05226_, _04377_);
  nand (_05228_, _05227_, _05224_);
  not (_05229_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_05230_, _04225_, _05229_);
  not (_05231_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_05232_, _04371_, _05231_);
  and (_05233_, _05232_, _04369_);
  nand (_05234_, _05233_, _05230_);
  nand (_05235_, _05234_, _05228_);
  nand (_05236_, _05235_, _03957_);
  not (_05237_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_05238_, _04371_, _05237_);
  not (_05239_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_05240_, _04225_, _05239_);
  and (_05241_, _05240_, _04377_);
  nand (_05242_, _05241_, _05238_);
  not (_05243_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_05244_, _04225_, _05243_);
  not (_05245_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05246_, _04371_, _05245_);
  and (_05247_, _05246_, _04369_);
  nand (_05248_, _05247_, _05244_);
  nand (_05249_, _05248_, _05242_);
  nand (_05250_, _05249_, _04385_);
  nand (_05251_, _05250_, _05236_);
  nand (_05252_, _05251_, _04402_);
  nand (_05253_, _05252_, _05222_);
  or (_05254_, _05253_, _03409_);
  and (_05255_, _03511_, _03409_);
  and (_05256_, _05255_, _03811_);
  and (_05257_, _05256_, _04257_);
  and (_05258_, _05257_, _03440_);
  nor (_05259_, _04292_, _03989_);
  and (_05260_, _05259_, _05005_);
  and (_05261_, _05260_, _05258_);
  and (_05262_, _05261_, \oc8051_golden_model_1.PCON [7]);
  not (_05263_, _05262_);
  and (_05264_, _04292_, _04139_);
  and (_05265_, _05264_, _03944_);
  and (_05266_, _05265_, _03513_);
  not (_05267_, _04257_);
  and (_05268_, _05267_, _03811_);
  and (_05269_, _05268_, _05255_);
  and (_05270_, _05269_, _05266_);
  and (_05271_, _05270_, \oc8051_golden_model_1.SBUF [7]);
  and (_05272_, _04292_, _03989_);
  and (_05273_, _05272_, _03944_);
  and (_05274_, _05273_, _03513_);
  not (_05275_, _03811_);
  and (_05276_, _04257_, _05275_);
  and (_05277_, _05276_, _05255_);
  and (_05278_, _05277_, _05274_);
  and (_05279_, _05278_, \oc8051_golden_model_1.IE [7]);
  nor (_05280_, _05279_, _05271_);
  and (_05281_, _05280_, _05263_);
  and (_05282_, _03944_, _03440_);
  and (_05283_, _05282_, _05272_);
  and (_05284_, _05283_, _05269_);
  and (_05285_, _05284_, \oc8051_golden_model_1.P1 [7]);
  and (_05286_, _05274_, _05257_);
  and (_05287_, _05286_, \oc8051_golden_model_1.TCON [7]);
  not (_05288_, _05287_);
  and (_05289_, _05283_, _05277_);
  and (_05290_, _05289_, \oc8051_golden_model_1.P2 [7]);
  nor (_05291_, _04257_, _03811_);
  and (_05292_, _05291_, _05255_);
  and (_05293_, _05292_, _05283_);
  and (_05294_, _05293_, \oc8051_golden_model_1.P3 [7]);
  nor (_05295_, _05294_, _05290_);
  nand (_05296_, _05295_, _05288_);
  nor (_05297_, _05296_, _05285_);
  and (_05298_, _05283_, _05257_);
  and (_05299_, _05298_, \oc8051_golden_model_1.P0 [7]);
  not (_05300_, _05299_);
  nor (_05301_, _03511_, _04493_);
  and (_05302_, _05301_, _05268_);
  and (_05303_, _05302_, _05283_);
  and (_05304_, _05303_, \oc8051_golden_model_1.PSW [7]);
  and (_05305_, _05301_, _05291_);
  and (_05306_, _05305_, _05283_);
  and (_05307_, _05306_, \oc8051_golden_model_1.B [7]);
  nor (_05308_, _05307_, _05304_);
  and (_05309_, _05292_, _05274_);
  and (_05310_, _05309_, \oc8051_golden_model_1.IP [7]);
  and (_05311_, _05301_, _05276_);
  and (_05312_, _05311_, _05283_);
  and (_05313_, _05312_, \oc8051_golden_model_1.ACC [7]);
  nor (_05314_, _05313_, _05310_);
  and (_05315_, _05314_, _05308_);
  and (_05316_, _05315_, _05300_);
  and (_05317_, _05316_, _05297_);
  nand (_05318_, _05317_, _05281_);
  and (_05319_, _05259_, _03944_);
  and (_05320_, _05319_, _05258_);
  and (_05321_, _05320_, \oc8051_golden_model_1.DPH [7]);
  not (_05322_, _05321_);
  and (_05323_, _05265_, _05258_);
  and (_05324_, _05323_, \oc8051_golden_model_1.SP [7]);
  nor (_05325_, _04292_, _04139_);
  and (_05326_, _05325_, _03944_);
  and (_05327_, _05326_, _05258_);
  and (_05328_, _05327_, \oc8051_golden_model_1.DPL [7]);
  nor (_05329_, _05328_, _05324_);
  and (_05330_, _05329_, _05322_);
  and (_05331_, _05266_, _05257_);
  and (_05332_, _05331_, \oc8051_golden_model_1.TMOD [7]);
  and (_05333_, _05274_, _05269_);
  and (_05334_, _05333_, \oc8051_golden_model_1.SCON [7]);
  nor (_05335_, _05334_, _05332_);
  not (_05336_, _05257_);
  nor (_05337_, _03944_, _03440_);
  nand (_05338_, _05337_, _05272_);
  nor (_05339_, _05338_, _05336_);
  and (_05340_, _05339_, \oc8051_golden_model_1.TH0 [7]);
  nand (_05341_, _05337_, _05264_);
  nor (_05342_, _05341_, _05336_);
  and (_05343_, _05342_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05344_, _05343_, _05340_);
  and (_05345_, _05344_, _05335_);
  nand (_05346_, _03944_, _03513_);
  nor (_05347_, _05346_, _05336_);
  and (_05348_, _05347_, _05325_);
  and (_05349_, _05348_, \oc8051_golden_model_1.TL0 [7]);
  and (_05350_, _05347_, _05259_);
  and (_05351_, _05350_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05352_, _05351_, _05349_);
  and (_05353_, _05352_, _05345_);
  and (_05354_, _05353_, _05330_);
  not (_05355_, _05354_);
  nor (_05356_, _05355_, _05318_);
  and (_05357_, _05356_, _05254_);
  not (_05358_, _05357_);
  not (_05359_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_05360_, _04225_, _05359_);
  not (_05361_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_05362_, _04371_, _05361_);
  and (_05363_, _05362_, _04369_);
  nand (_05364_, _05363_, _05360_);
  not (_05365_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_05366_, _04371_, _05365_);
  not (_05367_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_05368_, _04225_, _05367_);
  and (_05369_, _05368_, _04377_);
  nand (_05370_, _05369_, _05366_);
  nand (_05371_, _05370_, _05364_);
  nand (_05372_, _05371_, _03957_);
  not (_05373_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_05374_, _04371_, _05373_);
  not (_05375_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_05376_, _04225_, _05375_);
  and (_05377_, _05376_, _04377_);
  nand (_05378_, _05377_, _05374_);
  not (_05379_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_05380_, _04225_, _05379_);
  not (_05381_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_05382_, _04371_, _05381_);
  and (_05383_, _05382_, _04369_);
  nand (_05384_, _05383_, _05380_);
  nand (_05385_, _05384_, _05378_);
  nand (_05386_, _05385_, _04385_);
  nand (_05387_, _05386_, _05372_);
  nand (_05388_, _05387_, _03780_);
  nand (_05389_, _04225_, \oc8051_golden_model_1.IRAM[11] [6]);
  not (_05390_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05391_, _04225_, _05390_);
  and (_05392_, _05391_, _04377_);
  nand (_05393_, _05392_, _05389_);
  nand (_05394_, _04371_, \oc8051_golden_model_1.IRAM[8] [6]);
  not (_05395_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_05396_, _04371_, _05395_);
  and (_05397_, _05396_, _04369_);
  nand (_05398_, _05397_, _05394_);
  nand (_05399_, _05398_, _05393_);
  nand (_05400_, _05399_, _03957_);
  not (_05401_, \oc8051_golden_model_1.IRAM[15] [6]);
  or (_05402_, _04371_, _05401_);
  not (_05403_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05404_, _04225_, _05403_);
  and (_05405_, _05404_, _04377_);
  nand (_05406_, _05405_, _05402_);
  not (_05407_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_05408_, _04225_, _05407_);
  not (_05409_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_05410_, _04371_, _05409_);
  and (_05411_, _05410_, _04369_);
  nand (_05412_, _05411_, _05408_);
  nand (_05413_, _05412_, _05406_);
  nand (_05414_, _05413_, _04385_);
  nand (_05415_, _05414_, _05400_);
  nand (_05416_, _05415_, _04402_);
  nand (_05417_, _05416_, _05388_);
  or (_05418_, _05417_, _03409_);
  and (_05419_, _05261_, \oc8051_golden_model_1.PCON [6]);
  not (_05420_, _05419_);
  and (_05421_, _05270_, \oc8051_golden_model_1.SBUF [6]);
  and (_05422_, _05278_, \oc8051_golden_model_1.IE [6]);
  nor (_05423_, _05422_, _05421_);
  and (_05424_, _05423_, _05420_);
  and (_05425_, _05289_, \oc8051_golden_model_1.P2 [6]);
  and (_05426_, _05293_, \oc8051_golden_model_1.P3 [6]);
  nor (_05427_, _05426_, _05425_);
  and (_05428_, _05427_, _05424_);
  and (_05429_, _05309_, \oc8051_golden_model_1.IP [6]);
  not (_05430_, _05429_);
  and (_05431_, _05303_, \oc8051_golden_model_1.PSW [6]);
  not (_05432_, _05431_);
  and (_05433_, _05312_, \oc8051_golden_model_1.ACC [6]);
  and (_05434_, _05306_, \oc8051_golden_model_1.B [6]);
  nor (_05435_, _05434_, _05433_);
  and (_05436_, _05435_, _05432_);
  and (_05437_, _05436_, _05430_);
  and (_05438_, _05286_, \oc8051_golden_model_1.TCON [6]);
  and (_05439_, _05339_, \oc8051_golden_model_1.TH0 [6]);
  nor (_05440_, _05439_, _05438_);
  and (_05441_, _05284_, \oc8051_golden_model_1.P1 [6]);
  not (_05442_, _05259_);
  or (_05443_, _05346_, _05442_);
  nor (_05444_, _05443_, _05336_);
  and (_05445_, _05444_, \oc8051_golden_model_1.TL1 [6]);
  nor (_05446_, _05445_, _05441_);
  and (_05447_, _05446_, _05440_);
  and (_05448_, _05333_, \oc8051_golden_model_1.SCON [6]);
  and (_05449_, _05342_, \oc8051_golden_model_1.TH1 [6]);
  nor (_05450_, _05449_, _05448_);
  and (_05451_, _05331_, \oc8051_golden_model_1.TMOD [6]);
  and (_05452_, _05348_, \oc8051_golden_model_1.TL0 [6]);
  nor (_05453_, _05452_, _05451_);
  and (_05454_, _05453_, _05450_);
  and (_05455_, _05454_, _05447_);
  and (_05456_, _05455_, _05437_);
  and (_05457_, _05456_, _05428_);
  and (_05458_, _05298_, \oc8051_golden_model_1.P0 [6]);
  not (_05459_, _05458_);
  and (_05460_, _05320_, \oc8051_golden_model_1.DPH [6]);
  not (_05461_, _05460_);
  and (_05462_, _05323_, \oc8051_golden_model_1.SP [6]);
  and (_05463_, _05327_, \oc8051_golden_model_1.DPL [6]);
  nor (_05464_, _05463_, _05462_);
  and (_05465_, _05464_, _05461_);
  and (_05466_, _05465_, _05459_);
  and (_05467_, _05466_, _05457_);
  and (_05468_, _05467_, _05418_);
  not (_05469_, _05468_);
  not (_05470_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_05471_, _04225_, _05470_);
  not (_05472_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05473_, _04371_, _05472_);
  and (_05474_, _05473_, _04369_);
  nand (_05475_, _05474_, _05471_);
  not (_05476_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_05477_, _04371_, _05476_);
  not (_05478_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05479_, _04225_, _05478_);
  and (_05480_, _05479_, _04377_);
  nand (_05481_, _05480_, _05477_);
  nand (_05482_, _05481_, _05475_);
  nand (_05483_, _05482_, _03957_);
  not (_05484_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_05485_, _04371_, _05484_);
  not (_05486_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05487_, _04225_, _05486_);
  and (_05488_, _05487_, _04377_);
  nand (_05489_, _05488_, _05485_);
  not (_05490_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_05491_, _04225_, _05490_);
  not (_05492_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05493_, _04371_, _05492_);
  and (_05494_, _05493_, _04369_);
  nand (_05495_, _05494_, _05491_);
  nand (_05496_, _05495_, _05489_);
  nand (_05497_, _05496_, _04385_);
  nand (_05498_, _05497_, _05483_);
  nand (_05499_, _05498_, _03780_);
  nand (_05500_, _04225_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_05501_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05502_, _04225_, _05501_);
  and (_05503_, _05502_, _04377_);
  nand (_05504_, _05503_, _05500_);
  nand (_05505_, _04371_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_05506_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_05507_, _04371_, _05506_);
  and (_05508_, _05507_, _04369_);
  nand (_05509_, _05508_, _05505_);
  nand (_05510_, _05509_, _05504_);
  nand (_05511_, _05510_, _03957_);
  nand (_05512_, _04225_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_05513_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05514_, _04225_, _05513_);
  and (_05515_, _05514_, _04377_);
  nand (_05516_, _05515_, _05512_);
  nand (_05517_, _04371_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_05518_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_05519_, _04371_, _05518_);
  and (_05520_, _05519_, _04369_);
  nand (_05521_, _05520_, _05517_);
  nand (_05522_, _05521_, _05516_);
  nand (_05523_, _05522_, _04385_);
  nand (_05524_, _05523_, _05511_);
  nand (_05525_, _05524_, _04402_);
  nand (_05526_, _05525_, _05499_);
  or (_05527_, _05526_, _03409_);
  and (_05528_, _05320_, \oc8051_golden_model_1.DPH [5]);
  not (_05529_, _05528_);
  and (_05530_, _05323_, \oc8051_golden_model_1.SP [5]);
  and (_05531_, _05348_, \oc8051_golden_model_1.TL0 [5]);
  nor (_05532_, _05531_, _05530_);
  and (_05533_, _05532_, _05529_);
  and (_05534_, _05333_, \oc8051_golden_model_1.SCON [5]);
  not (_05535_, _05534_);
  and (_05536_, _05342_, \oc8051_golden_model_1.TH1 [5]);
  and (_05537_, _05270_, \oc8051_golden_model_1.SBUF [5]);
  nor (_05538_, _05537_, _05536_);
  and (_05539_, _05538_, _05535_);
  and (_05540_, _05327_, \oc8051_golden_model_1.DPL [5]);
  not (_05541_, _05540_);
  and (_05542_, _05331_, \oc8051_golden_model_1.TMOD [5]);
  and (_05543_, _05278_, \oc8051_golden_model_1.IE [5]);
  nor (_05544_, _05543_, _05542_);
  and (_05545_, _05544_, _05541_);
  and (_05546_, _05545_, _05539_);
  and (_05547_, _05546_, _05533_);
  not (_05548_, _05547_);
  and (_05549_, _05298_, \oc8051_golden_model_1.P0 [5]);
  not (_05550_, _05549_);
  and (_05551_, _05261_, \oc8051_golden_model_1.PCON [5]);
  not (_05552_, _05551_);
  and (_05553_, _05309_, \oc8051_golden_model_1.IP [5]);
  and (_05554_, _05306_, \oc8051_golden_model_1.B [5]);
  nor (_05555_, _05554_, _05553_);
  and (_05556_, _05303_, \oc8051_golden_model_1.PSW [5]);
  and (_05557_, _05312_, \oc8051_golden_model_1.ACC [5]);
  nor (_05558_, _05557_, _05556_);
  and (_05559_, _05558_, _05555_);
  and (_05560_, _05559_, _05552_);
  nand (_05561_, _05560_, _05550_);
  and (_05562_, _05339_, \oc8051_golden_model_1.TH0 [5]);
  and (_05563_, _05444_, \oc8051_golden_model_1.TL1 [5]);
  nor (_05564_, _05563_, _05562_);
  and (_05565_, _05284_, \oc8051_golden_model_1.P1 [5]);
  and (_05566_, _05286_, \oc8051_golden_model_1.TCON [5]);
  and (_05567_, _05289_, \oc8051_golden_model_1.P2 [5]);
  and (_05568_, _05293_, \oc8051_golden_model_1.P3 [5]);
  or (_05569_, _05568_, _05567_);
  or (_05570_, _05569_, _05566_);
  nor (_05571_, _05570_, _05565_);
  nand (_05572_, _05571_, _05564_);
  or (_05573_, _05572_, _05561_);
  nor (_05574_, _05573_, _05548_);
  and (_05575_, _05574_, _05527_);
  not (_05576_, _05575_);
  or (_05577_, _04885_, _03409_);
  and (_05578_, _05298_, \oc8051_golden_model_1.P0 [3]);
  not (_05579_, _05578_);
  and (_05580_, _05309_, \oc8051_golden_model_1.IP [3]);
  and (_05581_, _05306_, \oc8051_golden_model_1.B [3]);
  nor (_05582_, _05581_, _05580_);
  and (_05583_, _05303_, \oc8051_golden_model_1.PSW [3]);
  and (_05584_, _05312_, \oc8051_golden_model_1.ACC [3]);
  nor (_05585_, _05584_, _05583_);
  and (_05586_, _05585_, _05582_);
  and (_05587_, _05284_, \oc8051_golden_model_1.P1 [3]);
  not (_05588_, _05587_);
  and (_05589_, _05289_, \oc8051_golden_model_1.P2 [3]);
  and (_05590_, _05293_, \oc8051_golden_model_1.P3 [3]);
  nor (_05591_, _05590_, _05589_);
  and (_05592_, _05591_, _05588_);
  and (_05593_, _05592_, _05586_);
  and (_05594_, _05593_, _05579_);
  and (_05595_, _05323_, \oc8051_golden_model_1.SP [3]);
  and (_05596_, _05327_, \oc8051_golden_model_1.DPL [3]);
  nor (_05597_, _05596_, _05595_);
  and (_05598_, _05261_, \oc8051_golden_model_1.PCON [3]);
  not (_05599_, _05598_);
  and (_05600_, _05270_, \oc8051_golden_model_1.SBUF [3]);
  and (_05601_, _05278_, \oc8051_golden_model_1.IE [3]);
  nor (_05602_, _05601_, _05600_);
  and (_05603_, _05602_, _05599_);
  and (_05604_, _05603_, _05597_);
  and (_05605_, _05604_, _05594_);
  and (_05606_, _05348_, \oc8051_golden_model_1.TL0 [3]);
  not (_05607_, _05606_);
  and (_05608_, _05331_, \oc8051_golden_model_1.TMOD [3]);
  and (_05609_, _05333_, \oc8051_golden_model_1.SCON [3]);
  nor (_05610_, _05609_, _05608_);
  and (_05611_, _05286_, \oc8051_golden_model_1.TCON [3]);
  and (_05612_, _05342_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05613_, _05612_, _05611_);
  and (_05614_, _05613_, _05610_);
  and (_05615_, _05614_, _05607_);
  and (_05616_, _05350_, \oc8051_golden_model_1.TL1 [3]);
  not (_05617_, _05616_);
  and (_05618_, _05320_, \oc8051_golden_model_1.DPH [3]);
  and (_05619_, _05339_, \oc8051_golden_model_1.TH0 [3]);
  nor (_05620_, _05619_, _05618_);
  and (_05621_, _05620_, _05617_);
  and (_05622_, _05621_, _05615_);
  and (_05623_, _05622_, _05605_);
  and (_05624_, _05623_, _05577_);
  not (_05625_, _05624_);
  or (_05626_, _04635_, _03409_);
  and (_05627_, _05298_, \oc8051_golden_model_1.P0 [1]);
  not (_05628_, _05627_);
  and (_05629_, _05309_, \oc8051_golden_model_1.IP [1]);
  and (_05630_, _05312_, \oc8051_golden_model_1.ACC [1]);
  nor (_05631_, _05630_, _05629_);
  and (_05632_, _05303_, \oc8051_golden_model_1.PSW [1]);
  and (_05633_, _05306_, \oc8051_golden_model_1.B [1]);
  nor (_05634_, _05633_, _05632_);
  and (_05635_, _05634_, _05631_);
  and (_05636_, _05284_, \oc8051_golden_model_1.P1 [1]);
  not (_05637_, _05636_);
  and (_05638_, _05289_, \oc8051_golden_model_1.P2 [1]);
  and (_05639_, _05293_, \oc8051_golden_model_1.P3 [1]);
  nor (_05640_, _05639_, _05638_);
  and (_05641_, _05640_, _05637_);
  and (_05642_, _05641_, _05635_);
  and (_05643_, _05642_, _05628_);
  and (_05644_, _05323_, \oc8051_golden_model_1.SP [1]);
  and (_05645_, _05327_, \oc8051_golden_model_1.DPL [1]);
  nor (_05646_, _05645_, _05644_);
  and (_05647_, _05261_, \oc8051_golden_model_1.PCON [1]);
  not (_05648_, _05647_);
  and (_05649_, _05270_, \oc8051_golden_model_1.SBUF [1]);
  and (_05650_, _05278_, \oc8051_golden_model_1.IE [1]);
  nor (_05651_, _05650_, _05649_);
  and (_05652_, _05651_, _05648_);
  and (_05653_, _05652_, _05646_);
  and (_05654_, _05653_, _05643_);
  and (_05655_, _05348_, \oc8051_golden_model_1.TL0 [1]);
  not (_05656_, _05655_);
  and (_05657_, _05331_, \oc8051_golden_model_1.TMOD [1]);
  and (_05658_, _05333_, \oc8051_golden_model_1.SCON [1]);
  nor (_05659_, _05658_, _05657_);
  and (_05660_, _05286_, \oc8051_golden_model_1.TCON [1]);
  and (_05661_, _05342_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05662_, _05661_, _05660_);
  and (_05663_, _05662_, _05659_);
  and (_05664_, _05663_, _05656_);
  and (_05665_, _05350_, \oc8051_golden_model_1.TL1 [1]);
  not (_05666_, _05665_);
  and (_05667_, _05320_, \oc8051_golden_model_1.DPH [1]);
  and (_05668_, _05339_, \oc8051_golden_model_1.TH0 [1]);
  nor (_05669_, _05668_, _05667_);
  and (_05670_, _05669_, _05666_);
  and (_05671_, _05670_, _05664_);
  and (_05672_, _05671_, _05654_);
  and (_05673_, _05672_, _05626_);
  not (_05674_, _05673_);
  or (_05675_, _04462_, _03409_);
  and (_05676_, _05261_, \oc8051_golden_model_1.PCON [0]);
  not (_05677_, _05676_);
  and (_05678_, _05270_, \oc8051_golden_model_1.SBUF [0]);
  and (_05679_, _05278_, \oc8051_golden_model_1.IE [0]);
  nor (_05680_, _05679_, _05678_);
  and (_05681_, _05680_, _05677_);
  and (_05682_, _05286_, \oc8051_golden_model_1.TCON [0]);
  not (_05683_, _05682_);
  and (_05684_, _05284_, \oc8051_golden_model_1.P1 [0]);
  not (_05685_, _05684_);
  and (_05686_, _05289_, \oc8051_golden_model_1.P2 [0]);
  and (_05687_, _05293_, \oc8051_golden_model_1.P3 [0]);
  nor (_05688_, _05687_, _05686_);
  and (_05689_, _05688_, _05685_);
  and (_05690_, _05689_, _05683_);
  and (_05691_, _05298_, \oc8051_golden_model_1.P0 [0]);
  not (_05692_, _05691_);
  and (_05693_, _05309_, \oc8051_golden_model_1.IP [0]);
  and (_05694_, _05312_, \oc8051_golden_model_1.ACC [0]);
  nor (_05695_, _05694_, _05693_);
  and (_05696_, _05303_, \oc8051_golden_model_1.PSW [0]);
  and (_05697_, _05306_, \oc8051_golden_model_1.B [0]);
  nor (_05698_, _05697_, _05696_);
  and (_05699_, _05698_, _05695_);
  and (_05700_, _05699_, _05692_);
  and (_05701_, _05700_, _05690_);
  and (_05702_, _05701_, _05681_);
  and (_05703_, _05320_, \oc8051_golden_model_1.DPH [0]);
  not (_05704_, _05703_);
  and (_05705_, _05323_, \oc8051_golden_model_1.SP [0]);
  and (_05706_, _05327_, \oc8051_golden_model_1.DPL [0]);
  nor (_05707_, _05706_, _05705_);
  and (_05708_, _05707_, _05704_);
  and (_05709_, _05331_, \oc8051_golden_model_1.TMOD [0]);
  and (_05710_, _05333_, \oc8051_golden_model_1.SCON [0]);
  nor (_05711_, _05710_, _05709_);
  and (_05712_, _05339_, \oc8051_golden_model_1.TH0 [0]);
  and (_05713_, _05342_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05714_, _05713_, _05712_);
  and (_05715_, _05714_, _05711_);
  and (_05716_, _05348_, \oc8051_golden_model_1.TL0 [0]);
  and (_05717_, _05350_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05718_, _05717_, _05716_);
  and (_05719_, _05718_, _05715_);
  and (_05720_, _05719_, _05708_);
  and (_05721_, _05720_, _05702_);
  nand (_05722_, _05721_, _05675_);
  and (_05723_, _05722_, _05674_);
  or (_05724_, _05073_, _03409_);
  and (_05725_, _05261_, \oc8051_golden_model_1.PCON [2]);
  not (_05726_, _05725_);
  and (_05727_, _05270_, \oc8051_golden_model_1.SBUF [2]);
  and (_05728_, _05278_, \oc8051_golden_model_1.IE [2]);
  nor (_05729_, _05728_, _05727_);
  and (_05730_, _05729_, _05726_);
  and (_05731_, _05286_, \oc8051_golden_model_1.TCON [2]);
  not (_05732_, _05731_);
  and (_05733_, _05284_, \oc8051_golden_model_1.P1 [2]);
  not (_05734_, _05733_);
  and (_05735_, _05289_, \oc8051_golden_model_1.P2 [2]);
  and (_05736_, _05293_, \oc8051_golden_model_1.P3 [2]);
  nor (_05737_, _05736_, _05735_);
  and (_05738_, _05737_, _05734_);
  and (_05739_, _05738_, _05732_);
  and (_05740_, _05298_, \oc8051_golden_model_1.P0 [2]);
  not (_05741_, _05740_);
  and (_05742_, _05303_, \oc8051_golden_model_1.PSW [2]);
  and (_05743_, _05312_, \oc8051_golden_model_1.ACC [2]);
  nor (_05744_, _05743_, _05742_);
  and (_05745_, _05309_, \oc8051_golden_model_1.IP [2]);
  and (_05746_, _05306_, \oc8051_golden_model_1.B [2]);
  nor (_05747_, _05746_, _05745_);
  and (_05748_, _05747_, _05744_);
  and (_05749_, _05748_, _05741_);
  and (_05750_, _05749_, _05739_);
  and (_05751_, _05750_, _05730_);
  and (_05752_, _05320_, \oc8051_golden_model_1.DPH [2]);
  not (_05753_, _05752_);
  and (_05754_, _05323_, \oc8051_golden_model_1.SP [2]);
  and (_05755_, _05327_, \oc8051_golden_model_1.DPL [2]);
  nor (_05756_, _05755_, _05754_);
  and (_05757_, _05756_, _05753_);
  and (_05758_, _05331_, \oc8051_golden_model_1.TMOD [2]);
  and (_05759_, _05333_, \oc8051_golden_model_1.SCON [2]);
  nor (_05760_, _05759_, _05758_);
  and (_05761_, _05339_, \oc8051_golden_model_1.TH0 [2]);
  and (_05762_, _05342_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05763_, _05762_, _05761_);
  and (_05764_, _05763_, _05760_);
  and (_05765_, _05348_, \oc8051_golden_model_1.TL0 [2]);
  and (_05766_, _05350_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05767_, _05766_, _05765_);
  and (_05768_, _05767_, _05764_);
  and (_05769_, _05768_, _05757_);
  and (_05770_, _05769_, _05751_);
  and (_05771_, _05770_, _05724_);
  not (_05772_, _05771_);
  and (_05773_, _05772_, _05723_);
  and (_05774_, _05773_, _05625_);
  not (_05775_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_05776_, _04225_, _05775_);
  not (_05777_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05778_, _04371_, _05777_);
  and (_05779_, _05778_, _04369_);
  nand (_05780_, _05779_, _05776_);
  not (_05781_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_05782_, _04371_, _05781_);
  not (_05783_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05784_, _04225_, _05783_);
  and (_05785_, _05784_, _04377_);
  nand (_05786_, _05785_, _05782_);
  nand (_05787_, _05786_, _05780_);
  nand (_05788_, _05787_, _03957_);
  not (_05789_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05790_, _04371_, _05789_);
  not (_05791_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05792_, _04225_, _05791_);
  and (_05793_, _05792_, _04377_);
  nand (_05794_, _05793_, _05790_);
  not (_05795_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05796_, _04225_, _05795_);
  not (_05797_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05798_, _04371_, _05797_);
  and (_05799_, _05798_, _04369_);
  nand (_05800_, _05799_, _05796_);
  nand (_05801_, _05800_, _05794_);
  nand (_05802_, _05801_, _04385_);
  nand (_05803_, _05802_, _05788_);
  nand (_05804_, _05803_, _03780_);
  nand (_05805_, _04225_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_05806_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05807_, _04225_, _05806_);
  and (_05808_, _05807_, _04377_);
  nand (_05809_, _05808_, _05805_);
  nand (_05810_, _04371_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_05811_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05812_, _04371_, _05811_);
  and (_05813_, _05812_, _04369_);
  nand (_05814_, _05813_, _05810_);
  nand (_05815_, _05814_, _05809_);
  nand (_05816_, _05815_, _03957_);
  nand (_05817_, _04225_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_05818_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05819_, _04225_, _05818_);
  and (_05820_, _05819_, _04377_);
  nand (_05821_, _05820_, _05817_);
  nand (_05822_, _04371_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_05823_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05824_, _04371_, _05823_);
  and (_05825_, _05824_, _04369_);
  nand (_05826_, _05825_, _05822_);
  nand (_05827_, _05826_, _05821_);
  nand (_05828_, _05827_, _04385_);
  nand (_05829_, _05828_, _05816_);
  nand (_05830_, _05829_, _04402_);
  nand (_05831_, _05830_, _05804_);
  or (_05832_, _05831_, _03409_);
  and (_05833_, _05309_, \oc8051_golden_model_1.IP [4]);
  and (_05834_, _05306_, \oc8051_golden_model_1.B [4]);
  nor (_05835_, _05834_, _05833_);
  and (_05836_, _05303_, \oc8051_golden_model_1.PSW [4]);
  and (_05837_, _05312_, \oc8051_golden_model_1.ACC [4]);
  nor (_05838_, _05837_, _05836_);
  and (_05839_, _05838_, _05835_);
  and (_05840_, _05298_, \oc8051_golden_model_1.P0 [4]);
  not (_05841_, _05840_);
  and (_05842_, _05284_, \oc8051_golden_model_1.P1 [4]);
  not (_05843_, _05842_);
  and (_05844_, _05289_, \oc8051_golden_model_1.P2 [4]);
  and (_05845_, _05293_, \oc8051_golden_model_1.P3 [4]);
  nor (_05846_, _05845_, _05844_);
  and (_05847_, _05846_, _05843_);
  and (_05848_, _05847_, _05841_);
  and (_05849_, _05848_, _05839_);
  and (_05850_, _05323_, \oc8051_golden_model_1.SP [4]);
  and (_05851_, _05327_, \oc8051_golden_model_1.DPL [4]);
  nor (_05852_, _05851_, _05850_);
  and (_05853_, _05261_, \oc8051_golden_model_1.PCON [4]);
  not (_05854_, _05853_);
  and (_05855_, _05270_, \oc8051_golden_model_1.SBUF [4]);
  and (_05856_, _05278_, \oc8051_golden_model_1.IE [4]);
  nor (_05857_, _05856_, _05855_);
  and (_05858_, _05857_, _05854_);
  and (_05859_, _05858_, _05852_);
  and (_05860_, _05859_, _05849_);
  and (_05861_, _05348_, \oc8051_golden_model_1.TL0 [4]);
  not (_05862_, _05861_);
  and (_05863_, _05331_, \oc8051_golden_model_1.TMOD [4]);
  and (_05864_, _05333_, \oc8051_golden_model_1.SCON [4]);
  nor (_05865_, _05864_, _05863_);
  and (_05866_, _05286_, \oc8051_golden_model_1.TCON [4]);
  and (_05867_, _05342_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05868_, _05867_, _05866_);
  and (_05869_, _05868_, _05865_);
  and (_05870_, _05869_, _05862_);
  and (_05871_, _05350_, \oc8051_golden_model_1.TL1 [4]);
  not (_05872_, _05871_);
  and (_05873_, _05320_, \oc8051_golden_model_1.DPH [4]);
  and (_05874_, _05339_, \oc8051_golden_model_1.TH0 [4]);
  nor (_05875_, _05874_, _05873_);
  and (_05876_, _05875_, _05872_);
  and (_05877_, _05876_, _05870_);
  and (_05878_, _05877_, _05860_);
  and (_05879_, _05878_, _05832_);
  not (_05880_, _05879_);
  and (_05881_, _05880_, _05774_);
  and (_05882_, _05881_, _05576_);
  and (_05883_, _05882_, _05469_);
  nor (_05884_, _05883_, _05358_);
  and (_05885_, _05883_, _05358_);
  nor (_05886_, _05885_, _05884_);
  and (_05887_, _05886_, _04559_);
  not (_05888_, _05526_);
  not (_05889_, _05831_);
  nor (_05890_, _04635_, _04462_);
  nor (_05891_, _05073_, _04885_);
  and (_05892_, _05891_, _05890_);
  and (_05893_, _05892_, _05889_);
  and (_05894_, _05893_, _05888_);
  and (_05895_, _05417_, _05253_);
  nor (_05896_, _05417_, _05253_);
  nor (_05897_, _05896_, _05895_);
  and (_05898_, _05897_, _05894_);
  nor (_05899_, _05894_, _05253_);
  or (_05900_, _05899_, _05898_);
  and (_05901_, _05900_, _04737_);
  or (_05902_, _05901_, _04215_);
  and (_05903_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05904_, _05903_, \oc8051_golden_model_1.PC [6]);
  and (_05905_, _05904_, _02863_);
  and (_05906_, _05905_, \oc8051_golden_model_1.PC [7]);
  nor (_05907_, _05905_, \oc8051_golden_model_1.PC [7]);
  nor (_05908_, _05907_, _05906_);
  not (_05909_, _05908_);
  nand (_05910_, _05909_, _03168_);
  not (_05911_, _03167_);
  nor (_05912_, _04005_, _03561_);
  nor (_05913_, _05912_, _05911_);
  not (_05914_, _05913_);
  nor (_05915_, _04793_, _04778_);
  and (_05916_, _05915_, _05914_);
  and (_05917_, _05916_, _04509_);
  or (_05918_, _05917_, _03409_);
  not (_05919_, _03219_);
  not (_05920_, _03441_);
  nor (_05921_, _04258_, _05920_);
  nor (_05922_, _03812_, _03515_);
  and (_05923_, _05922_, _05921_);
  and (_05924_, _05923_, _05257_);
  and (_05925_, _05924_, \oc8051_golden_model_1.TCON [7]);
  not (_05926_, _03812_);
  and (_05927_, _05926_, _03515_);
  and (_05928_, _05927_, _05921_);
  and (_05929_, _05305_, _05928_);
  and (_05930_, _05929_, \oc8051_golden_model_1.B [7]);
  nor (_05931_, _05930_, _05925_);
  and (_05932_, _05302_, _05928_);
  and (_05933_, _05932_, \oc8051_golden_model_1.PSW [7]);
  not (_05934_, _05933_);
  and (_05935_, _05923_, _05292_);
  and (_05936_, _05935_, \oc8051_golden_model_1.IP [7]);
  and (_05937_, _05311_, _05928_);
  and (_05938_, _05937_, \oc8051_golden_model_1.ACC [7]);
  nor (_05939_, _05938_, _05936_);
  and (_05940_, _05939_, _05934_);
  and (_05941_, _05940_, _05931_);
  and (_05942_, _05923_, _05269_);
  and (_05943_, _05942_, \oc8051_golden_model_1.SCON [7]);
  and (_05944_, _05923_, _05277_);
  and (_05945_, _05944_, \oc8051_golden_model_1.IE [7]);
  nor (_05946_, _05945_, _05943_);
  and (_05947_, _05258_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05948_, _05277_, _05928_);
  and (_05949_, _05948_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05950_, _05949_, _05947_);
  and (_05951_, _05269_, _05928_);
  and (_05952_, _05951_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05953_, _05292_, _05928_);
  and (_05954_, _05953_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05955_, _05954_, _05952_);
  and (_05956_, _05955_, _05950_);
  and (_05957_, _05956_, _05946_);
  and (_05958_, _05957_, _05941_);
  and (_05959_, _05958_, _05254_);
  nor (_05960_, _05959_, _05260_);
  and (_05961_, _05260_, \oc8051_golden_model_1.PSW [7]);
  nor (_05962_, _05961_, _05960_);
  nor (_05963_, _05962_, _04946_);
  not (_05964_, _04466_);
  and (_05965_, _05948_, \oc8051_golden_model_1.P2 [7]);
  and (_05966_, _05953_, \oc8051_golden_model_1.P3 [7]);
  nor (_05967_, _05966_, _05965_);
  and (_05968_, _05258_, \oc8051_golden_model_1.P0 [7]);
  and (_05969_, _05951_, \oc8051_golden_model_1.P1 [7]);
  nor (_05970_, _05969_, _05968_);
  and (_05971_, _05970_, _05967_);
  and (_05972_, _05971_, _05946_);
  and (_05973_, _05972_, _05941_);
  and (_05974_, _05973_, _05254_);
  nor (_05975_, _05974_, _05260_);
  or (_05976_, _05975_, _05964_);
  not (_05977_, _03202_);
  not (_05978_, _03472_);
  not (_05979_, _05260_);
  nand (_05980_, _05974_, _05979_);
  or (_05981_, _05980_, _05978_);
  not (_05982_, _05253_);
  and (_05983_, _05831_, _05526_);
  and (_05984_, _04635_, _04462_);
  and (_05985_, _05073_, _04885_);
  and (_05986_, _05985_, _05984_);
  and (_05987_, _05986_, _05983_);
  and (_05988_, _05987_, _05417_);
  or (_05989_, _05988_, _05982_);
  nand (_05990_, _05988_, _05982_);
  and (_05991_, _05990_, _05989_);
  and (_05992_, _03561_, _03468_);
  not (_05993_, _05992_);
  nor (_05994_, _04327_, _03565_);
  nor (_05995_, _05994_, _03201_);
  nor (_05996_, _05995_, _04644_);
  and (_05997_, _05996_, _05993_);
  not (_05998_, _05997_);
  and (_05999_, _05998_, _05991_);
  nor (_06000_, _05909_, _03204_);
  and (_06001_, _03204_, \oc8051_golden_model_1.ACC [7]);
  or (_06002_, _06001_, _06000_);
  and (_06003_, _06002_, _05997_);
  or (_06005_, _06003_, _04012_);
  or (_06006_, _06005_, _05999_);
  not (_06008_, _04012_);
  nor (_06009_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_06011_, _06009_, _03857_);
  nor (_06012_, _06011_, _03526_);
  nor (_06014_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_06015_, _06014_, _03526_);
  and (_06017_, _06015_, _03455_);
  nor (_06018_, _06017_, _06012_);
  nor (_06020_, _06018_, _03858_);
  not (_06021_, _06020_);
  not (_06023_, _04885_);
  or (_06024_, _06023_, _04481_);
  and (_06026_, _04481_, _03440_);
  not (_06027_, _06026_);
  and (_06029_, _06027_, _03858_);
  nand (_06030_, _06029_, _06024_);
  and (_06032_, _06030_, _06021_);
  nor (_06033_, _06009_, _03857_);
  nor (_06035_, _06033_, _06011_);
  nor (_06036_, _06035_, _03858_);
  not (_06038_, _06036_);
  or (_06039_, _05074_, _04481_);
  and (_06041_, _04481_, _03944_);
  not (_06042_, _06041_);
  and (_06043_, _06042_, _03858_);
  nand (_06044_, _06043_, _06039_);
  and (_06045_, _06044_, _06038_);
  or (_06046_, _04429_, _04481_);
  not (_06047_, _03858_);
  and (_06048_, _04481_, _03989_);
  nor (_06049_, _06048_, _06047_);
  nand (_06050_, _06049_, _06046_);
  nor (_06051_, _03858_, \oc8051_golden_model_1.SP [0]);
  not (_06052_, _06051_);
  and (_06053_, _06052_, _06050_);
  nand (_06054_, _06053_, \oc8051_golden_model_1.IRAM[0] [7]);
  nor (_06055_, _04571_, _03858_);
  not (_06056_, _06055_);
  or (_06057_, _04635_, _04481_);
  nand (_06058_, _04566_, _04481_);
  and (_06059_, _06058_, _03858_);
  nand (_06060_, _06059_, _06057_);
  and (_06061_, _06060_, _06056_);
  not (_06062_, _06061_);
  or (_06063_, _06053_, _05195_);
  and (_06064_, _06063_, _06062_);
  nand (_06065_, _06064_, _06054_);
  nand (_06066_, _06053_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_06067_, _06053_, _05199_);
  and (_06068_, _06067_, _06061_);
  nand (_06069_, _06068_, _06066_);
  nand (_06070_, _06069_, _06065_);
  nand (_06071_, _06070_, _06045_);
  not (_06072_, _06045_);
  nand (_06073_, _06053_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_06074_, _06053_, _05215_);
  and (_06075_, _06074_, _06062_);
  nand (_06076_, _06075_, _06073_);
  nand (_06077_, _06053_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_06078_, _06053_, _05207_);
  and (_06079_, _06078_, _06061_);
  nand (_06080_, _06079_, _06077_);
  nand (_06081_, _06080_, _06076_);
  nand (_06082_, _06081_, _06072_);
  nand (_06083_, _06082_, _06071_);
  nand (_06084_, _06083_, _06032_);
  not (_06085_, _06032_);
  nand (_06086_, _06053_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_06087_, _06053_, _05223_);
  and (_06088_, _06087_, _06061_);
  nand (_06089_, _06088_, _06086_);
  nand (_06090_, _06053_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_06091_, _06053_, _05231_);
  and (_06092_, _06091_, _06062_);
  nand (_06093_, _06092_, _06090_);
  nand (_06094_, _06093_, _06089_);
  nand (_06095_, _06094_, _06045_);
  nand (_06096_, _06053_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_06097_, _06053_, _05245_);
  and (_06098_, _06097_, _06062_);
  nand (_06100_, _06098_, _06096_);
  nand (_06102_, _06053_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_06103_, _06053_, _05237_);
  and (_06105_, _06103_, _06061_);
  nand (_06106_, _06105_, _06102_);
  nand (_06108_, _06106_, _06100_);
  nand (_06109_, _06108_, _06072_);
  nand (_06111_, _06109_, _06095_);
  nand (_06112_, _06111_, _06085_);
  and (_06114_, _06112_, _06084_);
  or (_06115_, _06114_, _06008_);
  and (_06117_, _06115_, _06006_);
  or (_06118_, _06117_, _04433_);
  and (_06120_, _05879_, _05575_);
  not (_06121_, _05722_);
  and (_06123_, _06121_, _05673_);
  and (_06124_, _05771_, _05624_);
  and (_06126_, _06124_, _06123_);
  and (_06127_, _06126_, _06120_);
  and (_06129_, _06127_, _05468_);
  nor (_06130_, _06129_, _05358_);
  and (_06132_, _06129_, _05358_);
  nor (_06133_, _06132_, _06130_);
  or (_06134_, _06133_, _04434_);
  and (_06135_, _06134_, _06118_);
  or (_06136_, _06135_, _03472_);
  and (_06137_, _06136_, _05981_);
  or (_06138_, _06137_, _05977_);
  nor (_06139_, _05908_, _03202_);
  nor (_06140_, _06139_, _04458_);
  and (_06141_, _06140_, _06138_);
  nor (_06142_, _05253_, _04896_);
  or (_06143_, _06142_, _04466_);
  or (_06144_, _06143_, _06141_);
  and (_06145_, _06144_, _05976_);
  or (_06146_, _06145_, _03464_);
  and (_06147_, _05284_, \oc8051_golden_model_1.P1INREG [7]);
  not (_06148_, _06147_);
  and (_06149_, _05289_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06150_, _05293_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06151_, _06150_, _06149_);
  and (_06152_, _06151_, _05288_);
  and (_06153_, _06152_, _06148_);
  and (_06154_, _05298_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06155_, _06154_);
  and (_06156_, _06155_, _05315_);
  and (_06157_, _06156_, _06153_);
  and (_06158_, _06157_, _05281_);
  and (_06159_, _06158_, _05354_);
  and (_06160_, _06159_, _05254_);
  nand (_06161_, _06160_, _03464_);
  and (_06162_, _06161_, _03462_);
  and (_06163_, _06162_, _06146_);
  nor (_06164_, _05974_, _05979_);
  not (_06165_, _06164_);
  and (_06166_, _06165_, _05980_);
  and (_06167_, _06166_, _03461_);
  or (_06168_, _06167_, _06163_);
  and (_06169_, _06168_, _03207_);
  or (_06170_, _05909_, _03207_);
  nand (_06171_, _06170_, _03583_);
  or (_06172_, _06171_, _06169_);
  nand (_06173_, _06160_, _03584_);
  and (_06174_, _06173_, _06172_);
  or (_06175_, _06174_, _04481_);
  and (_06176_, _06114_, _04493_);
  nand (_06177_, _06159_, _04481_);
  or (_06178_, _06177_, _06176_);
  and (_06179_, _06178_, _04946_);
  and (_06180_, _06179_, _06175_);
  or (_06181_, _06180_, _05963_);
  and (_06182_, _06181_, _05919_);
  nand (_06183_, _05908_, _03219_);
  nand (_06184_, _06183_, _04499_);
  or (_06185_, _06184_, _06182_);
  or (_06186_, _05982_, _04499_);
  and (_06187_, _06186_, _06185_);
  or (_06188_, _06187_, _04501_);
  not (_06189_, _04501_);
  or (_06190_, _06114_, _06189_);
  and (_06191_, _06190_, _04754_);
  and (_06192_, _06191_, _06188_);
  not (_06193_, _05916_);
  nor (_06194_, _03409_, _03521_);
  not (_06195_, _06194_);
  and (_06196_, _03702_, _01685_);
  and (_06197_, _03720_, _01690_);
  nor (_06198_, _06197_, _06196_);
  and (_06199_, _03681_, _01696_);
  and (_06200_, _03684_, _01659_);
  nor (_06201_, _06200_, _06199_);
  and (_06202_, _06201_, _06198_);
  and (_06203_, _03696_, _01674_);
  and (_06204_, _03715_, _01671_);
  nor (_06205_, _06204_, _06203_);
  and (_06206_, _03690_, _01617_);
  and (_06207_, _03713_, _01653_);
  nor (_06208_, _06207_, _06206_);
  and (_06209_, _06208_, _06205_);
  and (_06210_, _06209_, _06202_);
  and (_06211_, _03709_, _01713_);
  and (_06212_, _03718_, _01681_);
  nor (_06213_, _06212_, _06211_);
  and (_06214_, _03671_, _01716_);
  and (_06215_, _03704_, _01701_);
  nor (_06216_, _06215_, _06214_);
  and (_06217_, _06216_, _06213_);
  and (_06218_, _03688_, _01647_);
  and (_06219_, _03694_, _01665_);
  nor (_06220_, _06219_, _06218_);
  and (_06221_, _03707_, _01709_);
  and (_06222_, _03674_, _01719_);
  nor (_06223_, _06222_, _06221_);
  and (_06224_, _06223_, _06220_);
  and (_06225_, _06224_, _06217_);
  and (_06226_, _06225_, _06210_);
  not (_06227_, _06226_);
  nor (_06228_, _06227_, _05253_);
  and (_06229_, _04325_, _04118_);
  and (_06230_, _03855_, _03725_);
  and (_06231_, _06230_, _06229_);
  and (_06232_, _03681_, _02197_);
  and (_06233_, _03684_, _02204_);
  nor (_06234_, _06233_, _06232_);
  and (_06235_, _03709_, _02212_);
  and (_06236_, _03704_, _02191_);
  nor (_06237_, _06236_, _06235_);
  and (_06238_, _06237_, _06234_);
  and (_06239_, _03696_, _02173_);
  and (_06240_, _03715_, _02171_);
  nor (_06241_, _06240_, _06239_);
  and (_06242_, _03690_, _02177_);
  and (_06243_, _03713_, _02220_);
  nor (_06244_, _06243_, _06242_);
  and (_06245_, _06244_, _06241_);
  and (_06246_, _06245_, _06238_);
  and (_06247_, _03718_, _02195_);
  and (_06248_, _03702_, _02184_);
  nor (_06249_, _06248_, _06247_);
  and (_06250_, _03671_, _02209_);
  and (_06251_, _03720_, _02186_);
  nor (_06252_, _06251_, _06250_);
  and (_06253_, _06252_, _06249_);
  and (_06254_, _03688_, _02217_);
  and (_06255_, _03694_, _02180_);
  nor (_06256_, _06255_, _06254_);
  and (_06257_, _03707_, _02201_);
  and (_06258_, _03674_, _02189_);
  nor (_06259_, _06258_, _06257_);
  and (_06260_, _06259_, _06256_);
  and (_06261_, _06260_, _06253_);
  and (_06262_, _06261_, _06246_);
  and (_06263_, _06262_, _06227_);
  and (_06264_, _03718_, _02140_);
  and (_06265_, _03715_, _02124_);
  nor (_06266_, _06265_, _06264_);
  and (_06267_, _03688_, _02161_);
  and (_06268_, _03713_, _02115_);
  nor (_06269_, _06268_, _06267_);
  and (_06270_, _06269_, _06266_);
  and (_06271_, _03702_, _02153_);
  and (_06272_, _03720_, _02131_);
  nor (_06273_, _06272_, _06271_);
  and (_06274_, _03671_, _02129_);
  and (_06275_, _03684_, _02147_);
  nor (_06276_, _06275_, _06274_);
  and (_06277_, _06276_, _06273_);
  and (_06278_, _06277_, _06270_);
  and (_06279_, _03707_, _02145_);
  and (_06280_, _03709_, _02136_);
  nor (_06281_, _06280_, _06279_);
  and (_06282_, _03681_, _02142_);
  and (_06283_, _03690_, _02121_);
  nor (_06284_, _06283_, _06282_);
  and (_06285_, _06284_, _06281_);
  and (_06286_, _03704_, _02156_);
  and (_06287_, _03696_, _02117_);
  nor (_06288_, _06287_, _06286_);
  and (_06289_, _03674_, _02134_);
  and (_06290_, _03694_, _02164_);
  nor (_06291_, _06290_, _06289_);
  and (_06292_, _06291_, _06288_);
  and (_06293_, _06292_, _06285_);
  and (_06294_, _06293_, _06278_);
  not (_06295_, _06294_);
  and (_06296_, _03684_, _02085_);
  and (_06297_, _03696_, _02061_);
  nor (_06298_, _06297_, _06296_);
  and (_06299_, _03713_, _02108_);
  and (_06300_, _03715_, _02068_);
  nor (_06301_, _06300_, _06299_);
  and (_06302_, _06301_, _06298_);
  and (_06303_, _03707_, _02090_);
  and (_06304_, _03671_, _02076_);
  nor (_06305_, _06304_, _06303_);
  and (_06306_, _03709_, _02100_);
  and (_06307_, _03702_, _02097_);
  nor (_06308_, _06307_, _06306_);
  and (_06309_, _06308_, _06305_);
  and (_06310_, _06309_, _06302_);
  and (_06311_, _03720_, _02079_);
  and (_06312_, _03690_, _02105_);
  nor (_06313_, _06312_, _06311_);
  and (_06314_, _03718_, _02087_);
  and (_06315_, _03694_, _02065_);
  nor (_06316_, _06315_, _06314_);
  and (_06317_, _06316_, _06313_);
  and (_06318_, _03704_, _02081_);
  and (_06319_, _03681_, _02092_);
  nor (_06320_, _06319_, _06318_);
  and (_06321_, _03674_, _02073_);
  and (_06322_, _03688_, _02059_);
  nor (_06323_, _06322_, _06321_);
  and (_06324_, _06323_, _06320_);
  and (_06325_, _06324_, _06317_);
  and (_06326_, _06325_, _06310_);
  and (_06327_, _06326_, _06295_);
  and (_06328_, _06327_, _06263_);
  and (_06329_, _06328_, _06231_);
  and (_06330_, _06329_, \oc8051_golden_model_1.P2INREG [7]);
  not (_06331_, _06330_);
  and (_06332_, _06326_, _06294_);
  and (_06333_, _06332_, _06263_);
  and (_06334_, _06333_, _06231_);
  and (_06335_, _06334_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06336_, _06335_);
  not (_06337_, _06326_);
  and (_06338_, _06337_, _06294_);
  and (_06339_, _06338_, _06263_);
  and (_06340_, _06339_, _06231_);
  and (_06341_, _06340_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_06342_, _06326_, _06294_);
  and (_06343_, _06342_, _06263_);
  and (_06344_, _06343_, _06231_);
  and (_06345_, _06344_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06346_, _06345_, _06341_);
  and (_06347_, _06346_, _06336_);
  and (_06348_, _06347_, _06331_);
  and (_06349_, _06333_, _06230_);
  not (_06350_, _04118_);
  and (_06351_, _04325_, _06350_);
  and (_06352_, _06351_, _06349_);
  and (_06353_, _06352_, \oc8051_golden_model_1.SP [7]);
  not (_06354_, _04325_);
  and (_06355_, _06354_, _04118_);
  not (_06356_, _03725_);
  and (_06357_, _03855_, _06356_);
  and (_06358_, _06357_, _06333_);
  and (_06359_, _06358_, _06355_);
  and (_06360_, _06359_, \oc8051_golden_model_1.TL0 [7]);
  nor (_06361_, _06360_, _06353_);
  and (_06362_, _06361_, _06348_);
  nor (_06363_, _06262_, _06226_);
  and (_06364_, _06363_, _06231_);
  and (_06365_, _06364_, _06338_);
  and (_06366_, _06365_, \oc8051_golden_model_1.PSW [7]);
  and (_06367_, _06364_, _06327_);
  and (_06368_, _06367_, \oc8051_golden_model_1.ACC [7]);
  nor (_06369_, _06368_, _06366_);
  and (_06370_, _06364_, _06342_);
  and (_06371_, _06370_, \oc8051_golden_model_1.B [7]);
  and (_06372_, _06357_, _06229_);
  and (_06373_, _06372_, _06263_);
  and (_06374_, _06373_, _06342_);
  and (_06375_, _06374_, \oc8051_golden_model_1.IP [7]);
  nor (_06376_, _06375_, _06371_);
  and (_06377_, _06376_, _06369_);
  and (_06378_, _06372_, _06328_);
  and (_06379_, _06378_, \oc8051_golden_model_1.IE [7]);
  not (_06380_, _06379_);
  and (_06381_, _06372_, _06339_);
  and (_06382_, _06381_, \oc8051_golden_model_1.SCON [7]);
  and (_06383_, _06357_, _06351_);
  and (_06384_, _06383_, _06339_);
  and (_06385_, _06384_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06386_, _06385_, _06382_);
  and (_06387_, _06386_, _06380_);
  and (_06388_, _06387_, _06377_);
  and (_06389_, _06388_, _06362_);
  nor (_06390_, _03855_, _03725_);
  and (_06391_, _06390_, _06333_);
  and (_06392_, _06391_, _06229_);
  and (_06393_, _06392_, \oc8051_golden_model_1.TH0 [7]);
  nor (_06394_, _04325_, _04118_);
  and (_06395_, _06394_, _06333_);
  and (_06396_, _06395_, _06357_);
  and (_06397_, _06396_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06398_, _06397_, _06393_);
  not (_06399_, _03855_);
  and (_06400_, _06399_, _03725_);
  and (_06401_, _06400_, _06395_);
  and (_06402_, _06401_, \oc8051_golden_model_1.PCON [7]);
  and (_06403_, _06358_, _06229_);
  and (_06404_, _06403_, \oc8051_golden_model_1.TCON [7]);
  nor (_06405_, _06404_, _06402_);
  and (_06406_, _06405_, _06398_);
  and (_06407_, _06395_, _06230_);
  and (_06408_, _06407_, \oc8051_golden_model_1.DPH [7]);
  and (_06409_, _06358_, _06351_);
  and (_06410_, _06409_, \oc8051_golden_model_1.TMOD [7]);
  nor (_06411_, _06410_, _06408_);
  and (_06412_, _06355_, _06349_);
  and (_06413_, _06412_, \oc8051_golden_model_1.DPL [7]);
  and (_06414_, _06391_, _06351_);
  and (_06415_, _06414_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06416_, _06415_, _06413_);
  and (_06417_, _06416_, _06411_);
  and (_06418_, _06417_, _06406_);
  and (_06419_, _06418_, _06389_);
  not (_06420_, _06419_);
  nor (_06421_, _06420_, _06228_);
  nor (_06422_, _06421_, _06195_);
  or (_06423_, _06422_, _06193_);
  or (_06424_, _06423_, _06192_);
  and (_06425_, _06424_, _05918_);
  not (_06426_, _04510_);
  nor (_06427_, _06226_, _06426_);
  or (_06428_, _06427_, _03168_);
  or (_06429_, _06428_, _06425_);
  and (_06430_, _06429_, _05910_);
  or (_06431_, _06430_, _04528_);
  not (_06432_, _04526_);
  not (_06433_, _04528_);
  and (_06434_, _06226_, _05357_);
  nor (_06435_, _06226_, _05357_);
  nor (_06436_, _06435_, _06434_);
  or (_06437_, _06436_, _06433_);
  and (_06438_, _06437_, _06432_);
  and (_06439_, _06438_, _06431_);
  not (_06440_, \oc8051_golden_model_1.ACC [7]);
  nor (_06441_, _05357_, _06440_);
  and (_06442_, _05357_, _06440_);
  nor (_06443_, _06442_, _06441_);
  and (_06444_, _06443_, _04526_);
  or (_06445_, _06444_, _04524_);
  or (_06446_, _06445_, _06439_);
  or (_06447_, _06435_, _04525_);
  and (_06448_, _06447_, _04522_);
  and (_06449_, _06448_, _06446_);
  and (_06450_, _06441_, _04521_);
  or (_06451_, _06450_, _03182_);
  or (_06452_, _06451_, _06449_);
  not (_06453_, _03618_);
  nor (_06454_, _06453_, _03409_);
  and (_06455_, _05909_, _03182_);
  nor (_06456_, _06455_, _06454_);
  and (_06457_, _06456_, _06452_);
  not (_06458_, _03741_);
  nor (_06459_, _06458_, _03409_);
  not (_06460_, _06454_);
  nor (_06461_, _06434_, _06460_);
  or (_06462_, _06461_, _06459_);
  or (_06463_, _06462_, _06457_);
  nand (_06464_, _06442_, _06459_);
  and (_06465_, _06464_, _04803_);
  and (_06466_, _06465_, _06463_);
  and (_06467_, _05908_, _03191_);
  nor (_06468_, _05994_, _05139_);
  or (_06469_, _06468_, _06467_);
  or (_06470_, _06469_, _06466_);
  not (_06471_, _06468_);
  or (_06472_, _06471_, _05991_);
  and (_06473_, _06472_, _04721_);
  and (_06474_, _06473_, _06470_);
  not (_06475_, _04721_);
  and (_06476_, _05991_, _06475_);
  or (_06477_, _06476_, _04544_);
  or (_06478_, _06477_, _06474_);
  not (_06479_, _04546_);
  not (_06480_, _04544_);
  not (_06481_, _06114_);
  nand (_06482_, _06053_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_06483_, _06053_, _05361_);
  and (_06484_, _06483_, _06062_);
  nand (_06485_, _06484_, _06482_);
  nand (_06486_, _06053_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_06487_, _06053_, _05365_);
  and (_06488_, _06487_, _06061_);
  nand (_06489_, _06488_, _06486_);
  nand (_06490_, _06489_, _06485_);
  nand (_06491_, _06490_, _06045_);
  nand (_06492_, _06053_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_06493_, _06053_, _05381_);
  and (_06494_, _06493_, _06062_);
  nand (_06495_, _06494_, _06492_);
  nand (_06496_, _06053_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_06497_, _06053_, _05373_);
  and (_06498_, _06497_, _06061_);
  nand (_06499_, _06498_, _06496_);
  nand (_06500_, _06499_, _06495_);
  nand (_06501_, _06500_, _06072_);
  and (_06502_, _06501_, _06032_);
  and (_06503_, _06502_, _06491_);
  nand (_06504_, _06053_, _05390_);
  or (_06505_, _06053_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_06506_, _06505_, _06504_);
  nand (_06507_, _06506_, _06061_);
  nand (_06508_, _06053_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_06509_, _06053_, _05395_);
  and (_06510_, _06509_, _06508_);
  nand (_06511_, _06510_, _06062_);
  nand (_06512_, _06511_, _06507_);
  nand (_06513_, _06512_, _06045_);
  nand (_06514_, _06053_, _05403_);
  or (_06515_, _06053_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_06516_, _06515_, _06514_);
  nand (_06517_, _06516_, _06061_);
  nand (_06518_, _06053_, _05407_);
  or (_06519_, _06053_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_06520_, _06519_, _06518_);
  nand (_06521_, _06520_, _06062_);
  nand (_06522_, _06521_, _06517_);
  nand (_06523_, _06522_, _06072_);
  and (_06524_, _06523_, _06085_);
  and (_06525_, _06524_, _06513_);
  or (_06526_, _06525_, _06503_);
  not (_06527_, _06526_);
  nand (_06528_, _06053_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_06529_, _06053_, _04580_);
  and (_06530_, _06529_, _06062_);
  nand (_06531_, _06530_, _06528_);
  nand (_06532_, _06053_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_06533_, _06053_, _04584_);
  and (_06534_, _06533_, _06061_);
  nand (_06535_, _06534_, _06532_);
  nand (_06536_, _06535_, _06531_);
  nand (_06537_, _06536_, _06045_);
  nand (_06538_, _06053_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_06539_, _06053_, _04601_);
  and (_06540_, _06539_, _06062_);
  nand (_06541_, _06540_, _06538_);
  nand (_06542_, _06053_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_06543_, _06053_, _04593_);
  and (_06544_, _06543_, _06061_);
  nand (_06545_, _06544_, _06542_);
  nand (_06546_, _06545_, _06541_);
  nand (_06547_, _06546_, _06072_);
  and (_06548_, _06547_, _06032_);
  and (_06549_, _06548_, _06537_);
  nand (_06550_, _06053_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_06551_, _06053_, _04609_);
  and (_06552_, _06551_, _06550_);
  nand (_06553_, _06552_, _06061_);
  nand (_06554_, _06053_, _04614_);
  or (_06555_, _06053_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_06556_, _06555_, _06554_);
  nand (_06557_, _06556_, _06062_);
  nand (_06558_, _06557_, _06553_);
  nand (_06559_, _06558_, _06045_);
  nand (_06560_, _06053_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_06561_, _06053_, _04621_);
  and (_06562_, _06561_, _06560_);
  nand (_06563_, _06562_, _06061_);
  nand (_06564_, _06053_, _04626_);
  or (_06565_, _06053_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_06566_, _06565_, _06564_);
  nand (_06567_, _06566_, _06062_);
  nand (_06568_, _06567_, _06563_);
  nand (_06569_, _06568_, _06072_);
  and (_06570_, _06569_, _06085_);
  and (_06571_, _06570_, _06559_);
  or (_06572_, _06571_, _06549_);
  nand (_06573_, _06053_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_06574_, _06053_, _04370_);
  and (_06575_, _06574_, _06062_);
  nand (_06576_, _06575_, _06573_);
  nand (_06577_, _06053_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_06578_, _06053_, _04375_);
  and (_06579_, _06578_, _06061_);
  nand (_06580_, _06579_, _06577_);
  nand (_06581_, _06580_, _06576_);
  nand (_06582_, _06581_, _06045_);
  nand (_06583_, _06053_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_06584_, _06053_, _04394_);
  and (_06585_, _06584_, _06062_);
  nand (_06586_, _06585_, _06583_);
  nand (_06587_, _06053_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_06588_, _06053_, _04386_);
  and (_06589_, _06588_, _06061_);
  nand (_06590_, _06589_, _06587_);
  nand (_06591_, _06590_, _06586_);
  nand (_06592_, _06591_, _06072_);
  and (_06593_, _06592_, _06032_);
  and (_06594_, _06593_, _06582_);
  nand (_06595_, _06053_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_06596_, _06053_, _04403_);
  and (_06597_, _06596_, _06595_);
  nand (_06598_, _06597_, _06061_);
  nand (_06599_, _06053_, _04408_);
  or (_06600_, _06053_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_06601_, _06600_, _06599_);
  nand (_06602_, _06601_, _06062_);
  nand (_06603_, _06602_, _06598_);
  nand (_06604_, _06603_, _06045_);
  nand (_06605_, _06053_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_06606_, _06053_, _04415_);
  and (_06607_, _06606_, _06605_);
  nand (_06608_, _06607_, _06061_);
  nand (_06609_, _06053_, _04420_);
  or (_06610_, _06053_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_06611_, _06610_, _06609_);
  nand (_06612_, _06611_, _06062_);
  nand (_06613_, _06612_, _06608_);
  nand (_06614_, _06613_, _06072_);
  and (_06615_, _06614_, _06085_);
  and (_06616_, _06615_, _06604_);
  or (_06617_, _06616_, _06594_);
  nor (_06618_, _06617_, _06572_);
  nand (_06619_, _06053_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_06620_, _06053_, _04831_);
  and (_06621_, _06620_, _06062_);
  nand (_06622_, _06621_, _06619_);
  nand (_06623_, _06053_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_06624_, _06053_, _04835_);
  and (_06625_, _06624_, _06061_);
  nand (_06626_, _06625_, _06623_);
  nand (_06627_, _06626_, _06622_);
  nand (_06628_, _06627_, _06045_);
  nand (_06629_, _06053_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_06630_, _06053_, _04851_);
  and (_06631_, _06630_, _06062_);
  nand (_06632_, _06631_, _06629_);
  nand (_06633_, _06053_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_06634_, _06053_, _04843_);
  and (_06635_, _06634_, _06061_);
  nand (_06636_, _06635_, _06633_);
  nand (_06637_, _06636_, _06632_);
  nand (_06638_, _06637_, _06072_);
  and (_06639_, _06638_, _06032_);
  and (_06640_, _06639_, _06628_);
  nand (_06641_, _06053_, _04861_);
  or (_06642_, _06053_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_06643_, _06642_, _06641_);
  nand (_06644_, _06643_, _06061_);
  nand (_06645_, _06053_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_06646_, _06053_, _04866_);
  and (_06647_, _06646_, _06645_);
  nand (_06648_, _06647_, _06062_);
  nand (_06649_, _06648_, _06644_);
  nand (_06650_, _06649_, _06045_);
  not (_06651_, _06053_);
  or (_06652_, _06651_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_06653_, _06053_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_06654_, _06653_, _06652_);
  nand (_06655_, _06654_, _06061_);
  nand (_06656_, _06053_, _04876_);
  or (_06657_, _06053_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_06658_, _06657_, _06656_);
  nand (_06659_, _06658_, _06062_);
  nand (_06660_, _06659_, _06655_);
  nand (_06661_, _06660_, _06072_);
  and (_06662_, _06661_, _06085_);
  and (_06663_, _06662_, _06650_);
  or (_06664_, _06663_, _06640_);
  nand (_06665_, _06053_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_06666_, _06053_, _05019_);
  and (_06667_, _06666_, _06062_);
  nand (_06668_, _06667_, _06665_);
  nand (_06669_, _06053_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_06670_, _06053_, _05023_);
  and (_06671_, _06670_, _06061_);
  nand (_06672_, _06671_, _06669_);
  nand (_06673_, _06672_, _06668_);
  nand (_06674_, _06673_, _06045_);
  nand (_06675_, _06053_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_06676_, _06053_, _05039_);
  and (_06677_, _06676_, _06062_);
  nand (_06678_, _06677_, _06675_);
  nand (_06679_, _06053_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_06680_, _06053_, _05031_);
  and (_06681_, _06680_, _06061_);
  nand (_06682_, _06681_, _06679_);
  nand (_06683_, _06682_, _06678_);
  nand (_06684_, _06683_, _06072_);
  and (_06685_, _06684_, _06032_);
  and (_06686_, _06685_, _06674_);
  nand (_06687_, _06053_, _05049_);
  or (_06688_, _06053_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_06689_, _06688_, _06687_);
  nand (_06690_, _06689_, _06061_);
  or (_06691_, _06651_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_06692_, _06053_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_06693_, _06692_, _06691_);
  nand (_06694_, _06693_, _06062_);
  nand (_06695_, _06694_, _06690_);
  nand (_06696_, _06695_, _06045_);
  nand (_06697_, _06053_, _05061_);
  or (_06698_, _06053_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_06699_, _06698_, _06697_);
  nand (_06700_, _06699_, _06061_);
  or (_06701_, _06651_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_06702_, _06053_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_06704_, _06702_, _06701_);
  nand (_06705_, _06704_, _06062_);
  nand (_06706_, _06705_, _06700_);
  nand (_06707_, _06706_, _06072_);
  and (_06708_, _06707_, _06085_);
  and (_06709_, _06708_, _06696_);
  or (_06710_, _06709_, _06686_);
  nor (_06711_, _06710_, _06664_);
  and (_06712_, _06711_, _06618_);
  nand (_06713_, _06053_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_06714_, _06053_, _05472_);
  and (_06715_, _06714_, _06062_);
  nand (_06716_, _06715_, _06713_);
  nand (_06717_, _06053_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_06718_, _06053_, _05476_);
  and (_06719_, _06718_, _06061_);
  nand (_06720_, _06719_, _06717_);
  nand (_06721_, _06720_, _06716_);
  nand (_06722_, _06721_, _06045_);
  nand (_06723_, _06053_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_06724_, _06053_, _05492_);
  and (_06725_, _06724_, _06062_);
  nand (_06726_, _06725_, _06723_);
  nand (_06727_, _06053_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_06728_, _06053_, _05484_);
  and (_06729_, _06728_, _06061_);
  nand (_06730_, _06729_, _06727_);
  nand (_06731_, _06730_, _06726_);
  nand (_06732_, _06731_, _06072_);
  and (_06733_, _06732_, _06032_);
  and (_06734_, _06733_, _06722_);
  nand (_06735_, _06053_, _05501_);
  or (_06736_, _06053_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_06737_, _06736_, _06735_);
  nand (_06738_, _06737_, _06061_);
  nand (_06739_, _06053_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_06740_, _06053_, _05506_);
  and (_06741_, _06740_, _06739_);
  nand (_06742_, _06741_, _06062_);
  nand (_06743_, _06742_, _06738_);
  nand (_06744_, _06743_, _06045_);
  nand (_06745_, _06053_, _05513_);
  or (_06746_, _06053_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_06747_, _06746_, _06745_);
  nand (_06748_, _06747_, _06061_);
  nand (_06749_, _06053_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_06750_, _06053_, _05518_);
  and (_06751_, _06750_, _06749_);
  nand (_06752_, _06751_, _06062_);
  nand (_06753_, _06752_, _06748_);
  nand (_06754_, _06753_, _06072_);
  and (_06755_, _06754_, _06085_);
  and (_06756_, _06755_, _06744_);
  or (_06757_, _06756_, _06734_);
  nand (_06758_, _06053_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_06759_, _06053_, _05777_);
  and (_06760_, _06759_, _06062_);
  nand (_06761_, _06760_, _06758_);
  nand (_06762_, _06053_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_06763_, _06053_, _05781_);
  and (_06764_, _06763_, _06061_);
  nand (_06765_, _06764_, _06762_);
  nand (_06766_, _06765_, _06761_);
  nand (_06767_, _06766_, _06045_);
  nand (_06768_, _06053_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_06769_, _06053_, _05797_);
  and (_06770_, _06769_, _06062_);
  nand (_06771_, _06770_, _06768_);
  nand (_06772_, _06053_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_06773_, _06053_, _05789_);
  and (_06774_, _06773_, _06061_);
  nand (_06775_, _06774_, _06772_);
  nand (_06776_, _06775_, _06771_);
  nand (_06777_, _06776_, _06072_);
  and (_06778_, _06777_, _06032_);
  and (_06779_, _06778_, _06767_);
  nand (_06780_, _06053_, _05806_);
  or (_06781_, _06053_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_06782_, _06781_, _06780_);
  nand (_06783_, _06782_, _06061_);
  nand (_06784_, _06053_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_06785_, _06053_, _05811_);
  and (_06786_, _06785_, _06784_);
  nand (_06787_, _06786_, _06062_);
  nand (_06788_, _06787_, _06783_);
  nand (_06789_, _06788_, _06045_);
  nand (_06790_, _06053_, _05818_);
  or (_06791_, _06053_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_06792_, _06791_, _06790_);
  nand (_06793_, _06792_, _06061_);
  nand (_06794_, _06053_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_06795_, _06053_, _05823_);
  and (_06796_, _06795_, _06794_);
  nand (_06797_, _06796_, _06062_);
  nand (_06798_, _06797_, _06793_);
  nand (_06799_, _06798_, _06072_);
  and (_06800_, _06799_, _06085_);
  and (_06801_, _06800_, _06789_);
  or (_06802_, _06801_, _06779_);
  nor (_06803_, _06802_, _06757_);
  and (_06804_, _06803_, _06712_);
  and (_06805_, _06804_, _06527_);
  nor (_06806_, _06805_, _06481_);
  and (_06807_, _06805_, _06481_);
  or (_06808_, _06807_, _06806_);
  or (_06809_, _06808_, _06480_);
  and (_06810_, _06809_, _06479_);
  and (_06811_, _06810_, _06478_);
  and (_06812_, _06133_, _04546_);
  or (_06813_, _06812_, _03645_);
  or (_06814_, _06813_, _06811_);
  and (_06815_, _02901_, \oc8051_golden_model_1.PC [2]);
  and (_06816_, _06815_, \oc8051_golden_model_1.PC [3]);
  and (_06817_, _06816_, _05904_);
  and (_06818_, _06817_, \oc8051_golden_model_1.PC [7]);
  nor (_06819_, _06817_, \oc8051_golden_model_1.PC [7]);
  nor (_06820_, _06819_, _06818_);
  not (_06821_, _06820_);
  nand (_06822_, _06821_, _03645_);
  and (_06823_, _06822_, _06814_);
  or (_06824_, _06823_, _03196_);
  and (_06825_, _05909_, _03196_);
  nor (_06826_, _06825_, _03448_);
  and (_06827_, _06826_, _06824_);
  and (_06828_, _05960_, _03448_);
  not (_06829_, _03193_);
  nor (_06830_, _05994_, _06829_);
  or (_06831_, _06830_, _06828_);
  or (_06832_, _06831_, _06827_);
  not (_06833_, _06830_);
  or (_06834_, _06833_, _05900_);
  and (_06835_, _06834_, _04736_);
  and (_06836_, _06835_, _06832_);
  or (_06837_, _06836_, _05902_);
  not (_06838_, _04215_);
  and (_06839_, _06617_, _06572_);
  and (_06840_, _06710_, _06664_);
  and (_06841_, _06840_, _06839_);
  and (_06842_, _06802_, _06757_);
  and (_06843_, _06842_, _06841_);
  and (_06844_, _06843_, _06526_);
  nor (_06845_, _06844_, _06481_);
  and (_06846_, _06844_, _06481_);
  or (_06847_, _06846_, _06845_);
  or (_06848_, _06847_, _06838_);
  and (_06849_, _06848_, _04746_);
  and (_06850_, _06849_, _06837_);
  or (_06851_, _06850_, _05887_);
  and (_06852_, _06851_, _05184_);
  or (_06853_, _06852_, _05192_);
  and (_06854_, _06853_, _05182_);
  not (_06855_, _03645_);
  and (_06856_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06857_, _06856_, \oc8051_golden_model_1.PC [10]);
  and (_06858_, _06857_, _06818_);
  and (_06859_, _06858_, \oc8051_golden_model_1.PC [11]);
  and (_06860_, _06859_, \oc8051_golden_model_1.PC [12]);
  and (_06861_, _06860_, \oc8051_golden_model_1.PC [13]);
  and (_06862_, _06861_, \oc8051_golden_model_1.PC [14]);
  nor (_06863_, _06862_, \oc8051_golden_model_1.PC [15]);
  and (_06864_, _06818_, \oc8051_golden_model_1.PC [8]);
  and (_06865_, _06864_, \oc8051_golden_model_1.PC [9]);
  and (_06866_, _06865_, \oc8051_golden_model_1.PC [10]);
  and (_06867_, _06866_, \oc8051_golden_model_1.PC [11]);
  and (_06868_, _06867_, \oc8051_golden_model_1.PC [12]);
  and (_06869_, _06868_, \oc8051_golden_model_1.PC [13]);
  and (_06870_, _06869_, \oc8051_golden_model_1.PC [14]);
  and (_06871_, _06870_, \oc8051_golden_model_1.PC [15]);
  nor (_06872_, _06871_, _06863_);
  or (_06873_, _06872_, _06855_);
  and (_06874_, _06857_, _05906_);
  and (_06875_, _06874_, \oc8051_golden_model_1.PC [11]);
  and (_06876_, _06875_, \oc8051_golden_model_1.PC [12]);
  and (_06877_, _06876_, \oc8051_golden_model_1.PC [13]);
  and (_06878_, _06877_, \oc8051_golden_model_1.PC [14]);
  nor (_06879_, _06878_, \oc8051_golden_model_1.PC [15]);
  and (_06880_, _05906_, \oc8051_golden_model_1.PC [8]);
  and (_06881_, _06880_, \oc8051_golden_model_1.PC [9]);
  and (_06882_, _06881_, \oc8051_golden_model_1.PC [10]);
  and (_06883_, _06882_, \oc8051_golden_model_1.PC [11]);
  and (_06884_, _06883_, \oc8051_golden_model_1.PC [12]);
  and (_06885_, _06884_, \oc8051_golden_model_1.PC [13]);
  and (_06886_, _06885_, \oc8051_golden_model_1.PC [14]);
  and (_06887_, _06886_, \oc8051_golden_model_1.PC [15]);
  nor (_06888_, _06887_, _06879_);
  or (_06889_, _06888_, _03645_);
  and (_06890_, _06889_, _06873_);
  and (_06891_, _06890_, _05177_);
  and (_06892_, _06891_, _05180_);
  or (_40769_, _06892_, _06854_);
  not (_06893_, \oc8051_golden_model_1.B [7]);
  nor (_06894_, _43189_, _06893_);
  nor (_06895_, _05306_, _06893_);
  not (_06896_, _05306_);
  nor (_06897_, _06896_, _05253_);
  or (_06898_, _06897_, _06895_);
  nor (_06899_, _03578_, _03565_);
  nor (_06900_, _06899_, _03261_);
  not (_06901_, _06900_);
  nor (_06902_, _04495_, _04076_);
  and (_06903_, _06902_, _06901_);
  or (_06904_, _06903_, _06898_);
  nor (_06905_, _05929_, _06893_);
  and (_06906_, _05975_, _05929_);
  or (_06907_, _06906_, _06905_);
  and (_06908_, _06907_, _03465_);
  and (_06909_, _06133_, _05306_);
  or (_06910_, _06909_, _06895_);
  or (_06911_, _06910_, _04432_);
  and (_06912_, _05306_, \oc8051_golden_model_1.ACC [7]);
  or (_06913_, _06912_, _06895_);
  and (_06914_, _06913_, _04436_);
  nor (_06915_, _04436_, _06893_);
  or (_06916_, _06915_, _03534_);
  or (_06917_, _06916_, _06914_);
  and (_06918_, _06917_, _03470_);
  and (_06919_, _06918_, _06911_);
  and (_06920_, _05980_, _05929_);
  or (_06921_, _06920_, _06905_);
  and (_06922_, _06921_, _03469_);
  or (_06923_, _06922_, _03527_);
  or (_06924_, _06923_, _06919_);
  or (_06925_, _06898_, _04457_);
  and (_06926_, _06925_, _06924_);
  or (_06927_, _06926_, _03530_);
  or (_06928_, _06913_, _03531_);
  and (_06929_, _06928_, _03466_);
  and (_06930_, _06929_, _06927_);
  or (_06931_, _06930_, _06908_);
  and (_06932_, _06931_, _03459_);
  and (_06933_, _03607_, _03558_);
  or (_06934_, _06905_, _06165_);
  and (_06935_, _06934_, _03458_);
  and (_06936_, _06935_, _06921_);
  or (_06937_, _06936_, _06933_);
  or (_06938_, _06937_, _06932_);
  and (_06939_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06940_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06941_, _06940_, _06939_);
  and (_06942_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06943_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_06944_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_06945_, _06944_, _06943_);
  nor (_06946_, _06945_, _06941_);
  and (_06947_, _06946_, _06942_);
  nor (_06948_, _06947_, _06941_);
  and (_06949_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06950_, _06949_, _06944_);
  and (_06951_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06952_, _06951_, _06939_);
  nor (_06953_, _06952_, _06950_);
  not (_06954_, _06953_);
  nor (_06955_, _06954_, _06948_);
  and (_06956_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06957_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06958_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06959_, _06958_, _06957_);
  nor (_06960_, _06958_, _06957_);
  nor (_06961_, _06960_, _06959_);
  and (_06962_, _06961_, _06956_);
  nor (_06963_, _06961_, _06956_);
  nor (_06964_, _06963_, _06962_);
  and (_06965_, _06954_, _06948_);
  nor (_06966_, _06965_, _06955_);
  and (_06967_, _06966_, _06964_);
  nor (_06968_, _06967_, _06955_);
  not (_06969_, _06944_);
  and (_06970_, _06949_, _06969_);
  and (_06971_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06972_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06973_, _06972_, _06957_);
  and (_06974_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06975_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06976_, _06975_, _06974_);
  nor (_06977_, _06976_, _06973_);
  and (_06978_, _06977_, _06971_);
  nor (_06979_, _06977_, _06971_);
  nor (_06980_, _06979_, _06978_);
  and (_06981_, _06980_, _06970_);
  nor (_06982_, _06980_, _06970_);
  nor (_06983_, _06982_, _06981_);
  not (_06984_, _06983_);
  nor (_06985_, _06984_, _06968_);
  and (_06986_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06987_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06988_, _06987_, _06986_);
  nor (_06989_, _06962_, _06959_);
  and (_06990_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06991_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06992_, _06991_, _06990_);
  nor (_06993_, _06991_, _06990_);
  nor (_06994_, _06993_, _06992_);
  not (_06995_, _06994_);
  nor (_06996_, _06995_, _06989_);
  and (_06997_, _06995_, _06989_);
  nor (_06998_, _06997_, _06996_);
  and (_06999_, _06998_, _06988_);
  nor (_07000_, _06998_, _06988_);
  nor (_07001_, _07000_, _06999_);
  and (_07002_, _06984_, _06968_);
  nor (_07003_, _07002_, _06985_);
  and (_07004_, _07003_, _07001_);
  nor (_07005_, _07004_, _06985_);
  nor (_07006_, _06978_, _06973_);
  and (_07007_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_07008_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_07009_, _07008_, _07007_);
  nor (_07010_, _07008_, _07007_);
  nor (_07011_, _07010_, _07009_);
  not (_07012_, _07011_);
  nor (_07013_, _07012_, _07006_);
  and (_07014_, _07012_, _07006_);
  nor (_07015_, _07014_, _07013_);
  and (_07016_, _07015_, _06992_);
  nor (_07017_, _07015_, _06992_);
  nor (_07018_, _07017_, _07016_);
  nor (_07019_, _06981_, _06950_);
  and (_07020_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_07021_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_07022_, _07021_, _06972_);
  nor (_07023_, _07021_, _06972_);
  nor (_07024_, _07023_, _07022_);
  and (_07025_, _07024_, _07020_);
  nor (_07026_, _07024_, _07020_);
  nor (_07027_, _07026_, _07025_);
  not (_07028_, _07027_);
  nor (_07029_, _07028_, _07019_);
  and (_07030_, _07028_, _07019_);
  nor (_07031_, _07030_, _07029_);
  and (_07032_, _07031_, _07018_);
  nor (_07033_, _07031_, _07018_);
  nor (_07034_, _07033_, _07032_);
  not (_07035_, _07034_);
  nor (_07036_, _07035_, _07005_);
  nor (_07037_, _06999_, _06996_);
  not (_07038_, _07037_);
  and (_07039_, _07035_, _07005_);
  nor (_07040_, _07039_, _07036_);
  and (_07041_, _07040_, _07038_);
  nor (_07042_, _07041_, _07036_);
  nor (_07043_, _07016_, _07013_);
  not (_07044_, _07043_);
  nor (_07045_, _07032_, _07029_);
  not (_07046_, _07045_);
  and (_07047_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_07048_, _07047_, _06972_);
  and (_07049_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_07050_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_07051_, _07050_, _07049_);
  nor (_07052_, _07051_, _07048_);
  nor (_07053_, _07025_, _07022_);
  and (_07054_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_07055_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_07056_, _07055_, _07054_);
  nor (_07057_, _07055_, _07054_);
  nor (_07058_, _07057_, _07056_);
  not (_07059_, _07058_);
  nor (_07060_, _07059_, _07053_);
  and (_07061_, _07059_, _07053_);
  nor (_07062_, _07061_, _07060_);
  and (_07063_, _07062_, _07009_);
  nor (_07064_, _07062_, _07009_);
  nor (_07065_, _07064_, _07063_);
  and (_07066_, _07065_, _07052_);
  nor (_07067_, _07065_, _07052_);
  nor (_07068_, _07067_, _07066_);
  and (_07069_, _07068_, _07046_);
  nor (_07070_, _07068_, _07046_);
  nor (_07071_, _07070_, _07069_);
  and (_07072_, _07071_, _07044_);
  nor (_07073_, _07071_, _07044_);
  nor (_07074_, _07073_, _07072_);
  not (_07075_, _07074_);
  nor (_07076_, _07075_, _07042_);
  nor (_07077_, _07072_, _07069_);
  nor (_07078_, _07063_, _07060_);
  not (_07079_, _07078_);
  and (_07080_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_07081_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_07082_, _07081_, _07080_);
  nor (_07083_, _07081_, _07080_);
  nor (_07084_, _07083_, _07082_);
  and (_07085_, _07084_, _07048_);
  nor (_07086_, _07084_, _07048_);
  nor (_07087_, _07086_, _07085_);
  and (_07088_, _07087_, _07056_);
  nor (_07089_, _07087_, _07056_);
  nor (_07090_, _07089_, _07088_);
  and (_07091_, _07090_, _07047_);
  nor (_07092_, _07090_, _07047_);
  nor (_07093_, _07092_, _07091_);
  and (_07094_, _07093_, _07066_);
  nor (_07095_, _07093_, _07066_);
  nor (_07096_, _07095_, _07094_);
  and (_07097_, _07096_, _07079_);
  nor (_07098_, _07096_, _07079_);
  nor (_07099_, _07098_, _07097_);
  not (_07100_, _07099_);
  nor (_07101_, _07100_, _07077_);
  and (_07102_, _07100_, _07077_);
  nor (_07103_, _07102_, _07101_);
  and (_07104_, _07103_, _07076_);
  nor (_07105_, _07097_, _07094_);
  nor (_07106_, _07088_, _07085_);
  not (_07107_, _07106_);
  and (_07108_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_07109_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_07110_, _07109_, _07108_);
  nor (_07111_, _07109_, _07108_);
  nor (_07112_, _07111_, _07110_);
  and (_07113_, _07112_, _07082_);
  nor (_07114_, _07112_, _07082_);
  nor (_07115_, _07114_, _07113_);
  and (_07116_, _07115_, _07091_);
  nor (_07117_, _07115_, _07091_);
  nor (_07118_, _07117_, _07116_);
  and (_07119_, _07118_, _07107_);
  nor (_07120_, _07118_, _07107_);
  nor (_07121_, _07120_, _07119_);
  not (_07122_, _07121_);
  nor (_07123_, _07122_, _07105_);
  and (_07124_, _07122_, _07105_);
  nor (_07125_, _07124_, _07123_);
  and (_07126_, _07125_, _07101_);
  nor (_07127_, _07125_, _07101_);
  nor (_07128_, _07127_, _07126_);
  and (_07129_, _07128_, _07104_);
  nor (_07130_, _07128_, _07104_);
  nor (_07131_, _07130_, _07129_);
  and (_07132_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_07133_, _07132_, _06944_);
  and (_07134_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_07135_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_07136_, _07135_, _06940_);
  nor (_07137_, _07136_, _07133_);
  and (_07138_, _07137_, _07134_);
  nor (_07139_, _07138_, _07133_);
  not (_07140_, _07139_);
  nor (_07141_, _06946_, _06942_);
  nor (_07142_, _07141_, _06947_);
  and (_07143_, _07142_, _07140_);
  and (_07144_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_07145_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_07146_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_07147_, _07146_, _07145_);
  nor (_07148_, _07146_, _07145_);
  nor (_07149_, _07148_, _07147_);
  and (_07150_, _07149_, _07144_);
  nor (_07151_, _07149_, _07144_);
  nor (_07152_, _07151_, _07150_);
  nor (_07153_, _07142_, _07140_);
  nor (_07154_, _07153_, _07143_);
  and (_07155_, _07154_, _07152_);
  nor (_07156_, _07155_, _07143_);
  nor (_07157_, _06966_, _06964_);
  nor (_07158_, _07157_, _06967_);
  not (_07159_, _07158_);
  nor (_07160_, _07159_, _07156_);
  and (_07161_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_07162_, _07161_, _06987_);
  nor (_07163_, _07150_, _07147_);
  nor (_07164_, _06987_, _06986_);
  nor (_07165_, _07164_, _06988_);
  not (_07166_, _07165_);
  nor (_07167_, _07166_, _07163_);
  and (_07168_, _07166_, _07163_);
  nor (_07169_, _07168_, _07167_);
  and (_07170_, _07169_, _07162_);
  nor (_07171_, _07169_, _07162_);
  nor (_07172_, _07171_, _07170_);
  and (_07173_, _07159_, _07156_);
  nor (_07174_, _07173_, _07160_);
  and (_07175_, _07174_, _07172_);
  nor (_07176_, _07175_, _07160_);
  nor (_07177_, _07003_, _07001_);
  nor (_07178_, _07177_, _07004_);
  not (_07179_, _07178_);
  nor (_07180_, _07179_, _07176_);
  nor (_07181_, _07170_, _07167_);
  not (_07182_, _07181_);
  and (_07183_, _07179_, _07176_);
  nor (_07184_, _07183_, _07180_);
  and (_07185_, _07184_, _07182_);
  nor (_07186_, _07185_, _07180_);
  nor (_07187_, _07040_, _07038_);
  nor (_07188_, _07187_, _07041_);
  not (_07189_, _07188_);
  nor (_07190_, _07189_, _07186_);
  and (_07191_, _07075_, _07042_);
  nor (_07192_, _07191_, _07076_);
  and (_07193_, _07192_, _07190_);
  nor (_07194_, _07103_, _07076_);
  nor (_07195_, _07194_, _07104_);
  and (_07196_, _07195_, _07193_);
  and (_07197_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_07198_, _07197_, _07132_);
  and (_07199_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_07200_, _07197_, _07132_);
  nor (_07201_, _07200_, _07198_);
  and (_07202_, _07201_, _07199_);
  nor (_07203_, _07202_, _07198_);
  not (_07204_, _07203_);
  nor (_07205_, _07137_, _07134_);
  nor (_07206_, _07205_, _07138_);
  and (_07207_, _07206_, _07204_);
  and (_07208_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_07209_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_07210_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_07211_, _07210_, _07209_);
  nor (_07212_, _07210_, _07209_);
  nor (_07213_, _07212_, _07211_);
  and (_07214_, _07213_, _07208_);
  nor (_07215_, _07213_, _07208_);
  nor (_07216_, _07215_, _07214_);
  nor (_07217_, _07206_, _07204_);
  nor (_07218_, _07217_, _07207_);
  and (_07219_, _07218_, _07216_);
  nor (_07220_, _07219_, _07207_);
  not (_07221_, _07220_);
  nor (_07222_, _07154_, _07152_);
  nor (_07223_, _07222_, _07155_);
  and (_07224_, _07223_, _07221_);
  nor (_07225_, _07214_, _07211_);
  and (_07226_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_07227_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_07228_, _07227_, _07226_);
  nor (_07229_, _07228_, _07162_);
  not (_07230_, _07229_);
  nor (_07231_, _07230_, _07225_);
  and (_07232_, _07230_, _07225_);
  nor (_07233_, _07232_, _07231_);
  nor (_07234_, _07223_, _07221_);
  nor (_07235_, _07234_, _07224_);
  and (_07236_, _07235_, _07233_);
  nor (_07237_, _07236_, _07224_);
  nor (_07238_, _07174_, _07172_);
  nor (_07239_, _07238_, _07175_);
  not (_07240_, _07239_);
  nor (_07241_, _07240_, _07237_);
  and (_07242_, _07240_, _07237_);
  nor (_07243_, _07242_, _07241_);
  and (_07244_, _07243_, _07231_);
  nor (_07245_, _07244_, _07241_);
  nor (_07246_, _07184_, _07182_);
  nor (_07247_, _07246_, _07185_);
  not (_07248_, _07247_);
  nor (_07249_, _07248_, _07245_);
  and (_07250_, _07189_, _07186_);
  nor (_07251_, _07250_, _07190_);
  and (_07252_, _07251_, _07249_);
  nor (_07253_, _07192_, _07190_);
  nor (_07254_, _07253_, _07193_);
  and (_07255_, _07254_, _07252_);
  nor (_07256_, _07254_, _07252_);
  nor (_07257_, _07256_, _07255_);
  and (_07258_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_07259_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_07260_, _07259_, _07258_);
  and (_07261_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_07262_, _07259_, _07258_);
  nor (_07263_, _07262_, _07260_);
  and (_07264_, _07263_, _07261_);
  nor (_07265_, _07264_, _07260_);
  not (_07266_, _07265_);
  nor (_07267_, _07201_, _07199_);
  nor (_07268_, _07267_, _07202_);
  and (_07269_, _07268_, _07266_);
  and (_07270_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_07271_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_07272_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_07273_, _07272_, _07271_);
  nor (_07274_, _07272_, _07271_);
  nor (_07275_, _07274_, _07273_);
  and (_07276_, _07275_, _07270_);
  nor (_07277_, _07275_, _07270_);
  nor (_07278_, _07277_, _07276_);
  nor (_07279_, _07268_, _07266_);
  nor (_07280_, _07279_, _07269_);
  and (_07281_, _07280_, _07278_);
  nor (_07282_, _07281_, _07269_);
  not (_07283_, _07282_);
  nor (_07284_, _07218_, _07216_);
  nor (_07285_, _07284_, _07219_);
  and (_07286_, _07285_, _07283_);
  not (_07287_, _07161_);
  nor (_07288_, _07276_, _07273_);
  nor (_07289_, _07288_, _07287_);
  and (_07290_, _07288_, _07287_);
  nor (_07291_, _07290_, _07289_);
  nor (_07292_, _07285_, _07283_);
  nor (_07293_, _07292_, _07286_);
  and (_07294_, _07293_, _07291_);
  nor (_07295_, _07294_, _07286_);
  not (_07296_, _07295_);
  nor (_07297_, _07235_, _07233_);
  nor (_07298_, _07297_, _07236_);
  and (_07299_, _07298_, _07296_);
  nor (_07300_, _07298_, _07296_);
  nor (_07301_, _07300_, _07299_);
  and (_07302_, _07301_, _07289_);
  nor (_07303_, _07302_, _07299_);
  nor (_07304_, _07243_, _07231_);
  nor (_07305_, _07304_, _07244_);
  not (_07306_, _07305_);
  nor (_07307_, _07306_, _07303_);
  and (_07308_, _07248_, _07245_);
  nor (_07309_, _07308_, _07249_);
  and (_07310_, _07309_, _07307_);
  nor (_07311_, _07251_, _07249_);
  nor (_07312_, _07311_, _07252_);
  and (_07313_, _07312_, _07310_);
  nor (_07314_, _07312_, _07310_);
  nor (_07315_, _07314_, _07313_);
  and (_07316_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_07317_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_07318_, _07317_, _07316_);
  and (_07319_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07320_, _07317_, _07316_);
  nor (_07321_, _07320_, _07318_);
  and (_07322_, _07321_, _07319_);
  nor (_07323_, _07322_, _07318_);
  not (_07324_, _07323_);
  nor (_07325_, _07263_, _07261_);
  nor (_07326_, _07325_, _07264_);
  and (_07327_, _07326_, _07324_);
  and (_07328_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_07329_, _07328_, _07272_);
  and (_07330_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_07331_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_07332_, _07331_, _07330_);
  nor (_07333_, _07332_, _07329_);
  nor (_07334_, _07326_, _07324_);
  nor (_07335_, _07334_, _07327_);
  and (_07336_, _07335_, _07333_);
  nor (_07337_, _07336_, _07327_);
  not (_07338_, _07337_);
  nor (_07339_, _07280_, _07278_);
  nor (_07340_, _07339_, _07281_);
  and (_07341_, _07340_, _07338_);
  nor (_07342_, _07340_, _07338_);
  nor (_07343_, _07342_, _07341_);
  and (_07344_, _07343_, _07329_);
  nor (_07345_, _07344_, _07341_);
  not (_07346_, _07345_);
  nor (_07347_, _07293_, _07291_);
  nor (_07348_, _07347_, _07294_);
  and (_07349_, _07348_, _07346_);
  nor (_07350_, _07301_, _07289_);
  nor (_07351_, _07350_, _07302_);
  and (_07352_, _07351_, _07349_);
  and (_07353_, _07306_, _07303_);
  nor (_07354_, _07353_, _07307_);
  and (_07355_, _07354_, _07352_);
  nor (_07356_, _07309_, _07307_);
  nor (_07357_, _07356_, _07310_);
  nor (_07358_, _07357_, _07355_);
  and (_07359_, _07357_, _07355_);
  not (_07360_, _07359_);
  and (_07361_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_07362_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_07363_, _07362_, _07361_);
  and (_07364_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_07365_, _07362_, _07361_);
  nor (_07366_, _07365_, _07363_);
  and (_07367_, _07366_, _07364_);
  nor (_07368_, _07367_, _07363_);
  not (_07369_, _07368_);
  nor (_07370_, _07321_, _07319_);
  nor (_07371_, _07370_, _07322_);
  and (_07372_, _07371_, _07369_);
  nor (_07373_, _07371_, _07369_);
  nor (_07374_, _07373_, _07372_);
  and (_07375_, _07374_, _07328_);
  nor (_07376_, _07375_, _07372_);
  not (_07377_, _07376_);
  nor (_07378_, _07335_, _07333_);
  nor (_07379_, _07378_, _07336_);
  and (_07380_, _07379_, _07377_);
  nor (_07381_, _07343_, _07329_);
  nor (_07382_, _07381_, _07344_);
  and (_07383_, _07382_, _07380_);
  nor (_07384_, _07348_, _07346_);
  nor (_07385_, _07384_, _07349_);
  and (_07386_, _07385_, _07383_);
  nor (_07387_, _07351_, _07349_);
  nor (_07388_, _07387_, _07352_);
  and (_07389_, _07388_, _07386_);
  nor (_07390_, _07354_, _07352_);
  nor (_07391_, _07390_, _07355_);
  and (_07392_, _07391_, _07389_);
  and (_07393_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_07394_, _07393_, _07362_);
  nor (_07395_, _07366_, _07364_);
  nor (_07396_, _07395_, _07367_);
  and (_07397_, _07396_, _07394_);
  nor (_07398_, _07374_, _07328_);
  nor (_07399_, _07398_, _07375_);
  and (_07400_, _07399_, _07397_);
  nor (_07401_, _07379_, _07377_);
  nor (_07402_, _07401_, _07380_);
  and (_07403_, _07402_, _07400_);
  nor (_07404_, _07382_, _07380_);
  nor (_07405_, _07404_, _07383_);
  and (_07406_, _07405_, _07403_);
  nor (_07407_, _07385_, _07383_);
  nor (_07408_, _07407_, _07386_);
  and (_07409_, _07408_, _07406_);
  nor (_07410_, _07388_, _07386_);
  nor (_07411_, _07410_, _07389_);
  and (_07412_, _07411_, _07409_);
  nor (_07413_, _07391_, _07389_);
  nor (_07414_, _07413_, _07392_);
  and (_07415_, _07414_, _07412_);
  nor (_07416_, _07415_, _07392_);
  and (_07417_, _07416_, _07360_);
  nor (_07418_, _07417_, _07358_);
  and (_07419_, _07418_, _07315_);
  nor (_07420_, _07419_, _07313_);
  not (_07421_, _07420_);
  and (_07422_, _07421_, _07257_);
  nor (_07423_, _07422_, _07255_);
  not (_07424_, _07423_);
  nor (_07425_, _07195_, _07193_);
  nor (_07426_, _07425_, _07196_);
  and (_07427_, _07426_, _07424_);
  nor (_07428_, _07427_, _07196_);
  not (_07429_, _07428_);
  and (_07430_, _07429_, _07131_);
  nor (_07431_, _07430_, _07129_);
  not (_07432_, _07431_);
  and (_07433_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_07434_, _07433_);
  nor (_07435_, _07434_, _07081_);
  nor (_07436_, _07435_, _07113_);
  nor (_07437_, _07119_, _07116_);
  nor (_07438_, _07437_, _07436_);
  and (_07439_, _07437_, _07436_);
  nor (_07440_, _07439_, _07438_);
  not (_07441_, _07440_);
  nor (_07442_, _07126_, _07123_);
  and (_07443_, _07442_, _07441_);
  nor (_07444_, _07442_, _07441_);
  nor (_07445_, _07444_, _07443_);
  and (_07446_, _07445_, _07432_);
  not (_07447_, _06933_);
  or (_07448_, _07438_, _07110_);
  or (_07449_, _07448_, _07444_);
  or (_07450_, _07449_, _07447_);
  or (_07451_, _07450_, _07446_);
  and (_07452_, _07451_, _03453_);
  and (_07453_, _07452_, _06938_);
  not (_07454_, _06903_);
  not (_07455_, _05929_);
  nor (_07456_, _05962_, _07455_);
  or (_07457_, _07456_, _06905_);
  and (_07458_, _07457_, _03452_);
  or (_07459_, _07458_, _07454_);
  or (_07460_, _07459_, _07453_);
  and (_07461_, _07460_, _06904_);
  or (_07462_, _07461_, _04082_);
  and (_07463_, _06114_, _05306_);
  or (_07464_, _06895_, _04500_);
  or (_07465_, _07464_, _07463_);
  and (_07466_, _07465_, _03521_);
  and (_07467_, _07466_, _07462_);
  and (_07468_, _03607_, _03158_);
  nor (_07469_, _06421_, _06896_);
  or (_07470_, _07469_, _06895_);
  and (_07471_, _07470_, _03224_);
  or (_07472_, _07471_, _07468_);
  or (_07473_, _07472_, _07467_);
  not (_07474_, _07468_);
  not (_07475_, \oc8051_golden_model_1.B [1]);
  nor (_07476_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_07477_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_07478_, _07477_, _07476_);
  and (_07479_, _07478_, _07475_);
  not (_07480_, \oc8051_golden_model_1.B [0]);
  and (_07481_, _07480_, \oc8051_golden_model_1.ACC [7]);
  nor (_07482_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_07483_, _07482_, _07481_);
  and (_07484_, _07483_, _07479_);
  not (_07485_, _07482_);
  and (_07486_, \oc8051_golden_model_1.B [0], _06440_);
  nor (_07487_, _07486_, _07485_);
  and (_07488_, _07487_, _07479_);
  or (_07489_, _07488_, _06440_);
  nor (_07490_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_07491_, _07490_, _07476_);
  nor (_07492_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.B [2]);
  and (_07493_, _07492_, _07491_);
  not (_07494_, _07493_);
  not (_07495_, \oc8051_golden_model_1.ACC [6]);
  and (_07496_, \oc8051_golden_model_1.B [0], _07495_);
  nor (_07497_, _07496_, _06440_);
  nor (_07498_, _07497_, _07475_);
  nor (_07499_, _07498_, _07494_);
  nor (_07500_, _07499_, _07489_);
  nor (_07501_, _07500_, _07484_);
  and (_07502_, _07499_, \oc8051_golden_model_1.B [0]);
  nor (_07503_, _07502_, _07495_);
  and (_07504_, _07503_, _07475_);
  nor (_07505_, _07503_, _07475_);
  nor (_07506_, _07505_, _07504_);
  nor (_07507_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07508_, _07507_, _07132_);
  nor (_07509_, _07508_, \oc8051_golden_model_1.ACC [4]);
  nor (_07510_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_07511_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_07512_, _07511_, _07480_);
  nor (_07513_, _07512_, _07510_);
  nor (_07514_, _07513_, _07509_);
  not (_07515_, _07514_);
  and (_07516_, _07515_, _07506_);
  nor (_07517_, _07501_, \oc8051_golden_model_1.B [2]);
  nor (_07518_, _07517_, _07504_);
  not (_07519_, _07518_);
  nor (_07520_, _07519_, _07516_);
  and (_07521_, \oc8051_golden_model_1.B [2], _06440_);
  nor (_07522_, _07521_, \oc8051_golden_model_1.B [7]);
  and (_07523_, _07522_, _07478_);
  not (_07524_, _07523_);
  nor (_07525_, _07524_, _07520_);
  nor (_07526_, _07525_, _07501_);
  nor (_07527_, _07526_, _07484_);
  not (_07528_, \oc8051_golden_model_1.B [2]);
  nor (_07529_, _07515_, _07506_);
  nor (_07530_, _07529_, _07516_);
  not (_07531_, _07530_);
  and (_07532_, _07531_, _07525_);
  nor (_07533_, _07525_, _07503_);
  nor (_07534_, _07533_, _07532_);
  and (_07535_, _07534_, _07528_);
  nor (_07536_, _07534_, _07528_);
  nor (_07537_, _07536_, _07535_);
  not (_07538_, _07537_);
  not (_07539_, \oc8051_golden_model_1.ACC [5]);
  nor (_07540_, _07525_, _07539_);
  and (_07541_, _07525_, _07508_);
  or (_07542_, _07541_, _07540_);
  and (_07543_, _07542_, _07475_);
  nor (_07544_, _07542_, _07475_);
  not (_07545_, \oc8051_golden_model_1.ACC [4]);
  and (_07546_, \oc8051_golden_model_1.B [0], _07545_);
  nor (_07547_, _07546_, _07544_);
  nor (_07548_, _07547_, _07543_);
  nor (_07549_, _07548_, _07538_);
  nor (_07550_, _07527_, \oc8051_golden_model_1.B [3]);
  nor (_07551_, _07550_, _07535_);
  not (_07552_, _07551_);
  nor (_07553_, _07552_, _07549_);
  not (_07554_, _07553_);
  and (_07555_, \oc8051_golden_model_1.B [3], _06440_);
  not (_07556_, _07555_);
  and (_07557_, _07556_, _07491_);
  and (_07558_, _07557_, _07554_);
  nor (_07559_, _07558_, _07527_);
  nor (_07560_, _07559_, _07484_);
  not (_07561_, \oc8051_golden_model_1.B [3]);
  not (_07562_, _07558_);
  and (_07563_, _07548_, _07538_);
  nor (_07564_, _07563_, _07549_);
  nor (_07565_, _07564_, _07562_);
  nor (_07566_, _07558_, _07534_);
  nor (_07567_, _07566_, _07565_);
  and (_07568_, _07567_, _07561_);
  nor (_07569_, _07567_, _07561_);
  nor (_07570_, _07569_, _07568_);
  not (_07571_, _07570_);
  nor (_07572_, _07558_, _07542_);
  nor (_07573_, _07544_, _07543_);
  and (_07574_, _07573_, _07546_);
  nor (_07575_, _07573_, _07546_);
  nor (_07576_, _07575_, _07574_);
  and (_07577_, _07576_, _07558_);
  or (_07578_, _07577_, _07572_);
  nor (_07579_, _07578_, \oc8051_golden_model_1.B [2]);
  and (_07580_, _07578_, \oc8051_golden_model_1.B [2]);
  nor (_07581_, _07558_, _07545_);
  nor (_07582_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07583_, _07582_, _07258_);
  and (_07584_, _07558_, _07583_);
  or (_07585_, _07584_, _07581_);
  and (_07586_, _07585_, _07475_);
  nor (_07587_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07588_, _07587_, _07316_);
  nor (_07589_, _07588_, \oc8051_golden_model_1.ACC [2]);
  nor (_07590_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_07591_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_07592_, _07591_, _07480_);
  nor (_07593_, _07592_, _07590_);
  nor (_07594_, _07593_, _07589_);
  not (_07595_, _07594_);
  nor (_07596_, _07585_, _07475_);
  nor (_07597_, _07596_, _07586_);
  and (_07598_, _07597_, _07595_);
  nor (_07599_, _07598_, _07586_);
  nor (_07600_, _07599_, _07580_);
  nor (_07601_, _07600_, _07579_);
  nor (_07602_, _07601_, _07571_);
  nor (_07603_, _07560_, \oc8051_golden_model_1.B [4]);
  nor (_07604_, _07603_, _07568_);
  not (_07605_, _07604_);
  nor (_07606_, _07605_, _07602_);
  not (_07607_, \oc8051_golden_model_1.B [5]);
  and (_07608_, _07490_, _07607_);
  and (_07609_, \oc8051_golden_model_1.B [4], _06440_);
  not (_07610_, _07609_);
  and (_07611_, _07610_, _07608_);
  not (_07612_, _07611_);
  nor (_07613_, _07612_, _07606_);
  nor (_07614_, _07613_, _07560_);
  nor (_07615_, _07614_, _07484_);
  not (_07616_, \oc8051_golden_model_1.B [4]);
  and (_07617_, _07601_, _07571_);
  nor (_07618_, _07617_, _07602_);
  not (_07619_, _07618_);
  and (_07620_, _07619_, _07613_);
  nor (_07621_, _07613_, _07567_);
  nor (_07622_, _07621_, _07620_);
  and (_07623_, _07622_, _07616_);
  nor (_07624_, _07622_, _07616_);
  nor (_07625_, _07624_, _07623_);
  not (_07626_, _07625_);
  nor (_07627_, _07613_, _07578_);
  nor (_07628_, _07580_, _07579_);
  and (_07629_, _07628_, _07599_);
  nor (_07630_, _07628_, _07599_);
  nor (_07631_, _07630_, _07629_);
  not (_07632_, _07631_);
  and (_07633_, _07632_, _07613_);
  nor (_07634_, _07633_, _07627_);
  nor (_07635_, _07634_, \oc8051_golden_model_1.B [3]);
  and (_07636_, _07634_, \oc8051_golden_model_1.B [3]);
  nor (_07637_, _07597_, _07595_);
  nor (_07638_, _07637_, _07598_);
  not (_07639_, _07638_);
  and (_07640_, _07639_, _07613_);
  nor (_07641_, _07613_, _07585_);
  nor (_07642_, _07641_, _07640_);
  and (_07643_, _07642_, _07528_);
  not (_07644_, \oc8051_golden_model_1.ACC [3]);
  nor (_07645_, _07613_, _07644_);
  and (_07646_, _07613_, _07588_);
  or (_07647_, _07646_, _07645_);
  and (_07648_, _07647_, _07475_);
  nor (_07649_, _07647_, _07475_);
  not (_07650_, \oc8051_golden_model_1.ACC [2]);
  and (_07651_, \oc8051_golden_model_1.B [0], _07650_);
  nor (_07652_, _07651_, _07649_);
  nor (_07653_, _07652_, _07648_);
  nor (_07654_, _07642_, _07528_);
  nor (_07655_, _07654_, _07643_);
  not (_07656_, _07655_);
  nor (_07657_, _07656_, _07653_);
  nor (_07658_, _07657_, _07643_);
  nor (_07659_, _07658_, _07636_);
  nor (_07660_, _07659_, _07635_);
  nor (_07661_, _07660_, _07626_);
  nor (_07662_, _07615_, \oc8051_golden_model_1.B [5]);
  nor (_07663_, _07662_, _07623_);
  not (_07664_, _07663_);
  nor (_07665_, _07664_, _07661_);
  not (_07666_, _07665_);
  not (_07667_, _07490_);
  and (_07668_, \oc8051_golden_model_1.B [5], _06440_);
  nor (_07669_, _07668_, _07667_);
  and (_07670_, _07669_, _07666_);
  nor (_07671_, _07670_, _07615_);
  nor (_07672_, _07671_, _07484_);
  nor (_07673_, _07672_, \oc8051_golden_model_1.B [6]);
  and (_07674_, \oc8051_golden_model_1.B [6], _06440_);
  not (_07675_, _07670_);
  and (_07676_, _07660_, _07626_);
  nor (_07677_, _07676_, _07661_);
  nor (_07678_, _07677_, _07675_);
  nor (_07679_, _07670_, _07622_);
  nor (_07680_, _07679_, _07678_);
  and (_07681_, _07680_, _07607_);
  nor (_07682_, _07680_, _07607_);
  nor (_07683_, _07682_, _07681_);
  not (_07684_, _07683_);
  nor (_07685_, _07636_, _07635_);
  nor (_07686_, _07685_, _07658_);
  and (_07687_, _07685_, _07658_);
  or (_07688_, _07687_, _07686_);
  nor (_07689_, _07688_, _07675_);
  and (_07690_, _07675_, _07634_);
  nor (_07691_, _07690_, _07689_);
  and (_07692_, _07691_, _07616_);
  nor (_07693_, _07691_, _07616_);
  and (_07694_, _07656_, _07653_);
  nor (_07695_, _07694_, _07657_);
  nor (_07696_, _07695_, _07675_);
  nor (_07697_, _07670_, _07642_);
  nor (_07698_, _07697_, _07696_);
  and (_07699_, _07698_, _07561_);
  nor (_07700_, _07649_, _07648_);
  nor (_07701_, _07700_, _07651_);
  and (_07702_, _07700_, _07651_);
  or (_07703_, _07702_, _07701_);
  nor (_07704_, _07703_, _07675_);
  nor (_07705_, _07670_, _07647_);
  nor (_07706_, _07705_, _07704_);
  and (_07707_, _07706_, _07528_);
  nor (_07708_, _07706_, _07528_);
  nor (_07709_, _07670_, \oc8051_golden_model_1.ACC [2]);
  nor (_07710_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07711_, _07710_, _07361_);
  nor (_07712_, _07675_, _07711_);
  nor (_07713_, _07712_, _07709_);
  and (_07714_, _07713_, _07475_);
  and (_07715_, \oc8051_golden_model_1.B [0], _03269_);
  not (_07716_, _07715_);
  nor (_07717_, _07713_, _07475_);
  nor (_07718_, _07717_, _07714_);
  and (_07719_, _07718_, _07716_);
  nor (_07720_, _07719_, _07714_);
  nor (_07721_, _07720_, _07708_);
  nor (_07722_, _07721_, _07707_);
  nor (_07723_, _07698_, _07561_);
  nor (_07724_, _07723_, _07699_);
  not (_07725_, _07724_);
  nor (_07726_, _07725_, _07722_);
  nor (_07727_, _07726_, _07699_);
  nor (_07728_, _07727_, _07693_);
  nor (_07729_, _07728_, _07692_);
  nor (_07730_, _07729_, _07684_);
  nor (_07731_, _07730_, _07681_);
  nor (_07732_, _07731_, _07674_);
  nor (_07733_, _07732_, _07673_);
  nor (_07734_, _07733_, \oc8051_golden_model_1.B [7]);
  nor (_07735_, _07734_, _07672_);
  or (_07736_, _07735_, _07484_);
  nor (_07737_, _07736_, \oc8051_golden_model_1.B [7]);
  nor (_07738_, _07737_, _07433_);
  not (_07739_, \oc8051_golden_model_1.B [6]);
  and (_07740_, _07729_, _07684_);
  nor (_07741_, _07740_, _07730_);
  not (_07742_, _07741_);
  and (_07743_, _07742_, _07734_);
  nor (_07744_, _07734_, _07680_);
  nor (_07745_, _07744_, _07743_);
  nor (_07746_, _07745_, _07739_);
  and (_07747_, _07745_, _07739_);
  nor (_07748_, _07747_, _07746_);
  not (_07749_, _07748_);
  nor (_07750_, _07749_, _07738_);
  and (_07751_, _07725_, _07722_);
  or (_07752_, _07751_, _07726_);
  and (_07753_, _07752_, _07734_);
  nor (_07754_, _07734_, _07698_);
  nor (_07755_, _07754_, _07753_);
  nor (_07756_, _07755_, _07616_);
  and (_07757_, _07755_, _07616_);
  nor (_07758_, _07757_, _07756_);
  nor (_07759_, _07693_, _07692_);
  nor (_07760_, _07759_, _07727_);
  and (_07761_, _07759_, _07727_);
  nor (_07762_, _07761_, _07760_);
  and (_07763_, _07762_, _07734_);
  nor (_07764_, _07734_, _07691_);
  or (_07765_, _07764_, _07763_);
  and (_07766_, _07765_, \oc8051_golden_model_1.B [5]);
  nor (_07767_, _07765_, \oc8051_golden_model_1.B [5]);
  nor (_07768_, _07767_, _07766_);
  and (_07769_, _07768_, _07758_);
  and (_07770_, _07769_, _07750_);
  nor (_07771_, _07708_, _07707_);
  nor (_07772_, _07771_, _07720_);
  and (_07773_, _07771_, _07720_);
  nor (_07774_, _07773_, _07772_);
  and (_07775_, _07774_, _07734_);
  nor (_07776_, _07734_, _07706_);
  or (_07777_, _07776_, _07775_);
  and (_07778_, _07777_, \oc8051_golden_model_1.B [3]);
  nor (_07779_, _07777_, \oc8051_golden_model_1.B [3]);
  nor (_07780_, _07779_, _07778_);
  nor (_07781_, _07718_, _07716_);
  nor (_07782_, _07781_, _07719_);
  and (_07783_, _07782_, _07734_);
  not (_07784_, _07713_);
  nor (_07785_, _07734_, _07784_);
  nor (_07786_, _07785_, _07783_);
  and (_07787_, _07786_, \oc8051_golden_model_1.B [2]);
  nor (_07788_, _07786_, \oc8051_golden_model_1.B [2]);
  nor (_07789_, _07788_, _07787_);
  and (_07790_, _07789_, _07780_);
  and (_07791_, _07480_, \oc8051_golden_model_1.ACC [0]);
  not (_07792_, _07791_);
  nor (_07793_, _07734_, \oc8051_golden_model_1.ACC [1]);
  and (_07794_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07795_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07796_, _07795_, _07794_);
  and (_07797_, _07734_, _07796_);
  nor (_07798_, _07797_, _07793_);
  and (_07799_, _07798_, _07475_);
  nor (_07800_, _07798_, _07475_);
  nor (_07801_, _07800_, _07799_);
  and (_07802_, \oc8051_golden_model_1.B [0], _03344_);
  not (_07803_, _07802_);
  and (_07804_, _07803_, _07801_);
  and (_07805_, _07804_, _07792_);
  and (_07806_, _07805_, _07790_);
  and (_07807_, _07806_, _07770_);
  not (_07808_, _07746_);
  nor (_07809_, _07808_, _07738_);
  not (_07810_, _07770_);
  nor (_07811_, _07792_, _07800_);
  nor (_07812_, _07811_, _07799_);
  and (_07813_, _07812_, _07790_);
  not (_07814_, _07813_);
  and (_07815_, _07787_, _07780_);
  nor (_07816_, _07815_, _07778_);
  and (_07817_, _07816_, _07814_);
  nor (_07818_, _07817_, _07810_);
  and (_07819_, _07768_, _07756_);
  nor (_07820_, _07819_, _07766_);
  not (_07821_, _07820_);
  and (_07822_, _07821_, _07750_);
  and (_07823_, _07672_, \oc8051_golden_model_1.B [7]);
  or (_07824_, _07823_, _07822_);
  or (_07825_, _07824_, _07818_);
  nor (_07826_, _07825_, _07809_);
  nor (_07827_, _07826_, _07807_);
  or (_07828_, _07827_, _07484_);
  and (_07829_, _07828_, _07736_);
  or (_07830_, _07829_, _07474_);
  and (_07831_, _07830_, _07473_);
  or (_07832_, _07831_, _03624_);
  and (_07833_, _06227_, _05306_);
  or (_07834_, _07833_, _06895_);
  or (_07835_, _07834_, _04509_);
  and (_07836_, _07835_, _04527_);
  and (_07837_, _07836_, _07832_);
  and (_07838_, _06436_, _05306_);
  or (_07839_, _07838_, _06895_);
  and (_07840_, _07839_, _03623_);
  or (_07841_, _07840_, _03744_);
  or (_07842_, _07841_, _07837_);
  and (_07843_, _06443_, _05306_);
  or (_07844_, _07843_, _06895_);
  or (_07845_, _07844_, _03745_);
  and (_07846_, _07845_, _04523_);
  and (_07847_, _07846_, _07842_);
  or (_07848_, _06895_, _05358_);
  and (_07849_, _07834_, _03611_);
  and (_07850_, _07849_, _07848_);
  or (_07851_, _07850_, _07847_);
  and (_07852_, _07851_, _03734_);
  and (_07853_, _06913_, _03733_);
  and (_07854_, _07853_, _07848_);
  or (_07855_, _07854_, _03618_);
  or (_07856_, _07855_, _07852_);
  nor (_07857_, _06434_, _06896_);
  or (_07858_, _06895_, _06453_);
  or (_07859_, _07858_, _07857_);
  and (_07860_, _07859_, _06458_);
  and (_07861_, _07860_, _07856_);
  nor (_07862_, _06442_, _06896_);
  or (_07863_, _07862_, _06895_);
  and (_07864_, _07863_, _03741_);
  or (_07865_, _07864_, _03767_);
  or (_07866_, _07865_, _07861_);
  or (_07867_, _06910_, _03948_);
  and (_07868_, _07867_, _03446_);
  and (_07869_, _07868_, _07866_);
  and (_07870_, _06907_, _03445_);
  or (_07871_, _07870_, _03473_);
  or (_07872_, _07871_, _07869_);
  and (_07873_, _05886_, _05306_);
  or (_07874_, _06895_, _03474_);
  or (_07875_, _07874_, _07873_);
  and (_07876_, _07875_, _43189_);
  and (_07877_, _07876_, _07872_);
  or (_07878_, _07877_, _06894_);
  and (_40770_, _07878_, _42003_);
  nor (_07879_, _43189_, _06440_);
  and (_07880_, _05253_, _06440_);
  nor (_07881_, _05253_, _06440_);
  nor (_07882_, _07881_, _07880_);
  nor (_07883_, _05417_, _07495_);
  and (_07884_, _05417_, _07495_);
  nor (_07885_, _07884_, _07883_);
  nor (_07886_, _05526_, _07539_);
  and (_07887_, _05526_, _07539_);
  nor (_07888_, _07887_, _07886_);
  not (_07889_, _07888_);
  nor (_07890_, _05831_, _07545_);
  and (_07891_, _05831_, _07545_);
  nor (_07892_, _07891_, _07890_);
  not (_07893_, _07892_);
  nor (_07894_, _04885_, _07644_);
  not (_07895_, _07894_);
  and (_07896_, _04885_, _07644_);
  nor (_07897_, _05073_, _07650_);
  and (_07898_, _05073_, _07650_);
  nor (_07899_, _07898_, _07897_);
  not (_07900_, _07899_);
  nor (_07901_, _04635_, _03269_);
  and (_07902_, _04635_, _03269_);
  nor (_07903_, _07902_, _07901_);
  and (_07904_, _04429_, \oc8051_golden_model_1.ACC [0]);
  and (_07905_, _07904_, _07903_);
  nor (_07906_, _07905_, _07901_);
  nor (_07907_, _07906_, _07900_);
  nor (_07908_, _07907_, _07897_);
  or (_07909_, _07908_, _07896_);
  and (_07910_, _07909_, _07895_);
  nor (_07911_, _07910_, _07893_);
  nor (_07912_, _07911_, _07890_);
  nor (_07913_, _07912_, _07889_);
  or (_07914_, _07913_, _07886_);
  and (_07915_, _07914_, _07885_);
  nor (_07916_, _07915_, _07883_);
  nor (_07917_, _07916_, _07882_);
  and (_07918_, _07916_, _07882_);
  or (_07919_, _07918_, _07917_);
  and (_07920_, _03188_, _02954_);
  not (_07921_, _07920_);
  or (_07922_, _07921_, _07919_);
  and (_07923_, _04005_, _03177_);
  nor (_07924_, _06114_, \oc8051_golden_model_1.ACC [7]);
  nand (_07925_, _07924_, _07923_);
  not (_07926_, _03177_);
  nor (_07927_, _06899_, _07926_);
  nand (_07928_, _07927_, _07880_);
  and (_07929_, _03607_, _03171_);
  not (_07930_, _07929_);
  and (_07931_, _03409_, \oc8051_golden_model_1.ACC [7]);
  nor (_07932_, _03409_, \oc8051_golden_model_1.ACC [7]);
  nor (_07933_, _07932_, _07931_);
  or (_07934_, _07933_, _07930_);
  nor (_07935_, _05312_, _06440_);
  not (_07936_, _05312_);
  nor (_07937_, _07936_, _05253_);
  nor (_07938_, _07937_, _07935_);
  nand (_07939_, _07938_, _07454_);
  and (_07940_, _03607_, _03218_);
  not (_07941_, _07940_);
  and (_07942_, _05259_, \oc8051_golden_model_1.PSW [7]);
  and (_07943_, _07942_, _05337_);
  and (_07944_, _07943_, _05291_);
  and (_07945_, _07944_, _04995_);
  nor (_07946_, _07945_, _04493_);
  and (_07947_, _07944_, _03512_);
  nor (_07948_, _07947_, _07946_);
  and (_07949_, _07948_, \oc8051_golden_model_1.ACC [7]);
  nor (_07950_, _07948_, \oc8051_golden_model_1.ACC [7]);
  nor (_07951_, _07950_, _07949_);
  not (_07952_, _07951_);
  nor (_07953_, _07944_, _04995_);
  nor (_07954_, _07953_, _07945_);
  nor (_07955_, _07954_, _07495_);
  and (_07956_, _07954_, _07495_);
  nor (_07957_, _07955_, _07956_);
  and (_07958_, _07943_, _05267_);
  nor (_07959_, _07958_, _05275_);
  nor (_07960_, _07959_, _07944_);
  nor (_07961_, _07960_, _07539_);
  and (_07962_, _07960_, _07539_);
  nor (_07963_, _07962_, _07961_);
  nor (_07964_, _07943_, _05267_);
  nor (_07965_, _07964_, _07958_);
  nor (_07966_, _07965_, _07545_);
  and (_07967_, _07965_, _07545_);
  nor (_07968_, _07967_, _07966_);
  and (_07969_, _07968_, _07963_);
  nor (_07970_, _05961_, _03513_);
  nor (_07971_, _07970_, _07943_);
  nor (_07972_, _07971_, _07644_);
  and (_07973_, _07971_, _07644_);
  nor (_07974_, _07973_, _07972_);
  nor (_07975_, _07942_, _05005_);
  nor (_07976_, _07975_, _05961_);
  nor (_07977_, _07976_, _07650_);
  and (_07978_, _07976_, _07650_);
  nor (_07979_, _07978_, _07977_);
  and (_07980_, _07979_, _07974_);
  not (_07981_, _07980_);
  not (_07982_, \oc8051_golden_model_1.PSW [7]);
  nor (_07983_, _03989_, _07982_);
  and (_07984_, _03989_, _07982_);
  nor (_07985_, _07984_, _07983_);
  and (_07986_, _07985_, _03344_);
  nor (_07987_, _07985_, _03344_);
  nor (_07988_, _07987_, _07986_);
  nor (_07989_, _04292_, _03269_);
  and (_07990_, _04292_, _03269_);
  nor (_07991_, _07990_, _07989_);
  and (_07992_, \oc8051_golden_model_1.PSW [7], _03344_);
  and (_07993_, _07982_, \oc8051_golden_model_1.ACC [0]);
  nor (_07994_, _07993_, _03989_);
  nor (_07995_, _07994_, _07992_);
  and (_07996_, _07995_, _07991_);
  nor (_07997_, _07995_, _07991_);
  nor (_07998_, _07997_, _07996_);
  nand (_07999_, _07998_, _07988_);
  nor (_08000_, _07999_, _07981_);
  nor (_08001_, _07983_, _04566_);
  nor (_08002_, _08001_, _07942_);
  and (_08003_, _08002_, _03269_);
  nor (_08004_, _08002_, _03269_);
  nor (_08005_, _07987_, _08004_);
  or (_08006_, _08005_, _08003_);
  and (_08007_, _08006_, _07980_);
  not (_08008_, _08007_);
  and (_08009_, _07978_, _07974_);
  nor (_08010_, _08009_, _07973_);
  and (_08011_, _08010_, _08008_);
  nor (_08012_, _08011_, _08000_);
  not (_08013_, _08012_);
  and (_08014_, _08013_, _07969_);
  nor (_08015_, _07966_, _07961_);
  nor (_08016_, _08015_, _07962_);
  or (_08017_, _08016_, _08014_);
  and (_08018_, _08017_, _07957_);
  or (_08019_, _08018_, _07955_);
  and (_08020_, _08019_, _07952_);
  nor (_08021_, _08019_, _07952_);
  or (_08022_, _08021_, _08020_);
  or (_08023_, _08022_, _07941_);
  not (_08024_, _04066_);
  and (_08025_, _06844_, \oc8051_golden_model_1.PSW [7]);
  nor (_08026_, _08025_, _06481_);
  and (_08027_, _08025_, _06481_);
  nor (_08028_, _08027_, _08026_);
  and (_08029_, _08028_, \oc8051_golden_model_1.ACC [7]);
  nor (_08030_, _08028_, \oc8051_golden_model_1.ACC [7]);
  nor (_08031_, _08030_, _08029_);
  and (_08032_, _06843_, \oc8051_golden_model_1.PSW [7]);
  nor (_08033_, _08032_, _06526_);
  nor (_08034_, _08033_, _08025_);
  nor (_08035_, _08034_, _07495_);
  and (_08036_, _08034_, _07495_);
  and (_08037_, _06839_, \oc8051_golden_model_1.PSW [7]);
  and (_08038_, _08037_, _06840_);
  and (_08039_, _08038_, _06802_);
  nor (_08040_, _08039_, _06757_);
  nor (_08041_, _08040_, _08032_);
  and (_08042_, _08041_, _07539_);
  nor (_08043_, _08041_, _07539_);
  nor (_08044_, _08038_, _06802_);
  nor (_08045_, _08044_, _08039_);
  nor (_08046_, _08045_, _07545_);
  nor (_08047_, _08046_, _08043_);
  nor (_08048_, _08047_, _08042_);
  nor (_08049_, _08043_, _08042_);
  and (_08050_, _08045_, _07545_);
  nor (_08051_, _08050_, _08046_);
  and (_08052_, _08051_, _08049_);
  not (_08053_, _08052_);
  and (_08054_, _06839_, _06710_);
  and (_08055_, _08054_, \oc8051_golden_model_1.PSW [7]);
  nor (_08056_, _08055_, _06664_);
  nor (_08057_, _08056_, _08038_);
  nor (_08058_, _08057_, _07644_);
  and (_08059_, _08057_, _07644_);
  nor (_08060_, _08059_, _08058_);
  nor (_08061_, _08037_, _06710_);
  nor (_08062_, _08061_, _08055_);
  nor (_08063_, _08062_, _07650_);
  and (_08064_, _08062_, _07650_);
  nor (_08065_, _08064_, _08063_);
  and (_08066_, _08065_, _08060_);
  and (_08067_, _06617_, \oc8051_golden_model_1.PSW [7]);
  nor (_08068_, _08067_, _06572_);
  nor (_08069_, _08068_, _08037_);
  and (_08070_, _08069_, _03269_);
  nor (_08071_, _08069_, _03269_);
  nor (_08072_, _06617_, \oc8051_golden_model_1.PSW [7]);
  nor (_08073_, _08072_, _08067_);
  nor (_08074_, _08073_, _03344_);
  nor (_08075_, _08074_, _08071_);
  nor (_08076_, _08075_, _08070_);
  not (_08077_, _08076_);
  and (_08078_, _08077_, _08066_);
  not (_08079_, _08078_);
  and (_08080_, _08064_, _08060_);
  nor (_08081_, _08080_, _08059_);
  and (_08082_, _08081_, _08079_);
  nor (_08083_, _08071_, _08070_);
  and (_08084_, _08073_, _03344_);
  nor (_08085_, _08074_, _08084_);
  and (_08086_, _08085_, _08083_);
  and (_08087_, _08086_, _08066_);
  nor (_08088_, _08087_, _08082_);
  nor (_08089_, _08088_, _08053_);
  nor (_08090_, _08089_, _08048_);
  nor (_08091_, _08090_, _08036_);
  or (_08092_, _08091_, _08035_);
  or (_08093_, _08092_, _08031_);
  nand (_08094_, _08092_, _08031_);
  and (_08095_, _08094_, _08093_);
  or (_08096_, _08095_, _08024_);
  nor (_08097_, _04775_, _03862_);
  and (_08098_, _08097_, _04663_);
  not (_08099_, _08098_);
  nand (_08100_, _08099_, _05253_);
  not (_08101_, _03536_);
  nor (_08102_, _06160_, _08101_);
  not (_08103_, _04007_);
  or (_08104_, _06114_, _08103_);
  nor (_08105_, _03208_, _03221_);
  not (_08106_, _08105_);
  nor (_08107_, _08106_, _05253_);
  and (_08108_, _03607_, _04003_);
  or (_08109_, _08108_, \oc8051_golden_model_1.ACC [7]);
  nand (_08110_, _08108_, \oc8051_golden_model_1.ACC [7]);
  and (_08111_, _08110_, _08109_);
  and (_08112_, _08111_, _08106_);
  or (_08113_, _08112_, _04007_);
  or (_08114_, _08113_, _08107_);
  and (_08115_, _08114_, _08101_);
  and (_08116_, _08115_, _08104_);
  or (_08117_, _08116_, _08102_);
  and (_08118_, _03607_, _03535_);
  nor (_08119_, _08118_, _03534_);
  and (_08120_, _08119_, _08117_);
  and (_08121_, _03607_, _03468_);
  and (_08122_, _06133_, _05312_);
  nor (_08123_, _08122_, _07935_);
  nor (_08124_, _08123_, _04432_);
  or (_08125_, _08124_, _08121_);
  or (_08126_, _08125_, _08120_);
  nor (_08127_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_08128_, _08127_, _07644_);
  and (_08129_, _08128_, _07511_);
  and (_08130_, _08129_, \oc8051_golden_model_1.ACC [6]);
  and (_08131_, _08130_, \oc8051_golden_model_1.ACC [7]);
  nor (_08132_, _08130_, \oc8051_golden_model_1.ACC [7]);
  nor (_08133_, _08132_, _08131_);
  and (_08134_, _08128_, \oc8051_golden_model_1.ACC [4]);
  nor (_08135_, _08134_, \oc8051_golden_model_1.ACC [5]);
  nor (_08136_, _08135_, _08129_);
  nor (_08137_, _08129_, \oc8051_golden_model_1.ACC [6]);
  nor (_08138_, _08137_, _08130_);
  nor (_08139_, _08138_, _08136_);
  not (_08140_, _08139_);
  and (_08141_, _08140_, _08133_);
  nor (_08142_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_08143_, _08142_, _08139_);
  nor (_08144_, _08143_, _08133_);
  nor (_08145_, _08144_, _08141_);
  not (_08146_, _08145_);
  nand (_08147_, _08146_, _08121_);
  and (_08148_, _08147_, _03532_);
  and (_08149_, _08148_, _08126_);
  nor (_08150_, _05937_, _06440_);
  and (_08151_, _05980_, _05937_);
  nor (_08152_, _08151_, _08150_);
  nor (_08153_, _08152_, _03470_);
  nor (_08154_, _07938_, _04457_);
  or (_08155_, _08154_, _08099_);
  or (_08156_, _08155_, _08153_);
  or (_08157_, _08156_, _08149_);
  and (_08158_, _08157_, _08100_);
  or (_08159_, _08158_, _04029_);
  not (_08160_, _04029_);
  or (_08161_, _06114_, _08160_);
  and (_08162_, _08161_, _03531_);
  and (_08163_, _08162_, _08159_);
  and (_08164_, _03607_, _03463_);
  nor (_08165_, _06160_, _03531_);
  or (_08166_, _08165_, _08164_);
  or (_08167_, _08166_, _08163_);
  nand (_08168_, _08164_, _07644_);
  and (_08169_, _08168_, _08167_);
  or (_08170_, _08169_, _03465_);
  and (_08171_, _05975_, _05937_);
  nor (_08172_, _08171_, _08150_);
  nand (_08173_, _08172_, _03465_);
  and (_08174_, _08173_, _03459_);
  and (_08175_, _08174_, _08170_);
  and (_08176_, _08151_, _06165_);
  nor (_08177_, _08176_, _08150_);
  nor (_08178_, _08177_, _03459_);
  or (_08179_, _08178_, _06933_);
  or (_08180_, _08179_, _08175_);
  nor (_08181_, _07411_, _07409_);
  nor (_08182_, _08181_, _07412_);
  or (_08183_, _08182_, _07447_);
  and (_08184_, _03561_, _03218_);
  not (_08185_, _08184_);
  nor (_08186_, _06899_, _03229_);
  and (_08187_, _03575_, _03218_);
  nor (_08188_, _08187_, _04063_);
  not (_08189_, _08188_);
  nor (_08190_, _08189_, _08186_);
  and (_08191_, _08190_, _08185_);
  and (_08192_, _08191_, _08183_);
  and (_08193_, _08192_, _08180_);
  not (_08194_, _08191_);
  not (_08195_, _05417_);
  and (_08196_, _05894_, \oc8051_golden_model_1.PSW [7]);
  and (_08197_, _08196_, _08195_);
  nor (_08198_, _08197_, _05253_);
  and (_08199_, _08197_, _05253_);
  nor (_08200_, _08199_, _08198_);
  and (_08201_, _08200_, \oc8051_golden_model_1.ACC [7]);
  nor (_08202_, _08200_, \oc8051_golden_model_1.ACC [7]);
  nor (_08203_, _08202_, _08201_);
  nor (_08204_, _08196_, _08195_);
  nor (_08205_, _08204_, _08197_);
  nor (_08206_, _08205_, _07495_);
  and (_08207_, _08205_, _07495_);
  and (_08208_, _05890_, \oc8051_golden_model_1.PSW [7]);
  and (_08209_, _08208_, _05891_);
  and (_08210_, _08209_, _05889_);
  nor (_08211_, _08210_, _05888_);
  nor (_08212_, _08211_, _08196_);
  and (_08213_, _08212_, _07539_);
  nor (_08214_, _08212_, _07539_);
  nor (_08215_, _08214_, _08213_);
  nor (_08216_, _08209_, _05889_);
  nor (_08217_, _08216_, _08210_);
  nor (_08218_, _08217_, _07545_);
  and (_08219_, _08217_, _07545_);
  nor (_08220_, _08219_, _08218_);
  and (_08221_, _08220_, _08215_);
  and (_08222_, _05890_, _05074_);
  and (_08223_, _08222_, \oc8051_golden_model_1.PSW [7]);
  nor (_08224_, _08223_, _06023_);
  nor (_08225_, _08224_, _08209_);
  nor (_08226_, _08225_, _07644_);
  and (_08227_, _08225_, _07644_);
  nor (_08228_, _08227_, _08226_);
  nor (_08229_, _08208_, _05074_);
  nor (_08230_, _08229_, _08223_);
  nor (_08231_, _08230_, _07650_);
  and (_08232_, _08230_, _07650_);
  nor (_08233_, _08232_, _08231_);
  and (_08234_, _08233_, _08228_);
  and (_08235_, _04429_, \oc8051_golden_model_1.PSW [7]);
  nor (_08236_, _08235_, _04636_);
  nor (_08237_, _08236_, _08208_);
  nor (_08238_, _08237_, _03269_);
  and (_08239_, _08237_, _03269_);
  and (_08240_, _04462_, _07982_);
  nor (_08241_, _08240_, _08235_);
  and (_08242_, _08241_, _03344_);
  nor (_08243_, _08242_, _08239_);
  or (_08244_, _08243_, _08238_);
  nand (_08245_, _08244_, _08234_);
  not (_08246_, _08226_);
  nand (_08247_, _08231_, _08228_);
  and (_08248_, _08247_, _08246_);
  and (_08249_, _08248_, _08245_);
  not (_08250_, _08249_);
  and (_08251_, _08250_, _08221_);
  not (_08252_, _08251_);
  and (_08253_, _08218_, _08215_);
  nor (_08254_, _08253_, _08214_);
  and (_08255_, _08254_, _08252_);
  nor (_08256_, _08255_, _08207_);
  or (_08257_, _08256_, _08206_);
  or (_08258_, _08257_, _08203_);
  nand (_08259_, _08257_, _08203_);
  and (_08260_, _08259_, _08258_);
  and (_08261_, _08260_, _08194_);
  or (_08262_, _08261_, _04066_);
  or (_08263_, _08262_, _08193_);
  and (_08264_, _08263_, _03599_);
  and (_08265_, _08264_, _08096_);
  nor (_08266_, _07940_, _03594_);
  not (_08267_, _08266_);
  and (_08268_, _06160_, _06440_);
  nor (_08269_, _06160_, _06440_);
  nor (_08270_, _08269_, _08268_);
  not (_08271_, _05438_);
  and (_08272_, _05465_, _08271_);
  nor (_08273_, _05445_, _05439_);
  and (_08274_, _08273_, _05453_);
  and (_08275_, _05289_, \oc8051_golden_model_1.P2INREG [6]);
  and (_08276_, _05293_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_08277_, _08276_, _08275_);
  and (_08278_, _05284_, \oc8051_golden_model_1.P1INREG [6]);
  and (_08279_, _05298_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_08280_, _08279_, _08278_);
  and (_08281_, _08280_, _08277_);
  and (_08282_, _08281_, _08274_);
  and (_08283_, _08282_, _08272_);
  and (_08284_, _05450_, _05424_);
  and (_08285_, _08284_, _05437_);
  and (_08286_, _08285_, _08283_);
  and (_08287_, _08286_, _05418_);
  and (_08288_, _08287_, \oc8051_golden_model_1.ACC [6]);
  nor (_08289_, _08287_, \oc8051_golden_model_1.ACC [6]);
  nor (_08290_, _08289_, _08288_);
  and (_08291_, _05298_, \oc8051_golden_model_1.P0INREG [5]);
  not (_08292_, _08291_);
  and (_08293_, _08292_, _05560_);
  and (_08294_, _05284_, \oc8051_golden_model_1.P1INREG [5]);
  not (_08295_, _08294_);
  not (_08296_, _05566_);
  and (_08297_, _05289_, \oc8051_golden_model_1.P2INREG [5]);
  and (_08298_, _05293_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_08299_, _08298_, _08297_);
  and (_08300_, _08299_, _08296_);
  and (_08301_, _08300_, _08295_);
  and (_08302_, _08301_, _05564_);
  and (_08303_, _08302_, _08293_);
  and (_08304_, _08303_, _05547_);
  and (_08305_, _08304_, _05527_);
  and (_08306_, _08305_, \oc8051_golden_model_1.ACC [5]);
  nor (_08307_, _08305_, \oc8051_golden_model_1.ACC [5]);
  and (_08308_, _05298_, \oc8051_golden_model_1.P0INREG [4]);
  not (_08309_, _08308_);
  and (_08310_, _05284_, \oc8051_golden_model_1.P1INREG [4]);
  not (_08311_, _08310_);
  and (_08312_, _05289_, \oc8051_golden_model_1.P2INREG [4]);
  and (_08313_, _05293_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08314_, _08313_, _08312_);
  and (_08315_, _08314_, _08311_);
  and (_08316_, _08315_, _05839_);
  and (_08317_, _08316_, _08309_);
  and (_08318_, _08317_, _05859_);
  and (_08319_, _08318_, _05877_);
  and (_08320_, _08319_, _05832_);
  and (_08321_, _08320_, \oc8051_golden_model_1.ACC [4]);
  and (_08322_, _05298_, \oc8051_golden_model_1.P0INREG [3]);
  not (_08323_, _08322_);
  and (_08324_, _05284_, \oc8051_golden_model_1.P1INREG [3]);
  not (_08325_, _08324_);
  and (_08326_, _05289_, \oc8051_golden_model_1.P2INREG [3]);
  and (_08327_, _05293_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08328_, _08327_, _08326_);
  and (_08329_, _08328_, _08325_);
  and (_08330_, _08329_, _05586_);
  and (_08331_, _08330_, _08323_);
  and (_08332_, _08331_, _05604_);
  and (_08333_, _08332_, _05622_);
  and (_08334_, _08333_, _05577_);
  and (_08335_, _08334_, \oc8051_golden_model_1.ACC [3]);
  nor (_08336_, _08334_, \oc8051_golden_model_1.ACC [3]);
  and (_08337_, _05284_, \oc8051_golden_model_1.P1INREG [2]);
  not (_08338_, _08337_);
  and (_08339_, _05289_, \oc8051_golden_model_1.P2INREG [2]);
  and (_08340_, _05293_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08341_, _08340_, _08339_);
  and (_08342_, _08341_, _05732_);
  and (_08343_, _08342_, _08338_);
  and (_08344_, _05298_, \oc8051_golden_model_1.P0INREG [2]);
  not (_08345_, _08344_);
  and (_08346_, _08345_, _05748_);
  and (_08347_, _08346_, _08343_);
  and (_08348_, _08347_, _05730_);
  and (_08349_, _08348_, _05769_);
  and (_08350_, _08349_, _05724_);
  and (_08351_, _08350_, \oc8051_golden_model_1.ACC [2]);
  and (_08352_, _05298_, \oc8051_golden_model_1.P0INREG [1]);
  not (_08353_, _08352_);
  and (_08354_, _05284_, \oc8051_golden_model_1.P1INREG [1]);
  not (_08355_, _08354_);
  and (_08356_, _05289_, \oc8051_golden_model_1.P2INREG [1]);
  and (_08357_, _05293_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_08358_, _08357_, _08356_);
  and (_08359_, _08358_, _08355_);
  and (_08360_, _08359_, _05635_);
  and (_08361_, _08360_, _08353_);
  and (_08362_, _08361_, _05653_);
  and (_08363_, _08362_, _05671_);
  and (_08364_, _08363_, _05626_);
  and (_08365_, _08364_, \oc8051_golden_model_1.ACC [1]);
  nor (_08366_, _08364_, \oc8051_golden_model_1.ACC [1]);
  and (_08367_, _05284_, \oc8051_golden_model_1.P1INREG [0]);
  not (_08368_, _08367_);
  and (_08369_, _05289_, \oc8051_golden_model_1.P2INREG [0]);
  and (_08370_, _05293_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_08371_, _08370_, _08369_);
  and (_08372_, _08371_, _05683_);
  and (_08373_, _08372_, _08368_);
  and (_08374_, _05298_, \oc8051_golden_model_1.P0INREG [0]);
  not (_08375_, _08374_);
  and (_08376_, _08375_, _05699_);
  and (_08377_, _08376_, _08373_);
  and (_08378_, _08377_, _05681_);
  and (_08379_, _08378_, _05720_);
  and (_08380_, _08379_, _05675_);
  nor (_08381_, _08380_, \oc8051_golden_model_1.ACC [0]);
  nor (_08382_, _08381_, _08366_);
  or (_08383_, _08382_, _08365_);
  nor (_08384_, _08350_, \oc8051_golden_model_1.ACC [2]);
  nor (_08385_, _08384_, _08351_);
  and (_08386_, _08385_, _08383_);
  nor (_08387_, _08386_, _08351_);
  nor (_08388_, _08387_, _08336_);
  or (_08389_, _08388_, _08335_);
  nor (_08390_, _08320_, \oc8051_golden_model_1.ACC [4]);
  nor (_08391_, _08390_, _08321_);
  and (_08392_, _08391_, _08389_);
  nor (_08393_, _08392_, _08321_);
  nor (_08394_, _08393_, _08307_);
  or (_08395_, _08394_, _08306_);
  and (_08396_, _08395_, _08290_);
  nor (_08397_, _08396_, _08288_);
  and (_08398_, _08397_, _08270_);
  nor (_08399_, _08397_, _08270_);
  nor (_08400_, _08399_, _08398_);
  not (_08401_, _08400_);
  nor (_08402_, _08395_, _08290_);
  nor (_08403_, _08402_, _08396_);
  nor (_08404_, _08306_, _08307_);
  not (_08405_, _08404_);
  and (_08406_, _08405_, _08393_);
  nor (_08407_, _08405_, _08393_);
  nor (_08408_, _08407_, _08406_);
  nor (_08409_, _08391_, _08389_);
  nor (_08410_, _08409_, _08392_);
  nor (_08411_, _08335_, _08336_);
  and (_08412_, _08411_, _08385_);
  nor (_08413_, _08365_, _08366_);
  and (_08414_, _08380_, \oc8051_golden_model_1.ACC [0]);
  nor (_08415_, _08414_, _08381_);
  and (_08416_, _08415_, _08413_);
  and (_08417_, _08416_, _08412_);
  and (_08418_, _08417_, \oc8051_golden_model_1.PSW [7]);
  not (_08419_, _08418_);
  nor (_08420_, _08419_, _08410_);
  not (_08421_, _08420_);
  nor (_08422_, _08421_, _08408_);
  not (_08423_, _08422_);
  nor (_08424_, _08423_, _08403_);
  nor (_08425_, _08424_, _08401_);
  and (_08426_, _08424_, _08401_);
  or (_08427_, _08426_, _07940_);
  or (_08428_, _08427_, _08425_);
  and (_08429_, _08428_, _08267_);
  or (_08430_, _08429_, _08265_);
  and (_08431_, _08430_, _08023_);
  or (_08432_, _08431_, _03334_);
  or (_08433_, _03409_, _03233_);
  and (_08434_, _08433_, _03453_);
  and (_08435_, _08434_, _08432_);
  not (_08436_, _05937_);
  nor (_08437_, _05962_, _08436_);
  nor (_08438_, _08437_, _08150_);
  nor (_08439_, _08438_, _03453_);
  or (_08440_, _08439_, _07454_);
  or (_08441_, _08440_, _08435_);
  and (_08442_, _08441_, _07939_);
  or (_08443_, _08442_, _04082_);
  and (_08444_, _06114_, _05312_);
  or (_08445_, _08444_, _07935_);
  or (_08446_, _08445_, _04500_);
  and (_08447_, _08446_, _03521_);
  and (_08448_, _08447_, _08443_);
  nor (_08449_, _06421_, _07936_);
  nor (_08450_, _08449_, _07935_);
  nor (_08451_, _08450_, _03521_);
  or (_08452_, _08451_, _07468_);
  or (_08453_, _08452_, _08448_);
  not (_08454_, _07488_);
  nand (_08455_, _08454_, _07468_);
  and (_08456_, _08455_, _08453_);
  or (_08457_, _08456_, _03262_);
  or (_08458_, _03409_, _03263_);
  and (_08459_, _08458_, _08457_);
  or (_08460_, _08459_, _03624_);
  and (_08461_, _03607_, _03167_);
  not (_08462_, _08461_);
  and (_08463_, _06227_, _05312_);
  nor (_08464_, _08463_, _07935_);
  nand (_08465_, _08464_, _03624_);
  and (_08466_, _08465_, _08462_);
  and (_08467_, _08466_, _08460_);
  and (_08468_, _08461_, _03409_);
  and (_08469_, _03572_, _03171_);
  or (_08470_, _08469_, _08468_);
  or (_08471_, _08470_, _08467_);
  not (_08472_, _08469_);
  or (_08473_, _08472_, _07882_);
  and (_08474_, _03566_, _03171_);
  nor (_08475_, _04330_, _08474_);
  and (_08476_, _03640_, _03171_);
  not (_08477_, _08476_);
  and (_08478_, _08477_, _08475_);
  and (_08479_, _08478_, _08473_);
  and (_08480_, _08479_, _08471_);
  and (_08481_, _04005_, _03171_);
  not (_08482_, _08478_);
  and (_08483_, _08482_, _07882_);
  or (_08484_, _08483_, _08481_);
  or (_08485_, _08484_, _08480_);
  not (_08486_, _03746_);
  not (_08487_, _08481_);
  and (_08488_, _06114_, \oc8051_golden_model_1.ACC [7]);
  nor (_08489_, _08488_, _07924_);
  or (_08490_, _08489_, _08487_);
  and (_08491_, _08490_, _08486_);
  and (_08492_, _08491_, _08485_);
  nor (_08493_, _07929_, _03746_);
  not (_08494_, _08493_);
  or (_08495_, _07929_, _06443_);
  and (_08496_, _08495_, _08494_);
  or (_08497_, _08496_, _08492_);
  and (_08498_, _08497_, _07934_);
  or (_08499_, _08498_, _03623_);
  and (_08500_, _06436_, _05312_);
  nor (_08501_, _08500_, _07935_);
  nand (_08502_, _08501_, _03623_);
  and (_08503_, _08502_, _03745_);
  and (_08504_, _08503_, _08499_);
  and (_08505_, _07935_, _03744_);
  nand (_08506_, _03181_, _02954_);
  not (_08507_, _08506_);
  or (_08508_, _08507_, _08505_);
  or (_08509_, _08508_, _08504_);
  not (_08510_, _04141_);
  or (_08511_, _08506_, _07881_);
  and (_08512_, _08511_, _08510_);
  and (_08513_, _08512_, _08509_);
  and (_08514_, _08488_, _04141_);
  or (_08515_, _08514_, _03735_);
  or (_08516_, _08515_, _08513_);
  and (_08517_, _03607_, _03181_);
  not (_08518_, _08517_);
  not (_08519_, _03735_);
  or (_08520_, _06441_, _08519_);
  and (_08521_, _08520_, _08518_);
  and (_08522_, _08521_, _08516_);
  and (_08523_, _08517_, _07931_);
  or (_08524_, _08523_, _08522_);
  and (_08525_, _08524_, _04523_);
  or (_08526_, _08464_, _06442_);
  nor (_08527_, _08526_, _04523_);
  or (_08528_, _08527_, _07927_);
  or (_08529_, _08528_, _08525_);
  and (_08530_, _08529_, _07928_);
  nor (_08531_, _05140_, _07926_);
  or (_08532_, _08531_, _08530_);
  not (_08533_, _04157_);
  nand (_08534_, _08531_, _07880_);
  and (_08535_, _08534_, _08533_);
  and (_08536_, _08535_, _08532_);
  nor (_08537_, _07880_, _08533_);
  or (_08538_, _08537_, _07923_);
  or (_08539_, _08538_, _08536_);
  and (_08540_, _08539_, _07925_);
  or (_08541_, _08540_, _03739_);
  and (_08542_, _03607_, _03177_);
  not (_08543_, _08542_);
  nand (_08544_, _06442_, _03739_);
  and (_08545_, _08544_, _08543_);
  and (_08546_, _08545_, _08541_);
  nor (_08547_, _08543_, _07932_);
  or (_08548_, _08547_, _08546_);
  and (_08549_, _08548_, _06453_);
  nor (_08550_, _06434_, _07936_);
  nor (_08551_, _08550_, _07935_);
  nor (_08552_, _08551_, _06453_);
  and (_08553_, _03572_, _03190_);
  and (_08554_, _03578_, _03190_);
  or (_08555_, _08554_, _04170_);
  or (_08556_, _08555_, _08553_);
  or (_08557_, _08556_, _08552_);
  or (_08558_, _08557_, _08549_);
  and (_08559_, _03561_, _03190_);
  not (_08560_, _08559_);
  nor (_08561_, _06899_, _04166_);
  nor (_08562_, _05140_, _04166_);
  nor (_08563_, _08562_, _08561_);
  and (_08564_, _08563_, _08560_);
  and (_08565_, _03640_, _03190_);
  not (_08566_, _08565_);
  and (_08567_, _08205_, \oc8051_golden_model_1.ACC [6]);
  nor (_08568_, _08206_, _08207_);
  and (_08569_, _08212_, \oc8051_golden_model_1.ACC [5]);
  and (_08570_, _08217_, \oc8051_golden_model_1.ACC [4]);
  and (_08571_, _08225_, \oc8051_golden_model_1.ACC [3]);
  and (_08572_, _08230_, \oc8051_golden_model_1.ACC [2]);
  and (_08573_, _08237_, \oc8051_golden_model_1.ACC [1]);
  nor (_08574_, _08239_, _08238_);
  and (_08575_, _08241_, \oc8051_golden_model_1.ACC [0]);
  not (_08576_, _08575_);
  nor (_08577_, _08576_, _08574_);
  nor (_08578_, _08577_, _08573_);
  nor (_08579_, _08578_, _08233_);
  nor (_08580_, _08579_, _08572_);
  nor (_08581_, _08580_, _08228_);
  nor (_08582_, _08581_, _08571_);
  nor (_08583_, _08582_, _08220_);
  nor (_08584_, _08583_, _08570_);
  nor (_08585_, _08584_, _08215_);
  nor (_08586_, _08585_, _08569_);
  nor (_08587_, _08586_, _08568_);
  nor (_08588_, _08587_, _08567_);
  nor (_08589_, _08588_, _08203_);
  and (_08590_, _08588_, _08203_);
  nor (_08591_, _08590_, _08589_);
  and (_08592_, _08591_, _08566_);
  or (_08593_, _08592_, _08564_);
  and (_08594_, _08593_, _08558_);
  and (_08595_, _04005_, _03190_);
  and (_08596_, _08591_, _08565_);
  or (_08597_, _08596_, _08595_);
  or (_08598_, _08597_, _08594_);
  not (_08599_, _08595_);
  and (_08600_, _08034_, \oc8051_golden_model_1.ACC [6]);
  nor (_08601_, _08035_, _08036_);
  and (_08602_, _08041_, \oc8051_golden_model_1.ACC [5]);
  and (_08603_, _08045_, \oc8051_golden_model_1.ACC [4]);
  and (_08604_, _08057_, \oc8051_golden_model_1.ACC [3]);
  and (_08605_, _08062_, \oc8051_golden_model_1.ACC [2]);
  and (_08606_, _08069_, \oc8051_golden_model_1.ACC [1]);
  and (_08607_, _08073_, \oc8051_golden_model_1.ACC [0]);
  not (_08608_, _08607_);
  nor (_08609_, _08608_, _08083_);
  nor (_08610_, _08609_, _08606_);
  nor (_08611_, _08610_, _08065_);
  nor (_08612_, _08611_, _08605_);
  nor (_08613_, _08612_, _08060_);
  nor (_08614_, _08613_, _08604_);
  nor (_08615_, _08614_, _08051_);
  nor (_08616_, _08615_, _08603_);
  nor (_08617_, _08616_, _08049_);
  nor (_08618_, _08617_, _08602_);
  nor (_08619_, _08618_, _08601_);
  nor (_08620_, _08619_, _08600_);
  nor (_08621_, _08620_, _08031_);
  and (_08622_, _08620_, _08031_);
  nor (_08623_, _08622_, _08621_);
  or (_08624_, _08623_, _08599_);
  and (_08625_, _08624_, _03732_);
  and (_08626_, _08625_, _08598_);
  and (_08627_, _03607_, _03190_);
  nor (_08628_, _08627_, _03731_);
  not (_08629_, _08628_);
  not (_08630_, _08287_);
  not (_08631_, _08305_);
  not (_08632_, _08320_);
  not (_08633_, _08334_);
  not (_08634_, _08350_);
  not (_08635_, _08364_);
  nor (_08636_, _08380_, _07982_);
  and (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _08634_);
  and (_08639_, _08638_, _08633_);
  and (_08640_, _08639_, _08632_);
  and (_08641_, _08640_, _08631_);
  and (_08642_, _08641_, _08630_);
  nor (_08643_, _08642_, _06160_);
  and (_08644_, _08642_, _06160_);
  nor (_08645_, _08644_, _08643_);
  and (_08646_, _08645_, \oc8051_golden_model_1.ACC [7]);
  nor (_08647_, _08645_, \oc8051_golden_model_1.ACC [7]);
  nor (_08648_, _08647_, _08646_);
  nor (_08649_, _08641_, _08630_);
  nor (_08650_, _08649_, _08642_);
  and (_08651_, _08650_, \oc8051_golden_model_1.ACC [6]);
  and (_08652_, _08650_, _07495_);
  nor (_08653_, _08650_, _07495_);
  nor (_08654_, _08653_, _08652_);
  nor (_08655_, _08640_, _08631_);
  nor (_08656_, _08655_, _08641_);
  and (_08657_, _08656_, \oc8051_golden_model_1.ACC [5]);
  nor (_08658_, _08656_, _07539_);
  and (_08659_, _08656_, _07539_);
  nor (_08660_, _08659_, _08658_);
  nor (_08661_, _08639_, _08632_);
  nor (_08662_, _08661_, _08640_);
  and (_08663_, _08662_, \oc8051_golden_model_1.ACC [4]);
  nor (_08664_, _08662_, _07545_);
  and (_08665_, _08662_, _07545_);
  nor (_08666_, _08665_, _08664_);
  nor (_08667_, _08638_, _08633_);
  nor (_08668_, _08667_, _08639_);
  and (_08669_, _08668_, \oc8051_golden_model_1.ACC [3]);
  nor (_08670_, _08668_, _07644_);
  and (_08671_, _08668_, _07644_);
  nor (_08672_, _08671_, _08670_);
  nor (_08673_, _08637_, _08634_);
  nor (_08674_, _08673_, _08638_);
  and (_08675_, _08674_, \oc8051_golden_model_1.ACC [2]);
  nor (_08676_, _08674_, _07650_);
  and (_08677_, _08674_, _07650_);
  nor (_08678_, _08677_, _08676_);
  nor (_08679_, _08636_, _08635_);
  nor (_08680_, _08679_, _08637_);
  and (_08681_, _08680_, \oc8051_golden_model_1.ACC [1]);
  and (_08682_, _08680_, _03269_);
  nor (_08683_, _08680_, _03269_);
  nor (_08684_, _08683_, _08682_);
  and (_08685_, _08380_, _07982_);
  nor (_08686_, _08685_, _08636_);
  and (_08687_, _08686_, \oc8051_golden_model_1.ACC [0]);
  not (_08688_, _08687_);
  nor (_08689_, _08688_, _08684_);
  nor (_08690_, _08689_, _08681_);
  nor (_08691_, _08690_, _08678_);
  nor (_08692_, _08691_, _08675_);
  nor (_08693_, _08692_, _08672_);
  nor (_08694_, _08693_, _08669_);
  nor (_08695_, _08694_, _08666_);
  nor (_08696_, _08695_, _08663_);
  nor (_08697_, _08696_, _08660_);
  nor (_08698_, _08697_, _08657_);
  nor (_08699_, _08698_, _08654_);
  nor (_08700_, _08699_, _08651_);
  nor (_08701_, _08700_, _08648_);
  and (_08702_, _08700_, _08648_);
  nor (_08703_, _08702_, _08701_);
  or (_08704_, _08703_, _08627_);
  and (_08705_, _08704_, _08629_);
  or (_08706_, _08705_, _08626_);
  and (_08707_, _03610_, _03190_);
  not (_08708_, _08707_);
  not (_08709_, _08627_);
  and (_08710_, _07954_, \oc8051_golden_model_1.ACC [6]);
  and (_08711_, _07960_, \oc8051_golden_model_1.ACC [5]);
  and (_08712_, _07965_, \oc8051_golden_model_1.ACC [4]);
  and (_08713_, _07971_, \oc8051_golden_model_1.ACC [3]);
  and (_08714_, _07976_, \oc8051_golden_model_1.ACC [2]);
  and (_08715_, _08002_, \oc8051_golden_model_1.ACC [1]);
  nor (_08716_, _08003_, _08004_);
  and (_08717_, _07985_, \oc8051_golden_model_1.ACC [0]);
  not (_08718_, _08717_);
  nor (_08719_, _08718_, _08716_);
  nor (_08720_, _08719_, _08715_);
  nor (_08721_, _08720_, _07979_);
  nor (_08722_, _08721_, _08714_);
  nor (_08723_, _08722_, _07974_);
  nor (_08724_, _08723_, _08713_);
  nor (_08725_, _08724_, _07968_);
  nor (_08726_, _08725_, _08712_);
  nor (_08727_, _08726_, _07963_);
  nor (_08728_, _08727_, _08711_);
  nor (_08729_, _08728_, _07957_);
  nor (_08730_, _08729_, _08710_);
  nor (_08731_, _08730_, _07951_);
  and (_08732_, _08730_, _07951_);
  nor (_08733_, _08732_, _08731_);
  or (_08734_, _08733_, _08709_);
  and (_08735_, _08734_, _08708_);
  and (_08736_, _08735_, _08706_);
  and (_08737_, _08707_, \oc8051_golden_model_1.ACC [6]);
  or (_08738_, _08737_, _07920_);
  or (_08739_, _08738_, _08736_);
  and (_08740_, _08739_, _07922_);
  or (_08741_, _08740_, _04184_);
  not (_08742_, _04184_);
  and (_08743_, _06526_, \oc8051_golden_model_1.ACC [6]);
  nor (_08744_, _06526_, \oc8051_golden_model_1.ACC [6]);
  nor (_08745_, _08744_, _08743_);
  nor (_08746_, _06757_, \oc8051_golden_model_1.ACC [5]);
  not (_08747_, _08746_);
  and (_08748_, _06757_, \oc8051_golden_model_1.ACC [5]);
  not (_08749_, _08748_);
  and (_08750_, _06802_, \oc8051_golden_model_1.ACC [4]);
  nor (_08751_, _06802_, \oc8051_golden_model_1.ACC [4]);
  nor (_08752_, _08751_, _08750_);
  nor (_08753_, _06664_, \oc8051_golden_model_1.ACC [3]);
  not (_08754_, _08753_);
  and (_08755_, _06664_, \oc8051_golden_model_1.ACC [3]);
  not (_08756_, _08755_);
  and (_08757_, _06710_, \oc8051_golden_model_1.ACC [2]);
  nor (_08758_, _06710_, \oc8051_golden_model_1.ACC [2]);
  nor (_08759_, _08758_, _08757_);
  not (_08760_, _08759_);
  and (_08761_, _06572_, \oc8051_golden_model_1.ACC [1]);
  nor (_08762_, _06572_, \oc8051_golden_model_1.ACC [1]);
  nor (_08763_, _08762_, _08761_);
  and (_08764_, _06617_, \oc8051_golden_model_1.ACC [0]);
  and (_08765_, _08764_, _08763_);
  nor (_08766_, _08765_, _08761_);
  nor (_08767_, _08766_, _08760_);
  nor (_08768_, _08767_, _08757_);
  nand (_08769_, _08768_, _08756_);
  and (_08770_, _08769_, _08754_);
  and (_08771_, _08770_, _08752_);
  nor (_08772_, _08771_, _08750_);
  nand (_08773_, _08772_, _08749_);
  and (_08774_, _08773_, _08747_);
  and (_08775_, _08774_, _08745_);
  nor (_08776_, _08775_, _08743_);
  nor (_08777_, _08776_, _08489_);
  and (_08778_, _08776_, _08489_);
  or (_08779_, _08778_, _08777_);
  or (_08780_, _08779_, _08742_);
  and (_08781_, _08780_, _03480_);
  and (_08782_, _08781_, _08741_);
  and (_08783_, _03607_, _03188_);
  nor (_08784_, _08783_, _03478_);
  not (_08785_, _08784_);
  not (_08786_, _08783_);
  nor (_08787_, _08287_, _07495_);
  nor (_08788_, _08305_, _07539_);
  nor (_08789_, _08320_, _07545_);
  not (_08790_, _08391_);
  nor (_08791_, _08350_, _07650_);
  nor (_08792_, _08364_, _03269_);
  nor (_08793_, _08380_, _03344_);
  not (_08794_, _08793_);
  nor (_08795_, _08794_, _08413_);
  nor (_08796_, _08795_, _08792_);
  nor (_08797_, _08796_, _08385_);
  nor (_08798_, _08797_, _08791_);
  nor (_08799_, _08798_, _08334_);
  or (_08800_, _08799_, \oc8051_golden_model_1.ACC [3]);
  nand (_08801_, _08798_, _08334_);
  and (_08802_, _08801_, _08800_);
  and (_08803_, _08802_, _08790_);
  nor (_08804_, _08803_, _08789_);
  nor (_08805_, _08804_, _08404_);
  nor (_08806_, _08805_, _08788_);
  nor (_08807_, _08806_, _08290_);
  nor (_08808_, _08807_, _08787_);
  nor (_08809_, _08808_, _08270_);
  and (_08810_, _08808_, _08270_);
  nor (_08811_, _08810_, _08809_);
  nand (_08812_, _08811_, _08786_);
  and (_08813_, _08812_, _08785_);
  or (_08814_, _08813_, _08782_);
  and (_08815_, _03610_, _03188_);
  not (_08816_, _08815_);
  nor (_08817_, _03511_, _07495_);
  and (_08818_, _03511_, _07495_);
  nor (_08819_, _08818_, _08817_);
  nor (_08820_, _03811_, _07539_);
  and (_08821_, _03811_, _07539_);
  nor (_08822_, _04257_, _07545_);
  and (_08823_, _04257_, _07545_);
  nor (_08824_, _08823_, _08822_);
  nor (_08825_, _03440_, _07644_);
  and (_08826_, _03440_, _07644_);
  nor (_08827_, _03944_, _07650_);
  and (_08828_, _03944_, _07650_);
  nor (_08829_, _08828_, _08827_);
  not (_08830_, _08829_);
  nor (_08831_, _03989_, _03344_);
  and (_08832_, _08831_, _07991_);
  nor (_08833_, _08832_, _07989_);
  nor (_08834_, _08833_, _08830_);
  nor (_08835_, _08834_, _08827_);
  nor (_08836_, _08835_, _08826_);
  or (_08837_, _08836_, _08825_);
  and (_08838_, _08837_, _08824_);
  nor (_08839_, _08838_, _08822_);
  nor (_08840_, _08839_, _08821_);
  or (_08841_, _08840_, _08820_);
  and (_08842_, _08841_, _08819_);
  nor (_08843_, _08842_, _08817_);
  nor (_08844_, _08843_, _07933_);
  and (_08845_, _08843_, _07933_);
  or (_08846_, _08845_, _08844_);
  or (_08847_, _08846_, _08786_);
  and (_08848_, _08847_, _08816_);
  and (_08849_, _08848_, _08814_);
  and (_08850_, _08815_, \oc8051_golden_model_1.ACC [6]);
  or (_08851_, _08850_, _03767_);
  or (_08852_, _08851_, _08849_);
  and (_08853_, _03607_, _03195_);
  not (_08854_, _08853_);
  nand (_08855_, _08123_, _03767_);
  and (_08856_, _08855_, _08854_);
  and (_08857_, _08856_, _08852_);
  and (_08858_, _03610_, _03195_);
  nor (_08859_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08860_, _08859_, _07590_);
  and (_08861_, _08860_, _07510_);
  and (_08862_, _08861_, _07495_);
  nor (_08863_, _08862_, _06440_);
  and (_08864_, _08862_, _06440_);
  nor (_08865_, _08864_, _08863_);
  nor (_08866_, _08865_, _08854_);
  or (_08867_, _08866_, _08858_);
  or (_08868_, _08867_, _08857_);
  nand (_08869_, _08858_, _07982_);
  and (_08870_, _08869_, _03446_);
  and (_08871_, _08870_, _08868_);
  nor (_08872_, _08172_, _03446_);
  or (_08873_, _08872_, _03473_);
  or (_08874_, _08873_, _08871_);
  and (_08875_, _03607_, _03193_);
  not (_08876_, _08875_);
  and (_08877_, _05886_, _05312_);
  nor (_08878_, _08877_, _07935_);
  nand (_08879_, _08878_, _03473_);
  and (_08880_, _08879_, _08876_);
  and (_08881_, _08880_, _08874_);
  and (_08882_, _03610_, _03193_);
  and (_08883_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08884_, _08883_, _07591_);
  nor (_08885_, _08884_, _07545_);
  and (_08886_, _08885_, \oc8051_golden_model_1.ACC [5]);
  and (_08887_, _08886_, \oc8051_golden_model_1.ACC [6]);
  nor (_08888_, _08887_, \oc8051_golden_model_1.ACC [7]);
  and (_08889_, _08887_, \oc8051_golden_model_1.ACC [7]);
  nor (_08890_, _08889_, _08888_);
  and (_08891_, _08890_, _08875_);
  or (_08892_, _08891_, _08882_);
  or (_08893_, _08892_, _08881_);
  nand (_08894_, _08882_, _03344_);
  and (_08895_, _08894_, _43189_);
  and (_08896_, _08895_, _08893_);
  or (_08897_, _08896_, _07879_);
  and (_40772_, _08897_, _42003_);
  not (_08898_, \oc8051_golden_model_1.DPL [7]);
  nor (_08899_, _43189_, _08898_);
  nor (_08900_, _05327_, _08898_);
  not (_08901_, _05327_);
  nor (_08902_, _06442_, _08901_);
  or (_08903_, _08902_, _08900_);
  and (_08904_, _08903_, _03741_);
  not (_08905_, _03625_);
  nor (_08906_, _08901_, _05253_);
  or (_08907_, _08906_, _08900_);
  or (_08908_, _08907_, _06903_);
  and (_08909_, _06133_, _05327_);
  or (_08910_, _08909_, _08900_);
  or (_08911_, _08910_, _04432_);
  and (_08912_, _05327_, \oc8051_golden_model_1.ACC [7]);
  or (_08913_, _08912_, _08900_);
  and (_08914_, _08913_, _04436_);
  nor (_08915_, _04436_, _08898_);
  or (_08916_, _08915_, _03534_);
  or (_08917_, _08916_, _08914_);
  and (_08918_, _08917_, _04457_);
  and (_08919_, _08918_, _08911_);
  and (_08920_, _08907_, _03527_);
  or (_08921_, _08920_, _03530_);
  or (_08922_, _08921_, _08919_);
  nor (_08923_, _03232_, _03213_);
  not (_08924_, _08923_);
  or (_08925_, _08913_, _03531_);
  and (_08926_, _08925_, _08924_);
  and (_08927_, _08926_, _08922_);
  and (_08928_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08929_, _08928_, \oc8051_golden_model_1.DPL [2]);
  and (_08930_, _08929_, \oc8051_golden_model_1.DPL [3]);
  and (_08931_, _08930_, \oc8051_golden_model_1.DPL [4]);
  and (_08932_, _08931_, \oc8051_golden_model_1.DPL [5]);
  and (_08933_, _08932_, \oc8051_golden_model_1.DPL [6]);
  nor (_08934_, _08933_, \oc8051_golden_model_1.DPL [7]);
  and (_08935_, _08933_, \oc8051_golden_model_1.DPL [7]);
  nor (_08936_, _08935_, _08934_);
  and (_08937_, _08936_, _08923_);
  or (_08938_, _08937_, _08927_);
  and (_08939_, _08938_, _03622_);
  nor (_08940_, _06226_, _03622_);
  or (_08942_, _08940_, _07454_);
  or (_08943_, _08942_, _08939_);
  and (_08944_, _08943_, _08908_);
  or (_08945_, _08944_, _04082_);
  and (_08946_, _06114_, _05327_);
  or (_08947_, _08900_, _04500_);
  or (_08948_, _08947_, _08946_);
  and (_08949_, _08948_, _03521_);
  and (_08950_, _08949_, _08945_);
  nor (_08951_, _06421_, _08901_);
  or (_08953_, _08951_, _08900_);
  and (_08954_, _08953_, _03224_);
  or (_08955_, _08954_, _08950_);
  or (_08956_, _08955_, _08905_);
  and (_08957_, _06436_, _05327_);
  or (_08958_, _08900_, _04527_);
  or (_08959_, _08958_, _08957_);
  and (_08960_, _06227_, _05327_);
  or (_08961_, _08960_, _08900_);
  or (_08962_, _08961_, _04509_);
  and (_08964_, _08962_, _03745_);
  and (_08965_, _08964_, _08959_);
  and (_08966_, _08965_, _08956_);
  and (_08967_, _06443_, _05327_);
  or (_08968_, _08967_, _08900_);
  and (_08969_, _08968_, _03744_);
  or (_08970_, _08969_, _08966_);
  and (_08971_, _08970_, _04523_);
  or (_08972_, _08900_, _05358_);
  and (_08973_, _08961_, _03611_);
  and (_08975_, _08973_, _08972_);
  or (_08976_, _08975_, _08971_);
  and (_08977_, _08976_, _03734_);
  and (_08978_, _08913_, _03733_);
  and (_08979_, _08978_, _08972_);
  or (_08980_, _08979_, _03618_);
  or (_08981_, _08980_, _08977_);
  nor (_08982_, _06434_, _08901_);
  or (_08983_, _08900_, _06453_);
  or (_08984_, _08983_, _08982_);
  and (_08986_, _08984_, _06458_);
  and (_08987_, _08986_, _08981_);
  or (_08988_, _08987_, _08904_);
  and (_08989_, _08988_, _03948_);
  and (_08990_, _08910_, _03767_);
  or (_08991_, _08990_, _03473_);
  or (_08992_, _08991_, _08989_);
  and (_08993_, _05886_, _05327_);
  or (_08994_, _08900_, _03474_);
  or (_08995_, _08994_, _08993_);
  and (_08997_, _08995_, _43189_);
  and (_08998_, _08997_, _08992_);
  or (_08999_, _08998_, _08899_);
  and (_40773_, _08999_, _42003_);
  not (_09000_, \oc8051_golden_model_1.DPH [7]);
  nor (_09001_, _43189_, _09000_);
  nor (_09002_, _05320_, _09000_);
  not (_09003_, _05320_);
  nor (_09004_, _06442_, _09003_);
  or (_09005_, _09004_, _09002_);
  and (_09007_, _09005_, _03741_);
  nor (_09008_, _09003_, _05253_);
  or (_09009_, _09008_, _09002_);
  or (_09010_, _09009_, _06903_);
  and (_09011_, _06133_, _05320_);
  or (_09012_, _09011_, _09002_);
  or (_09013_, _09012_, _04432_);
  and (_09014_, _05320_, \oc8051_golden_model_1.ACC [7]);
  or (_09015_, _09014_, _09002_);
  and (_09016_, _09015_, _04436_);
  nor (_09017_, _04436_, _09000_);
  or (_09018_, _09017_, _03534_);
  or (_09019_, _09018_, _09016_);
  and (_09020_, _09019_, _04457_);
  and (_09021_, _09020_, _09013_);
  and (_09022_, _09009_, _03527_);
  or (_09023_, _09022_, _03530_);
  or (_09024_, _09023_, _09021_);
  or (_09025_, _09015_, _03531_);
  and (_09026_, _09025_, _08924_);
  and (_09027_, _09026_, _09024_);
  and (_09028_, _08935_, \oc8051_golden_model_1.DPH [0]);
  and (_09029_, _09028_, \oc8051_golden_model_1.DPH [1]);
  and (_09030_, _09029_, \oc8051_golden_model_1.DPH [2]);
  and (_09031_, _09030_, \oc8051_golden_model_1.DPH [3]);
  and (_09032_, _09031_, \oc8051_golden_model_1.DPH [4]);
  and (_09033_, _09032_, \oc8051_golden_model_1.DPH [5]);
  nand (_09034_, _09033_, \oc8051_golden_model_1.DPH [6]);
  or (_09035_, _09034_, _09000_);
  nand (_09036_, _09034_, _09000_);
  and (_09037_, _09036_, _08923_);
  and (_09038_, _09037_, _09035_);
  or (_09039_, _09038_, _09027_);
  and (_09040_, _09039_, _03622_);
  and (_09041_, _03621_, _03409_);
  or (_09042_, _09041_, _07454_);
  or (_09043_, _09042_, _09040_);
  and (_09044_, _09043_, _09010_);
  or (_09045_, _09044_, _04082_);
  and (_09046_, _06114_, _05320_);
  or (_09047_, _09002_, _04500_);
  or (_09048_, _09047_, _09046_);
  and (_09049_, _09048_, _03521_);
  and (_09050_, _09049_, _09045_);
  nor (_09051_, _06421_, _09003_);
  or (_09052_, _09051_, _09002_);
  and (_09053_, _09052_, _03224_);
  or (_09054_, _09053_, _09050_);
  or (_09055_, _09054_, _08905_);
  and (_09056_, _06436_, _05320_);
  or (_09057_, _09002_, _04527_);
  or (_09058_, _09057_, _09056_);
  and (_09059_, _06227_, _05320_);
  or (_09060_, _09059_, _09002_);
  or (_09061_, _09060_, _04509_);
  and (_09062_, _09061_, _03745_);
  and (_09063_, _09062_, _09058_);
  and (_09064_, _09063_, _09055_);
  and (_09065_, _06443_, _05320_);
  or (_09066_, _09065_, _09002_);
  and (_09067_, _09066_, _03744_);
  or (_09068_, _09067_, _09064_);
  and (_09069_, _09068_, _04523_);
  or (_09070_, _09002_, _05358_);
  and (_09071_, _09060_, _03611_);
  and (_09072_, _09071_, _09070_);
  or (_09073_, _09072_, _09069_);
  and (_09074_, _09073_, _03734_);
  and (_09075_, _09015_, _03733_);
  and (_09076_, _09075_, _09070_);
  or (_09077_, _09076_, _03618_);
  or (_09078_, _09077_, _09074_);
  nor (_09079_, _06434_, _09003_);
  or (_09080_, _09002_, _06453_);
  or (_09081_, _09080_, _09079_);
  and (_09082_, _09081_, _06458_);
  and (_09083_, _09082_, _09078_);
  or (_09084_, _09083_, _09007_);
  and (_09085_, _09084_, _03948_);
  and (_09086_, _09012_, _03767_);
  or (_09087_, _09086_, _03473_);
  or (_09088_, _09087_, _09085_);
  and (_09089_, _05886_, _05320_);
  or (_09090_, _09002_, _03474_);
  or (_09091_, _09090_, _09089_);
  and (_09092_, _09091_, _43189_);
  and (_09093_, _09092_, _09088_);
  or (_09094_, _09093_, _09001_);
  and (_40774_, _09094_, _42003_);
  not (_09095_, \oc8051_golden_model_1.IE [7]);
  nor (_09096_, _05278_, _09095_);
  not (_09097_, _05278_);
  nor (_09098_, _09097_, _05253_);
  nor (_09099_, _09098_, _09096_);
  and (_09100_, _09099_, _07454_);
  nor (_09101_, _05944_, _09095_);
  and (_09102_, _05975_, _05944_);
  nor (_09103_, _09102_, _09101_);
  nor (_09104_, _09103_, _03466_);
  and (_09105_, _05278_, \oc8051_golden_model_1.ACC [7]);
  nor (_09106_, _09105_, _09096_);
  nor (_09107_, _09106_, _04437_);
  nor (_09108_, _04436_, _09095_);
  or (_09109_, _09108_, _09107_);
  and (_09110_, _09109_, _04432_);
  and (_09111_, _06133_, _05278_);
  nor (_09112_, _09111_, _09096_);
  nor (_09113_, _09112_, _04432_);
  or (_09114_, _09113_, _09110_);
  and (_09115_, _09114_, _03470_);
  and (_09116_, _05980_, _05944_);
  nor (_09117_, _09116_, _09101_);
  nor (_09118_, _09117_, _03470_);
  or (_09119_, _09118_, _03527_);
  or (_09120_, _09119_, _09115_);
  nand (_09121_, _09099_, _03527_);
  and (_09122_, _09121_, _09120_);
  and (_09123_, _09122_, _03531_);
  nor (_09124_, _09106_, _03531_);
  or (_09125_, _09124_, _09123_);
  and (_09126_, _09125_, _03466_);
  nor (_09127_, _09126_, _09104_);
  nor (_09128_, _09127_, _03458_);
  nor (_09129_, _09101_, _06165_);
  or (_09130_, _09117_, _03459_);
  nor (_09131_, _09130_, _09129_);
  nor (_09132_, _09131_, _09128_);
  nor (_09133_, _09132_, _03452_);
  not (_09134_, _05944_);
  nor (_09135_, _05962_, _09134_);
  nor (_09136_, _09135_, _09101_);
  nor (_09137_, _09136_, _03453_);
  nor (_09138_, _09137_, _07454_);
  not (_09139_, _09138_);
  nor (_09140_, _09139_, _09133_);
  nor (_09141_, _09140_, _09100_);
  nor (_09142_, _09141_, _04082_);
  and (_09143_, _06114_, _05278_);
  nor (_09144_, _09096_, _04500_);
  not (_09145_, _09144_);
  nor (_09146_, _09145_, _09143_);
  nor (_09147_, _09146_, _03224_);
  not (_09148_, _09147_);
  nor (_09149_, _09148_, _09142_);
  nor (_09150_, _06421_, _09097_);
  nor (_09151_, _09150_, _09096_);
  nor (_09152_, _09151_, _03521_);
  or (_09153_, _09152_, _08905_);
  or (_09154_, _09153_, _09149_);
  and (_09155_, _06436_, _05278_);
  or (_09156_, _09096_, _04527_);
  or (_09157_, _09156_, _09155_);
  and (_09158_, _06227_, _05278_);
  nor (_09159_, _09158_, _09096_);
  and (_09160_, _09159_, _03624_);
  nor (_09161_, _09160_, _03744_);
  and (_09162_, _09161_, _09157_);
  and (_09163_, _09162_, _09154_);
  and (_09164_, _06443_, _05278_);
  nor (_09165_, _09164_, _09096_);
  nor (_09166_, _09165_, _03745_);
  nor (_09167_, _09166_, _09163_);
  nor (_09168_, _09167_, _03611_);
  nor (_09169_, _09096_, _05358_);
  not (_09170_, _09169_);
  nor (_09171_, _09159_, _04523_);
  and (_09172_, _09171_, _09170_);
  nor (_09173_, _09172_, _09168_);
  nor (_09174_, _09173_, _03733_);
  nor (_09175_, _09106_, _03734_);
  and (_09176_, _09175_, _09170_);
  or (_09177_, _09176_, _09174_);
  and (_09178_, _09177_, _06453_);
  nor (_09179_, _06434_, _09097_);
  nor (_09180_, _09179_, _09096_);
  nor (_09181_, _09180_, _06453_);
  or (_09182_, _09181_, _09178_);
  and (_09183_, _09182_, _06458_);
  nor (_09184_, _06442_, _09097_);
  nor (_09185_, _09184_, _09096_);
  nor (_09186_, _09185_, _06458_);
  or (_09187_, _09186_, _09183_);
  and (_09188_, _09187_, _03948_);
  nor (_09189_, _09112_, _03948_);
  or (_09190_, _09189_, _09188_);
  and (_09191_, _09190_, _03446_);
  nor (_09192_, _09103_, _03446_);
  or (_09193_, _09192_, _09191_);
  and (_09194_, _09193_, _03474_);
  and (_09195_, _05886_, _05278_);
  nor (_09196_, _09195_, _09096_);
  nor (_09197_, _09196_, _03474_);
  or (_09198_, _09197_, _09194_);
  or (_09199_, _09198_, _43193_);
  or (_09200_, _43189_, \oc8051_golden_model_1.IE [7]);
  and (_09201_, _09200_, _42003_);
  and (_40775_, _09201_, _09199_);
  not (_09202_, \oc8051_golden_model_1.IP [7]);
  nor (_09203_, _05309_, _09202_);
  not (_09204_, _05309_);
  nor (_09205_, _09204_, _05253_);
  nor (_09206_, _09205_, _09203_);
  and (_09207_, _09206_, _07454_);
  nor (_09208_, _05935_, _09202_);
  and (_09209_, _05975_, _05935_);
  nor (_09210_, _09209_, _09208_);
  nor (_09211_, _09210_, _03466_);
  and (_09212_, _05309_, \oc8051_golden_model_1.ACC [7]);
  nor (_09213_, _09212_, _09203_);
  nor (_09214_, _09213_, _04437_);
  nor (_09215_, _04436_, _09202_);
  or (_09216_, _09215_, _09214_);
  and (_09217_, _09216_, _04432_);
  and (_09218_, _06133_, _05309_);
  nor (_09219_, _09218_, _09203_);
  nor (_09220_, _09219_, _04432_);
  or (_09221_, _09220_, _09217_);
  and (_09222_, _09221_, _03470_);
  and (_09223_, _05980_, _05935_);
  nor (_09224_, _09223_, _09208_);
  nor (_09225_, _09224_, _03470_);
  or (_09226_, _09225_, _03527_);
  or (_09227_, _09226_, _09222_);
  nand (_09228_, _09206_, _03527_);
  and (_09229_, _09228_, _09227_);
  and (_09230_, _09229_, _03531_);
  nor (_09231_, _09213_, _03531_);
  or (_09232_, _09231_, _09230_);
  and (_09233_, _09232_, _03466_);
  nor (_09234_, _09233_, _09211_);
  nor (_09235_, _09234_, _03458_);
  nor (_09236_, _09208_, _06165_);
  or (_09237_, _09224_, _03459_);
  nor (_09238_, _09237_, _09236_);
  nor (_09239_, _09238_, _09235_);
  nor (_09240_, _09239_, _03452_);
  not (_09241_, _05935_);
  nor (_09242_, _05962_, _09241_);
  nor (_09243_, _09242_, _09208_);
  nor (_09244_, _09243_, _03453_);
  nor (_09245_, _09244_, _07454_);
  not (_09246_, _09245_);
  nor (_09247_, _09246_, _09240_);
  nor (_09248_, _09247_, _09207_);
  nor (_09249_, _09248_, _04082_);
  and (_09250_, _06114_, _05309_);
  nor (_09251_, _09203_, _04500_);
  not (_09252_, _09251_);
  nor (_09253_, _09252_, _09250_);
  nor (_09254_, _09253_, _03224_);
  not (_09255_, _09254_);
  nor (_09256_, _09255_, _09249_);
  nor (_09257_, _06421_, _09204_);
  nor (_09258_, _09257_, _09203_);
  nor (_09259_, _09258_, _03521_);
  or (_09260_, _09259_, _08905_);
  or (_09261_, _09260_, _09256_);
  and (_09262_, _06436_, _05309_);
  or (_09263_, _09203_, _04527_);
  or (_09264_, _09263_, _09262_);
  and (_09265_, _06227_, _05309_);
  nor (_09266_, _09265_, _09203_);
  and (_09267_, _09266_, _03624_);
  nor (_09268_, _09267_, _03744_);
  and (_09269_, _09268_, _09264_);
  and (_09270_, _09269_, _09261_);
  and (_09271_, _06443_, _05309_);
  nor (_09272_, _09271_, _09203_);
  nor (_09273_, _09272_, _03745_);
  nor (_09274_, _09273_, _09270_);
  nor (_09275_, _09274_, _03611_);
  nor (_09276_, _09203_, _05358_);
  not (_09277_, _09276_);
  nor (_09278_, _09266_, _04523_);
  and (_09279_, _09278_, _09277_);
  nor (_09280_, _09279_, _09275_);
  nor (_09281_, _09280_, _03733_);
  nor (_09282_, _09213_, _03734_);
  and (_09283_, _09282_, _09277_);
  or (_09284_, _09283_, _09281_);
  and (_09285_, _09284_, _06453_);
  nor (_09286_, _06434_, _09204_);
  nor (_09287_, _09286_, _09203_);
  nor (_09288_, _09287_, _06453_);
  or (_09289_, _09288_, _09285_);
  and (_09290_, _09289_, _06458_);
  nor (_09291_, _06442_, _09204_);
  nor (_09292_, _09291_, _09203_);
  nor (_09293_, _09292_, _06458_);
  or (_09294_, _09293_, _09290_);
  and (_09295_, _09294_, _03948_);
  nor (_09296_, _09219_, _03948_);
  or (_09297_, _09296_, _09295_);
  and (_09298_, _09297_, _03446_);
  nor (_09299_, _09210_, _03446_);
  or (_09300_, _09299_, _09298_);
  and (_09301_, _09300_, _03474_);
  and (_09302_, _05886_, _05309_);
  nor (_09303_, _09302_, _09203_);
  nor (_09304_, _09303_, _03474_);
  or (_09305_, _09304_, _09301_);
  or (_09306_, _09305_, _43193_);
  or (_09307_, _43189_, \oc8051_golden_model_1.IP [7]);
  and (_09308_, _09307_, _42003_);
  and (_40776_, _09308_, _09306_);
  not (_09309_, \oc8051_golden_model_1.P0 [7]);
  nor (_09310_, _05298_, _09309_);
  not (_09311_, _05298_);
  nor (_09312_, _09311_, _05253_);
  or (_09313_, _09312_, _09310_);
  or (_09314_, _09313_, _06903_);
  nor (_09315_, _05258_, _09309_);
  and (_09316_, _05975_, _05258_);
  or (_09317_, _09316_, _09315_);
  and (_09318_, _09317_, _03465_);
  and (_09319_, _06133_, _05298_);
  or (_09320_, _09319_, _09310_);
  or (_09321_, _09320_, _04432_);
  and (_09322_, _05298_, \oc8051_golden_model_1.ACC [7]);
  or (_09323_, _09322_, _09310_);
  and (_09324_, _09323_, _04436_);
  nor (_09325_, _04436_, _09309_);
  or (_09326_, _09325_, _03534_);
  or (_09327_, _09326_, _09324_);
  and (_09328_, _09327_, _03470_);
  and (_09329_, _09328_, _09321_);
  and (_09330_, _05980_, _05258_);
  or (_09331_, _09330_, _09315_);
  and (_09332_, _09331_, _03469_);
  or (_09333_, _09332_, _03527_);
  or (_09334_, _09333_, _09329_);
  or (_09335_, _09313_, _04457_);
  and (_09336_, _09335_, _09334_);
  or (_09337_, _09336_, _03530_);
  or (_09338_, _09323_, _03531_);
  and (_09339_, _09338_, _03466_);
  and (_09340_, _09339_, _09337_);
  or (_09341_, _09340_, _09318_);
  and (_09342_, _09341_, _03459_);
  or (_09343_, _09315_, _06165_);
  and (_09344_, _09343_, _03458_);
  and (_09345_, _09344_, _09331_);
  or (_09346_, _09345_, _09342_);
  and (_09347_, _09346_, _03453_);
  or (_09348_, _05975_, _05961_);
  and (_09349_, _09348_, _05258_);
  or (_09350_, _09349_, _09315_);
  and (_09351_, _09350_, _03452_);
  or (_09352_, _09351_, _07454_);
  or (_09353_, _09352_, _09347_);
  and (_09354_, _09353_, _09314_);
  or (_09355_, _09354_, _04082_);
  and (_09356_, _06114_, _05298_);
  or (_09357_, _09310_, _04500_);
  or (_09358_, _09357_, _09356_);
  and (_09359_, _09358_, _03521_);
  and (_09360_, _09359_, _09355_);
  and (_09361_, _06334_, \oc8051_golden_model_1.P0 [7]);
  and (_09362_, _06329_, \oc8051_golden_model_1.P2 [7]);
  and (_09363_, _06340_, \oc8051_golden_model_1.P1 [7]);
  and (_09364_, _06344_, \oc8051_golden_model_1.P3 [7]);
  or (_09365_, _09364_, _09363_);
  or (_09366_, _09365_, _09362_);
  nor (_09367_, _09366_, _09361_);
  and (_09368_, _09367_, _06361_);
  and (_09369_, _09368_, _06388_);
  nand (_09370_, _09369_, _06418_);
  or (_09371_, _09370_, _06228_);
  and (_09372_, _09371_, _05298_);
  or (_09373_, _09372_, _09310_);
  and (_09374_, _09373_, _03224_);
  or (_09375_, _09374_, _08905_);
  or (_09376_, _09375_, _09360_);
  and (_09377_, _06436_, _05298_);
  or (_09378_, _09310_, _04527_);
  or (_09379_, _09378_, _09377_);
  and (_09380_, _06227_, _05298_);
  or (_09381_, _09380_, _09310_);
  or (_09382_, _09381_, _04509_);
  and (_09383_, _09382_, _03745_);
  and (_09384_, _09383_, _09379_);
  and (_09385_, _09384_, _09376_);
  and (_09386_, _06443_, _05298_);
  or (_09387_, _09386_, _09310_);
  and (_09388_, _09387_, _03744_);
  or (_09389_, _09388_, _09385_);
  and (_09390_, _09389_, _04523_);
  or (_09391_, _09310_, _05358_);
  and (_09392_, _09381_, _03611_);
  and (_09393_, _09392_, _09391_);
  or (_09394_, _09393_, _09390_);
  and (_09395_, _09394_, _03734_);
  and (_09396_, _09323_, _03733_);
  and (_09397_, _09396_, _09391_);
  or (_09398_, _09397_, _03618_);
  or (_09399_, _09398_, _09395_);
  nor (_09400_, _06434_, _09311_);
  or (_09401_, _09310_, _06453_);
  or (_09402_, _09401_, _09400_);
  and (_09403_, _09402_, _06458_);
  and (_09404_, _09403_, _09399_);
  nor (_09405_, _06442_, _09311_);
  or (_09406_, _09405_, _09310_);
  and (_09407_, _09406_, _03741_);
  or (_09408_, _09407_, _03767_);
  or (_09409_, _09408_, _09404_);
  or (_09410_, _09320_, _03948_);
  and (_09411_, _09410_, _03446_);
  and (_09412_, _09411_, _09409_);
  and (_09413_, _09317_, _03445_);
  or (_09414_, _09413_, _03473_);
  or (_09415_, _09414_, _09412_);
  and (_09416_, _05886_, _05298_);
  or (_09417_, _09310_, _03474_);
  or (_09418_, _09417_, _09416_);
  and (_09419_, _09418_, _43189_);
  and (_09420_, _09419_, _09415_);
  nor (_09421_, _43189_, _09309_);
  or (_09422_, _09421_, rst);
  or (_40778_, _09422_, _09420_);
  not (_09423_, \oc8051_golden_model_1.P1 [7]);
  nor (_09424_, _43189_, _09423_);
  or (_09425_, _09424_, rst);
  nor (_09426_, _05284_, _09423_);
  not (_09427_, _05284_);
  nor (_09428_, _09427_, _05253_);
  or (_09429_, _09428_, _09426_);
  or (_09430_, _09429_, _06903_);
  nor (_09431_, _05951_, _09423_);
  and (_09432_, _05975_, _05951_);
  or (_09433_, _09432_, _09431_);
  and (_09434_, _09433_, _03465_);
  and (_09435_, _06133_, _05284_);
  or (_09436_, _09435_, _09426_);
  or (_09437_, _09436_, _04432_);
  and (_09438_, _05284_, \oc8051_golden_model_1.ACC [7]);
  or (_09439_, _09438_, _09426_);
  and (_09440_, _09439_, _04436_);
  nor (_09441_, _04436_, _09423_);
  or (_09442_, _09441_, _03534_);
  or (_09443_, _09442_, _09440_);
  and (_09444_, _09443_, _03470_);
  and (_09445_, _09444_, _09437_);
  and (_09446_, _05980_, _05951_);
  or (_09447_, _09446_, _09431_);
  and (_09448_, _09447_, _03469_);
  or (_09449_, _09448_, _03527_);
  or (_09450_, _09449_, _09445_);
  or (_09451_, _09429_, _04457_);
  and (_09452_, _09451_, _09450_);
  or (_09453_, _09452_, _03530_);
  or (_09454_, _09439_, _03531_);
  and (_09455_, _09454_, _03466_);
  and (_09456_, _09455_, _09453_);
  or (_09457_, _09456_, _09434_);
  and (_09458_, _09457_, _03459_);
  and (_09459_, _06166_, _05951_);
  or (_09460_, _09459_, _09431_);
  and (_09461_, _09460_, _03458_);
  or (_09462_, _09461_, _09458_);
  and (_09463_, _09462_, _03453_);
  and (_09464_, _09348_, _05951_);
  or (_09465_, _09464_, _09431_);
  and (_09466_, _09465_, _03452_);
  or (_09467_, _09466_, _07454_);
  or (_09468_, _09467_, _09463_);
  and (_09469_, _09468_, _09430_);
  or (_09470_, _09469_, _04082_);
  and (_09471_, _06114_, _05284_);
  or (_09472_, _09426_, _04500_);
  or (_09473_, _09472_, _09471_);
  and (_09474_, _09473_, _03521_);
  and (_09475_, _09474_, _09470_);
  and (_09476_, _09371_, _05284_);
  or (_09477_, _09476_, _09426_);
  and (_09478_, _09477_, _03224_);
  or (_09479_, _09478_, _08905_);
  or (_09480_, _09479_, _09475_);
  and (_09481_, _06436_, _05284_);
  or (_09482_, _09426_, _04527_);
  or (_09483_, _09482_, _09481_);
  and (_09484_, _06227_, _05284_);
  or (_09485_, _09484_, _09426_);
  or (_09486_, _09485_, _04509_);
  and (_09487_, _09486_, _03745_);
  and (_09488_, _09487_, _09483_);
  and (_09489_, _09488_, _09480_);
  and (_09490_, _06443_, _05284_);
  or (_09491_, _09490_, _09426_);
  and (_09492_, _09491_, _03744_);
  or (_09493_, _09492_, _09489_);
  and (_09494_, _09493_, _04523_);
  or (_09495_, _09426_, _05358_);
  and (_09496_, _09485_, _03611_);
  and (_09497_, _09496_, _09495_);
  or (_09498_, _09497_, _09494_);
  and (_09499_, _09498_, _03734_);
  and (_09500_, _09439_, _03733_);
  and (_09501_, _09500_, _09495_);
  or (_09502_, _09501_, _03618_);
  or (_09503_, _09502_, _09499_);
  nor (_09504_, _06434_, _09427_);
  or (_09505_, _09426_, _06453_);
  or (_09506_, _09505_, _09504_);
  and (_09507_, _09506_, _06458_);
  and (_09508_, _09507_, _09503_);
  nor (_09509_, _06442_, _09427_);
  or (_09510_, _09509_, _09426_);
  and (_09511_, _09510_, _03741_);
  or (_09512_, _09511_, _03767_);
  or (_09513_, _09512_, _09508_);
  or (_09514_, _09436_, _03948_);
  and (_09515_, _09514_, _03446_);
  and (_09516_, _09515_, _09513_);
  and (_09517_, _09433_, _03445_);
  or (_09518_, _09517_, _03473_);
  or (_09519_, _09518_, _09516_);
  and (_09520_, _05886_, _05284_);
  or (_09521_, _09426_, _03474_);
  or (_09522_, _09521_, _09520_);
  and (_09523_, _09522_, _43189_);
  and (_09524_, _09523_, _09519_);
  or (_40779_, _09524_, _09425_);
  not (_09525_, \oc8051_golden_model_1.P2 [7]);
  nor (_09526_, _43189_, _09525_);
  or (_09527_, _09526_, rst);
  nor (_09528_, _05289_, _09525_);
  not (_09529_, _05289_);
  nor (_09530_, _09529_, _05253_);
  or (_09531_, _09530_, _09528_);
  or (_09532_, _09531_, _06903_);
  nor (_09533_, _05948_, _09525_);
  and (_09534_, _05975_, _05948_);
  or (_09535_, _09534_, _09533_);
  and (_09536_, _09535_, _03465_);
  and (_09537_, _06133_, _05289_);
  or (_09538_, _09537_, _09528_);
  or (_09539_, _09538_, _04432_);
  and (_09540_, _05289_, \oc8051_golden_model_1.ACC [7]);
  or (_09541_, _09540_, _09528_);
  and (_09542_, _09541_, _04436_);
  nor (_09543_, _04436_, _09525_);
  or (_09544_, _09543_, _03534_);
  or (_09545_, _09544_, _09542_);
  and (_09546_, _09545_, _03470_);
  and (_09547_, _09546_, _09539_);
  and (_09548_, _05980_, _05948_);
  or (_09549_, _09548_, _09533_);
  and (_09550_, _09549_, _03469_);
  or (_09551_, _09550_, _03527_);
  or (_09553_, _09551_, _09547_);
  or (_09554_, _09531_, _04457_);
  and (_09555_, _09554_, _09553_);
  or (_09556_, _09555_, _03530_);
  or (_09557_, _09541_, _03531_);
  and (_09558_, _09557_, _03466_);
  and (_09559_, _09558_, _09556_);
  or (_09560_, _09559_, _09536_);
  and (_09561_, _09560_, _03459_);
  and (_09562_, _06166_, _05948_);
  or (_09563_, _09562_, _09533_);
  and (_09564_, _09563_, _03458_);
  or (_09565_, _09564_, _09561_);
  and (_09566_, _09565_, _03453_);
  and (_09567_, _09348_, _05948_);
  or (_09568_, _09567_, _09533_);
  and (_09569_, _09568_, _03452_);
  or (_09570_, _09569_, _07454_);
  or (_09571_, _09570_, _09566_);
  and (_09572_, _09571_, _09532_);
  or (_09574_, _09572_, _04082_);
  and (_09575_, _06114_, _05289_);
  or (_09576_, _09528_, _04500_);
  or (_09577_, _09576_, _09575_);
  and (_09578_, _09577_, _03521_);
  and (_09579_, _09578_, _09574_);
  and (_09580_, _09371_, _05289_);
  or (_09581_, _09580_, _09528_);
  and (_09582_, _09581_, _03224_);
  or (_09583_, _09582_, _08905_);
  or (_09584_, _09583_, _09579_);
  and (_09585_, _06436_, _05289_);
  or (_09586_, _09528_, _04527_);
  or (_09587_, _09586_, _09585_);
  and (_09588_, _06227_, _05289_);
  or (_09589_, _09588_, _09528_);
  or (_09590_, _09589_, _04509_);
  and (_09591_, _09590_, _03745_);
  and (_09592_, _09591_, _09587_);
  and (_09593_, _09592_, _09584_);
  and (_09594_, _06443_, _05289_);
  or (_09595_, _09594_, _09528_);
  and (_09596_, _09595_, _03744_);
  or (_09597_, _09596_, _09593_);
  and (_09598_, _09597_, _04523_);
  or (_09599_, _09528_, _05358_);
  and (_09600_, _09589_, _03611_);
  and (_09601_, _09600_, _09599_);
  or (_09602_, _09601_, _09598_);
  and (_09603_, _09602_, _03734_);
  and (_09604_, _09541_, _03733_);
  and (_09605_, _09604_, _09599_);
  or (_09606_, _09605_, _03618_);
  or (_09607_, _09606_, _09603_);
  nor (_09608_, _06434_, _09529_);
  or (_09609_, _09528_, _06453_);
  or (_09610_, _09609_, _09608_);
  and (_09611_, _09610_, _06458_);
  and (_09612_, _09611_, _09607_);
  nor (_09613_, _06442_, _09529_);
  or (_09614_, _09613_, _09528_);
  and (_09615_, _09614_, _03741_);
  or (_09616_, _09615_, _03767_);
  or (_09617_, _09616_, _09612_);
  or (_09618_, _09538_, _03948_);
  and (_09619_, _09618_, _03446_);
  and (_09620_, _09619_, _09617_);
  and (_09621_, _09535_, _03445_);
  or (_09622_, _09621_, _03473_);
  or (_09623_, _09622_, _09620_);
  and (_09624_, _05886_, _05289_);
  or (_09625_, _09528_, _03474_);
  or (_09626_, _09625_, _09624_);
  and (_09627_, _09626_, _43189_);
  and (_09628_, _09627_, _09623_);
  or (_40780_, _09628_, _09527_);
  not (_09629_, \oc8051_golden_model_1.P3 [7]);
  nor (_09630_, _43189_, _09629_);
  or (_09631_, _09630_, rst);
  nor (_09632_, _05293_, _09629_);
  not (_09633_, _05293_);
  nor (_09634_, _09633_, _05253_);
  or (_09635_, _09634_, _09632_);
  or (_09636_, _09635_, _06903_);
  nor (_09637_, _05953_, _09629_);
  and (_09638_, _05975_, _05953_);
  or (_09639_, _09638_, _09637_);
  and (_09640_, _09639_, _03465_);
  and (_09641_, _06133_, _05293_);
  or (_09642_, _09641_, _09632_);
  or (_09643_, _09642_, _04432_);
  and (_09644_, _05293_, \oc8051_golden_model_1.ACC [7]);
  or (_09645_, _09644_, _09632_);
  and (_09646_, _09645_, _04436_);
  nor (_09647_, _04436_, _09629_);
  or (_09648_, _09647_, _03534_);
  or (_09649_, _09648_, _09646_);
  and (_09650_, _09649_, _03470_);
  and (_09651_, _09650_, _09643_);
  and (_09652_, _05980_, _05953_);
  or (_09653_, _09652_, _09637_);
  and (_09654_, _09653_, _03469_);
  or (_09655_, _09654_, _03527_);
  or (_09656_, _09655_, _09651_);
  or (_09657_, _09635_, _04457_);
  and (_09658_, _09657_, _09656_);
  or (_09659_, _09658_, _03530_);
  or (_09660_, _09645_, _03531_);
  and (_09661_, _09660_, _03466_);
  and (_09662_, _09661_, _09659_);
  or (_09663_, _09662_, _09640_);
  and (_09664_, _09663_, _03459_);
  and (_09665_, _06166_, _05953_);
  or (_09666_, _09665_, _09637_);
  and (_09667_, _09666_, _03458_);
  or (_09668_, _09667_, _09664_);
  and (_09669_, _09668_, _03453_);
  and (_09670_, _09348_, _05953_);
  or (_09671_, _09670_, _09637_);
  and (_09672_, _09671_, _03452_);
  or (_09673_, _09672_, _07454_);
  or (_09674_, _09673_, _09669_);
  and (_09675_, _09674_, _09636_);
  or (_09676_, _09675_, _04082_);
  and (_09677_, _06114_, _05293_);
  or (_09678_, _09632_, _04500_);
  or (_09679_, _09678_, _09677_);
  and (_09680_, _09679_, _03521_);
  and (_09681_, _09680_, _09676_);
  and (_09682_, _09371_, _05293_);
  or (_09683_, _09682_, _09632_);
  and (_09684_, _09683_, _03224_);
  or (_09685_, _09684_, _08905_);
  or (_09686_, _09685_, _09681_);
  and (_09687_, _06436_, _05293_);
  or (_09688_, _09632_, _04527_);
  or (_09689_, _09688_, _09687_);
  and (_09690_, _06227_, _05293_);
  or (_09691_, _09690_, _09632_);
  or (_09692_, _09691_, _04509_);
  and (_09693_, _09692_, _03745_);
  and (_09694_, _09693_, _09689_);
  and (_09695_, _09694_, _09686_);
  and (_09696_, _06443_, _05293_);
  or (_09697_, _09696_, _09632_);
  and (_09698_, _09697_, _03744_);
  or (_09699_, _09698_, _09695_);
  and (_09700_, _09699_, _04523_);
  or (_09701_, _09632_, _05358_);
  and (_09702_, _09691_, _03611_);
  and (_09703_, _09702_, _09701_);
  or (_09704_, _09703_, _09700_);
  and (_09705_, _09704_, _03734_);
  and (_09706_, _09645_, _03733_);
  and (_09707_, _09706_, _09701_);
  or (_09708_, _09707_, _03618_);
  or (_09709_, _09708_, _09705_);
  nor (_09710_, _06434_, _09633_);
  or (_09711_, _09632_, _06453_);
  or (_09712_, _09711_, _09710_);
  and (_09713_, _09712_, _06458_);
  and (_09714_, _09713_, _09709_);
  nor (_09715_, _06442_, _09633_);
  or (_09716_, _09715_, _09632_);
  and (_09717_, _09716_, _03741_);
  or (_09718_, _09717_, _03767_);
  or (_09719_, _09718_, _09714_);
  or (_09720_, _09642_, _03948_);
  and (_09721_, _09720_, _03446_);
  and (_09722_, _09721_, _09719_);
  and (_09723_, _09639_, _03445_);
  or (_09724_, _09723_, _03473_);
  or (_09725_, _09724_, _09722_);
  and (_09726_, _05886_, _05293_);
  or (_09727_, _09632_, _03474_);
  or (_09728_, _09727_, _09726_);
  and (_09729_, _09728_, _43189_);
  and (_09730_, _09729_, _09725_);
  or (_40781_, _09730_, _09631_);
  not (_09731_, _07931_);
  nor (_09732_, _08843_, _07932_);
  nor (_09733_, _09732_, _08786_);
  nand (_09734_, _09733_, _09731_);
  nor (_09735_, _07948_, _06440_);
  or (_09736_, _09735_, _08731_);
  and (_09737_, _07958_, _05275_);
  and (_09738_, _09737_, _05301_);
  or (_09739_, _09738_, _09736_);
  and (_09740_, _09739_, _08627_);
  nor (_09741_, _08028_, _06440_);
  nor (_09742_, _09741_, _08621_);
  and (_09743_, _08039_, _06757_);
  nand (_09744_, _09743_, _06526_);
  or (_09745_, _09744_, _06481_);
  and (_09746_, _09745_, _08595_);
  and (_09747_, _09746_, _09742_);
  nor (_09748_, _05303_, _07982_);
  not (_09749_, _09748_);
  nand (_09750_, _06443_, _05303_);
  and (_09751_, _09750_, _09749_);
  or (_09752_, _09751_, _03745_);
  not (_09753_, _05303_);
  or (_09754_, _06421_, _09753_);
  and (_09755_, _09754_, _09749_);
  or (_09756_, _09755_, _03521_);
  or (_09757_, _09753_, _05253_);
  and (_09758_, _09757_, _09749_);
  and (_09759_, _09758_, _07454_);
  and (_09760_, _08035_, _08031_);
  nor (_09761_, _09760_, _08029_);
  not (_09762_, _09761_);
  and (_09763_, _08601_, _08031_);
  not (_09764_, _09763_);
  nor (_09765_, _09764_, _08090_);
  nor (_09766_, _09765_, _09762_);
  nand (_09767_, _09745_, _04066_);
  nor (_09768_, _09767_, _09766_);
  not (_09769_, _03587_);
  not (_09770_, _05326_);
  and (_09771_, _05942_, \oc8051_golden_model_1.SCON [2]);
  and (_09772_, _05944_, \oc8051_golden_model_1.IE [2]);
  nor (_09773_, _09772_, _09771_);
  and (_09774_, _05924_, \oc8051_golden_model_1.TCON [2]);
  and (_09775_, _05953_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_09776_, _09775_, _09774_);
  and (_09777_, _09776_, _09773_);
  and (_09778_, _05932_, \oc8051_golden_model_1.PSW [2]);
  and (_09779_, _05937_, \oc8051_golden_model_1.ACC [2]);
  nor (_09780_, _09779_, _09778_);
  and (_09781_, _05935_, \oc8051_golden_model_1.IP [2]);
  and (_09782_, _05929_, \oc8051_golden_model_1.B [2]);
  nor (_09783_, _09782_, _09781_);
  and (_09784_, _09783_, _09780_);
  and (_09785_, _05951_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09786_, _05948_, \oc8051_golden_model_1.P2INREG [2]);
  and (_09787_, _05258_, \oc8051_golden_model_1.P0INREG [2]);
  or (_09788_, _09787_, _09786_);
  nor (_09789_, _09788_, _09785_);
  and (_09790_, _09789_, _09784_);
  and (_09791_, _09790_, _09777_);
  and (_09792_, _09791_, _05724_);
  nor (_09793_, _09792_, _09770_);
  not (_09794_, _05265_);
  and (_09795_, _05924_, \oc8051_golden_model_1.TCON [1]);
  and (_09796_, _05929_, \oc8051_golden_model_1.B [1]);
  nor (_09797_, _09796_, _09795_);
  and (_09798_, _05932_, \oc8051_golden_model_1.PSW [1]);
  not (_09799_, _09798_);
  and (_09800_, _05935_, \oc8051_golden_model_1.IP [1]);
  and (_09801_, _05937_, \oc8051_golden_model_1.ACC [1]);
  nor (_09802_, _09801_, _09800_);
  and (_09803_, _09802_, _09799_);
  and (_09804_, _09803_, _09797_);
  and (_09805_, _05942_, \oc8051_golden_model_1.SCON [1]);
  and (_09806_, _05944_, \oc8051_golden_model_1.IE [1]);
  nor (_09807_, _09806_, _09805_);
  and (_09808_, _05258_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09809_, _05948_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09810_, _09809_, _09808_);
  and (_09811_, _05951_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09812_, _05953_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09813_, _09812_, _09811_);
  and (_09814_, _09813_, _09810_);
  and (_09815_, _09814_, _09807_);
  and (_09816_, _09815_, _09804_);
  and (_09817_, _09816_, _05626_);
  nor (_09818_, _09817_, _09794_);
  nor (_09819_, _09818_, _09793_);
  and (_09820_, _05272_, _05005_);
  not (_09821_, _09820_);
  and (_09822_, _05924_, \oc8051_golden_model_1.TCON [4]);
  and (_09823_, _05929_, \oc8051_golden_model_1.B [4]);
  nor (_09824_, _09823_, _09822_);
  and (_09825_, _05932_, \oc8051_golden_model_1.PSW [4]);
  not (_09826_, _09825_);
  and (_09827_, _05935_, \oc8051_golden_model_1.IP [4]);
  and (_09828_, _05937_, \oc8051_golden_model_1.ACC [4]);
  nor (_09829_, _09828_, _09827_);
  and (_09830_, _09829_, _09826_);
  and (_09831_, _09830_, _09824_);
  and (_09832_, _05942_, \oc8051_golden_model_1.SCON [4]);
  and (_09833_, _05944_, \oc8051_golden_model_1.IE [4]);
  nor (_09834_, _09833_, _09832_);
  and (_09835_, _05258_, \oc8051_golden_model_1.P0INREG [4]);
  and (_09836_, _05948_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_09837_, _09836_, _09835_);
  and (_09838_, _05951_, \oc8051_golden_model_1.P1INREG [4]);
  and (_09839_, _05953_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09840_, _09839_, _09838_);
  and (_09841_, _09840_, _09837_);
  and (_09842_, _09841_, _09834_);
  and (_09843_, _09842_, _09831_);
  and (_09844_, _09843_, _05832_);
  nor (_09845_, _09844_, _09821_);
  nor (_09846_, _05959_, _05979_);
  nor (_09847_, _09846_, _09845_);
  and (_09848_, _09847_, _09819_);
  not (_09849_, _05273_);
  and (_09850_, _05942_, \oc8051_golden_model_1.SCON [0]);
  not (_09851_, _09850_);
  and (_09852_, _05944_, \oc8051_golden_model_1.IE [0]);
  and (_09853_, _05937_, \oc8051_golden_model_1.ACC [0]);
  nor (_09854_, _09853_, _09852_);
  and (_09855_, _09854_, _09851_);
  and (_09856_, _05932_, \oc8051_golden_model_1.PSW [0]);
  and (_09857_, _05929_, \oc8051_golden_model_1.B [0]);
  nor (_09858_, _09857_, _09856_);
  and (_09859_, _05924_, \oc8051_golden_model_1.TCON [0]);
  and (_09860_, _05935_, \oc8051_golden_model_1.IP [0]);
  nor (_09861_, _09860_, _09859_);
  and (_09862_, _09861_, _09858_);
  and (_09863_, _09862_, _09855_);
  and (_09864_, _05258_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09865_, _05948_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09866_, _09865_, _09864_);
  and (_09867_, _05951_, \oc8051_golden_model_1.P1INREG [0]);
  and (_09868_, _05953_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09869_, _09868_, _09867_);
  and (_09870_, _09869_, _09866_);
  and (_09871_, _09870_, _09863_);
  and (_09872_, _09871_, _05675_);
  nor (_09873_, _09872_, _09849_);
  and (_09874_, _05325_, _05005_);
  not (_09875_, _09874_);
  and (_09876_, _05935_, \oc8051_golden_model_1.IP [6]);
  and (_09877_, _05929_, \oc8051_golden_model_1.B [6]);
  nor (_09878_, _09877_, _09876_);
  and (_09879_, _05942_, \oc8051_golden_model_1.SCON [6]);
  and (_09880_, _05944_, \oc8051_golden_model_1.IE [6]);
  nor (_09881_, _09880_, _09879_);
  and (_09882_, _05932_, \oc8051_golden_model_1.PSW [6]);
  and (_09883_, _05937_, \oc8051_golden_model_1.ACC [6]);
  nor (_09884_, _09883_, _09882_);
  and (_09885_, _09884_, _09881_);
  and (_09886_, _09885_, _09878_);
  and (_09887_, _05924_, \oc8051_golden_model_1.TCON [6]);
  and (_09888_, _05953_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09889_, _09888_, _09887_);
  and (_09890_, _05951_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09891_, _05948_, \oc8051_golden_model_1.P2INREG [6]);
  and (_09892_, _05258_, \oc8051_golden_model_1.P0INREG [6]);
  or (_09893_, _09892_, _09891_);
  nor (_09894_, _09893_, _09890_);
  and (_09895_, _09894_, _09889_);
  and (_09896_, _09895_, _09886_);
  and (_09897_, _09896_, _05418_);
  nor (_09898_, _09897_, _09875_);
  nor (_09899_, _09898_, _09873_);
  not (_09900_, _05319_);
  and (_09901_, _05924_, \oc8051_golden_model_1.TCON [3]);
  and (_09902_, _05937_, \oc8051_golden_model_1.ACC [3]);
  nor (_09903_, _09902_, _09901_);
  and (_09904_, _05935_, \oc8051_golden_model_1.IP [3]);
  not (_09905_, _09904_);
  and (_09906_, _05932_, \oc8051_golden_model_1.PSW [3]);
  and (_09907_, _05929_, \oc8051_golden_model_1.B [3]);
  nor (_09908_, _09907_, _09906_);
  and (_09909_, _09908_, _09905_);
  and (_09910_, _09909_, _09903_);
  and (_09911_, _05942_, \oc8051_golden_model_1.SCON [3]);
  and (_09912_, _05944_, \oc8051_golden_model_1.IE [3]);
  nor (_09913_, _09912_, _09911_);
  and (_09914_, _05258_, \oc8051_golden_model_1.P0INREG [3]);
  and (_09915_, _05948_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09916_, _09915_, _09914_);
  and (_09917_, _05951_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09918_, _05953_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_09919_, _09918_, _09917_);
  and (_09920_, _09919_, _09916_);
  and (_09921_, _09920_, _09913_);
  and (_09922_, _09921_, _09910_);
  and (_09923_, _09922_, _05577_);
  nor (_09924_, _09923_, _09900_);
  and (_09925_, _05264_, _05005_);
  not (_09926_, _09925_);
  and (_09927_, _05935_, \oc8051_golden_model_1.IP [5]);
  and (_09928_, _05929_, \oc8051_golden_model_1.B [5]);
  nor (_09929_, _09928_, _09927_);
  and (_09930_, _05932_, \oc8051_golden_model_1.PSW [5]);
  and (_09931_, _05937_, \oc8051_golden_model_1.ACC [5]);
  nor (_09932_, _09931_, _09930_);
  and (_09933_, _09932_, _09929_);
  and (_09934_, _05944_, \oc8051_golden_model_1.IE [5]);
  not (_09935_, _09934_);
  and (_09936_, _05924_, \oc8051_golden_model_1.TCON [5]);
  and (_09937_, _05942_, \oc8051_golden_model_1.SCON [5]);
  nor (_09938_, _09937_, _09936_);
  and (_09939_, _09938_, _09935_);
  and (_09940_, _05258_, \oc8051_golden_model_1.P0INREG [5]);
  and (_09941_, _05953_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09942_, _09941_, _09940_);
  and (_09943_, _05951_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09944_, _05948_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_09945_, _09944_, _09943_);
  and (_09946_, _09945_, _09942_);
  and (_09947_, _09946_, _09939_);
  and (_09948_, _09947_, _09933_);
  and (_09949_, _09948_, _05527_);
  nor (_09950_, _09949_, _09926_);
  nor (_09951_, _09950_, _09924_);
  and (_09952_, _09951_, _09899_);
  and (_09953_, _09952_, _09848_);
  or (_09954_, _09953_, _09769_);
  not (_09955_, _08413_);
  nor (_09956_, _08414_, _09955_);
  or (_09957_, _09956_, _08366_);
  nand (_09958_, _09957_, _08412_);
  and (_09959_, _08411_, _08384_);
  nor (_09960_, _09959_, _08336_);
  nand (_09961_, _09960_, _09958_);
  and (_09962_, _08404_, _08391_);
  not (_09963_, _08270_);
  and (_09964_, _08290_, _09963_);
  and (_09965_, _09964_, _09962_);
  nand (_09966_, _09965_, _09961_);
  nor (_09967_, _08390_, _08307_);
  nor (_09968_, _09967_, _08306_);
  nand (_09969_, _09964_, _09968_);
  or (_09970_, _06160_, \oc8051_golden_model_1.ACC [7]);
  nand (_09971_, _08289_, _09963_);
  and (_09972_, _09971_, _09970_);
  and (_09973_, _09972_, _09969_);
  and (_09974_, _09973_, _09966_);
  and (_09975_, _09965_, _08417_);
  or (_09976_, _09975_, _03994_);
  or (_09977_, _09976_, _09974_);
  and (_09978_, _06133_, _05303_);
  nor (_09979_, _09978_, _09748_);
  and (_09980_, _09979_, _03534_);
  and (_09981_, _05303_, \oc8051_golden_model_1.ACC [7]);
  nor (_09982_, _09981_, _09748_);
  or (_09983_, _09982_, _04437_);
  or (_09984_, _04436_, _07982_);
  and (_09985_, _09984_, _04432_);
  and (_09986_, _09985_, _09983_);
  or (_09987_, _09986_, _08121_);
  or (_09988_, _09987_, _09980_);
  nor (_09989_, _08131_, \oc8051_golden_model_1.PSW [7]);
  not (_09990_, _09989_);
  nor (_09991_, _09990_, _08141_);
  not (_09992_, _09991_);
  nand (_09993_, _09992_, _08121_);
  nor (_09994_, _03232_, _03201_);
  nor (_09995_, _09994_, _03533_);
  and (_09996_, _09995_, _09993_);
  and (_09997_, _09996_, _09988_);
  nor (_09998_, _05932_, _07982_);
  not (_09999_, _09998_);
  nand (_10000_, _05980_, _05932_);
  and (_10001_, _10000_, _09999_);
  and (_10002_, _10001_, _03469_);
  and (_10003_, _09758_, _03527_);
  or (_10004_, _10003_, _10002_);
  or (_10005_, _10004_, _09997_);
  and (_10006_, _10005_, _03531_);
  and (_10007_, _09982_, _03530_);
  nor (_10008_, _03232_, _03211_);
  or (_10009_, _10008_, _03465_);
  or (_10010_, _10009_, _10007_);
  or (_10011_, _10010_, _10006_);
  and (_10012_, _05975_, _05932_);
  nor (_10013_, _10012_, _09998_);
  or (_10014_, _10013_, _03466_);
  and (_10015_, _06899_, _05140_);
  nor (_10016_, _10015_, _03206_);
  nor (_10017_, _10016_, _04040_);
  and (_10018_, _10017_, _10014_);
  and (_10019_, _10018_, _10011_);
  and (_10020_, _04005_, _03457_);
  not (_10021_, _10017_);
  not (_10022_, _05254_);
  and (_10023_, _05417_, _04995_);
  nor (_10024_, _10023_, _10022_);
  nor (_10025_, _05417_, _04995_);
  not (_10026_, _10025_);
  and (_10027_, _05253_, _03409_);
  nor (_10028_, _05526_, _05275_);
  nor (_10029_, _10028_, _10027_);
  and (_10030_, _10029_, _10026_);
  and (_10031_, _10030_, _10024_);
  and (_10032_, _05526_, _05275_);
  not (_10033_, _10032_);
  nor (_10034_, _05831_, _05267_);
  and (_10035_, _05831_, _05267_);
  nor (_10036_, _10035_, _10034_);
  and (_10037_, _10036_, _10033_);
  and (_10038_, _10037_, _10031_);
  nor (_10039_, _04635_, _04566_);
  and (_10040_, _04635_, _04566_);
  and (_10041_, _04429_, _03989_);
  or (_10042_, _10041_, _10040_);
  nor (_10043_, _10042_, _10039_);
  and (_10044_, _04462_, _04139_);
  not (_10045_, _10044_);
  and (_10046_, _04885_, _03513_);
  nor (_10047_, _04885_, _03513_);
  nor (_10048_, _10047_, _10046_);
  and (_10049_, _05073_, _05005_);
  nor (_10050_, _05073_, _05005_);
  nor (_10051_, _10050_, _10049_);
  and (_10052_, _10051_, _10048_);
  and (_10053_, _10052_, _10045_);
  and (_10054_, _10053_, _10043_);
  and (_10055_, _10054_, _10038_);
  or (_10056_, _10043_, _10040_);
  nand (_10057_, _10056_, _10052_);
  and (_10058_, _10049_, _10048_);
  nor (_10059_, _10058_, _10046_);
  nand (_10060_, _10059_, _10057_);
  nand (_10061_, _10060_, _10038_);
  nor (_10062_, _10027_, _10023_);
  or (_10063_, _10062_, _10022_);
  or (_10064_, _10032_, _10035_);
  nand (_10065_, _10064_, _10031_);
  and (_10066_, _10065_, _10063_);
  and (_10067_, _10066_, _10061_);
  or (_10068_, _10067_, _10055_);
  and (_10069_, _10068_, _10021_);
  or (_10070_, _10069_, _10020_);
  or (_10071_, _10070_, _10019_);
  and (_10072_, _06757_, _03811_);
  nor (_10073_, _10072_, _06176_);
  nor (_10074_, _06114_, _04493_);
  nor (_10075_, _06526_, _03511_);
  nor (_10076_, _10075_, _10074_);
  nand (_10077_, _06526_, _03511_);
  and (_10078_, _10077_, _10076_);
  and (_10079_, _10078_, _10073_);
  nand (_10080_, _06802_, _04257_);
  or (_10081_, _06757_, _03811_);
  or (_10082_, _06802_, _04257_);
  and (_10083_, _10082_, _10081_);
  and (_10084_, _10083_, _10080_);
  and (_10085_, _10084_, _10079_);
  and (_10086_, _06664_, _03440_);
  not (_10087_, _10086_);
  or (_10088_, _06664_, _03440_);
  and (_10089_, _10088_, _10087_);
  or (_10090_, _06710_, _03944_);
  nand (_10091_, _06710_, _03944_);
  and (_10092_, _10091_, _10090_);
  and (_10093_, _10092_, _10089_);
  or (_10094_, _06572_, _04292_);
  nand (_10095_, _06617_, _03989_);
  or (_10096_, _06572_, _04566_);
  nand (_10097_, _06572_, _04566_);
  nand (_10098_, _10097_, _10096_);
  and (_10099_, _10098_, _10095_);
  not (_10100_, _10099_);
  nand (_10101_, _10100_, _10094_);
  nand (_10102_, _10101_, _10093_);
  or (_10103_, _10090_, _10086_);
  and (_10104_, _10103_, _10088_);
  nand (_10105_, _10104_, _10102_);
  nand (_10106_, _10105_, _10085_);
  or (_10107_, _10076_, _06176_);
  not (_10108_, _10079_);
  or (_10109_, _10083_, _10108_);
  and (_10110_, _10109_, _10107_);
  and (_10111_, _10110_, _10106_);
  not (_10112_, _10020_);
  or (_10113_, _06617_, _03989_);
  and (_10114_, _10099_, _10113_);
  and (_10115_, _10114_, _10093_);
  and (_10116_, _10115_, _10085_);
  or (_10117_, _10116_, _10112_);
  or (_10118_, _10117_, _10111_);
  and (_10119_, _10118_, _10071_);
  or (_10120_, _10119_, _03547_);
  and (_10121_, _10120_, _09977_);
  nor (_10122_, _03232_, _03206_);
  nor (_10123_, _10122_, _03608_);
  not (_10124_, _10123_);
  or (_10125_, _10124_, _10121_);
  nand (_10126_, _10122_, _07982_);
  nor (_10127_, _08825_, _08826_);
  nor (_10128_, _10127_, _08829_);
  or (_10129_, _04292_, \oc8051_golden_model_1.ACC [1]);
  and (_10130_, _04292_, \oc8051_golden_model_1.ACC [1]);
  and (_10131_, _03989_, \oc8051_golden_model_1.ACC [0]);
  or (_10132_, _10131_, _10130_);
  nand (_10133_, _10132_, _10129_);
  nand (_10134_, _10133_, _10128_);
  and (_10135_, _03440_, \oc8051_golden_model_1.ACC [3]);
  nor (_10136_, _03440_, \oc8051_golden_model_1.ACC [3]);
  nor (_10137_, _03944_, \oc8051_golden_model_1.ACC [2]);
  nor (_10138_, _10137_, _10136_);
  or (_10139_, _10138_, _10135_);
  nand (_10140_, _10139_, _10134_);
  nor (_10141_, _08821_, _08820_);
  nor (_10142_, _10141_, _08824_);
  nor (_10143_, _08819_, _07933_);
  and (_10144_, _10143_, _10142_);
  nand (_10145_, _10144_, _10140_);
  and (_10146_, _03811_, \oc8051_golden_model_1.ACC [5]);
  nor (_10147_, _03811_, \oc8051_golden_model_1.ACC [5]);
  nor (_10148_, _04257_, \oc8051_golden_model_1.ACC [4]);
  nor (_10149_, _10148_, _10147_);
  nor (_10150_, _10149_, _10146_);
  nand (_10151_, _10143_, _10150_);
  nand (_10152_, _03409_, _06440_);
  or (_10153_, _03511_, \oc8051_golden_model_1.ACC [6]);
  or (_10154_, _10153_, _07933_);
  and (_10155_, _10154_, _10152_);
  and (_10156_, _10155_, _10151_);
  and (_10157_, _10156_, _10145_);
  not (_10158_, _03608_);
  and (_10159_, _03989_, _03344_);
  nor (_10160_, _10159_, _08831_);
  nor (_10161_, _10160_, _07991_);
  and (_10162_, _10161_, _10128_);
  and (_10163_, _10162_, _10144_);
  or (_10164_, _10163_, _10158_);
  or (_10165_, _10164_, _10157_);
  and (_10166_, _10165_, _10126_);
  and (_10167_, _10166_, _10125_);
  or (_10168_, _10167_, _03553_);
  and (_10169_, _05258_, \oc8051_golden_model_1.P0 [2]);
  and (_10170_, _05951_, \oc8051_golden_model_1.P1 [2]);
  nor (_10171_, _10170_, _10169_);
  and (_10172_, _05953_, \oc8051_golden_model_1.P3 [2]);
  and (_10173_, _05948_, \oc8051_golden_model_1.P2 [2]);
  or (_10174_, _10173_, _10172_);
  nor (_10175_, _10174_, _09774_);
  and (_10176_, _10175_, _09784_);
  and (_10177_, _10176_, _09773_);
  and (_10178_, _10177_, _10171_);
  and (_10179_, _10178_, _05724_);
  nor (_10180_, _10179_, _09770_);
  and (_10181_, _05948_, \oc8051_golden_model_1.P2 [1]);
  and (_10182_, _05953_, \oc8051_golden_model_1.P3 [1]);
  nor (_10183_, _10182_, _10181_);
  and (_10184_, _05258_, \oc8051_golden_model_1.P0 [1]);
  and (_10185_, _05951_, \oc8051_golden_model_1.P1 [1]);
  nor (_10186_, _10185_, _10184_);
  and (_10187_, _10186_, _10183_);
  and (_10188_, _10187_, _09807_);
  and (_10189_, _10188_, _09804_);
  and (_10190_, _10189_, _05626_);
  nor (_10191_, _10190_, _09794_);
  nor (_10192_, _10191_, _10180_);
  and (_10193_, _05948_, \oc8051_golden_model_1.P2 [4]);
  and (_10194_, _05953_, \oc8051_golden_model_1.P3 [4]);
  nor (_10195_, _10194_, _10193_);
  and (_10196_, _05258_, \oc8051_golden_model_1.P0 [4]);
  and (_10197_, _05951_, \oc8051_golden_model_1.P1 [4]);
  nor (_10198_, _10197_, _10196_);
  and (_10199_, _10198_, _10195_);
  and (_10200_, _10199_, _09834_);
  and (_10201_, _10200_, _09831_);
  and (_10202_, _10201_, _05832_);
  nor (_10203_, _09821_, _10202_);
  nor (_10204_, _10203_, _06164_);
  and (_10205_, _10204_, _10192_);
  and (_10206_, _05258_, \oc8051_golden_model_1.P0 [0]);
  and (_10207_, _05953_, \oc8051_golden_model_1.P3 [0]);
  nor (_10208_, _10207_, _10206_);
  and (_10209_, _05951_, \oc8051_golden_model_1.P1 [0]);
  and (_10210_, _05948_, \oc8051_golden_model_1.P2 [0]);
  nor (_10211_, _10210_, _10209_);
  and (_10212_, _10211_, _10208_);
  and (_10213_, _10212_, _09863_);
  and (_10214_, _10213_, _05675_);
  nor (_10215_, _10214_, _09849_);
  and (_10216_, _05258_, \oc8051_golden_model_1.P0 [6]);
  and (_10217_, _05953_, \oc8051_golden_model_1.P3 [6]);
  nor (_10218_, _10217_, _10216_);
  not (_10219_, _09887_);
  and (_10220_, _05951_, \oc8051_golden_model_1.P1 [6]);
  and (_10221_, _05948_, \oc8051_golden_model_1.P2 [6]);
  nor (_10222_, _10221_, _10220_);
  and (_10223_, _10222_, _10219_);
  and (_10224_, _10223_, _10218_);
  and (_10225_, _10224_, _09886_);
  and (_10226_, _10225_, _05418_);
  nor (_10227_, _09875_, _10226_);
  nor (_10228_, _10227_, _10215_);
  and (_10229_, _05948_, \oc8051_golden_model_1.P2 [3]);
  and (_10230_, _05953_, \oc8051_golden_model_1.P3 [3]);
  nor (_10231_, _10230_, _10229_);
  and (_10232_, _05258_, \oc8051_golden_model_1.P0 [3]);
  and (_10233_, _05951_, \oc8051_golden_model_1.P1 [3]);
  nor (_10234_, _10233_, _10232_);
  and (_10235_, _10234_, _10231_);
  and (_10236_, _10235_, _09913_);
  and (_10237_, _10236_, _09910_);
  and (_10238_, _10237_, _05577_);
  nor (_10239_, _10238_, _09900_);
  and (_10240_, _05258_, \oc8051_golden_model_1.P0 [5]);
  and (_10241_, _05953_, \oc8051_golden_model_1.P3 [5]);
  nor (_10242_, _10241_, _10240_);
  and (_10243_, _05951_, \oc8051_golden_model_1.P1 [5]);
  and (_10244_, _05948_, \oc8051_golden_model_1.P2 [5]);
  nor (_10245_, _10244_, _10243_);
  and (_10246_, _10245_, _10242_);
  and (_10247_, _10246_, _09939_);
  and (_10248_, _10247_, _09933_);
  and (_10249_, _10248_, _05527_);
  nor (_10250_, _09926_, _10249_);
  nor (_10251_, _10250_, _10239_);
  and (_10252_, _10251_, _10228_);
  and (_10253_, _10252_, _10205_);
  and (_10254_, _10253_, \oc8051_golden_model_1.PSW [7]);
  nand (_10255_, _10254_, _03522_);
  and (_10256_, _09999_, _06164_);
  or (_10257_, _10256_, _03459_);
  or (_10258_, _10257_, _10001_);
  and (_10259_, _10258_, _10255_);
  and (_10260_, _10259_, _10168_);
  or (_10261_, _06933_, _03587_);
  or (_10262_, _10261_, _10260_);
  and (_10263_, _10262_, _09954_);
  or (_10264_, _10263_, _03586_);
  not (_10265_, _03586_);
  nor (_10266_, _10253_, \oc8051_golden_model_1.PSW [7]);
  or (_10267_, _10266_, _10265_);
  and (_10268_, _10267_, _08190_);
  and (_10269_, _10268_, _10264_);
  and (_10270_, _08210_, _05888_);
  and (_10271_, _10270_, _05896_);
  and (_10272_, _08206_, _08203_);
  nor (_10273_, _10272_, _08201_);
  not (_10274_, _10273_);
  and (_10275_, _08568_, _08203_);
  not (_10276_, _10275_);
  nor (_10277_, _10276_, _08255_);
  nor (_10278_, _10277_, _10274_);
  nor (_10279_, _10278_, _10271_);
  nor (_10280_, _10279_, _08184_);
  nor (_10281_, _10280_, _08191_);
  or (_10282_, _10281_, _10269_);
  or (_10283_, _10279_, _08185_);
  and (_10284_, _10283_, _08024_);
  and (_10285_, _10284_, _10282_);
  or (_10286_, _10285_, _09768_);
  and (_10287_, _10286_, _03599_);
  not (_10288_, _06160_);
  and (_10289_, _08642_, _10288_);
  and (_10290_, _08653_, _08648_);
  nor (_10291_, _10290_, _08646_);
  not (_10292_, _10291_);
  and (_10293_, _08666_, _08660_);
  not (_10294_, _10293_);
  and (_10295_, _08678_, _08672_);
  not (_10296_, _10295_);
  nor (_10297_, _08686_, _03344_);
  nor (_10298_, _10297_, _08683_);
  nor (_10299_, _10298_, _08682_);
  nor (_10300_, _10299_, _10296_);
  nor (_10301_, _08677_, _08671_);
  or (_10302_, _10301_, _08670_);
  not (_10303_, _10302_);
  nor (_10304_, _10303_, _10300_);
  and (_10305_, _08686_, _03344_);
  nor (_10306_, _10297_, _10305_);
  nor (_10307_, _08380_, _07993_);
  nor (_10308_, _10307_, _07992_);
  and (_10309_, _10308_, _08413_);
  nor (_10310_, _10308_, _08413_);
  or (_10311_, _10310_, _10309_);
  nand (_10312_, _10311_, _10306_);
  nor (_10313_, _10312_, _10296_);
  nor (_10314_, _10313_, _10304_);
  nor (_10315_, _10314_, _10294_);
  not (_10316_, _10315_);
  nor (_10317_, _08664_, _08658_);
  or (_10318_, _10317_, _08659_);
  and (_10319_, _10318_, _10316_);
  and (_10320_, _08654_, _08648_);
  not (_10321_, _10320_);
  nor (_10322_, _10321_, _10319_);
  nor (_10323_, _10322_, _10292_);
  nor (_10324_, _10323_, _10289_);
  and (_10325_, _10324_, _03594_);
  or (_10326_, _10325_, _07940_);
  or (_10327_, _10326_, _10287_);
  and (_10328_, _07957_, _07951_);
  and (_10329_, _10328_, _08014_);
  and (_10330_, _10328_, _08016_);
  not (_10331_, _10330_);
  and (_10332_, _07955_, _07951_);
  nor (_10333_, _10332_, _07949_);
  and (_10334_, _10333_, _10331_);
  not (_10335_, _10334_);
  nor (_10336_, _10335_, _10329_);
  nor (_10337_, _10336_, _09738_);
  or (_10338_, _10337_, _07941_);
  and (_10339_, _10338_, _06903_);
  and (_10340_, _10339_, _10327_);
  or (_10341_, _10340_, _09759_);
  and (_10342_, _10341_, _04500_);
  nand (_10343_, _06114_, _05303_);
  nor (_10344_, _09748_, _04500_);
  and (_10345_, _10344_, _10343_);
  or (_10346_, _10345_, _03224_);
  or (_10347_, _10346_, _10342_);
  and (_10348_, _10347_, _09756_);
  or (_10349_, _07468_, _03517_);
  or (_10350_, _10349_, _10348_);
  not (_10351_, _03517_);
  or (_10352_, _10253_, _07982_);
  or (_10353_, _10352_, _10351_);
  and (_10354_, _10353_, _04509_);
  and (_10355_, _10354_, _10350_);
  and (_10356_, _06227_, _05303_);
  nor (_10357_, _10356_, _09748_);
  and (_10358_, _10357_, _03624_);
  or (_10359_, _10358_, _10355_);
  and (_10360_, _10359_, _04121_);
  and (_10361_, _10253_, _07982_);
  and (_10362_, _10361_, _03516_);
  or (_10363_, _10362_, _10360_);
  and (_10364_, _10363_, _04527_);
  nand (_10365_, _06436_, _05303_);
  and (_10366_, _10365_, _09749_);
  and (_10367_, _10366_, _03623_);
  or (_10368_, _10367_, _03744_);
  or (_10369_, _10368_, _10364_);
  and (_10370_, _10369_, _09752_);
  or (_10371_, _10370_, _03611_);
  and (_10372_, _09749_, _05357_);
  or (_10373_, _10357_, _04523_);
  or (_10374_, _10373_, _10372_);
  and (_10375_, _10374_, _10371_);
  or (_10376_, _10375_, _03733_);
  or (_10377_, _09982_, _03734_);
  or (_10378_, _10377_, _10372_);
  and (_10379_, _10378_, _06453_);
  and (_10380_, _10379_, _10376_);
  or (_10381_, _06434_, _09753_);
  nor (_10382_, _09748_, _06453_);
  and (_10383_, _10382_, _10381_);
  or (_10384_, _10383_, _03741_);
  or (_10385_, _10384_, _10380_);
  or (_10386_, _06442_, _09753_);
  and (_10387_, _10386_, _09749_);
  or (_10388_, _10387_, _06458_);
  and (_10389_, _10388_, _08563_);
  and (_10390_, _10389_, _10385_);
  not (_10391_, _10271_);
  nor (_10392_, _08200_, _06440_);
  nor (_10393_, _10392_, _08589_);
  and (_10394_, _10393_, _10391_);
  nor (_10395_, _10394_, _08559_);
  nor (_10396_, _10395_, _08564_);
  or (_10397_, _10396_, _10390_);
  or (_10398_, _10394_, _08560_);
  and (_10399_, _10398_, _08599_);
  and (_10400_, _10399_, _10397_);
  or (_10401_, _10400_, _09747_);
  nand (_10402_, _10401_, _03732_);
  nor (_10403_, _08645_, _06440_);
  or (_10404_, _10403_, _08701_);
  or (_10405_, _10289_, _03732_);
  or (_10406_, _10405_, _10404_);
  and (_10407_, _10406_, _08709_);
  and (_10408_, _10407_, _10402_);
  or (_10409_, _10408_, _09740_);
  and (_10410_, _10409_, _08708_);
  and (_10411_, _08707_, \oc8051_golden_model_1.ACC [7]);
  or (_10412_, _10411_, _07920_);
  or (_10413_, _10412_, _10410_);
  and (_10414_, _07915_, _07882_);
  not (_10415_, _07880_);
  or (_10416_, _07883_, _07881_);
  and (_10417_, _10416_, _10415_);
  or (_10418_, _10417_, _07921_);
  or (_10419_, _10418_, _10414_);
  and (_10420_, _10419_, _10413_);
  or (_10421_, _10420_, _04184_);
  not (_10422_, _08488_);
  nor (_10423_, _08776_, _07924_);
  nor (_10424_, _10423_, _08742_);
  nand (_10425_, _10424_, _10422_);
  and (_10426_, _10425_, _03480_);
  and (_10427_, _10426_, _10421_);
  not (_10428_, _08268_);
  not (_10429_, _08269_);
  nand (_10430_, _08808_, _10429_);
  and (_10431_, _10430_, _03478_);
  and (_10432_, _10431_, _10428_);
  or (_10433_, _10432_, _08783_);
  or (_10434_, _10433_, _10427_);
  and (_10435_, _10434_, _09734_);
  nor (_10436_, _10435_, _03767_);
  and (_10437_, _09979_, _03767_);
  nor (_10438_, _10437_, _08858_);
  not (_10439_, _10438_);
  nor (_10440_, _10439_, _10436_);
  and (_10441_, _08858_, \oc8051_golden_model_1.ACC [0]);
  or (_10442_, _10441_, _10440_);
  and (_10443_, _10442_, _03446_);
  nor (_10444_, _10013_, _03446_);
  or (_10445_, _10444_, _10443_);
  and (_10446_, _10445_, _03474_);
  and (_10447_, _05886_, _05303_);
  nor (_10448_, _10447_, _09748_);
  nor (_10449_, _10448_, _03474_);
  or (_10450_, _10449_, _10446_);
  or (_10451_, _10450_, _43193_);
  or (_10452_, _43189_, \oc8051_golden_model_1.PSW [7]);
  and (_10453_, _10452_, _42003_);
  and (_40782_, _10453_, _10451_);
  not (_10454_, \oc8051_golden_model_1.PCON [7]);
  nor (_10455_, _05261_, _10454_);
  not (_10456_, _05261_);
  nor (_10457_, _06442_, _10456_);
  nor (_10458_, _10457_, _10455_);
  nor (_10459_, _10458_, _06458_);
  and (_10460_, _06227_, _05261_);
  nor (_10461_, _10460_, _10455_);
  and (_10462_, _10461_, _03624_);
  and (_10463_, _05261_, \oc8051_golden_model_1.ACC [7]);
  nor (_10464_, _10463_, _10455_);
  nor (_10465_, _10464_, _03531_);
  nor (_10466_, _10464_, _04437_);
  nor (_10467_, _04436_, _10454_);
  or (_10468_, _10467_, _10466_);
  and (_10469_, _10468_, _04432_);
  and (_10470_, _06133_, _05261_);
  nor (_10471_, _10470_, _10455_);
  nor (_10472_, _10471_, _04432_);
  or (_10473_, _10472_, _10469_);
  and (_10474_, _10473_, _04457_);
  nor (_10475_, _10456_, _05253_);
  nor (_10476_, _10475_, _10455_);
  nor (_10477_, _10476_, _04457_);
  nor (_10478_, _10477_, _10474_);
  nor (_10479_, _10478_, _03530_);
  or (_10480_, _10479_, _07454_);
  nor (_10481_, _10480_, _10465_);
  and (_10482_, _10476_, _07454_);
  nor (_10483_, _10482_, _10481_);
  nor (_10484_, _10483_, _04082_);
  and (_10485_, _06114_, _05261_);
  nor (_10486_, _10455_, _04500_);
  not (_10487_, _10486_);
  nor (_10488_, _10487_, _10485_);
  or (_10489_, _10488_, _03224_);
  nor (_10490_, _10489_, _10484_);
  nor (_10491_, _06421_, _10456_);
  nor (_10492_, _10491_, _10455_);
  nor (_10493_, _10492_, _03521_);
  or (_10494_, _10493_, _03624_);
  nor (_10495_, _10494_, _10490_);
  nor (_10496_, _10495_, _10462_);
  or (_10497_, _10496_, _03623_);
  and (_10498_, _06436_, _05261_);
  or (_10499_, _10498_, _10455_);
  or (_10500_, _10499_, _04527_);
  and (_10501_, _10500_, _03745_);
  and (_10502_, _10501_, _10497_);
  and (_10503_, _06443_, _05261_);
  nor (_10504_, _10503_, _10455_);
  nor (_10505_, _10504_, _03745_);
  nor (_10506_, _10505_, _10502_);
  nor (_10507_, _10506_, _03611_);
  nor (_10508_, _10455_, _05358_);
  not (_10509_, _10508_);
  nor (_10510_, _10461_, _04523_);
  and (_10511_, _10510_, _10509_);
  nor (_10512_, _10511_, _10507_);
  nor (_10513_, _10512_, _03733_);
  nor (_10514_, _10464_, _03734_);
  and (_10515_, _10514_, _10509_);
  or (_10516_, _10515_, _10513_);
  and (_10517_, _10516_, _06453_);
  nor (_10518_, _06434_, _10456_);
  nor (_10519_, _10518_, _10455_);
  nor (_10520_, _10519_, _06453_);
  or (_10521_, _10520_, _10517_);
  and (_10522_, _10521_, _06458_);
  nor (_10523_, _10522_, _10459_);
  nor (_10524_, _10523_, _03767_);
  nor (_10525_, _10471_, _03948_);
  or (_10526_, _10525_, _03473_);
  nor (_10527_, _10526_, _10524_);
  and (_10528_, _05886_, _05261_);
  or (_10529_, _10455_, _03474_);
  nor (_10530_, _10529_, _10528_);
  nor (_10531_, _10530_, _10527_);
  or (_10532_, _10531_, _43193_);
  or (_10533_, _43189_, \oc8051_golden_model_1.PCON [7]);
  and (_10534_, _10533_, _42003_);
  and (_40784_, _10534_, _10532_);
  not (_10535_, \oc8051_golden_model_1.SBUF [7]);
  nor (_10536_, _05270_, _10535_);
  not (_10537_, _05270_);
  nor (_10538_, _06442_, _10537_);
  nor (_10539_, _10538_, _10536_);
  nor (_10540_, _10539_, _06458_);
  and (_10541_, _06227_, _05270_);
  nor (_10542_, _10541_, _10536_);
  and (_10543_, _10542_, _03624_);
  and (_10544_, _05270_, \oc8051_golden_model_1.ACC [7]);
  nor (_10545_, _10544_, _10536_);
  nor (_10546_, _10545_, _03531_);
  nor (_10547_, _10545_, _04437_);
  nor (_10548_, _04436_, _10535_);
  or (_10549_, _10548_, _10547_);
  and (_10550_, _10549_, _04432_);
  and (_10551_, _06133_, _05270_);
  nor (_10552_, _10551_, _10536_);
  nor (_10553_, _10552_, _04432_);
  or (_10554_, _10553_, _10550_);
  and (_10555_, _10554_, _04457_);
  nor (_10556_, _10537_, _05253_);
  nor (_10557_, _10556_, _10536_);
  nor (_10558_, _10557_, _04457_);
  nor (_10559_, _10558_, _10555_);
  nor (_10560_, _10559_, _03530_);
  or (_10561_, _10560_, _07454_);
  nor (_10562_, _10561_, _10546_);
  and (_10563_, _10557_, _07454_);
  nor (_10564_, _10563_, _10562_);
  nor (_10565_, _10564_, _04082_);
  and (_10566_, _06114_, _05270_);
  nor (_10567_, _10536_, _04500_);
  not (_10568_, _10567_);
  nor (_10569_, _10568_, _10566_);
  or (_10570_, _10569_, _03224_);
  nor (_10571_, _10570_, _10565_);
  nor (_10572_, _06421_, _10537_);
  nor (_10573_, _10572_, _10536_);
  nor (_10574_, _10573_, _03521_);
  or (_10575_, _10574_, _03624_);
  nor (_10576_, _10575_, _10571_);
  nor (_10577_, _10576_, _10543_);
  or (_10578_, _10577_, _03623_);
  and (_10579_, _06436_, _05270_);
  or (_10580_, _10579_, _10536_);
  or (_10581_, _10580_, _04527_);
  and (_10582_, _10581_, _03745_);
  and (_10583_, _10582_, _10578_);
  and (_10584_, _06443_, _05270_);
  nor (_10585_, _10584_, _10536_);
  nor (_10586_, _10585_, _03745_);
  nor (_10587_, _10586_, _10583_);
  nor (_10588_, _10587_, _03611_);
  nor (_10589_, _10536_, _05358_);
  not (_10590_, _10589_);
  nor (_10591_, _10542_, _04523_);
  and (_10592_, _10591_, _10590_);
  nor (_10593_, _10592_, _10588_);
  nor (_10594_, _10593_, _03733_);
  nor (_10595_, _10545_, _03734_);
  and (_10596_, _10595_, _10590_);
  or (_10597_, _10596_, _10594_);
  and (_10598_, _10597_, _06453_);
  nor (_10599_, _06434_, _10537_);
  nor (_10600_, _10599_, _10536_);
  nor (_10601_, _10600_, _06453_);
  or (_10602_, _10601_, _10598_);
  and (_10603_, _10602_, _06458_);
  nor (_10604_, _10603_, _10540_);
  nor (_10605_, _10604_, _03767_);
  nor (_10606_, _10552_, _03948_);
  or (_10607_, _10606_, _03473_);
  nor (_10608_, _10607_, _10605_);
  and (_10609_, _05886_, _05270_);
  or (_10610_, _10536_, _03474_);
  nor (_10611_, _10610_, _10609_);
  nor (_10612_, _10611_, _10608_);
  or (_10613_, _10612_, _43193_);
  or (_10614_, _43189_, \oc8051_golden_model_1.SBUF [7]);
  and (_10615_, _10614_, _42003_);
  and (_40785_, _10615_, _10613_);
  not (_10616_, \oc8051_golden_model_1.SCON [7]);
  nor (_10617_, _05333_, _10616_);
  not (_10618_, _05333_);
  nor (_10619_, _10618_, _05253_);
  nor (_10620_, _10619_, _10617_);
  and (_10621_, _10620_, _07454_);
  nor (_10622_, _05942_, _10616_);
  and (_10623_, _05975_, _05942_);
  nor (_10624_, _10623_, _10622_);
  nor (_10625_, _10624_, _03466_);
  and (_10626_, _05333_, \oc8051_golden_model_1.ACC [7]);
  nor (_10627_, _10626_, _10617_);
  nor (_10628_, _10627_, _04437_);
  nor (_10629_, _04436_, _10616_);
  or (_10630_, _10629_, _10628_);
  and (_10631_, _10630_, _04432_);
  and (_10632_, _06133_, _05333_);
  nor (_10633_, _10632_, _10617_);
  nor (_10634_, _10633_, _04432_);
  or (_10635_, _10634_, _10631_);
  and (_10636_, _10635_, _03470_);
  and (_10637_, _05980_, _05942_);
  nor (_10638_, _10637_, _10622_);
  nor (_10639_, _10638_, _03470_);
  or (_10640_, _10639_, _03527_);
  or (_10641_, _10640_, _10636_);
  nand (_10642_, _10620_, _03527_);
  and (_10643_, _10642_, _10641_);
  and (_10644_, _10643_, _03531_);
  nor (_10645_, _10627_, _03531_);
  or (_10646_, _10645_, _10644_);
  and (_10647_, _10646_, _03466_);
  nor (_10648_, _10647_, _10625_);
  nor (_10649_, _10648_, _03458_);
  nor (_10650_, _10622_, _06165_);
  or (_10651_, _10638_, _03459_);
  nor (_10652_, _10651_, _10650_);
  nor (_10653_, _10652_, _10649_);
  nor (_10654_, _10653_, _03452_);
  not (_10655_, _05942_);
  nor (_10656_, _05962_, _10655_);
  nor (_10657_, _10656_, _10622_);
  nor (_10658_, _10657_, _03453_);
  nor (_10659_, _10658_, _07454_);
  not (_10660_, _10659_);
  nor (_10661_, _10660_, _10654_);
  nor (_10662_, _10661_, _10621_);
  nor (_10663_, _10662_, _04082_);
  and (_10664_, _06114_, _05333_);
  nor (_10665_, _10617_, _04500_);
  not (_10666_, _10665_);
  nor (_10667_, _10666_, _10664_);
  nor (_10668_, _10667_, _03224_);
  not (_10669_, _10668_);
  nor (_10670_, _10669_, _10663_);
  nor (_10671_, _06421_, _10618_);
  nor (_10672_, _10671_, _10617_);
  nor (_10673_, _10672_, _03521_);
  or (_10674_, _10673_, _08905_);
  or (_10675_, _10674_, _10670_);
  and (_10676_, _06436_, _05333_);
  or (_10677_, _10617_, _04527_);
  or (_10678_, _10677_, _10676_);
  and (_10679_, _06227_, _05333_);
  nor (_10680_, _10679_, _10617_);
  and (_10681_, _10680_, _03624_);
  nor (_10682_, _10681_, _03744_);
  and (_10683_, _10682_, _10678_);
  and (_10684_, _10683_, _10675_);
  and (_10685_, _06443_, _05333_);
  nor (_10686_, _10685_, _10617_);
  nor (_10687_, _10686_, _03745_);
  nor (_10688_, _10687_, _10684_);
  nor (_10689_, _10688_, _03611_);
  nor (_10690_, _10617_, _05358_);
  not (_10691_, _10690_);
  nor (_10692_, _10680_, _04523_);
  and (_10693_, _10692_, _10691_);
  nor (_10694_, _10693_, _10689_);
  nor (_10695_, _10694_, _03733_);
  nor (_10696_, _10627_, _03734_);
  and (_10697_, _10696_, _10691_);
  nor (_10698_, _10697_, _03618_);
  not (_10700_, _10698_);
  nor (_10701_, _10700_, _10695_);
  nor (_10702_, _06434_, _10618_);
  or (_10703_, _10617_, _06453_);
  nor (_10704_, _10703_, _10702_);
  or (_10705_, _10704_, _03741_);
  nor (_10706_, _10705_, _10701_);
  nor (_10707_, _06442_, _10618_);
  nor (_10708_, _10707_, _10617_);
  nor (_10709_, _10708_, _06458_);
  or (_10711_, _10709_, _10706_);
  and (_10712_, _10711_, _03948_);
  nor (_10713_, _10633_, _03948_);
  or (_10714_, _10713_, _10712_);
  and (_10715_, _10714_, _03446_);
  nor (_10716_, _10624_, _03446_);
  or (_10717_, _10716_, _10715_);
  and (_10718_, _10717_, _03474_);
  and (_10719_, _05886_, _05333_);
  nor (_10720_, _10719_, _10617_);
  nor (_10722_, _10720_, _03474_);
  or (_10723_, _10722_, _10718_);
  or (_10724_, _10723_, _43193_);
  or (_10725_, _43189_, \oc8051_golden_model_1.SCON [7]);
  and (_10726_, _10725_, _42003_);
  and (_40786_, _10726_, _10724_);
  and (_10727_, _04891_, \oc8051_golden_model_1.SP [4]);
  and (_10728_, _10727_, \oc8051_golden_model_1.SP [5]);
  and (_10729_, _10728_, \oc8051_golden_model_1.SP [6]);
  nor (_10730_, _10729_, \oc8051_golden_model_1.SP [7]);
  and (_10732_, _10729_, \oc8051_golden_model_1.SP [7]);
  nor (_10733_, _10732_, _10730_);
  nor (_10734_, _10733_, _04553_);
  not (_10735_, _03752_);
  not (_10736_, \oc8051_golden_model_1.SP [7]);
  nor (_10737_, _05323_, _10736_);
  and (_10738_, _06443_, _05323_);
  nor (_10739_, _10738_, _10737_);
  nor (_10740_, _10739_, _03745_);
  not (_10741_, _05323_);
  nor (_10743_, _10741_, _05253_);
  nor (_10744_, _10743_, _10737_);
  nor (_10745_, _10744_, _06903_);
  or (_10746_, _10745_, _04082_);
  and (_10747_, _06133_, _05323_);
  nor (_10748_, _10747_, _10737_);
  and (_10749_, _10748_, _03534_);
  and (_10750_, _05323_, \oc8051_golden_model_1.ACC [7]);
  nor (_10751_, _10750_, _10737_);
  or (_10752_, _10751_, _04437_);
  nor (_10754_, _04436_, _04435_);
  nand (_10755_, _10754_, \oc8051_golden_model_1.SP [7]);
  not (_10756_, _10733_);
  nor (_10757_, _10756_, _03204_);
  nor (_10758_, _10757_, _03534_);
  and (_10759_, _10758_, _10755_);
  and (_10760_, _10759_, _10752_);
  nor (_10761_, _10760_, _05977_);
  not (_10762_, _10761_);
  nor (_10763_, _10762_, _10749_);
  nor (_10765_, _10756_, _03202_);
  or (_10766_, _10765_, _03527_);
  nor (_10767_, _10766_, _10763_);
  not (_10768_, \oc8051_golden_model_1.SP [6]);
  not (_10769_, \oc8051_golden_model_1.SP [5]);
  not (_10770_, \oc8051_golden_model_1.SP [4]);
  and (_10771_, _06015_, _10770_);
  and (_10772_, _10771_, _10769_);
  and (_10773_, _10772_, _10768_);
  and (_10774_, _10773_, _03455_);
  nor (_10775_, _10774_, _10736_);
  and (_10776_, _10774_, _10736_);
  nor (_10777_, _10776_, _10775_);
  and (_10778_, _10777_, _03527_);
  nor (_10779_, _10778_, _10767_);
  and (_10780_, _10779_, _03531_);
  nor (_10781_, _10751_, _03531_);
  or (_10782_, _10781_, _10780_);
  and (_10783_, _10782_, _04577_);
  and (_10784_, _10729_, \oc8051_golden_model_1.SP [0]);
  nor (_10785_, _10784_, _10736_);
  and (_10786_, _10784_, _10736_);
  nor (_10787_, _10786_, _10785_);
  nor (_10788_, _10787_, _04577_);
  nor (_10789_, _10788_, _04756_);
  not (_10790_, _10789_);
  nor (_10791_, _10790_, _10783_);
  and (_10792_, _10756_, _04756_);
  or (_10793_, _10792_, _07454_);
  nor (_10794_, _10793_, _10791_);
  nor (_10795_, _10794_, _10746_);
  and (_10796_, _06114_, _05323_);
  nor (_10797_, _10737_, _04500_);
  not (_10798_, _10797_);
  nor (_10799_, _10798_, _10796_);
  nor (_10800_, _10799_, _03224_);
  not (_10801_, _10800_);
  nor (_10802_, _10801_, _10795_);
  nor (_10803_, _06421_, _10741_);
  nor (_10804_, _10803_, _10737_);
  nor (_10805_, _10804_, _03521_);
  or (_10806_, _10805_, _03624_);
  or (_10807_, _10806_, _10802_);
  and (_10808_, _06227_, _05323_);
  nor (_10809_, _10808_, _10737_);
  nand (_10810_, _10809_, _03624_);
  and (_10811_, _10810_, _10807_);
  nor (_10812_, _10811_, _03168_);
  and (_10813_, _10756_, _03168_);
  nor (_10814_, _10813_, _10812_);
  nor (_10815_, _10814_, _03623_);
  and (_10816_, _06436_, _05323_);
  or (_10817_, _10737_, _04527_);
  nor (_10818_, _10817_, _10816_);
  or (_10819_, _10818_, _03744_);
  nor (_10820_, _10819_, _10815_);
  nor (_10821_, _10820_, _10740_);
  nor (_10822_, _10821_, _03611_);
  nor (_10823_, _10737_, _05358_);
  not (_10824_, _10823_);
  nor (_10825_, _10809_, _04523_);
  and (_10826_, _10825_, _10824_);
  nor (_10827_, _10826_, _10822_);
  nor (_10828_, _03733_, _03182_);
  not (_10829_, _10828_);
  nor (_10830_, _10829_, _10827_);
  and (_10831_, _10733_, _03182_);
  or (_10832_, _10823_, _03734_);
  nor (_10833_, _10832_, _10751_);
  nor (_10834_, _10833_, _10831_);
  and (_10835_, _10834_, _06453_);
  not (_10836_, _10835_);
  nor (_10837_, _10836_, _10830_);
  nor (_10838_, _06434_, _10741_);
  nor (_10839_, _10838_, _10737_);
  and (_10840_, _10839_, _03618_);
  nor (_10841_, _10840_, _10837_);
  and (_10842_, _10841_, _06458_);
  nor (_10843_, _06442_, _10741_);
  nor (_10844_, _10843_, _10737_);
  nor (_10845_, _10844_, _06458_);
  or (_10846_, _10845_, _10842_);
  and (_10847_, _10846_, _10735_);
  nor (_10848_, _03752_, _03191_);
  nor (_10849_, _10773_, \oc8051_golden_model_1.SP [7]);
  and (_10850_, _10773_, \oc8051_golden_model_1.SP [7]);
  nor (_10851_, _10850_, _10849_);
  nor (_10852_, _10851_, _03191_);
  nor (_10853_, _10852_, _10848_);
  nor (_10854_, _10853_, _10847_);
  and (_10855_, _10756_, _03191_);
  nor (_10856_, _10855_, _10854_);
  and (_10857_, _10856_, _03476_);
  and (_10858_, _10851_, _03475_);
  or (_10859_, _10858_, _10857_);
  and (_10860_, _10859_, _03948_);
  nor (_10861_, _10748_, _03948_);
  nor (_10862_, _10861_, _04986_);
  not (_10863_, _10862_);
  nor (_10864_, _10863_, _10860_);
  nor (_10865_, _10864_, _10734_);
  and (_10866_, _10865_, _03474_);
  and (_10867_, _05886_, _05323_);
  nor (_10868_, _10867_, _10737_);
  nor (_10869_, _10868_, _03474_);
  or (_10870_, _10869_, _10866_);
  or (_10871_, _10870_, _43193_);
  or (_10872_, _43189_, \oc8051_golden_model_1.SP [7]);
  and (_10873_, _10872_, _42003_);
  and (_40787_, _10873_, _10871_);
  not (_10874_, \oc8051_golden_model_1.TCON [7]);
  nor (_10875_, _05286_, _10874_);
  not (_10876_, _05286_);
  nor (_10877_, _10876_, _05253_);
  nor (_10878_, _10877_, _10875_);
  and (_10879_, _10878_, _07454_);
  nor (_10880_, _05924_, _10874_);
  and (_10881_, _05975_, _05924_);
  nor (_10882_, _10881_, _10880_);
  nor (_10883_, _10882_, _03466_);
  and (_10884_, _05286_, \oc8051_golden_model_1.ACC [7]);
  nor (_10885_, _10884_, _10875_);
  nor (_10886_, _10885_, _04437_);
  nor (_10887_, _04436_, _10874_);
  or (_10888_, _10887_, _10886_);
  and (_10889_, _10888_, _04432_);
  and (_10890_, _06133_, _05286_);
  nor (_10891_, _10890_, _10875_);
  nor (_10892_, _10891_, _04432_);
  or (_10893_, _10892_, _10889_);
  and (_10894_, _10893_, _03470_);
  and (_10895_, _05980_, _05924_);
  nor (_10896_, _10895_, _10880_);
  nor (_10897_, _10896_, _03470_);
  or (_10898_, _10897_, _03527_);
  or (_10899_, _10898_, _10894_);
  nand (_10900_, _10878_, _03527_);
  and (_10901_, _10900_, _10899_);
  and (_10902_, _10901_, _03531_);
  nor (_10903_, _10885_, _03531_);
  or (_10904_, _10903_, _10902_);
  and (_10905_, _10904_, _03466_);
  nor (_10906_, _10905_, _10883_);
  nor (_10907_, _10906_, _03458_);
  and (_10908_, _06166_, _05924_);
  nor (_10909_, _10908_, _10880_);
  nor (_10910_, _10909_, _03459_);
  nor (_10911_, _10910_, _10907_);
  nor (_10912_, _10911_, _03452_);
  not (_10913_, _05924_);
  nor (_10914_, _05962_, _10913_);
  nor (_10915_, _10914_, _10880_);
  nor (_10916_, _10915_, _03453_);
  nor (_10917_, _10916_, _07454_);
  not (_10918_, _10917_);
  nor (_10919_, _10918_, _10912_);
  nor (_10920_, _10919_, _10879_);
  nor (_10921_, _10920_, _04082_);
  and (_10922_, _06114_, _05286_);
  nor (_10923_, _10875_, _04500_);
  not (_10924_, _10923_);
  nor (_10925_, _10924_, _10922_);
  nor (_10926_, _10925_, _03224_);
  not (_10927_, _10926_);
  nor (_10928_, _10927_, _10921_);
  nor (_10929_, _06421_, _10876_);
  nor (_10930_, _10929_, _10875_);
  nor (_10931_, _10930_, _03521_);
  or (_10932_, _10931_, _08905_);
  or (_10933_, _10932_, _10928_);
  and (_10934_, _06436_, _05286_);
  or (_10935_, _10875_, _04527_);
  or (_10936_, _10935_, _10934_);
  and (_10937_, _06227_, _05286_);
  nor (_10938_, _10937_, _10875_);
  and (_10939_, _10938_, _03624_);
  nor (_10940_, _10939_, _03744_);
  and (_10941_, _10940_, _10936_);
  and (_10942_, _10941_, _10933_);
  and (_10943_, _06443_, _05286_);
  nor (_10944_, _10943_, _10875_);
  nor (_10945_, _10944_, _03745_);
  nor (_10946_, _10945_, _10942_);
  nor (_10947_, _10946_, _03611_);
  nor (_10948_, _10875_, _05358_);
  not (_10949_, _10948_);
  nor (_10950_, _10938_, _04523_);
  and (_10951_, _10950_, _10949_);
  nor (_10952_, _10951_, _10947_);
  nor (_10953_, _10952_, _03733_);
  nor (_10954_, _10885_, _03734_);
  and (_10955_, _10954_, _10949_);
  or (_10956_, _10955_, _10953_);
  and (_10957_, _10956_, _06453_);
  nor (_10958_, _06434_, _10876_);
  nor (_10959_, _10958_, _10875_);
  nor (_10960_, _10959_, _06453_);
  or (_10961_, _10960_, _10957_);
  and (_10962_, _10961_, _06458_);
  nor (_10963_, _06442_, _10876_);
  nor (_10964_, _10963_, _10875_);
  nor (_10965_, _10964_, _06458_);
  or (_10966_, _10965_, _10962_);
  and (_10967_, _10966_, _03948_);
  nor (_10968_, _10891_, _03948_);
  or (_10969_, _10968_, _10967_);
  and (_10970_, _10969_, _03446_);
  nor (_10971_, _10882_, _03446_);
  or (_10972_, _10971_, _10970_);
  and (_10973_, _10972_, _03474_);
  and (_10974_, _05886_, _05286_);
  nor (_10975_, _10974_, _10875_);
  nor (_10976_, _10975_, _03474_);
  or (_10977_, _10976_, _10973_);
  or (_10978_, _10977_, _43193_);
  or (_10979_, _43189_, \oc8051_golden_model_1.TCON [7]);
  and (_10980_, _10979_, _42003_);
  and (_40788_, _10980_, _10978_);
  not (_10981_, \oc8051_golden_model_1.TH0 [7]);
  nor (_10982_, _05339_, _10981_);
  not (_10983_, _05339_);
  nor (_10984_, _06442_, _10983_);
  nor (_10985_, _10984_, _10982_);
  nor (_10986_, _10985_, _06458_);
  and (_10987_, _06227_, _05339_);
  nor (_10988_, _10987_, _10982_);
  and (_10989_, _10988_, _03624_);
  nor (_10990_, _10983_, _05253_);
  nor (_10991_, _10990_, _10982_);
  and (_10992_, _10991_, _07454_);
  and (_10993_, _05339_, \oc8051_golden_model_1.ACC [7]);
  nor (_10994_, _10993_, _10982_);
  nor (_10995_, _10994_, _04437_);
  nor (_10996_, _04436_, _10981_);
  or (_10997_, _10996_, _10995_);
  and (_10998_, _10997_, _04432_);
  and (_10999_, _06133_, _05339_);
  nor (_11000_, _10999_, _10982_);
  nor (_11001_, _11000_, _04432_);
  or (_11002_, _11001_, _10998_);
  and (_11003_, _11002_, _04457_);
  nor (_11004_, _10991_, _04457_);
  nor (_11005_, _11004_, _11003_);
  nor (_11006_, _11005_, _03530_);
  nor (_11007_, _10994_, _03531_);
  nor (_11008_, _11007_, _07454_);
  not (_11009_, _11008_);
  nor (_11010_, _11009_, _11006_);
  nor (_11011_, _11010_, _10992_);
  nor (_11012_, _11011_, _04082_);
  and (_11013_, _06114_, _05339_);
  nor (_11014_, _10982_, _04500_);
  not (_11015_, _11014_);
  nor (_11016_, _11015_, _11013_);
  or (_11017_, _11016_, _03224_);
  nor (_11018_, _11017_, _11012_);
  nor (_11019_, _06421_, _10983_);
  nor (_11020_, _11019_, _10982_);
  nor (_11021_, _11020_, _03521_);
  or (_11022_, _11021_, _03624_);
  nor (_11023_, _11022_, _11018_);
  nor (_11024_, _11023_, _10989_);
  or (_11025_, _11024_, _03623_);
  and (_11026_, _06436_, _05339_);
  or (_11027_, _11026_, _10982_);
  or (_11028_, _11027_, _04527_);
  and (_11029_, _11028_, _03745_);
  and (_11030_, _11029_, _11025_);
  and (_11031_, _06443_, _05339_);
  nor (_11032_, _11031_, _10982_);
  nor (_11033_, _11032_, _03745_);
  nor (_11034_, _11033_, _11030_);
  nor (_11035_, _11034_, _03611_);
  nor (_11036_, _10982_, _05358_);
  not (_11037_, _11036_);
  nor (_11038_, _10988_, _04523_);
  and (_11039_, _11038_, _11037_);
  nor (_11040_, _11039_, _11035_);
  nor (_11041_, _11040_, _03733_);
  nor (_11042_, _10994_, _03734_);
  and (_11043_, _11042_, _11037_);
  nor (_11044_, _11043_, _03618_);
  not (_11045_, _11044_);
  nor (_11046_, _11045_, _11041_);
  nor (_11047_, _06434_, _10983_);
  or (_11048_, _10982_, _06453_);
  nor (_11049_, _11048_, _11047_);
  or (_11050_, _11049_, _03741_);
  nor (_11051_, _11050_, _11046_);
  nor (_11052_, _11051_, _10986_);
  nor (_11053_, _11052_, _03767_);
  nor (_11054_, _11000_, _03948_);
  or (_11055_, _11054_, _03473_);
  nor (_11056_, _11055_, _11053_);
  and (_11057_, _05886_, _05339_);
  or (_11058_, _10982_, _03474_);
  nor (_11059_, _11058_, _11057_);
  nor (_11060_, _11059_, _11056_);
  or (_11061_, _11060_, _43193_);
  or (_11062_, _43189_, \oc8051_golden_model_1.TH0 [7]);
  and (_11063_, _11062_, _42003_);
  and (_40790_, _11063_, _11061_);
  not (_11064_, \oc8051_golden_model_1.TH1 [7]);
  nor (_11065_, _05342_, _11064_);
  not (_11066_, _05342_);
  nor (_11067_, _06442_, _11066_);
  nor (_11068_, _11067_, _11065_);
  nor (_11069_, _11068_, _06458_);
  and (_11070_, _06227_, _05342_);
  nor (_11071_, _11070_, _11065_);
  and (_11072_, _11071_, _03624_);
  and (_11073_, _05342_, \oc8051_golden_model_1.ACC [7]);
  nor (_11074_, _11073_, _11065_);
  nor (_11075_, _11074_, _03531_);
  nor (_11076_, _11074_, _04437_);
  nor (_11077_, _04436_, _11064_);
  or (_11078_, _11077_, _11076_);
  and (_11079_, _11078_, _04432_);
  and (_11080_, _06133_, _05342_);
  nor (_11081_, _11080_, _11065_);
  nor (_11082_, _11081_, _04432_);
  or (_11083_, _11082_, _11079_);
  and (_11084_, _11083_, _04457_);
  nor (_11085_, _11066_, _05253_);
  nor (_11086_, _11085_, _11065_);
  nor (_11087_, _11086_, _04457_);
  nor (_11088_, _11087_, _11084_);
  nor (_11089_, _11088_, _03530_);
  or (_11090_, _11089_, _07454_);
  nor (_11091_, _11090_, _11075_);
  and (_11092_, _11086_, _07454_);
  nor (_11093_, _11092_, _11091_);
  nor (_11094_, _11093_, _04082_);
  and (_11095_, _06114_, _05342_);
  nor (_11096_, _11065_, _04500_);
  not (_11097_, _11096_);
  nor (_11098_, _11097_, _11095_);
  or (_11099_, _11098_, _03224_);
  nor (_11100_, _11099_, _11094_);
  nor (_11101_, _06421_, _11066_);
  nor (_11102_, _11101_, _11065_);
  nor (_11103_, _11102_, _03521_);
  or (_11104_, _11103_, _03624_);
  nor (_11105_, _11104_, _11100_);
  nor (_11106_, _11105_, _11072_);
  or (_11107_, _11106_, _03623_);
  and (_11108_, _06436_, _05342_);
  or (_11109_, _11108_, _11065_);
  or (_11110_, _11109_, _04527_);
  and (_11111_, _11110_, _03745_);
  and (_11112_, _11111_, _11107_);
  and (_11113_, _06443_, _05342_);
  nor (_11114_, _11113_, _11065_);
  nor (_11115_, _11114_, _03745_);
  nor (_11116_, _11115_, _11112_);
  nor (_11117_, _11116_, _03611_);
  nor (_11118_, _11065_, _05358_);
  not (_11119_, _11118_);
  nor (_11120_, _11071_, _04523_);
  and (_11121_, _11120_, _11119_);
  nor (_11122_, _11121_, _11117_);
  nor (_11123_, _11122_, _03733_);
  nor (_11124_, _11074_, _03734_);
  and (_11125_, _11124_, _11119_);
  or (_11126_, _11125_, _11123_);
  and (_11127_, _11126_, _06453_);
  nor (_11128_, _06434_, _11066_);
  nor (_11129_, _11128_, _11065_);
  nor (_11130_, _11129_, _06453_);
  or (_11131_, _11130_, _11127_);
  and (_11132_, _11131_, _06458_);
  nor (_11133_, _11132_, _11069_);
  nor (_11134_, _11133_, _03767_);
  nor (_11135_, _11081_, _03948_);
  or (_11136_, _11135_, _03473_);
  nor (_11137_, _11136_, _11134_);
  and (_11138_, _05886_, _05342_);
  or (_11139_, _11065_, _03474_);
  nor (_11140_, _11139_, _11138_);
  nor (_11141_, _11140_, _11137_);
  or (_11142_, _11141_, _43193_);
  or (_11143_, _43189_, \oc8051_golden_model_1.TH1 [7]);
  and (_11144_, _11143_, _42003_);
  and (_40791_, _11144_, _11142_);
  not (_11145_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11146_, _05348_, _11145_);
  not (_11147_, _05348_);
  nor (_11148_, _06442_, _11147_);
  nor (_11149_, _11148_, _11146_);
  nor (_11150_, _11149_, _06458_);
  and (_11151_, _06227_, _05348_);
  nor (_11152_, _11151_, _11146_);
  and (_11153_, _11152_, _03624_);
  and (_11154_, _05348_, \oc8051_golden_model_1.ACC [7]);
  nor (_11155_, _11154_, _11146_);
  nor (_11156_, _11155_, _03531_);
  nor (_11157_, _11155_, _04437_);
  nor (_11158_, _04436_, _11145_);
  or (_11159_, _11158_, _11157_);
  and (_11160_, _11159_, _04432_);
  and (_11161_, _06133_, _05348_);
  nor (_11162_, _11161_, _11146_);
  nor (_11163_, _11162_, _04432_);
  or (_11164_, _11163_, _11160_);
  and (_11165_, _11164_, _04457_);
  nor (_11166_, _11147_, _05253_);
  nor (_11167_, _11166_, _11146_);
  nor (_11168_, _11167_, _04457_);
  nor (_11169_, _11168_, _11165_);
  nor (_11170_, _11169_, _03530_);
  or (_11171_, _11170_, _07454_);
  nor (_11172_, _11171_, _11156_);
  and (_11173_, _11167_, _07454_);
  nor (_11174_, _11173_, _11172_);
  nor (_11175_, _11174_, _04082_);
  and (_11176_, _06114_, _05348_);
  nor (_11177_, _11146_, _04500_);
  not (_11178_, _11177_);
  nor (_11179_, _11178_, _11176_);
  or (_11180_, _11179_, _03224_);
  nor (_11181_, _11180_, _11175_);
  nor (_11182_, _06421_, _11147_);
  nor (_11183_, _11182_, _11146_);
  nor (_11184_, _11183_, _03521_);
  or (_11185_, _11184_, _03624_);
  nor (_11186_, _11185_, _11181_);
  nor (_11187_, _11186_, _11153_);
  or (_11188_, _11187_, _03623_);
  and (_11189_, _06436_, _05348_);
  or (_11190_, _11189_, _11146_);
  or (_11191_, _11190_, _04527_);
  and (_11192_, _11191_, _03745_);
  and (_11193_, _11192_, _11188_);
  and (_11194_, _06443_, _05348_);
  nor (_11195_, _11194_, _11146_);
  nor (_11196_, _11195_, _03745_);
  nor (_11197_, _11196_, _11193_);
  nor (_11198_, _11197_, _03611_);
  nor (_11199_, _11146_, _05358_);
  not (_11200_, _11199_);
  nor (_11201_, _11152_, _04523_);
  and (_11202_, _11201_, _11200_);
  nor (_11203_, _11202_, _11198_);
  nor (_11204_, _11203_, _03733_);
  nor (_11205_, _11155_, _03734_);
  and (_11206_, _11205_, _11200_);
  nor (_11207_, _11206_, _03618_);
  not (_11208_, _11207_);
  nor (_11209_, _11208_, _11204_);
  nor (_11210_, _06434_, _11147_);
  or (_11211_, _11146_, _06453_);
  nor (_11212_, _11211_, _11210_);
  or (_11213_, _11212_, _03741_);
  nor (_11214_, _11213_, _11209_);
  nor (_11215_, _11214_, _11150_);
  nor (_11216_, _11215_, _03767_);
  nor (_11217_, _11162_, _03948_);
  or (_11218_, _11217_, _03473_);
  nor (_11219_, _11218_, _11216_);
  and (_11220_, _05886_, _05348_);
  nor (_11221_, _11220_, _11146_);
  and (_11222_, _11221_, _03473_);
  nor (_11223_, _11222_, _11219_);
  or (_11224_, _11223_, _43193_);
  or (_11225_, _43189_, \oc8051_golden_model_1.TL0 [7]);
  and (_11226_, _11225_, _42003_);
  and (_40792_, _11226_, _11224_);
  not (_11227_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11228_, _05444_, _11227_);
  not (_11229_, _05350_);
  nor (_11230_, _06442_, _11229_);
  nor (_11231_, _11230_, _11228_);
  nor (_11232_, _11231_, _06458_);
  and (_11233_, _06227_, _05444_);
  nor (_11234_, _11233_, _11228_);
  and (_11235_, _11234_, _03624_);
  and (_11236_, _05444_, \oc8051_golden_model_1.ACC [7]);
  nor (_11237_, _11236_, _11228_);
  nor (_11238_, _11237_, _03531_);
  nor (_11239_, _11237_, _04437_);
  nor (_11240_, _04436_, _11227_);
  or (_11241_, _11240_, _11239_);
  and (_11242_, _11241_, _04432_);
  and (_11243_, _06133_, _05350_);
  nor (_11244_, _11243_, _11228_);
  nor (_11245_, _11244_, _04432_);
  or (_11246_, _11245_, _11242_);
  and (_11247_, _11246_, _04457_);
  nor (_11248_, _11229_, _05253_);
  nor (_11249_, _11248_, _11228_);
  nor (_11250_, _11249_, _04457_);
  nor (_11251_, _11250_, _11247_);
  nor (_11252_, _11251_, _03530_);
  or (_11253_, _11252_, _07454_);
  nor (_11254_, _11253_, _11238_);
  and (_11255_, _11249_, _07454_);
  nor (_11256_, _11255_, _11254_);
  nor (_11257_, _11256_, _04082_);
  nor (_11258_, _11228_, _04500_);
  nand (_11259_, _06114_, _05444_);
  and (_11260_, _11259_, _11258_);
  or (_11261_, _11260_, _03224_);
  nor (_11262_, _11261_, _11257_);
  not (_11263_, _05444_);
  nor (_11264_, _06421_, _11263_);
  nor (_11265_, _11264_, _11228_);
  nor (_11266_, _11265_, _03521_);
  or (_11267_, _11266_, _03624_);
  nor (_11268_, _11267_, _11262_);
  nor (_11269_, _11268_, _11235_);
  or (_11270_, _11269_, _03623_);
  and (_11271_, _06436_, _05444_);
  or (_11272_, _11271_, _11228_);
  or (_11273_, _11272_, _04527_);
  and (_11274_, _11273_, _03745_);
  and (_11275_, _11274_, _11270_);
  and (_11276_, _06443_, _05350_);
  nor (_11277_, _11276_, _11228_);
  nor (_11278_, _11277_, _03745_);
  nor (_11279_, _11278_, _11275_);
  nor (_11280_, _11279_, _03611_);
  nor (_11281_, _11228_, _05358_);
  not (_11282_, _11281_);
  nor (_11283_, _11234_, _04523_);
  and (_11284_, _11283_, _11282_);
  nor (_11285_, _11284_, _11280_);
  nor (_11286_, _11285_, _03733_);
  nor (_11287_, _11237_, _03734_);
  and (_11288_, _11287_, _11282_);
  nor (_11289_, _11288_, _03618_);
  not (_11290_, _11289_);
  nor (_11291_, _11290_, _11286_);
  or (_11292_, _06434_, _11229_);
  nor (_11293_, _11228_, _06453_);
  and (_11294_, _11293_, _11292_);
  or (_11295_, _11294_, _03741_);
  nor (_11296_, _11295_, _11291_);
  nor (_11297_, _11296_, _11232_);
  nor (_11298_, _11297_, _03767_);
  nor (_11299_, _11244_, _03948_);
  or (_11300_, _11299_, _03473_);
  nor (_11301_, _11300_, _11298_);
  nand (_11302_, _05886_, _05350_);
  nor (_11303_, _11228_, _03474_);
  and (_11304_, _11303_, _11302_);
  nor (_11305_, _11304_, _11301_);
  or (_11306_, _11305_, _43193_);
  or (_11307_, _43189_, \oc8051_golden_model_1.TL1 [7]);
  and (_11308_, _11307_, _42003_);
  and (_40793_, _11308_, _11306_);
  not (_11309_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11310_, _05331_, _11309_);
  not (_11311_, _05331_);
  nor (_11312_, _06442_, _11311_);
  nor (_11313_, _11312_, _11310_);
  nor (_11314_, _11313_, _06458_);
  and (_11315_, _06227_, _05331_);
  nor (_11316_, _11315_, _11310_);
  and (_11317_, _11316_, _03624_);
  nor (_11318_, _11311_, _05253_);
  nor (_11319_, _11318_, _11310_);
  and (_11320_, _11319_, _07454_);
  and (_11321_, _05331_, \oc8051_golden_model_1.ACC [7]);
  nor (_11322_, _11321_, _11310_);
  nor (_11323_, _11322_, _04437_);
  nor (_11324_, _04436_, _11309_);
  or (_11325_, _11324_, _11323_);
  and (_11326_, _11325_, _04432_);
  and (_11327_, _06133_, _05331_);
  nor (_11328_, _11327_, _11310_);
  nor (_11329_, _11328_, _04432_);
  or (_11330_, _11329_, _11326_);
  and (_11331_, _11330_, _04457_);
  nor (_11332_, _11319_, _04457_);
  nor (_11333_, _11332_, _11331_);
  nor (_11334_, _11333_, _03530_);
  nor (_11335_, _11322_, _03531_);
  nor (_11336_, _11335_, _07454_);
  not (_11337_, _11336_);
  nor (_11338_, _11337_, _11334_);
  nor (_11339_, _11338_, _11320_);
  nor (_11340_, _11339_, _04082_);
  and (_11341_, _06114_, _05331_);
  nor (_11342_, _11310_, _04500_);
  not (_11343_, _11342_);
  nor (_11344_, _11343_, _11341_);
  or (_11345_, _11344_, _03224_);
  nor (_11346_, _11345_, _11340_);
  nor (_11347_, _06421_, _11311_);
  nor (_11348_, _11347_, _11310_);
  nor (_11349_, _11348_, _03521_);
  or (_11350_, _11349_, _03624_);
  nor (_11351_, _11350_, _11346_);
  nor (_11352_, _11351_, _11317_);
  or (_11353_, _11352_, _03623_);
  and (_11354_, _06436_, _05331_);
  or (_11355_, _11354_, _11310_);
  or (_11356_, _11355_, _04527_);
  and (_11357_, _11356_, _03745_);
  and (_11358_, _11357_, _11353_);
  and (_11359_, _06443_, _05331_);
  nor (_11360_, _11359_, _11310_);
  nor (_11361_, _11360_, _03745_);
  nor (_11362_, _11361_, _11358_);
  nor (_11363_, _11362_, _03611_);
  nor (_11364_, _11310_, _05358_);
  not (_11365_, _11364_);
  nor (_11366_, _11316_, _04523_);
  and (_11367_, _11366_, _11365_);
  nor (_11368_, _11367_, _11363_);
  nor (_11369_, _11368_, _03733_);
  nor (_11370_, _11322_, _03734_);
  and (_11371_, _11370_, _11365_);
  or (_11372_, _11371_, _11369_);
  and (_11373_, _11372_, _06453_);
  nor (_11374_, _06434_, _11311_);
  nor (_11375_, _11374_, _11310_);
  nor (_11376_, _11375_, _06453_);
  or (_11377_, _11376_, _11373_);
  and (_11378_, _11377_, _06458_);
  nor (_11379_, _11378_, _11314_);
  nor (_11380_, _11379_, _03767_);
  nor (_11381_, _11328_, _03948_);
  or (_11382_, _11381_, _03473_);
  nor (_11383_, _11382_, _11380_);
  and (_11384_, _05886_, _05331_);
  or (_11385_, _11310_, _03474_);
  nor (_11386_, _11385_, _11384_);
  nor (_11387_, _11386_, _11383_);
  or (_11388_, _11387_, _43193_);
  or (_11389_, _43189_, \oc8051_golden_model_1.TMOD [7]);
  and (_11390_, _11389_, _42003_);
  and (_40794_, _11390_, _11388_);
  not (_11391_, _03615_);
  nor (_11392_, _08882_, _08875_);
  not (_11393_, _02884_);
  and (_11394_, _05904_, _11393_);
  and (_11395_, _11394_, \oc8051_golden_model_1.PC [7]);
  and (_11396_, _11395_, _06857_);
  and (_11397_, _11396_, \oc8051_golden_model_1.PC [11]);
  and (_11398_, _11397_, \oc8051_golden_model_1.PC [12]);
  and (_11399_, _11398_, \oc8051_golden_model_1.PC [13]);
  and (_11400_, _11399_, \oc8051_golden_model_1.PC [14]);
  nor (_11401_, _11400_, \oc8051_golden_model_1.PC [15]);
  and (_11402_, _11400_, \oc8051_golden_model_1.PC [15]);
  nor (_11403_, _11402_, _11401_);
  nor (_11404_, _11403_, _11392_);
  not (_11405_, _03189_);
  nor (_11406_, _07920_, _04184_);
  nor (_11407_, _11406_, _11403_);
  and (_11408_, _08564_, _08599_);
  nor (_11409_, _11408_, _11403_);
  nor (_11410_, _08542_, _03739_);
  not (_11411_, _07923_);
  nand (_11412_, _03177_, _02954_);
  and (_11413_, _11412_, _11411_);
  nor (_11414_, _11413_, _11403_);
  and (_11415_, _08478_, _08472_);
  and (_11416_, _11415_, _08487_);
  nor (_11417_, _11416_, _11403_);
  and (_11418_, _06872_, _03224_);
  and (_11419_, _08191_, _08024_);
  nor (_11420_, _11419_, _11403_);
  and (_11421_, _03223_, _03558_);
  not (_11422_, _11421_);
  nor (_11423_, _08923_, _06933_);
  and (_11424_, _11423_, _11422_);
  not (_11425_, _11424_);
  and (_11426_, _11425_, _11403_);
  and (_11427_, _06888_, _03530_);
  and (_11428_, _03532_, _03202_);
  nor (_11429_, _11428_, _06888_);
  nor (_11430_, _09994_, _08121_);
  not (_11431_, _11430_);
  not (_11432_, _06872_);
  and (_11433_, _05722_, _05673_);
  and (_11434_, _06124_, _11433_);
  and (_11435_, _05468_, _05357_);
  and (_11436_, _11435_, _06120_);
  and (_11437_, _11436_, _11434_);
  and (_11438_, _11437_, _11432_);
  nand (_11439_, _11436_, _11434_);
  nor (_11440_, _06861_, \oc8051_golden_model_1.PC [14]);
  nor (_11441_, _11440_, _06862_);
  not (_11442_, _11441_);
  nor (_11443_, _11442_, _06226_);
  and (_11444_, _11442_, _06226_);
  nor (_11445_, _11444_, _11443_);
  not (_11446_, _11445_);
  nor (_11447_, _06860_, \oc8051_golden_model_1.PC [13]);
  nor (_11448_, _11447_, _06861_);
  and (_11449_, _11448_, _06227_);
  nor (_11450_, _11448_, _06227_);
  nor (_11451_, _06859_, \oc8051_golden_model_1.PC [12]);
  nor (_11452_, _11451_, _06860_);
  not (_11453_, _11452_);
  nor (_11454_, _11453_, _06226_);
  nor (_11455_, _06865_, \oc8051_golden_model_1.PC [10]);
  nor (_11456_, _11455_, _06858_);
  not (_11457_, _11456_);
  nor (_11458_, _11457_, _06226_);
  not (_11459_, _11458_);
  not (_11460_, \oc8051_golden_model_1.PC [11]);
  nor (_11461_, _06858_, _11460_);
  and (_11462_, _06858_, _11460_);
  or (_11463_, _11462_, _11461_);
  not (_11464_, _11463_);
  nor (_11465_, _11464_, _06226_);
  and (_11466_, _11464_, _06226_);
  nor (_11467_, _11466_, _11465_);
  and (_11468_, _11457_, _06226_);
  nor (_11469_, _11468_, _11458_);
  and (_11470_, _11469_, _11467_);
  nor (_11471_, _06864_, \oc8051_golden_model_1.PC [9]);
  nor (_11472_, _11471_, _06865_);
  not (_11473_, _11472_);
  nor (_11474_, _11473_, _06226_);
  and (_11475_, _11473_, _06226_);
  nor (_11476_, _11475_, _11474_);
  nor (_11477_, _06821_, _06226_);
  and (_11478_, _06821_, _06226_);
  and (_11479_, _06816_, _05903_);
  nor (_11480_, _11479_, \oc8051_golden_model_1.PC [6]);
  nor (_11481_, _11480_, _06817_);
  not (_11482_, _11481_);
  nor (_11483_, _11482_, _06262_);
  and (_11484_, _11482_, _06262_);
  nor (_11485_, _11484_, _11483_);
  not (_11486_, _11485_);
  and (_11487_, _06816_, \oc8051_golden_model_1.PC [4]);
  nor (_11488_, _11487_, \oc8051_golden_model_1.PC [5]);
  nor (_11489_, _11488_, _11479_);
  not (_11490_, _11489_);
  nor (_11491_, _11490_, _06294_);
  and (_11492_, _11490_, _06294_);
  nor (_11493_, _06816_, \oc8051_golden_model_1.PC [4]);
  nor (_11494_, _11493_, _11487_);
  not (_11495_, _11494_);
  nor (_11496_, _11495_, _06326_);
  nor (_11497_, _06815_, \oc8051_golden_model_1.PC [3]);
  nor (_11498_, _11497_, _06816_);
  not (_11499_, _11498_);
  nor (_11500_, _11499_, _03725_);
  and (_11501_, _11499_, _03725_);
  nor (_11502_, _02901_, \oc8051_golden_model_1.PC [2]);
  nor (_11503_, _11502_, _06815_);
  not (_11504_, _11503_);
  nor (_11505_, _11504_, _03855_);
  nor (_11506_, _04325_, _03313_);
  nor (_11507_, _04118_, \oc8051_golden_model_1.PC [0]);
  and (_11508_, _04325_, _03313_);
  nor (_11509_, _11508_, _11506_);
  and (_11510_, _11509_, _11507_);
  nor (_11511_, _11510_, _11506_);
  and (_11512_, _11504_, _03855_);
  nor (_11513_, _11512_, _11505_);
  not (_11514_, _11513_);
  nor (_11515_, _11514_, _11511_);
  nor (_11516_, _11515_, _11505_);
  nor (_11517_, _11516_, _11501_);
  nor (_11518_, _11517_, _11500_);
  and (_11519_, _11495_, _06326_);
  nor (_11520_, _11519_, _11496_);
  not (_11521_, _11520_);
  nor (_11522_, _11521_, _11518_);
  nor (_11523_, _11522_, _11496_);
  nor (_11524_, _11523_, _11492_);
  nor (_11525_, _11524_, _11491_);
  nor (_11526_, _11525_, _11486_);
  nor (_11527_, _11526_, _11483_);
  nor (_11528_, _11527_, _11478_);
  or (_11529_, _11528_, _11477_);
  nor (_11530_, _06818_, \oc8051_golden_model_1.PC [8]);
  nor (_11531_, _11530_, _06864_);
  not (_11532_, _11531_);
  nor (_11533_, _11532_, _06226_);
  and (_11534_, _11532_, _06226_);
  nor (_11535_, _11534_, _11533_);
  and (_11536_, _11535_, _11529_);
  and (_11537_, _11536_, _11476_);
  and (_11538_, _11537_, _11470_);
  nor (_11539_, _11533_, _11474_);
  not (_11540_, _11539_);
  and (_11541_, _11540_, _11470_);
  or (_11542_, _11541_, _11465_);
  nor (_11543_, _11542_, _11538_);
  and (_11544_, _11543_, _11459_);
  and (_11545_, _11453_, _06226_);
  nor (_11546_, _11545_, _11454_);
  not (_11547_, _11546_);
  nor (_11548_, _11547_, _11544_);
  nor (_11549_, _11548_, _11454_);
  nor (_11550_, _11549_, _11450_);
  nor (_11551_, _11550_, _11449_);
  nor (_11552_, _11551_, _11446_);
  nor (_11553_, _11552_, _11443_);
  and (_11554_, _11432_, _06226_);
  nor (_11555_, _11432_, _06226_);
  nor (_11556_, _11555_, _11554_);
  and (_11557_, _11556_, _11553_);
  nor (_11558_, _11556_, _11553_);
  nor (_11559_, _11558_, _11557_);
  and (_11560_, _11559_, _11439_);
  or (_11561_, _11560_, _04432_);
  or (_11562_, _11561_, _11438_);
  and (_11563_, _05985_, _05983_);
  and (_11564_, _04635_, _04429_);
  and (_11565_, _11564_, _05895_);
  and (_11566_, _11565_, _11563_);
  and (_11567_, _11566_, _06888_);
  nor (_11568_, _06877_, \oc8051_golden_model_1.PC [14]);
  nor (_11569_, _11568_, _06878_);
  and (_11570_, _11569_, _03409_);
  nor (_11571_, _11569_, _03409_);
  nor (_11572_, _11571_, _11570_);
  nor (_11573_, _06876_, \oc8051_golden_model_1.PC [13]);
  nor (_11574_, _11573_, _06877_);
  and (_11575_, _11574_, _03409_);
  nor (_11576_, _11574_, _03409_);
  nor (_11577_, _06875_, \oc8051_golden_model_1.PC [12]);
  nor (_11578_, _11577_, _06876_);
  and (_11579_, _11578_, _03409_);
  nor (_11580_, _06882_, \oc8051_golden_model_1.PC [11]);
  nor (_11581_, _11580_, _06883_);
  and (_11582_, _11581_, _03409_);
  nor (_11583_, _11581_, _03409_);
  nor (_11584_, _11583_, _11582_);
  nor (_11585_, _06881_, \oc8051_golden_model_1.PC [10]);
  nor (_11586_, _11585_, _06874_);
  and (_11587_, _11586_, _03409_);
  nor (_11588_, _11586_, _03409_);
  nor (_11589_, _11588_, _11587_);
  and (_11590_, _11589_, _11584_);
  nor (_11591_, _06880_, \oc8051_golden_model_1.PC [9]);
  nor (_11592_, _11591_, _06881_);
  and (_11593_, _11592_, _03409_);
  nor (_11594_, _11592_, _03409_);
  nor (_11595_, _11594_, _11593_);
  and (_11596_, _05908_, _03409_);
  nor (_11597_, _05908_, _03409_);
  and (_11598_, _05903_, _02863_);
  nor (_11599_, _11598_, \oc8051_golden_model_1.PC [6]);
  nor (_11600_, _11599_, _05905_);
  not (_11601_, _11600_);
  nor (_11602_, _11601_, _03511_);
  and (_11603_, _11601_, _03511_);
  nor (_11604_, _11603_, _11602_);
  not (_11605_, _11604_);
  and (_11606_, _02863_, \oc8051_golden_model_1.PC [4]);
  nor (_11607_, _11606_, \oc8051_golden_model_1.PC [5]);
  nor (_11608_, _11607_, _11598_);
  not (_11609_, _11608_);
  nor (_11610_, _11609_, _03811_);
  and (_11611_, _11609_, _03811_);
  nor (_11612_, _02863_, \oc8051_golden_model_1.PC [4]);
  nor (_11613_, _11612_, _11606_);
  not (_11614_, _11613_);
  nor (_11615_, _11614_, _04257_);
  nor (_11616_, _03440_, _03665_);
  and (_11617_, _03440_, _03665_);
  not (_11618_, _03294_);
  nor (_11619_, _03944_, _11618_);
  nor (_11620_, _04292_, \oc8051_golden_model_1.PC [1]);
  nor (_11621_, _03989_, _02897_);
  and (_11622_, _04292_, \oc8051_golden_model_1.PC [1]);
  nor (_11623_, _11622_, _11620_);
  and (_11624_, _11623_, _11621_);
  nor (_11625_, _11624_, _11620_);
  and (_11626_, _03944_, _11618_);
  nor (_11627_, _11626_, _11619_);
  not (_11628_, _11627_);
  nor (_11629_, _11628_, _11625_);
  nor (_11630_, _11629_, _11619_);
  nor (_11631_, _11630_, _11617_);
  nor (_11632_, _11631_, _11616_);
  and (_11633_, _11614_, _04257_);
  nor (_11634_, _11633_, _11615_);
  not (_11635_, _11634_);
  nor (_11636_, _11635_, _11632_);
  nor (_11637_, _11636_, _11615_);
  nor (_11638_, _11637_, _11611_);
  nor (_11639_, _11638_, _11610_);
  nor (_11640_, _11639_, _11605_);
  nor (_11641_, _11640_, _11602_);
  nor (_11642_, _11641_, _11597_);
  or (_11643_, _11642_, _11596_);
  nor (_11644_, _05906_, \oc8051_golden_model_1.PC [8]);
  nor (_11645_, _11644_, _06880_);
  and (_11646_, _11645_, _03409_);
  nor (_11647_, _11645_, _03409_);
  nor (_11648_, _11647_, _11646_);
  and (_11649_, _11648_, _11643_);
  and (_11650_, _11649_, _11595_);
  and (_11651_, _11650_, _11590_);
  nor (_11652_, _11646_, _11593_);
  not (_11653_, _11652_);
  and (_11654_, _11653_, _11590_);
  or (_11655_, _11654_, _11587_);
  or (_11656_, _11655_, _11651_);
  nor (_11657_, _11656_, _11582_);
  nor (_11658_, _11578_, _03409_);
  nor (_11659_, _11658_, _11579_);
  not (_11660_, _11659_);
  nor (_11661_, _11660_, _11657_);
  nor (_11662_, _11661_, _11579_);
  nor (_11663_, _11662_, _11576_);
  nor (_11664_, _11663_, _11575_);
  not (_11665_, _11664_);
  and (_11666_, _11665_, _11572_);
  nor (_11667_, _11666_, _11570_);
  nor (_11668_, _06888_, _03409_);
  and (_11669_, _06888_, _03409_);
  nor (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _11667_);
  nor (_11672_, _11670_, _11667_);
  nor (_11673_, _11672_, _11671_);
  nor (_11674_, _11566_, _11673_);
  or (_11675_, _11674_, _05997_);
  nor (_11676_, _11675_, _11567_);
  not (_11677_, _03209_);
  nand (_11678_, _11403_, _08118_);
  not (_11679_, _11403_);
  nor (_11680_, _08105_, _04007_);
  nor (_11681_, _04005_, _02954_);
  nor (_11682_, _11681_, _03203_);
  nor (_11683_, _11682_, _08108_);
  and (_11684_, _11683_, _11680_);
  or (_11685_, _11684_, _11679_);
  not (_11686_, _08118_);
  and (_11687_, _11680_, _11686_);
  not (_11688_, _11682_);
  and (_11689_, _03204_, \oc8051_golden_model_1.PC [15]);
  nor (_11690_, _08108_, _04436_);
  and (_11691_, _11690_, _11689_);
  and (_11692_, _11691_, _11688_);
  nand (_11693_, _11692_, _11687_);
  and (_11694_, _11693_, _11685_);
  or (_11695_, _11694_, _03536_);
  and (_11696_, _11695_, _11678_);
  or (_11697_, _11696_, _11677_);
  not (_11698_, _06888_);
  nand (_11699_, _10754_, _08101_);
  nor (_11700_, _11699_, _11677_);
  or (_11701_, _11700_, _11698_);
  and (_11702_, _11701_, _05997_);
  and (_11703_, _11702_, _11697_);
  not (_11704_, _11703_);
  nor (_11705_, _04012_, _03534_);
  nand (_11706_, _11705_, _11704_);
  or (_11707_, _11706_, _11676_);
  and (_11708_, _11707_, _11562_);
  or (_11709_, _11708_, _11431_);
  nand (_11710_, _11430_, _06008_);
  nand (_11711_, _11710_, _11403_);
  and (_11712_, _11711_, _11428_);
  and (_11713_, _11712_, _11709_);
  nor (_11714_, _11713_, _11429_);
  and (_11715_, _08098_, _08160_);
  not (_11716_, _11715_);
  nor (_11717_, _11716_, _11714_);
  nor (_11718_, _11715_, _11403_);
  nor (_11719_, _11718_, _03530_);
  not (_11720_, _11719_);
  nor (_11721_, _11720_, _11717_);
  nor (_11722_, _11721_, _11427_);
  nor (_11723_, _10008_, _08164_);
  not (_11724_, _11723_);
  nor (_11725_, _11724_, _11722_);
  nor (_11726_, _11723_, _11679_);
  not (_11727_, _03212_);
  nor (_11728_, _03464_, _11727_);
  and (_11729_, _11728_, _03466_);
  not (_11730_, _11729_);
  nor (_11731_, _11730_, _11726_);
  not (_11732_, _11731_);
  nor (_11733_, _11732_, _11725_);
  nor (_11734_, _11729_, _06888_);
  nor (_11735_, _11734_, _11733_);
  nor (_11736_, _11735_, _10021_);
  and (_11737_, _10055_, _06872_);
  nor (_11738_, _11559_, _10055_);
  or (_11739_, _11738_, _11737_);
  nor (_11740_, _11739_, _10017_);
  or (_11741_, _11740_, _10020_);
  nor (_11742_, _11741_, _11736_);
  nand (_11743_, _10115_, _10085_);
  not (_11744_, _11559_);
  and (_11745_, _11744_, _11743_);
  and (_11746_, _10116_, _06872_);
  nor (_11747_, _11746_, _11745_);
  nor (_11748_, _11747_, _10112_);
  or (_11749_, _11748_, _03547_);
  or (_11750_, _11749_, _11742_);
  and (_11751_, _09975_, _06872_);
  nor (_11752_, _11559_, _09975_);
  or (_11753_, _11752_, _03994_);
  or (_11754_, _11753_, _11751_);
  and (_11755_, _11754_, _10123_);
  and (_11756_, _11755_, _11750_);
  and (_11757_, _11403_, _10122_);
  not (_11758_, _11757_);
  nor (_11759_, _04481_, _04755_);
  and (_11760_, _11759_, _03523_);
  and (_11761_, _11760_, _03583_);
  and (_11762_, _11761_, _11758_);
  and (_11763_, _10163_, _11432_);
  not (_11764_, _10163_);
  and (_11765_, _11559_, _11764_);
  or (_11766_, _11765_, _10158_);
  or (_11767_, _11766_, _11763_);
  and (_11768_, _11767_, _11762_);
  not (_11769_, _11768_);
  nor (_11770_, _11769_, _11756_);
  nor (_11771_, _11761_, _06888_);
  nor (_11772_, _11771_, _11425_);
  not (_11773_, _11772_);
  nor (_11774_, _11773_, _11770_);
  or (_11775_, _11774_, _11426_);
  not (_11776_, _03214_);
  nor (_11777_, _03587_, _11776_);
  and (_11778_, _11777_, _10265_);
  nand (_11779_, _11778_, _11775_);
  not (_11780_, _11419_);
  nor (_11781_, _11778_, _11698_);
  nor (_11782_, _11781_, _11780_);
  and (_11783_, _11782_, _11779_);
  or (_11784_, _11783_, _11420_);
  nand (_11785_, _11784_, _08266_);
  nor (_11786_, _08266_, _06888_);
  nor (_11787_, _11786_, _03334_);
  nand (_11788_, _11787_, _11785_);
  and (_11789_, _11403_, _03334_);
  nor (_11790_, _03452_, _03219_);
  not (_11791_, _11790_);
  nor (_11792_, _11791_, _11789_);
  nand (_11793_, _11792_, _11788_);
  nor (_11794_, _11790_, _06888_);
  nor (_11795_, _11794_, _03621_);
  nand (_11796_, _11795_, _11793_);
  and (_11797_, _06903_, _04500_);
  and (_11798_, _06872_, _03621_);
  not (_11799_, _11798_);
  and (_11800_, _11799_, _11797_);
  nand (_11801_, _11800_, _11796_);
  nor (_11802_, _11797_, _06888_);
  nor (_11803_, _11802_, _03224_);
  and (_11804_, _11803_, _11801_);
  or (_11805_, _11804_, _11418_);
  nor (_11806_, _07468_, _03262_);
  nand (_11807_, _11806_, _11805_);
  nor (_11808_, _03517_, _03159_);
  not (_11809_, _11808_);
  nor (_11810_, _11806_, _11679_);
  nor (_11811_, _11810_, _11809_);
  and (_11812_, _11811_, _11807_);
  and (_11813_, _03444_, _03158_);
  not (_11814_, _11813_);
  and (_11815_, _11814_, _11808_);
  and (_11816_, _11814_, _06888_);
  nor (_11817_, _11816_, _11815_);
  or (_11818_, _11817_, _11812_);
  nor (_11819_, _11814_, _11673_);
  nor (_11820_, _11819_, _06193_);
  nand (_11821_, _11820_, _11818_);
  nor (_11822_, _06888_, _05916_);
  nor (_11823_, _11822_, _03624_);
  nand (_11824_, _11823_, _11821_);
  and (_11825_, _06872_, _03624_);
  nor (_11826_, _11825_, _08461_);
  nand (_11827_, _11826_, _11824_);
  and (_11828_, _03610_, _03167_);
  nor (_11829_, _08462_, _06888_);
  nor (_11830_, _11829_, _11828_);
  nand (_11831_, _11830_, _11827_);
  and (_11832_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_11833_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_11834_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11835_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11836_, _11835_, _11834_);
  not (_11837_, _11836_);
  and (_11838_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_11839_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  and (_11840_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11841_, _03250_, _03246_);
  nor (_11842_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11843_, _11842_, _11840_);
  not (_11844_, _11843_);
  nor (_11845_, _11844_, _11841_);
  nor (_11846_, _11845_, _11840_);
  nor (_11847_, _11846_, _11839_);
  nor (_11848_, _11847_, _11838_);
  nor (_11849_, _11848_, _11837_);
  nor (_11850_, _11849_, _11834_);
  nor (_11851_, _11850_, _11833_);
  or (_11852_, _11851_, _11832_);
  and (_11853_, _11852_, \oc8051_golden_model_1.DPH [0]);
  and (_11854_, _11853_, \oc8051_golden_model_1.DPH [1]);
  and (_11855_, _11854_, \oc8051_golden_model_1.DPH [2]);
  and (_11856_, _11855_, \oc8051_golden_model_1.DPH [3]);
  and (_11857_, _11856_, \oc8051_golden_model_1.DPH [4]);
  and (_11858_, _11857_, \oc8051_golden_model_1.DPH [5]);
  and (_11859_, _11858_, \oc8051_golden_model_1.DPH [6]);
  and (_11860_, _11859_, \oc8051_golden_model_1.DPH [7]);
  nor (_11861_, _11859_, \oc8051_golden_model_1.DPH [7]);
  nor (_11862_, _11861_, _11860_);
  and (_11863_, _11862_, _11828_);
  nor (_11864_, _03516_, _03168_);
  not (_11865_, _11864_);
  nor (_11866_, _11865_, _11863_);
  nand (_11867_, _11866_, _11831_);
  and (_11868_, _03444_, _03167_);
  nor (_11869_, _11864_, _06888_);
  nor (_11870_, _11869_, _11868_);
  nand (_11871_, _11870_, _11867_);
  not (_11872_, _11416_);
  and (_11873_, _08864_, _06888_);
  nor (_11874_, _11673_, _08864_);
  or (_11875_, _11874_, _11873_);
  and (_11876_, _11875_, _11868_);
  nor (_11877_, _11876_, _11872_);
  and (_11878_, _11877_, _11871_);
  or (_11879_, _11878_, _11417_);
  nand (_11880_, _11879_, _08493_);
  nor (_11881_, _08493_, _06888_);
  nor (_11882_, _11881_, _03623_);
  nand (_11883_, _11882_, _11880_);
  and (_11884_, _06872_, _03623_);
  nor (_11885_, _03744_, _03172_);
  not (_11886_, _11885_);
  nor (_11887_, _11886_, _11884_);
  nand (_11888_, _11887_, _11883_);
  and (_11889_, _03444_, _03171_);
  nor (_11890_, _11885_, _06888_);
  nor (_11891_, _11890_, _11889_);
  nand (_11892_, _11891_, _11888_);
  not (_11893_, _11889_);
  not (_11894_, _08864_);
  nand (_11895_, _11894_, _06888_);
  or (_11896_, _11673_, _11894_);
  and (_11897_, _11896_, _11895_);
  or (_11898_, _11897_, _11893_);
  nand (_11899_, _11898_, _11892_);
  not (_11900_, _03181_);
  nor (_11901_, _11681_, _11900_);
  not (_11902_, _11901_);
  nand (_11903_, _11902_, _11899_);
  nor (_11904_, _08517_, _03735_);
  not (_11905_, _11904_);
  and (_11906_, _11901_, _11403_);
  nor (_11907_, _11906_, _11905_);
  nand (_11908_, _11907_, _11903_);
  nor (_11909_, _11904_, _06888_);
  nor (_11910_, _11909_, _03611_);
  nand (_11911_, _11910_, _11908_);
  and (_11912_, _06872_, _03611_);
  nor (_11913_, _11912_, _10829_);
  and (_11914_, _11913_, _11911_);
  and (_11915_, _03444_, _03181_);
  nor (_11916_, _10828_, _06888_);
  or (_11917_, _11916_, _11915_);
  or (_11918_, _11917_, _11914_);
  not (_11919_, _11413_);
  and (_11920_, _06888_, \oc8051_golden_model_1.PSW [7]);
  nor (_11921_, _11673_, \oc8051_golden_model_1.PSW [7]);
  or (_11922_, _11921_, _11920_);
  and (_11923_, _11922_, _11915_);
  nor (_11924_, _11923_, _11919_);
  and (_11925_, _11924_, _11918_);
  or (_11926_, _11925_, _11414_);
  nand (_11927_, _11926_, _11410_);
  nor (_11928_, _11410_, _06888_);
  nor (_11929_, _11928_, _03618_);
  nand (_11930_, _11929_, _11927_);
  and (_11931_, _06872_, _03618_);
  nor (_11932_, _03741_, _03178_);
  not (_11933_, _11932_);
  nor (_11934_, _11933_, _11931_);
  nand (_11935_, _11934_, _11930_);
  and (_11936_, _03444_, _03177_);
  nor (_11937_, _11932_, _06888_);
  nor (_11938_, _11937_, _11936_);
  nand (_11939_, _11938_, _11935_);
  not (_11940_, _11408_);
  and (_11941_, _11673_, \oc8051_golden_model_1.PSW [7]);
  not (_11942_, _11936_);
  nor (_11943_, _06888_, \oc8051_golden_model_1.PSW [7]);
  nor (_11944_, _11943_, _11942_);
  not (_11945_, _11944_);
  nor (_11946_, _11945_, _11941_);
  nor (_11947_, _11946_, _11940_);
  and (_11948_, _11947_, _11939_);
  or (_11949_, _11948_, _11409_);
  nand (_11950_, _11949_, _08628_);
  nor (_11951_, _08628_, _06888_);
  nor (_11952_, _11951_, _08707_);
  nand (_11953_, _11952_, _11950_);
  and (_11954_, _11403_, _08707_);
  nor (_11955_, _11954_, _03752_);
  and (_11956_, _11955_, _11953_);
  and (_11957_, _05253_, _03752_);
  or (_11958_, _11957_, _11956_);
  nand (_11959_, _11958_, _04803_);
  nor (_11960_, _06888_, _04803_);
  nor (_11961_, _11960_, _03617_);
  nand (_11962_, _11961_, _11959_);
  not (_11963_, _11406_);
  and (_11964_, _11559_, _09953_);
  nor (_11965_, _09953_, _06872_);
  or (_11966_, _11965_, _03814_);
  nor (_11967_, _11966_, _11964_);
  nor (_11968_, _11967_, _11963_);
  and (_11969_, _11968_, _11962_);
  or (_11970_, _11969_, _11407_);
  nand (_11971_, _11970_, _08784_);
  nor (_11972_, _08784_, _06888_);
  nor (_11973_, _11972_, _08815_);
  nand (_11974_, _11973_, _11971_);
  and (_11975_, _11403_, _08815_);
  nor (_11976_, _11975_, _03475_);
  and (_11977_, _11976_, _11974_);
  and (_11978_, _05253_, _03475_);
  or (_11979_, _11978_, _11977_);
  nand (_11980_, _11979_, _11405_);
  nor (_11981_, _06888_, _11405_);
  nor (_11982_, _11981_, _03644_);
  nand (_11983_, _11982_, _11980_);
  nor (_11984_, _11744_, _09953_);
  and (_11985_, _09953_, _11432_);
  nor (_11986_, _11985_, _11984_);
  and (_11987_, _11986_, _03644_);
  nor (_11988_, _06899_, _05139_);
  nor (_11989_, _11988_, _05141_);
  and (_11990_, _11989_, _05137_);
  and (_11991_, _11990_, _06480_);
  not (_11992_, _11991_);
  nor (_11993_, _11992_, _11987_);
  nand (_11994_, _11993_, _11983_);
  nor (_11995_, _11991_, _11403_);
  nor (_11996_, _11995_, _03767_);
  nand (_11997_, _11996_, _11994_);
  nor (_11998_, _08858_, _08853_);
  not (_11999_, _11998_);
  and (_12000_, _06888_, _03767_);
  nor (_12001_, _12000_, _11999_);
  nand (_12002_, _12001_, _11997_);
  nor (_12003_, _11403_, _11998_);
  nor (_12004_, _12003_, _03645_);
  nand (_12005_, _12004_, _12002_);
  and (_12006_, _03645_, _03409_);
  nor (_12007_, _12006_, _03196_);
  nand (_12008_, _12007_, _12005_);
  not (_12009_, _03196_);
  nor (_12010_, _06888_, _12009_);
  nor (_12011_, _12010_, _03445_);
  nand (_12012_, _12011_, _12008_);
  and (_12013_, _11986_, _03445_);
  and (_12014_, _03193_, _02954_);
  nor (_12015_, _12014_, _04215_);
  not (_12016_, _12015_);
  nor (_12017_, _12016_, _12013_);
  nand (_12018_, _12017_, _12012_);
  nor (_12019_, _12015_, _11403_);
  nor (_12020_, _12019_, _03473_);
  nand (_12021_, _12020_, _12018_);
  not (_12022_, _11392_);
  and (_12023_, _06888_, _03473_);
  nor (_12024_, _12023_, _12022_);
  and (_12025_, _12024_, _12021_);
  or (_12026_, _12025_, _11404_);
  nand (_12027_, _12026_, _11391_);
  nor (_12028_, _11391_, _03409_);
  nor (_12029_, _12028_, _03194_);
  nand (_12030_, _12029_, _12027_);
  and (_12031_, _03444_, _03193_);
  and (_12032_, _06888_, _03194_);
  nor (_12033_, _12032_, _12031_);
  and (_12034_, _12033_, _12030_);
  not (_12035_, _12031_);
  nor (_12036_, _12035_, _11403_);
  nor (_12037_, _12036_, _12034_);
  or (_12038_, _12037_, _43193_);
  or (_12039_, _43189_, \oc8051_golden_model_1.PC [15]);
  and (_12040_, _12039_, _42003_);
  and (_40796_, _12040_, _12038_);
  and (_12041_, _43193_, \oc8051_golden_model_1.P0INREG [7]);
  or (_12042_, _12041_, _01087_);
  and (_40797_, _12042_, _42003_);
  and (_12043_, _43193_, \oc8051_golden_model_1.P1INREG [7]);
  or (_12044_, _12043_, _01008_);
  and (_40798_, _12044_, _42003_);
  and (_12045_, _43193_, \oc8051_golden_model_1.P2INREG [7]);
  or (_12046_, _12045_, _00917_);
  and (_40799_, _12046_, _42003_);
  and (_12047_, _43193_, \oc8051_golden_model_1.P3INREG [7]);
  or (_12048_, _12047_, _01187_);
  and (_40800_, _12048_, _42003_);
  nor (_12049_, _05185_, _04744_);
  nor (_12050_, _12049_, _05186_);
  nor (_12051_, _05185_, _05161_);
  nor (_12052_, _12051_, _05189_);
  and (_12053_, _12052_, _05184_);
  nand (_12054_, _12053_, _12050_);
  nand (_12055_, _03196_, _02897_);
  not (_12056_, _06459_);
  nor (_12057_, _05722_, _06350_);
  nor (_12058_, _12057_, _06460_);
  and (_12059_, _05722_, _06350_);
  and (_12060_, _12059_, _04524_);
  or (_12061_, _04499_, _04429_);
  nand (_12062_, _08380_, _03584_);
  nor (_12063_, _10214_, _05273_);
  or (_12064_, _12063_, _05964_);
  nor (_12065_, _05722_, _04434_);
  or (_12066_, _05997_, _04462_);
  nor (_12067_, _03204_, _02897_);
  and (_12068_, _03204_, \oc8051_golden_model_1.ACC [0]);
  nor (_12069_, _12068_, _12067_);
  and (_12070_, _12069_, _05997_);
  nor (_12071_, _12070_, _04433_);
  and (_12072_, _12071_, _12066_);
  or (_12073_, _12072_, _12065_);
  and (_12074_, _12073_, _05978_);
  nand (_12075_, _10214_, _09849_);
  and (_12076_, _12075_, _03472_);
  or (_12077_, _12076_, _05977_);
  or (_12078_, _12077_, _12074_);
  nor (_12079_, _03202_, \oc8051_golden_model_1.PC [0]);
  nor (_12080_, _12079_, _04458_);
  and (_12081_, _12080_, _12078_);
  and (_12082_, _04458_, _04429_);
  or (_12083_, _12082_, _12081_);
  or (_12084_, _12083_, _04466_);
  and (_12085_, _12084_, _12064_);
  or (_12086_, _12085_, _03464_);
  nand (_12087_, _08380_, _03464_);
  and (_12088_, _12087_, _03462_);
  and (_12089_, _12088_, _12086_);
  nand (_12090_, _12075_, _03461_);
  nor (_12091_, _12090_, _10215_);
  or (_12092_, _12091_, _12089_);
  and (_12093_, _12092_, _03207_);
  or (_12094_, _03207_, _02897_);
  nand (_12095_, _03583_, _12094_);
  or (_12096_, _12095_, _12093_);
  and (_12097_, _12096_, _12062_);
  or (_12098_, _12097_, _04481_);
  and (_12099_, _06617_, _04493_);
  nand (_12100_, _08379_, _04481_);
  or (_12101_, _12100_, _12099_);
  and (_12102_, _12101_, _12098_);
  or (_12103_, _12102_, _04480_);
  nor (_12104_, _09872_, _05273_);
  and (_12105_, _05273_, \oc8051_golden_model_1.PSW [7]);
  nor (_12106_, _12105_, _12104_);
  nand (_12107_, _12106_, _04480_);
  and (_12108_, _12107_, _05919_);
  and (_12109_, _12108_, _12103_);
  nand (_12110_, _03219_, \oc8051_golden_model_1.PC [0]);
  nand (_12111_, _04499_, _12110_);
  or (_12112_, _12111_, _12109_);
  and (_12113_, _12112_, _12061_);
  or (_12114_, _12113_, _04501_);
  or (_12115_, _06617_, _06189_);
  and (_12116_, _12115_, _04754_);
  and (_12117_, _12116_, _12114_);
  and (_12118_, _06226_, _04429_);
  and (_12119_, _06407_, \oc8051_golden_model_1.DPH [0]);
  and (_12120_, _06414_, \oc8051_golden_model_1.TH1 [0]);
  nor (_12121_, _12120_, _12119_);
  and (_12122_, _06329_, \oc8051_golden_model_1.P2INREG [0]);
  not (_12123_, _12122_);
  and (_12124_, _06334_, \oc8051_golden_model_1.P0INREG [0]);
  not (_12125_, _12124_);
  and (_12126_, _06340_, \oc8051_golden_model_1.P1INREG [0]);
  and (_12127_, _06344_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_12128_, _12127_, _12126_);
  and (_12129_, _12128_, _12125_);
  and (_12130_, _12129_, _12123_);
  and (_12131_, _12130_, _12121_);
  and (_12132_, _06378_, \oc8051_golden_model_1.IE [0]);
  not (_12133_, _12132_);
  and (_12134_, _06381_, \oc8051_golden_model_1.SCON [0]);
  and (_12135_, _06384_, \oc8051_golden_model_1.SBUF [0]);
  nor (_12136_, _12135_, _12134_);
  and (_12137_, _12136_, _12133_);
  and (_12138_, _06365_, \oc8051_golden_model_1.PSW [0]);
  and (_12139_, _06367_, \oc8051_golden_model_1.ACC [0]);
  nor (_12140_, _12139_, _12138_);
  and (_12141_, _06370_, \oc8051_golden_model_1.B [0]);
  and (_12142_, _06374_, \oc8051_golden_model_1.IP [0]);
  nor (_12143_, _12142_, _12141_);
  and (_12144_, _12143_, _12140_);
  and (_12145_, _12144_, _12137_);
  and (_12146_, _12145_, _12131_);
  and (_12147_, _06392_, \oc8051_golden_model_1.TH0 [0]);
  and (_12148_, _06396_, \oc8051_golden_model_1.TL1 [0]);
  nor (_12149_, _12148_, _12147_);
  and (_12150_, _06401_, \oc8051_golden_model_1.PCON [0]);
  and (_12151_, _06403_, \oc8051_golden_model_1.TCON [0]);
  nor (_12152_, _12151_, _12150_);
  and (_12153_, _12152_, _12149_);
  and (_12154_, _06352_, \oc8051_golden_model_1.SP [0]);
  and (_12155_, _06412_, \oc8051_golden_model_1.DPL [0]);
  nor (_12156_, _12155_, _12154_);
  and (_12157_, _06359_, \oc8051_golden_model_1.TL0 [0]);
  and (_12158_, _06409_, \oc8051_golden_model_1.TMOD [0]);
  nor (_12159_, _12158_, _12157_);
  and (_12160_, _12159_, _12156_);
  and (_12161_, _12160_, _12153_);
  and (_12162_, _12161_, _12146_);
  not (_12163_, _12162_);
  nor (_12164_, _12163_, _12118_);
  nor (_12165_, _12164_, _06195_);
  or (_12166_, _12165_, _06193_);
  or (_12167_, _12166_, _12117_);
  and (_12168_, _06193_, _03989_);
  nor (_12169_, _12168_, _04510_);
  and (_12170_, _12169_, _12167_);
  nor (_12171_, _06426_, _04118_);
  or (_12172_, _12171_, _03168_);
  or (_12173_, _12172_, _12170_);
  and (_12174_, _03168_, _02897_);
  nor (_12175_, _12174_, _04528_);
  and (_12176_, _12175_, _12173_);
  nor (_12177_, _12059_, _12057_);
  nor (_12178_, _12177_, _04526_);
  nor (_12179_, _12178_, _04529_);
  or (_12180_, _12179_, _12176_);
  nor (_12181_, _05722_, \oc8051_golden_model_1.ACC [0]);
  and (_12182_, _05722_, \oc8051_golden_model_1.ACC [0]);
  nor (_12183_, _12182_, _12181_);
  or (_12184_, _12183_, _06432_);
  and (_12185_, _12184_, _04525_);
  and (_12186_, _12185_, _12180_);
  or (_12187_, _12186_, _12060_);
  and (_12188_, _12187_, _04522_);
  and (_12189_, _12182_, _04521_);
  or (_12190_, _12189_, _03182_);
  or (_12191_, _12190_, _12188_);
  and (_12192_, _03182_, _02897_);
  nor (_12193_, _12192_, _06454_);
  and (_12194_, _12193_, _12191_);
  or (_12195_, _12194_, _12058_);
  and (_12196_, _12195_, _12056_);
  nor (_12197_, _12181_, _12056_);
  or (_12198_, _12197_, _03191_);
  or (_12199_, _12198_, _12196_);
  nand (_12200_, _03191_, _02897_);
  and (_12201_, _12200_, _11990_);
  and (_12202_, _12201_, _12199_);
  nor (_12203_, _11990_, _04429_);
  or (_12204_, _12203_, _12202_);
  and (_12205_, _12204_, _06480_);
  nor (_12206_, _06617_, _06480_);
  or (_12207_, _12206_, _04546_);
  or (_12208_, _12207_, _12205_);
  nand (_12209_, _05722_, _04546_);
  and (_12210_, _12209_, _06855_);
  and (_12211_, _12210_, _12208_);
  and (_12212_, _03645_, _02897_);
  or (_12213_, _12212_, _03196_);
  or (_12214_, _12213_, _12211_);
  and (_12215_, _12214_, _12055_);
  or (_12216_, _12215_, _03448_);
  not (_12217_, _12014_);
  or (_12218_, _12104_, _03449_);
  and (_12219_, _12218_, _12217_);
  and (_12220_, _12219_, _12216_);
  or (_12221_, _04462_, _04215_);
  and (_12222_, _12221_, _12016_);
  or (_12223_, _12222_, _12220_);
  nand (_12224_, _06617_, _04215_);
  and (_12225_, _12224_, _12223_);
  or (_12226_, _12225_, _04559_);
  nand (_12227_, _05722_, _04559_);
  and (_12228_, _12227_, _05184_);
  and (_12229_, _12228_, _12226_);
  or (_12230_, _12229_, _12054_);
  and (_12231_, _05177_, _05169_);
  nor (_12232_, _12231_, _05178_);
  and (_12233_, _05177_, _04570_);
  and (_12234_, _12233_, _12232_);
  and (_12235_, _12054_, _03958_);
  nor (_12236_, _12235_, _12234_);
  and (_12237_, _12236_, _12230_);
  nand (_12238_, _11532_, _03645_);
  or (_12239_, _11645_, _03645_);
  and (_12240_, _12239_, _12238_);
  and (_12241_, _12240_, _05177_);
  and (_12242_, _12241_, _12234_);
  or (_40839_, _12242_, _12237_);
  nor (_12243_, _05176_, _04745_);
  and (_12244_, _12243_, _05169_);
  and (_12245_, _12243_, _05172_);
  or (_12246_, _12245_, _12244_);
  nand (_12247_, _12243_, _04570_);
  or (_12248_, _12247_, _12246_);
  nand (_12249_, _12054_, _04578_);
  and (_12250_, _12249_, _12248_);
  nor (_12251_, _05984_, _05890_);
  and (_12252_, _12251_, _12014_);
  and (_12253_, _03191_, _02860_);
  or (_12254_, _04636_, _04499_);
  nand (_12255_, _08364_, _03584_);
  nor (_12256_, _10190_, _05265_);
  or (_12257_, _12256_, _05964_);
  nand (_12258_, _12251_, _05998_);
  nor (_12259_, _03204_, \oc8051_golden_model_1.PC [1]);
  and (_12260_, _03204_, \oc8051_golden_model_1.ACC [1]);
  nor (_12261_, _12260_, _12259_);
  nand (_12262_, _12261_, _05997_);
  and (_12263_, _12262_, _12258_);
  or (_12264_, _12263_, _04433_);
  nor (_12265_, _06123_, _05723_);
  nand (_12266_, _12265_, _04433_);
  and (_12267_, _12266_, _12264_);
  or (_12268_, _12267_, _03472_);
  nand (_12269_, _10190_, _09794_);
  or (_12270_, _12269_, _05978_);
  and (_12271_, _12270_, _12268_);
  or (_12272_, _12271_, _05977_);
  nor (_12273_, _03202_, _02860_);
  nor (_12274_, _12273_, _04458_);
  and (_12275_, _12274_, _12272_);
  nor (_12276_, _04635_, _04896_);
  or (_12277_, _12276_, _04466_);
  or (_12278_, _12277_, _12275_);
  and (_12279_, _12278_, _12257_);
  or (_12280_, _12279_, _03464_);
  nand (_12281_, _08364_, _03464_);
  and (_12282_, _12281_, _03462_);
  and (_12283_, _12282_, _12280_);
  not (_12284_, _10191_);
  and (_12285_, _12269_, _12284_);
  and (_12286_, _12285_, _03461_);
  or (_12287_, _12286_, _12283_);
  and (_12288_, _12287_, _03207_);
  or (_12289_, _03207_, \oc8051_golden_model_1.PC [1]);
  nand (_12290_, _03583_, _12289_);
  or (_12291_, _12290_, _12288_);
  and (_12292_, _12291_, _12255_);
  or (_12293_, _12292_, _04481_);
  and (_12294_, _06572_, _04493_);
  nand (_12295_, _08363_, _04481_);
  or (_12296_, _12295_, _12294_);
  and (_12297_, _12296_, _12293_);
  or (_12298_, _12297_, _04480_);
  nor (_12299_, _09817_, _05265_);
  and (_12300_, _05265_, \oc8051_golden_model_1.PSW [7]);
  nor (_12301_, _12300_, _12299_);
  nand (_12302_, _12301_, _04480_);
  and (_12303_, _12302_, _05919_);
  and (_12304_, _12303_, _12298_);
  nand (_12305_, _03219_, _02860_);
  nand (_12306_, _04499_, _12305_);
  or (_12307_, _12306_, _12304_);
  and (_12308_, _12307_, _12254_);
  or (_12309_, _12308_, _04501_);
  nand (_12310_, _04490_, _04005_);
  or (_12311_, _06572_, _12310_);
  and (_12312_, _12311_, _06195_);
  and (_12313_, _12312_, _12309_);
  nor (_12314_, _06227_, _04635_);
  and (_12315_, _06329_, \oc8051_golden_model_1.P2INREG [1]);
  not (_12316_, _12315_);
  and (_12317_, _06334_, \oc8051_golden_model_1.P0INREG [1]);
  not (_12318_, _12317_);
  and (_12319_, _06340_, \oc8051_golden_model_1.P1INREG [1]);
  and (_12320_, _06344_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_12321_, _12320_, _12319_);
  and (_12322_, _12321_, _12318_);
  and (_12323_, _12322_, _12316_);
  and (_12324_, _06352_, \oc8051_golden_model_1.SP [1]);
  and (_12325_, _06359_, \oc8051_golden_model_1.TL0 [1]);
  nor (_12326_, _12325_, _12324_);
  and (_12327_, _12326_, _12323_);
  and (_12328_, _06378_, \oc8051_golden_model_1.IE [1]);
  not (_12329_, _12328_);
  and (_12330_, _06381_, \oc8051_golden_model_1.SCON [1]);
  and (_12331_, _06384_, \oc8051_golden_model_1.SBUF [1]);
  nor (_12332_, _12331_, _12330_);
  and (_12333_, _12332_, _12329_);
  and (_12334_, _06365_, \oc8051_golden_model_1.PSW [1]);
  and (_12335_, _06370_, \oc8051_golden_model_1.B [1]);
  nor (_12336_, _12335_, _12334_);
  and (_12337_, _06367_, \oc8051_golden_model_1.ACC [1]);
  and (_12338_, _06374_, \oc8051_golden_model_1.IP [1]);
  nor (_12339_, _12338_, _12337_);
  and (_12340_, _12339_, _12336_);
  and (_12341_, _12340_, _12333_);
  and (_12342_, _12341_, _12327_);
  and (_12343_, _06392_, \oc8051_golden_model_1.TH0 [1]);
  and (_12344_, _06396_, \oc8051_golden_model_1.TL1 [1]);
  nor (_12345_, _12344_, _12343_);
  and (_12346_, _06401_, \oc8051_golden_model_1.PCON [1]);
  and (_12347_, _06403_, \oc8051_golden_model_1.TCON [1]);
  nor (_12348_, _12347_, _12346_);
  and (_12349_, _12348_, _12345_);
  and (_12350_, _06407_, \oc8051_golden_model_1.DPH [1]);
  and (_12351_, _06409_, \oc8051_golden_model_1.TMOD [1]);
  nor (_12352_, _12351_, _12350_);
  and (_12353_, _06412_, \oc8051_golden_model_1.DPL [1]);
  and (_12354_, _06414_, \oc8051_golden_model_1.TH1 [1]);
  nor (_12355_, _12354_, _12353_);
  and (_12356_, _12355_, _12352_);
  and (_12357_, _12356_, _12349_);
  and (_12358_, _12357_, _12342_);
  not (_12359_, _12358_);
  nor (_12360_, _12359_, _12314_);
  nor (_12361_, _12360_, _06195_);
  or (_12362_, _12361_, _06193_);
  or (_12363_, _12362_, _12313_);
  and (_12364_, _06193_, _04292_);
  nor (_12365_, _12364_, _04510_);
  and (_12366_, _12365_, _12363_);
  nor (_12367_, _06426_, _04325_);
  or (_12368_, _12367_, _03168_);
  or (_12369_, _12368_, _12366_);
  and (_12370_, _03168_, \oc8051_golden_model_1.PC [1]);
  nor (_12371_, _12370_, _04528_);
  and (_12372_, _12371_, _12369_);
  and (_12373_, _05673_, _04325_);
  nor (_12374_, _05673_, _04325_);
  nor (_12375_, _12374_, _12373_);
  and (_12376_, _12375_, _04528_);
  or (_12377_, _12376_, _12372_);
  and (_12378_, _12377_, _06432_);
  nor (_12379_, _05673_, _03269_);
  and (_12380_, _05673_, _03269_);
  nor (_12381_, _12380_, _12379_);
  and (_12382_, _12381_, _04526_);
  or (_12383_, _12382_, _12378_);
  and (_12384_, _12383_, _04525_);
  and (_12385_, _12374_, _04524_);
  or (_12386_, _12385_, _12384_);
  and (_12387_, _12386_, _04522_);
  and (_12388_, _12379_, _04521_);
  or (_12389_, _12388_, _03182_);
  or (_12390_, _12389_, _12387_);
  and (_12391_, _03182_, \oc8051_golden_model_1.PC [1]);
  nor (_12392_, _12391_, _06454_);
  and (_12393_, _12392_, _12390_);
  nor (_12394_, _12373_, _06460_);
  or (_12395_, _12394_, _06459_);
  or (_12396_, _12395_, _12393_);
  nand (_12397_, _12380_, _06459_);
  and (_12398_, _12397_, _04803_);
  and (_12399_, _12398_, _12396_);
  nor (_12400_, _12399_, _12253_);
  nor (_12401_, _12400_, _03861_);
  and (_12402_, _03565_, _03195_);
  nand (_12403_, _12251_, _03017_);
  and (_12404_, _12403_, _12402_);
  or (_12405_, _12404_, _05144_);
  or (_12406_, _12405_, _12401_);
  nand (_12407_, _05143_, _04718_);
  nand (_12408_, _12407_, _12251_);
  and (_12409_, _12408_, _06480_);
  and (_12410_, _12409_, _12406_);
  nor (_12411_, _06839_, _06618_);
  nor (_12412_, _12411_, _06480_);
  or (_12413_, _12412_, _12410_);
  and (_12414_, _12413_, _06479_);
  nor (_12415_, _12265_, _06479_);
  or (_12416_, _12415_, _03645_);
  or (_12417_, _12416_, _12414_);
  nand (_12418_, _03645_, _03313_);
  and (_12419_, _12418_, _12009_);
  and (_12420_, _12419_, _12417_);
  and (_12421_, _03196_, _02860_);
  or (_12422_, _03448_, _12421_);
  or (_12423_, _12422_, _12420_);
  or (_12424_, _12299_, _03449_);
  and (_12425_, _12424_, _12217_);
  and (_12426_, _12425_, _12423_);
  or (_12427_, _12426_, _12252_);
  and (_12428_, _12427_, _06838_);
  and (_12429_, _12411_, _04215_);
  or (_12430_, _12429_, _04559_);
  or (_12431_, _12430_, _12428_);
  or (_12432_, _12265_, _04746_);
  and (_12433_, _12432_, _05184_);
  and (_12434_, _12433_, _12431_);
  or (_12435_, _12434_, _12054_);
  and (_12436_, _12435_, _12250_);
  nand (_12437_, _11473_, _03645_);
  or (_12438_, _11592_, _03645_);
  and (_12439_, _12438_, _12437_);
  and (_12440_, _12439_, _05177_);
  and (_12441_, _12440_, _12234_);
  or (_40840_, _12441_, _12436_);
  nand (_12442_, _12054_, _05017_);
  and (_12443_, _12442_, _12248_);
  or (_12444_, _05890_, _05074_);
  nor (_12445_, _12217_, _08222_);
  and (_12446_, _12445_, _12444_);
  not (_12447_, _06710_);
  and (_12448_, _06618_, _12447_);
  nor (_12449_, _06618_, _12447_);
  or (_12450_, _12449_, _12448_);
  and (_12451_, _12450_, _04201_);
  and (_12452_, _05984_, _05073_);
  nor (_12453_, _05984_, _05073_);
  or (_12454_, _12453_, _12452_);
  or (_12455_, _12454_, _04721_);
  and (_12456_, _03629_, _03195_);
  or (_12457_, _12454_, _06471_);
  nor (_12458_, _05771_, _03855_);
  and (_12459_, _12458_, _04524_);
  nor (_12460_, _10179_, _05326_);
  or (_12461_, _12460_, _05964_);
  nand (_12462_, _10179_, _09770_);
  or (_12463_, _12462_, _05978_);
  and (_12464_, _05771_, _05673_);
  and (_12465_, _12464_, _06121_);
  nor (_12466_, _06123_, _05771_);
  nor (_12467_, _12466_, _12465_);
  nor (_12468_, _12467_, _04434_);
  or (_12469_, _12454_, _05997_);
  nor (_12470_, _11618_, _03204_);
  and (_12471_, _03204_, \oc8051_golden_model_1.ACC [2]);
  nor (_12472_, _12471_, _12470_);
  and (_12473_, _12472_, _05997_);
  nor (_12474_, _12473_, _04433_);
  and (_12475_, _12474_, _12469_);
  or (_12476_, _12475_, _03472_);
  or (_12477_, _12476_, _12468_);
  and (_12478_, _12477_, _12463_);
  or (_12479_, _12478_, _05977_);
  nor (_12480_, _03294_, _03202_);
  nor (_12481_, _12480_, _04458_);
  and (_12482_, _12481_, _12479_);
  nor (_12483_, _05073_, _04896_);
  or (_12484_, _12483_, _04466_);
  or (_12485_, _12484_, _12482_);
  and (_12486_, _12485_, _12461_);
  or (_12487_, _12486_, _03464_);
  nand (_12488_, _08350_, _03464_);
  and (_12489_, _12488_, _03462_);
  and (_12490_, _12489_, _12487_);
  not (_12491_, _10180_);
  and (_12492_, _12462_, _12491_);
  and (_12493_, _12492_, _03461_);
  or (_12494_, _12493_, _12490_);
  and (_12495_, _12494_, _03207_);
  or (_12496_, _11618_, _03207_);
  nand (_12497_, _03583_, _12496_);
  or (_12498_, _12497_, _12495_);
  nand (_12499_, _08350_, _03584_);
  and (_12500_, _12499_, _12498_);
  or (_12501_, _12500_, _04481_);
  and (_12502_, _06710_, _04493_);
  nand (_12503_, _08349_, _04481_);
  or (_12504_, _12503_, _12502_);
  and (_12505_, _12504_, _12501_);
  or (_12506_, _12505_, _04480_);
  nor (_12507_, _09792_, _05326_);
  and (_12508_, _05326_, \oc8051_golden_model_1.PSW [7]);
  nor (_12509_, _12508_, _12507_);
  nand (_12510_, _12509_, _04480_);
  and (_12511_, _12510_, _05919_);
  and (_12512_, _12511_, _12506_);
  nand (_12513_, _03294_, _03219_);
  nand (_12514_, _04499_, _12513_);
  or (_12515_, _12514_, _12512_);
  or (_12516_, _05074_, _04499_);
  and (_12517_, _12516_, _12515_);
  or (_12518_, _12517_, _04501_);
  or (_12519_, _06710_, _06189_);
  and (_12520_, _12519_, _04754_);
  and (_12521_, _12520_, _12518_);
  nor (_12522_, _06227_, _05073_);
  and (_12523_, _06329_, \oc8051_golden_model_1.P2INREG [2]);
  not (_12524_, _12523_);
  and (_12525_, _06334_, \oc8051_golden_model_1.P0INREG [2]);
  not (_12526_, _12525_);
  and (_12527_, _06340_, \oc8051_golden_model_1.P1INREG [2]);
  and (_12528_, _06344_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_12529_, _12528_, _12527_);
  and (_12530_, _12529_, _12526_);
  and (_12531_, _12530_, _12524_);
  and (_12532_, _06359_, \oc8051_golden_model_1.TL0 [2]);
  and (_12533_, _06409_, \oc8051_golden_model_1.TMOD [2]);
  nor (_12534_, _12533_, _12532_);
  and (_12535_, _12534_, _12531_);
  and (_12536_, _06378_, \oc8051_golden_model_1.IE [2]);
  not (_12537_, _12536_);
  and (_12538_, _06381_, \oc8051_golden_model_1.SCON [2]);
  and (_12539_, _06384_, \oc8051_golden_model_1.SBUF [2]);
  nor (_12540_, _12539_, _12538_);
  and (_12541_, _12540_, _12537_);
  and (_12542_, _06407_, \oc8051_golden_model_1.DPH [2]);
  and (_12543_, _06414_, \oc8051_golden_model_1.TH1 [2]);
  nor (_12544_, _12543_, _12542_);
  and (_12545_, _12544_, _12541_);
  and (_12546_, _12545_, _12535_);
  and (_12547_, _06392_, \oc8051_golden_model_1.TH0 [2]);
  and (_12548_, _06396_, \oc8051_golden_model_1.TL1 [2]);
  nor (_12549_, _12548_, _12547_);
  and (_12550_, _06401_, \oc8051_golden_model_1.PCON [2]);
  and (_12551_, _06403_, \oc8051_golden_model_1.TCON [2]);
  nor (_12552_, _12551_, _12550_);
  and (_12553_, _12552_, _12549_);
  and (_12554_, _06370_, \oc8051_golden_model_1.B [2]);
  and (_12555_, _06374_, \oc8051_golden_model_1.IP [2]);
  nor (_12556_, _12555_, _12554_);
  and (_12557_, _06365_, \oc8051_golden_model_1.PSW [2]);
  and (_12558_, _06367_, \oc8051_golden_model_1.ACC [2]);
  nor (_12559_, _12558_, _12557_);
  and (_12560_, _12559_, _12556_);
  and (_12561_, _06352_, \oc8051_golden_model_1.SP [2]);
  and (_12562_, _06412_, \oc8051_golden_model_1.DPL [2]);
  nor (_12563_, _12562_, _12561_);
  and (_12564_, _12563_, _12560_);
  and (_12565_, _12564_, _12553_);
  and (_12566_, _12565_, _12546_);
  not (_12567_, _12566_);
  nor (_12568_, _12567_, _12522_);
  nor (_12569_, _12568_, _06195_);
  or (_12570_, _12569_, _06193_);
  or (_12571_, _12570_, _12521_);
  and (_12572_, _06193_, _03944_);
  nor (_12573_, _12572_, _04510_);
  and (_12574_, _12573_, _12571_);
  nor (_12575_, _06426_, _03855_);
  or (_12576_, _12575_, _03168_);
  or (_12577_, _12576_, _12574_);
  and (_12578_, _11618_, _03168_);
  nor (_12579_, _12578_, _04528_);
  and (_12580_, _12579_, _12577_);
  and (_12581_, _05771_, _03855_);
  nor (_12582_, _12581_, _12458_);
  nor (_12583_, _12582_, _04526_);
  nor (_12584_, _12583_, _04529_);
  or (_12585_, _12584_, _12580_);
  nor (_12586_, _05771_, _07650_);
  and (_12587_, _05771_, _07650_);
  nor (_12588_, _12587_, _12586_);
  or (_12589_, _12588_, _06432_);
  and (_12590_, _12589_, _04525_);
  and (_12591_, _12590_, _12585_);
  or (_12592_, _12591_, _12459_);
  and (_12593_, _12592_, _04522_);
  and (_12594_, _12586_, _04521_);
  or (_12595_, _12594_, _03182_);
  or (_12596_, _12595_, _12593_);
  and (_12597_, _11618_, _03182_);
  nor (_12598_, _12597_, _06454_);
  and (_12599_, _12598_, _12596_);
  nor (_12600_, _12581_, _06460_);
  or (_12601_, _12600_, _06459_);
  or (_12602_, _12601_, _12599_);
  nand (_12603_, _12587_, _06459_);
  and (_12604_, _12603_, _04803_);
  and (_12605_, _12604_, _12602_);
  and (_12606_, _03294_, _03191_);
  or (_12607_, _06468_, _12606_);
  or (_12608_, _12607_, _12605_);
  and (_12609_, _12608_, _12457_);
  nor (_12610_, _12609_, _06475_);
  nor (_12611_, _12610_, _12456_);
  and (_12612_, _12611_, _12455_);
  and (_12613_, _12450_, _12456_);
  nor (_12614_, _12613_, _12612_);
  nor (_12615_, _12614_, _04201_);
  or (_12616_, _12615_, _12451_);
  and (_12617_, _12616_, _06479_);
  nor (_12618_, _12467_, _06479_);
  or (_12619_, _12618_, _03645_);
  or (_12620_, _12619_, _12617_);
  nand (_12621_, _11504_, _03645_);
  and (_12622_, _12621_, _12009_);
  and (_12623_, _12622_, _12620_);
  and (_12624_, _03294_, _03196_);
  or (_12625_, _03448_, _12624_);
  or (_12626_, _12625_, _12623_);
  or (_12627_, _12507_, _03449_);
  and (_12628_, _12627_, _12217_);
  and (_12629_, _12628_, _12626_);
  or (_12630_, _12629_, _12446_);
  and (_12631_, _12630_, _06838_);
  or (_12632_, _06839_, _06710_);
  nor (_12633_, _08054_, _06838_);
  and (_12634_, _12633_, _12632_);
  or (_12635_, _12634_, _04559_);
  or (_12636_, _12635_, _12631_);
  nor (_12637_, _05772_, _05723_);
  nor (_12638_, _12637_, _05773_);
  or (_12639_, _12638_, _04746_);
  and (_12640_, _12639_, _05184_);
  and (_12641_, _12640_, _12636_);
  or (_12642_, _12641_, _12054_);
  and (_12643_, _12642_, _12443_);
  nand (_12644_, _11457_, _03645_);
  or (_12645_, _11586_, _03645_);
  and (_12646_, _12645_, _12644_);
  and (_12647_, _12646_, _05177_);
  and (_12648_, _12647_, _12234_);
  or (_40841_, _12648_, _12643_);
  nand (_12649_, _12054_, _04829_);
  and (_12650_, _12649_, _12248_);
  nor (_12651_, _12465_, _05624_);
  nor (_12652_, _12651_, _06126_);
  nor (_12653_, _12652_, _06479_);
  not (_12654_, _06664_);
  nor (_12655_, _12448_, _12654_);
  or (_12656_, _12655_, _06712_);
  and (_12657_, _12656_, _04544_);
  and (_12658_, _03191_, _02866_);
  nor (_12659_, _05624_, _03725_);
  and (_12660_, _12659_, _04524_);
  or (_12661_, _06023_, _04499_);
  nor (_12662_, _10238_, _05319_);
  or (_12663_, _12662_, _05964_);
  nand (_12664_, _10238_, _09900_);
  or (_12665_, _12664_, _05978_);
  nor (_12666_, _12652_, _04434_);
  nor (_12667_, _12452_, _04885_);
  or (_12668_, _12667_, _05986_);
  or (_12669_, _12668_, _05997_);
  nor (_12670_, _03204_, _03665_);
  and (_12671_, _03204_, \oc8051_golden_model_1.ACC [3]);
  nor (_12672_, _12671_, _12670_);
  and (_12673_, _12672_, _05997_);
  nor (_12674_, _12673_, _04433_);
  and (_12675_, _12674_, _12669_);
  or (_12676_, _12675_, _03472_);
  or (_12677_, _12676_, _12666_);
  and (_12678_, _12677_, _12665_);
  or (_12679_, _12678_, _05977_);
  nor (_12680_, _03202_, _02866_);
  nor (_12681_, _12680_, _04458_);
  and (_12682_, _12681_, _12679_);
  nor (_12683_, _04885_, _04896_);
  or (_12684_, _12683_, _04466_);
  or (_12685_, _12684_, _12682_);
  and (_12686_, _12685_, _12663_);
  or (_12687_, _12686_, _03464_);
  nand (_12688_, _08334_, _03464_);
  and (_12689_, _12688_, _03462_);
  and (_12690_, _12689_, _12687_);
  not (_12691_, _10239_);
  and (_12692_, _12664_, _12691_);
  and (_12693_, _12692_, _03461_);
  or (_12694_, _12693_, _12690_);
  and (_12695_, _12694_, _03207_);
  or (_12696_, _03207_, _03665_);
  nand (_12697_, _03583_, _12696_);
  or (_12698_, _12697_, _12695_);
  nand (_12699_, _08334_, _03584_);
  and (_12700_, _12699_, _12698_);
  or (_12701_, _12700_, _04481_);
  and (_12702_, _06664_, _04493_);
  nand (_12703_, _08333_, _04481_);
  or (_12704_, _12703_, _12702_);
  and (_12705_, _12704_, _12701_);
  or (_12706_, _12705_, _04480_);
  and (_12707_, _05319_, \oc8051_golden_model_1.PSW [7]);
  nor (_12708_, _09923_, _05319_);
  nor (_12709_, _12708_, _12707_);
  nand (_12711_, _12709_, _04480_);
  and (_12712_, _12711_, _05919_);
  and (_12713_, _12712_, _12706_);
  nand (_12714_, _02866_, _03219_);
  nand (_12715_, _04499_, _12714_);
  or (_12716_, _12715_, _12713_);
  and (_12717_, _12716_, _12661_);
  or (_12718_, _12717_, _04501_);
  or (_12719_, _06664_, _06189_);
  and (_12720_, _12719_, _04754_);
  and (_12721_, _12720_, _12718_);
  nor (_12722_, _06227_, _04885_);
  and (_12723_, _06365_, \oc8051_golden_model_1.PSW [3]);
  not (_12724_, _12723_);
  and (_12725_, _06372_, _06343_);
  and (_12726_, _12725_, \oc8051_golden_model_1.IP [3]);
  not (_12727_, _12726_);
  and (_12728_, _06367_, \oc8051_golden_model_1.ACC [3]);
  and (_12729_, _06342_, _06231_);
  and (_12730_, _06363_, _12729_);
  and (_12732_, _12730_, \oc8051_golden_model_1.B [3]);
  nor (_12733_, _12732_, _12728_);
  and (_12734_, _12733_, _12727_);
  and (_12735_, _12734_, _12724_);
  and (_12736_, _06352_, \oc8051_golden_model_1.SP [3]);
  not (_12737_, _12736_);
  and (_12738_, _06412_, \oc8051_golden_model_1.DPL [3]);
  and (_12739_, _06334_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_12740_, _12739_, _12738_);
  and (_12741_, _12740_, _12737_);
  and (_12742_, _12741_, _12735_);
  and (_12743_, _06378_, \oc8051_golden_model_1.IE [3]);
  not (_12744_, _12743_);
  and (_12745_, _06381_, \oc8051_golden_model_1.SCON [3]);
  and (_12746_, _06384_, \oc8051_golden_model_1.SBUF [3]);
  nor (_12747_, _12746_, _12745_);
  and (_12748_, _12747_, _12744_);
  and (_12749_, _06344_, \oc8051_golden_model_1.P3INREG [3]);
  and (_12750_, _06329_, \oc8051_golden_model_1.P2INREG [3]);
  and (_12751_, _06340_, \oc8051_golden_model_1.P1INREG [3]);
  or (_12752_, _12751_, _12750_);
  nor (_12753_, _12752_, _12749_);
  and (_12754_, _12753_, _12748_);
  and (_12755_, _06392_, \oc8051_golden_model_1.TH0 [3]);
  and (_12756_, _06396_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12757_, _12756_, _12755_);
  and (_12758_, _06401_, \oc8051_golden_model_1.PCON [3]);
  and (_12759_, _06403_, \oc8051_golden_model_1.TCON [3]);
  nor (_12760_, _12759_, _12758_);
  and (_12761_, _12760_, _12757_);
  and (_12762_, _06407_, \oc8051_golden_model_1.DPH [3]);
  and (_12763_, _06409_, \oc8051_golden_model_1.TMOD [3]);
  nor (_12764_, _12763_, _12762_);
  and (_12765_, _06414_, \oc8051_golden_model_1.TH1 [3]);
  and (_12766_, _06359_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12767_, _12766_, _12765_);
  and (_12768_, _12767_, _12764_);
  and (_12769_, _12768_, _12761_);
  and (_12770_, _12769_, _12754_);
  and (_12771_, _12770_, _12742_);
  not (_12772_, _12771_);
  nor (_12773_, _12772_, _12722_);
  nor (_12774_, _12773_, _06195_);
  or (_12775_, _12774_, _06193_);
  or (_12776_, _12775_, _12721_);
  and (_12777_, _06193_, _03440_);
  nor (_12778_, _12777_, _04510_);
  and (_12779_, _12778_, _12776_);
  nor (_12780_, _06426_, _03725_);
  or (_12781_, _12780_, _03168_);
  or (_12782_, _12781_, _12779_);
  and (_12783_, _03665_, _03168_);
  nor (_12784_, _12783_, _04528_);
  and (_12785_, _12784_, _12782_);
  and (_12786_, _05624_, _03725_);
  nor (_12787_, _12786_, _12659_);
  nor (_12788_, _12787_, _04526_);
  nor (_12789_, _12788_, _04529_);
  or (_12790_, _12789_, _12785_);
  nor (_12791_, _05624_, _07644_);
  and (_12792_, _05624_, _07644_);
  nor (_12793_, _12792_, _12791_);
  or (_12794_, _12793_, _06432_);
  and (_12795_, _12794_, _04525_);
  and (_12796_, _12795_, _12790_);
  or (_12797_, _12796_, _12660_);
  and (_12798_, _12797_, _04522_);
  and (_12799_, _12791_, _04521_);
  or (_12800_, _12799_, _03182_);
  or (_12801_, _12800_, _12798_);
  and (_12802_, _03182_, _03665_);
  nor (_12803_, _12802_, _06454_);
  and (_12804_, _12803_, _12801_);
  nor (_12805_, _12786_, _06460_);
  or (_12806_, _12805_, _06459_);
  or (_12807_, _12806_, _12804_);
  nand (_12808_, _12792_, _06459_);
  and (_12809_, _12808_, _04803_);
  and (_12810_, _12809_, _12807_);
  nor (_12811_, _12810_, _12658_);
  or (_12812_, _12811_, _11988_);
  nor (_12813_, _04720_, _04205_);
  nand (_12814_, _12668_, _11988_);
  and (_12815_, _12814_, _12813_);
  nand (_12816_, _12815_, _12812_);
  or (_12817_, _12813_, _12668_);
  and (_12818_, _12817_, _06480_);
  and (_12819_, _12818_, _12816_);
  or (_12820_, _12819_, _12657_);
  and (_12821_, _12820_, _06479_);
  or (_12822_, _12821_, _12653_);
  and (_12823_, _12822_, _06855_);
  and (_12824_, _11498_, _03645_);
  or (_12825_, _12824_, _03196_);
  or (_12826_, _12825_, _12823_);
  and (_12827_, _03196_, _03665_);
  nor (_12828_, _12827_, _03448_);
  and (_12829_, _12828_, _12826_);
  and (_12830_, _12708_, _03448_);
  or (_12831_, _12830_, _12829_);
  and (_12832_, _12831_, _12015_);
  or (_12833_, _08054_, _06664_);
  nor (_12834_, _06841_, _06838_);
  and (_12835_, _12834_, _12833_);
  or (_12836_, _08222_, _06023_);
  nor (_12837_, _12217_, _05892_);
  and (_12838_, _12837_, _12836_);
  or (_12839_, _12838_, _04559_);
  or (_12840_, _12839_, _12835_);
  or (_12841_, _12840_, _12832_);
  nor (_12842_, _05773_, _05625_);
  nor (_12843_, _12842_, _05774_);
  or (_12844_, _12843_, _04746_);
  and (_12845_, _12844_, _05184_);
  and (_12846_, _12845_, _12841_);
  or (_12847_, _12846_, _12054_);
  and (_12848_, _12847_, _12650_);
  nand (_12849_, _11464_, _03645_);
  or (_12850_, _11581_, _03645_);
  and (_12851_, _12850_, _12849_);
  and (_12852_, _12851_, _05177_);
  and (_12853_, _12852_, _12234_);
  or (_40843_, _12853_, _12848_);
  and (_12854_, _06126_, _05879_);
  nor (_12855_, _06126_, _05879_);
  nor (_12856_, _12855_, _12854_);
  nand (_12857_, _12856_, _04546_);
  nor (_12858_, _05986_, _05831_);
  and (_12859_, _05986_, _05831_);
  or (_12860_, _12859_, _12858_);
  or (_12861_, _12860_, _06471_);
  nor (_12862_, _06326_, _05879_);
  and (_12863_, _12862_, _04524_);
  nor (_12864_, _09820_, _10202_);
  or (_12865_, _12864_, _05964_);
  nand (_12866_, _09821_, _10202_);
  or (_12867_, _12866_, _05978_);
  and (_12868_, _12860_, _05998_);
  nor (_12869_, _11614_, _03204_);
  and (_12870_, _03204_, \oc8051_golden_model_1.ACC [4]);
  or (_12871_, _12870_, _12869_);
  and (_12872_, _12871_, _05997_);
  or (_12873_, _12872_, _04012_);
  or (_12874_, _12873_, _12868_);
  or (_12875_, _06802_, _06008_);
  and (_12876_, _12875_, _12874_);
  or (_12877_, _12876_, _04433_);
  nand (_12878_, _12856_, _04433_);
  and (_12879_, _12878_, _12877_);
  or (_12880_, _12879_, _03472_);
  and (_12881_, _12880_, _12867_);
  or (_12882_, _12881_, _05977_);
  nor (_12883_, _11613_, _03202_);
  nor (_12884_, _12883_, _04458_);
  and (_12885_, _12884_, _12882_);
  nor (_12886_, _05831_, _04896_);
  or (_12887_, _12886_, _04466_);
  or (_12888_, _12887_, _12885_);
  and (_12889_, _12888_, _12865_);
  or (_12890_, _12889_, _03464_);
  nand (_12891_, _08320_, _03464_);
  and (_12892_, _12891_, _03462_);
  and (_12893_, _12892_, _12890_);
  not (_12894_, _10203_);
  and (_12895_, _12866_, _12894_);
  and (_12896_, _12895_, _03461_);
  or (_12897_, _12896_, _12893_);
  and (_12898_, _12897_, _03207_);
  or (_12899_, _11614_, _03207_);
  nand (_12900_, _12899_, _03583_);
  or (_12901_, _12900_, _12898_);
  nand (_12902_, _08320_, _03584_);
  and (_12903_, _12902_, _12901_);
  or (_12904_, _12903_, _04481_);
  and (_12905_, _06802_, _04493_);
  nand (_12906_, _08319_, _04481_);
  or (_12907_, _12906_, _12905_);
  and (_12908_, _12907_, _12904_);
  or (_12909_, _12908_, _04480_);
  nor (_12910_, _09844_, _09820_);
  and (_12911_, _09820_, \oc8051_golden_model_1.PSW [7]);
  nor (_12912_, _12911_, _12910_);
  nand (_12913_, _12912_, _04480_);
  and (_12914_, _12913_, _05919_);
  and (_12915_, _12914_, _12909_);
  nand (_12916_, _11613_, _03219_);
  nand (_12917_, _12916_, _04499_);
  or (_12918_, _12917_, _12915_);
  or (_12919_, _05889_, _04499_);
  and (_12920_, _12919_, _12918_);
  or (_12921_, _12920_, _04501_);
  or (_12922_, _06802_, _06189_);
  and (_12923_, _12922_, _04754_);
  and (_12924_, _12923_, _12921_);
  nor (_12925_, _06227_, _05831_);
  and (_12926_, _06329_, \oc8051_golden_model_1.P2INREG [4]);
  not (_12927_, _12926_);
  and (_12928_, _06334_, \oc8051_golden_model_1.P0INREG [4]);
  not (_12929_, _12928_);
  and (_12930_, _06340_, \oc8051_golden_model_1.P1INREG [4]);
  and (_12931_, _06344_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_12932_, _12931_, _12930_);
  and (_12933_, _12932_, _12929_);
  and (_12934_, _12933_, _12927_);
  and (_12935_, _06352_, \oc8051_golden_model_1.SP [4]);
  and (_12936_, _06359_, \oc8051_golden_model_1.TL0 [4]);
  nor (_12937_, _12936_, _12935_);
  and (_12938_, _12937_, _12934_);
  and (_12939_, _06378_, \oc8051_golden_model_1.IE [4]);
  not (_12940_, _12939_);
  and (_12941_, _06381_, \oc8051_golden_model_1.SCON [4]);
  and (_12942_, _06384_, \oc8051_golden_model_1.SBUF [4]);
  nor (_12943_, _12942_, _12941_);
  and (_12944_, _12943_, _12940_);
  and (_12945_, _06370_, \oc8051_golden_model_1.B [4]);
  and (_12946_, _06374_, \oc8051_golden_model_1.IP [4]);
  nor (_12947_, _12946_, _12945_);
  and (_12948_, _06365_, \oc8051_golden_model_1.PSW [4]);
  and (_12949_, _06367_, \oc8051_golden_model_1.ACC [4]);
  nor (_12950_, _12949_, _12948_);
  and (_12951_, _12950_, _12947_);
  and (_12952_, _12951_, _12944_);
  and (_12953_, _12952_, _12938_);
  and (_12954_, _06407_, \oc8051_golden_model_1.DPH [4]);
  and (_12955_, _06409_, \oc8051_golden_model_1.TMOD [4]);
  nor (_12956_, _12955_, _12954_);
  and (_12957_, _06412_, \oc8051_golden_model_1.DPL [4]);
  and (_12958_, _06414_, \oc8051_golden_model_1.TH1 [4]);
  nor (_12959_, _12958_, _12957_);
  and (_12960_, _12959_, _12956_);
  and (_12961_, _06372_, _06333_);
  and (_12962_, _12961_, \oc8051_golden_model_1.TCON [4]);
  and (_12963_, _06392_, \oc8051_golden_model_1.TH0 [4]);
  nor (_12964_, _12963_, _12962_);
  and (_12965_, _06401_, \oc8051_golden_model_1.PCON [4]);
  and (_12966_, _06396_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12967_, _12966_, _12965_);
  and (_12968_, _12967_, _12964_);
  and (_12969_, _12968_, _12960_);
  and (_12970_, _12969_, _12953_);
  not (_12971_, _12970_);
  nor (_12972_, _12971_, _12925_);
  nor (_12973_, _12972_, _06195_);
  or (_12974_, _12973_, _06193_);
  or (_12975_, _12974_, _12924_);
  and (_12976_, _06193_, _04257_);
  nor (_12977_, _12976_, _04510_);
  and (_12978_, _12977_, _12975_);
  nor (_12979_, _06326_, _06426_);
  or (_12980_, _12979_, _03168_);
  or (_12981_, _12980_, _12978_);
  and (_12982_, _11614_, _03168_);
  nor (_12983_, _12982_, _04528_);
  and (_12984_, _12983_, _12981_);
  and (_12985_, _06326_, _05879_);
  nor (_12986_, _12985_, _12862_);
  nor (_12987_, _12986_, _04526_);
  nor (_12988_, _12987_, _04529_);
  or (_12989_, _12988_, _12984_);
  nor (_12990_, _05879_, _07545_);
  and (_12991_, _05879_, _07545_);
  nor (_12992_, _12991_, _12990_);
  or (_12993_, _12992_, _06432_);
  and (_12994_, _12993_, _04525_);
  and (_12995_, _12994_, _12989_);
  or (_12996_, _12995_, _12863_);
  and (_12997_, _12996_, _04522_);
  and (_12998_, _12990_, _04521_);
  or (_12999_, _12998_, _03182_);
  or (_13000_, _12999_, _12997_);
  and (_13001_, _11614_, _03182_);
  nor (_13002_, _13001_, _06454_);
  and (_13003_, _13002_, _13000_);
  nor (_13004_, _12985_, _06460_);
  or (_13005_, _13004_, _06459_);
  or (_13006_, _13005_, _13003_);
  nand (_13007_, _12991_, _06459_);
  and (_13008_, _13007_, _04803_);
  and (_13009_, _13008_, _13006_);
  and (_13010_, _11613_, _03191_);
  or (_13011_, _13010_, _06468_);
  or (_13012_, _13011_, _13009_);
  and (_13013_, _13012_, _12861_);
  or (_13014_, _13013_, _06475_);
  or (_13015_, _12860_, _04721_);
  and (_13016_, _13015_, _06480_);
  and (_13017_, _13016_, _13014_);
  not (_13018_, _06802_);
  and (_13019_, _06712_, _13018_);
  nor (_13020_, _06712_, _13018_);
  or (_13021_, _13020_, _13019_);
  and (_13022_, _13021_, _04544_);
  or (_13023_, _13022_, _04546_);
  or (_13024_, _13023_, _13017_);
  and (_13025_, _13024_, _12857_);
  or (_13026_, _13025_, _03645_);
  nand (_13027_, _11495_, _03645_);
  and (_13028_, _13027_, _12009_);
  and (_13029_, _13028_, _13026_);
  and (_13030_, _11613_, _03196_);
  or (_13031_, _13030_, _03448_);
  or (_13032_, _13031_, _13029_);
  or (_13033_, _12910_, _03449_);
  and (_13034_, _13033_, _06833_);
  and (_13035_, _13034_, _13032_);
  nor (_13036_, _05892_, _05889_);
  nor (_13037_, _13036_, _05893_);
  and (_13038_, _13037_, _06830_);
  or (_13039_, _13038_, _04737_);
  or (_13040_, _13039_, _13035_);
  or (_13041_, _13037_, _04736_);
  and (_13042_, _13041_, _06838_);
  and (_13043_, _13042_, _13040_);
  or (_13044_, _06841_, _06802_);
  and (_13045_, _06841_, _06802_);
  nor (_13046_, _13045_, _06838_);
  and (_13047_, _13046_, _13044_);
  or (_13048_, _13047_, _04559_);
  or (_13049_, _13048_, _13043_);
  nor (_13050_, _05880_, _05774_);
  nor (_13051_, _13050_, _05881_);
  or (_13052_, _13051_, _04746_);
  and (_13053_, _13052_, _05184_);
  and (_13054_, _13053_, _13049_);
  or (_13055_, _13054_, _12054_);
  nand (_13056_, _12054_, _05775_);
  and (_13057_, _13056_, _12248_);
  and (_13058_, _13057_, _13055_);
  nand (_13059_, _11453_, _03645_);
  or (_13060_, _11578_, _03645_);
  and (_13061_, _13060_, _13059_);
  and (_13062_, _13061_, _05177_);
  and (_13063_, _13062_, _12234_);
  or (_40844_, _13063_, _13058_);
  nand (_13064_, _12054_, _05470_);
  and (_13065_, _13064_, _12248_);
  nor (_13066_, _05893_, _05888_);
  nor (_13067_, _13066_, _05894_);
  and (_13068_, _13067_, _12014_);
  nor (_13069_, _12854_, _05575_);
  nor (_13070_, _13069_, _06127_);
  nand (_13071_, _13070_, _04546_);
  nor (_13072_, _06294_, _05575_);
  and (_13073_, _13072_, _04524_);
  nor (_13074_, _09949_, _09925_);
  and (_13075_, _09925_, \oc8051_golden_model_1.PSW [7]);
  nor (_13076_, _13075_, _13074_);
  nor (_13077_, _13076_, _04946_);
  nor (_13078_, _09925_, _10249_);
  or (_13079_, _13078_, _05964_);
  nor (_13080_, _13070_, _04434_);
  or (_13081_, _06757_, _06008_);
  nor (_13082_, _12859_, _05526_);
  or (_13083_, _13082_, _05987_);
  and (_13084_, _13083_, _05998_);
  or (_13085_, _11608_, _03204_);
  nand (_13086_, _03204_, _07539_);
  and (_13087_, _13086_, _13085_);
  and (_13088_, _13087_, _05997_);
  or (_13089_, _13088_, _04012_);
  or (_13090_, _13089_, _13084_);
  and (_13091_, _13090_, _04434_);
  and (_13092_, _13091_, _13081_);
  or (_13093_, _13092_, _13080_);
  and (_13094_, _13093_, _05978_);
  nand (_13095_, _09926_, _10249_);
  and (_13096_, _13095_, _03472_);
  or (_13097_, _13096_, _05977_);
  or (_13098_, _13097_, _13094_);
  nor (_13099_, _11608_, _03202_);
  nor (_13100_, _13099_, _04458_);
  and (_13101_, _13100_, _13098_);
  nor (_13102_, _05526_, _04896_);
  or (_13103_, _13102_, _04466_);
  or (_13104_, _13103_, _13101_);
  and (_13105_, _13104_, _13079_);
  or (_13106_, _13105_, _03464_);
  nand (_13107_, _08305_, _03464_);
  and (_13108_, _13107_, _03462_);
  and (_13109_, _13108_, _13106_);
  not (_13110_, _10250_);
  and (_13111_, _13095_, _13110_);
  and (_13112_, _13111_, _03461_);
  or (_13113_, _13112_, _13109_);
  and (_13114_, _13113_, _03207_);
  or (_13115_, _11609_, _03207_);
  nand (_13116_, _13115_, _03583_);
  or (_13117_, _13116_, _13114_);
  nand (_13118_, _08305_, _03584_);
  and (_13119_, _13118_, _13117_);
  or (_13120_, _13119_, _04481_);
  and (_13121_, _06757_, _04493_);
  nand (_13122_, _08304_, _04481_);
  or (_13123_, _13122_, _13121_);
  and (_13124_, _13123_, _04946_);
  and (_13125_, _13124_, _13120_);
  or (_13126_, _13125_, _13077_);
  and (_13127_, _13126_, _05919_);
  nand (_13128_, _11608_, _03219_);
  nand (_13129_, _13128_, _04499_);
  or (_13130_, _13129_, _13127_);
  or (_13131_, _05888_, _04499_);
  and (_13132_, _13131_, _13130_);
  or (_13133_, _13132_, _04501_);
  or (_13134_, _06757_, _06189_);
  and (_13135_, _13134_, _04754_);
  and (_13136_, _13135_, _13133_);
  nor (_13137_, _06227_, _05526_);
  and (_13138_, _12725_, \oc8051_golden_model_1.IP [5]);
  not (_13139_, _13138_);
  and (_13140_, _06365_, \oc8051_golden_model_1.PSW [5]);
  not (_13141_, _13140_);
  and (_13142_, _06367_, \oc8051_golden_model_1.ACC [5]);
  and (_13143_, _12730_, \oc8051_golden_model_1.B [5]);
  nor (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _13141_);
  and (_13146_, _13145_, _13139_);
  and (_13147_, _06352_, \oc8051_golden_model_1.SP [5]);
  not (_13148_, _13147_);
  and (_13149_, _06412_, \oc8051_golden_model_1.DPL [5]);
  and (_13150_, _06334_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_13151_, _13150_, _13149_);
  and (_13152_, _13151_, _13148_);
  and (_13153_, _13152_, _13146_);
  and (_13154_, _06378_, \oc8051_golden_model_1.IE [5]);
  not (_13155_, _13154_);
  and (_13156_, _06381_, \oc8051_golden_model_1.SCON [5]);
  and (_13157_, _06384_, \oc8051_golden_model_1.SBUF [5]);
  nor (_13158_, _13157_, _13156_);
  and (_13159_, _13158_, _13155_);
  and (_13160_, _06344_, \oc8051_golden_model_1.P3INREG [5]);
  and (_13161_, _06329_, \oc8051_golden_model_1.P2INREG [5]);
  and (_13162_, _06340_, \oc8051_golden_model_1.P1INREG [5]);
  or (_13163_, _13162_, _13161_);
  nor (_13164_, _13163_, _13160_);
  and (_13165_, _13164_, _13159_);
  and (_13166_, _06392_, \oc8051_golden_model_1.TH0 [5]);
  and (_13167_, _06396_, \oc8051_golden_model_1.TL1 [5]);
  nor (_13168_, _13167_, _13166_);
  and (_13169_, _06401_, \oc8051_golden_model_1.PCON [5]);
  and (_13170_, _06403_, \oc8051_golden_model_1.TCON [5]);
  nor (_13171_, _13170_, _13169_);
  and (_13172_, _13171_, _13168_);
  and (_13173_, _06407_, \oc8051_golden_model_1.DPH [5]);
  and (_13174_, _06409_, \oc8051_golden_model_1.TMOD [5]);
  nor (_13175_, _13174_, _13173_);
  and (_13176_, _06414_, \oc8051_golden_model_1.TH1 [5]);
  and (_13177_, _06359_, \oc8051_golden_model_1.TL0 [5]);
  nor (_13178_, _13177_, _13176_);
  and (_13179_, _13178_, _13175_);
  and (_13180_, _13179_, _13172_);
  and (_13181_, _13180_, _13165_);
  and (_13182_, _13181_, _13153_);
  not (_13183_, _13182_);
  nor (_13184_, _13183_, _13137_);
  nor (_13185_, _13184_, _06195_);
  or (_13186_, _13185_, _06193_);
  or (_13187_, _13186_, _13136_);
  and (_13188_, _06193_, _03811_);
  nor (_13189_, _13188_, _04510_);
  and (_13190_, _13189_, _13187_);
  nor (_13191_, _06294_, _06426_);
  or (_13192_, _13191_, _03168_);
  or (_13193_, _13192_, _13190_);
  and (_13194_, _11609_, _03168_);
  nor (_13195_, _13194_, _04528_);
  and (_13196_, _13195_, _13193_);
  and (_13197_, _06294_, _05575_);
  nor (_13198_, _13197_, _13072_);
  nor (_13199_, _13198_, _04526_);
  nor (_13200_, _13199_, _04529_);
  or (_13201_, _13200_, _13196_);
  nor (_13202_, _05575_, _07539_);
  and (_13203_, _05575_, _07539_);
  nor (_13204_, _13203_, _13202_);
  or (_13205_, _13204_, _06432_);
  and (_13206_, _13205_, _04525_);
  and (_13207_, _13206_, _13201_);
  or (_13208_, _13207_, _13073_);
  and (_13209_, _13208_, _04522_);
  and (_13210_, _13202_, _04521_);
  or (_13211_, _13210_, _03182_);
  or (_13212_, _13211_, _13209_);
  and (_13213_, _11609_, _03182_);
  nor (_13214_, _13213_, _06454_);
  and (_13215_, _13214_, _13212_);
  nor (_13216_, _13197_, _06460_);
  or (_13217_, _13216_, _06459_);
  or (_13218_, _13217_, _13215_);
  nand (_13219_, _13203_, _06459_);
  and (_13220_, _13219_, _04803_);
  and (_13221_, _13220_, _13218_);
  nand (_13222_, _11608_, _03191_);
  nand (_13223_, _13222_, _11990_);
  or (_13224_, _13223_, _13221_);
  or (_13225_, _13083_, _11990_);
  and (_13226_, _13225_, _06480_);
  and (_13227_, _13226_, _13224_);
  not (_13228_, _06757_);
  nor (_13229_, _13019_, _13228_);
  or (_13230_, _13229_, _06804_);
  and (_13231_, _13230_, _04544_);
  or (_13232_, _13231_, _04546_);
  or (_13233_, _13232_, _13227_);
  and (_13234_, _13233_, _13071_);
  or (_13235_, _13234_, _03645_);
  nand (_13236_, _11490_, _03645_);
  and (_13237_, _13236_, _12009_);
  and (_13238_, _13237_, _13235_);
  and (_13239_, _11608_, _03196_);
  or (_13240_, _13239_, _03448_);
  or (_13241_, _13240_, _13238_);
  or (_13242_, _13074_, _03449_);
  and (_13243_, _13242_, _12217_);
  and (_13244_, _13243_, _13241_);
  or (_13245_, _13244_, _13068_);
  and (_13246_, _13245_, _06838_);
  or (_13247_, _13045_, _06757_);
  nor (_13248_, _06843_, _06838_);
  and (_13249_, _13248_, _13247_);
  or (_13250_, _13249_, _04559_);
  or (_13251_, _13250_, _13246_);
  nor (_13252_, _05881_, _05576_);
  nor (_13253_, _13252_, _05882_);
  or (_13254_, _13253_, _04746_);
  and (_13255_, _13254_, _05184_);
  and (_13256_, _13255_, _13251_);
  or (_13257_, _13256_, _12054_);
  and (_13258_, _13257_, _13065_);
  not (_13259_, _11574_);
  nor (_13260_, _13259_, _03645_);
  and (_13261_, _11448_, _03645_);
  or (_13262_, _13261_, _13260_);
  and (_13263_, _13262_, _05177_);
  and (_13264_, _13263_, _12234_);
  or (_40846_, _13264_, _13258_);
  nand (_13265_, _12054_, _05359_);
  and (_13266_, _13265_, _12248_);
  nor (_13267_, _06843_, _06526_);
  nor (_13268_, _13267_, _06844_);
  or (_13269_, _13268_, _06838_);
  nor (_13270_, _06804_, _06527_);
  or (_13271_, _13270_, _06805_);
  and (_13272_, _13271_, _04544_);
  nor (_13273_, _05987_, _05417_);
  or (_13274_, _13273_, _05988_);
  or (_13275_, _13274_, _06471_);
  nor (_13276_, _05468_, _07495_);
  or (_13277_, _13276_, _04522_);
  and (_13278_, _11600_, _03219_);
  nor (_13279_, _05417_, _04896_);
  nand (_13280_, _09875_, _10226_);
  or (_13281_, _13280_, _05978_);
  or (_13282_, _06526_, _06008_);
  and (_13283_, _13274_, _05998_);
  nor (_13284_, _11601_, _03204_);
  and (_13285_, _03204_, \oc8051_golden_model_1.ACC [6]);
  or (_13286_, _13285_, _13284_);
  and (_13287_, _13286_, _05997_);
  or (_13288_, _13287_, _04012_);
  or (_13289_, _13288_, _13283_);
  and (_13290_, _13289_, _13282_);
  or (_13291_, _13290_, _04433_);
  nor (_13292_, _06127_, _05468_);
  nor (_13293_, _13292_, _06129_);
  nand (_13294_, _13293_, _04433_);
  and (_13295_, _13294_, _13291_);
  or (_13296_, _13295_, _03472_);
  and (_13297_, _13296_, _13281_);
  or (_13298_, _13297_, _05977_);
  nor (_13299_, _11600_, _03202_);
  nor (_13300_, _13299_, _04458_);
  and (_13301_, _13300_, _13298_);
  or (_13302_, _13301_, _13279_);
  and (_13303_, _13302_, _05964_);
  nor (_13304_, _09874_, _10226_);
  and (_13305_, _13304_, _04466_);
  or (_13306_, _13305_, _03464_);
  or (_13307_, _13306_, _13303_);
  nand (_13308_, _08287_, _03464_);
  and (_13309_, _13308_, _03462_);
  and (_13310_, _13309_, _13307_);
  not (_13311_, _10227_);
  and (_13312_, _13280_, _13311_);
  and (_13313_, _13312_, _03461_);
  or (_13314_, _13313_, _13310_);
  and (_13315_, _13314_, _03207_);
  or (_13316_, _11601_, _03207_);
  nand (_13317_, _13316_, _03583_);
  or (_13318_, _13317_, _13315_);
  nand (_13319_, _08287_, _03584_);
  and (_13320_, _13319_, _13318_);
  or (_13321_, _13320_, _04481_);
  and (_13322_, _06526_, _04493_);
  nand (_13323_, _08286_, _04481_);
  or (_13324_, _13323_, _13322_);
  and (_13325_, _13324_, _13321_);
  or (_13326_, _13325_, _04480_);
  nor (_13327_, _09897_, _09874_);
  and (_13328_, _09874_, \oc8051_golden_model_1.PSW [7]);
  nor (_13329_, _13328_, _13327_);
  nand (_13330_, _13329_, _04480_);
  and (_13331_, _13330_, _05919_);
  and (_13332_, _13331_, _13326_);
  or (_13333_, _13332_, _13278_);
  and (_13334_, _13333_, _04499_);
  nor (_13335_, _05417_, _04499_);
  or (_13336_, _13335_, _04501_);
  or (_13337_, _13336_, _13334_);
  or (_13338_, _06526_, _12310_);
  and (_13339_, _13338_, _06195_);
  and (_13340_, _13339_, _13337_);
  nor (_13341_, _06227_, _05417_);
  and (_13342_, _06365_, \oc8051_golden_model_1.PSW [6]);
  and (_13343_, _06370_, \oc8051_golden_model_1.B [6]);
  nor (_13344_, _13343_, _13342_);
  and (_13345_, _06367_, \oc8051_golden_model_1.ACC [6]);
  and (_13346_, _06374_, \oc8051_golden_model_1.IP [6]);
  nor (_13347_, _13346_, _13345_);
  and (_13348_, _13347_, _13344_);
  and (_13349_, _06329_, \oc8051_golden_model_1.P2INREG [6]);
  not (_13350_, _13349_);
  and (_13351_, _06334_, \oc8051_golden_model_1.P0INREG [6]);
  not (_13352_, _13351_);
  and (_13353_, _06340_, \oc8051_golden_model_1.P1INREG [6]);
  and (_13354_, _06344_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _13352_);
  and (_13357_, _13356_, _13350_);
  and (_13358_, _13357_, _13348_);
  and (_13359_, _06378_, \oc8051_golden_model_1.IE [6]);
  not (_13360_, _13359_);
  and (_13361_, _06381_, \oc8051_golden_model_1.SCON [6]);
  and (_13362_, _06384_, \oc8051_golden_model_1.SBUF [6]);
  nor (_13363_, _13362_, _13361_);
  and (_13364_, _13363_, _13360_);
  and (_13365_, _06407_, \oc8051_golden_model_1.DPH [6]);
  and (_13366_, _06414_, \oc8051_golden_model_1.TH1 [6]);
  nor (_13367_, _13366_, _13365_);
  and (_13368_, _13367_, _13364_);
  and (_13369_, _13368_, _13358_);
  and (_13370_, _06392_, \oc8051_golden_model_1.TH0 [6]);
  and (_13371_, _06396_, \oc8051_golden_model_1.TL1 [6]);
  nor (_13372_, _13371_, _13370_);
  and (_13373_, _06401_, \oc8051_golden_model_1.PCON [6]);
  and (_13374_, _06403_, \oc8051_golden_model_1.TCON [6]);
  nor (_13375_, _13374_, _13373_);
  and (_13376_, _13375_, _13372_);
  and (_13377_, _06412_, \oc8051_golden_model_1.DPL [6]);
  and (_13378_, _06359_, \oc8051_golden_model_1.TL0 [6]);
  nor (_13379_, _13378_, _13377_);
  and (_13380_, _06352_, \oc8051_golden_model_1.SP [6]);
  and (_13381_, _06409_, \oc8051_golden_model_1.TMOD [6]);
  nor (_13382_, _13381_, _13380_);
  and (_13383_, _13382_, _13379_);
  and (_13384_, _13383_, _13376_);
  and (_13385_, _13384_, _13369_);
  not (_13386_, _13385_);
  nor (_13387_, _13386_, _13341_);
  nor (_13388_, _13387_, _06195_);
  or (_13389_, _13388_, _06193_);
  or (_13390_, _13389_, _13340_);
  and (_13391_, _06193_, _03511_);
  nor (_13392_, _13391_, _04510_);
  and (_13393_, _13392_, _13390_);
  nor (_13394_, _06262_, _06426_);
  or (_13395_, _13394_, _03168_);
  or (_13396_, _13395_, _13393_);
  and (_13397_, _11601_, _03168_);
  nor (_13398_, _13397_, _04528_);
  and (_13399_, _13398_, _13396_);
  and (_13400_, _06262_, _05468_);
  nor (_13401_, _06262_, _05468_);
  nor (_13402_, _13401_, _13400_);
  and (_13403_, _13402_, _04528_);
  or (_13404_, _13403_, _04526_);
  or (_13405_, _13404_, _13399_);
  and (_13406_, _05468_, _07495_);
  nor (_13407_, _13406_, _13276_);
  or (_13408_, _13407_, _06432_);
  and (_13409_, _13408_, _04525_);
  and (_13410_, _13409_, _13405_);
  and (_13411_, _13401_, _04524_);
  or (_13412_, _13411_, _04521_);
  or (_13413_, _13412_, _13410_);
  and (_13414_, _13413_, _13277_);
  or (_13415_, _13414_, _03182_);
  and (_13416_, _11601_, _03182_);
  nor (_13417_, _13416_, _06454_);
  and (_13418_, _13417_, _13415_);
  nor (_13419_, _13400_, _06460_);
  or (_13420_, _13419_, _06459_);
  or (_13421_, _13420_, _13418_);
  nand (_13422_, _13406_, _06459_);
  and (_13423_, _13422_, _04803_);
  and (_13424_, _13423_, _13421_);
  and (_13425_, _11600_, _03191_);
  or (_13426_, _13425_, _06468_);
  or (_13427_, _13426_, _13424_);
  and (_13428_, _13427_, _13275_);
  or (_13429_, _13428_, _06475_);
  or (_13430_, _13274_, _04721_);
  and (_13431_, _13430_, _06480_);
  and (_13432_, _13431_, _13429_);
  or (_13433_, _13432_, _13272_);
  and (_13434_, _13433_, _06479_);
  nor (_13435_, _13293_, _06479_);
  or (_13436_, _13435_, _03645_);
  or (_13437_, _13436_, _13434_);
  nand (_13438_, _11482_, _03645_);
  and (_13439_, _13438_, _12009_);
  and (_13440_, _13439_, _13437_);
  and (_13441_, _11600_, _03196_);
  or (_13442_, _13441_, _03448_);
  or (_13443_, _13442_, _13440_);
  or (_13444_, _13327_, _03449_);
  and (_13445_, _13444_, _12217_);
  and (_13446_, _13445_, _13443_);
  nor (_13447_, _05894_, _05417_);
  and (_13448_, _05894_, _05417_);
  or (_13449_, _13448_, _13447_);
  and (_13450_, _13449_, _12014_);
  or (_13451_, _13450_, _04215_);
  or (_13452_, _13451_, _13446_);
  and (_13453_, _13452_, _13269_);
  or (_13454_, _13453_, _04559_);
  nor (_13455_, _05882_, _05469_);
  nor (_13456_, _13455_, _05883_);
  or (_13457_, _13456_, _04746_);
  and (_13458_, _13457_, _05184_);
  and (_13459_, _13458_, _13454_);
  or (_13460_, _13459_, _12054_);
  and (_13461_, _13460_, _13266_);
  nand (_13462_, _11442_, _03645_);
  or (_13463_, _11569_, _03645_);
  and (_13464_, _13463_, _13462_);
  and (_13465_, _13464_, _05177_);
  and (_13466_, _13465_, _12234_);
  or (_40847_, _13466_, _13461_);
  nand (_13467_, _12054_, _05193_);
  and (_13468_, _13467_, _12248_);
  or (_13469_, _12054_, _06852_);
  and (_13470_, _13469_, _13468_);
  and (_13471_, _12234_, _06891_);
  or (_40848_, _13471_, _13470_);
  and (_13472_, _05186_, _04744_);
  and (_13473_, _13472_, _12052_);
  or (_13474_, _13473_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_13475_, _12243_, _04887_);
  or (_13476_, _13475_, _12246_);
  and (_13477_, _13476_, _13474_);
  not (_13478_, _13473_);
  or (_13479_, _13478_, _12229_);
  and (_13480_, _13479_, _13477_);
  and (_13481_, _05177_, _04887_);
  and (_13482_, _13481_, _12232_);
  and (_13483_, _13482_, _12241_);
  or (_40853_, _13483_, _13480_);
  or (_13484_, _13473_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_13485_, _13484_, _13476_);
  or (_13486_, _13478_, _12434_);
  and (_13487_, _13486_, _13485_);
  and (_13488_, _13482_, _12440_);
  or (_40854_, _13488_, _13487_);
  or (_13489_, _13473_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_13490_, _13489_, _13476_);
  or (_13491_, _13478_, _12641_);
  and (_13492_, _13491_, _13490_);
  and (_13493_, _13482_, _12647_);
  or (_40855_, _13493_, _13492_);
  or (_13494_, _13473_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_13495_, _13494_, _13476_);
  or (_13496_, _13478_, _12846_);
  and (_13497_, _13496_, _13495_);
  and (_13498_, _13482_, _12852_);
  or (_40856_, _13498_, _13497_);
  or (_13499_, _13473_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_13500_, _13499_, _13476_);
  or (_13501_, _13478_, _13054_);
  and (_13502_, _13501_, _13500_);
  and (_13503_, _13482_, _13062_);
  or (_40857_, _13503_, _13502_);
  or (_13504_, _13473_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_13505_, _13504_, _13476_);
  or (_13506_, _13478_, _13256_);
  and (_13507_, _13506_, _13505_);
  and (_13508_, _13482_, _13263_);
  or (_40859_, _13508_, _13507_);
  or (_13509_, _13473_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_13510_, _13509_, _13476_);
  or (_13511_, _13478_, _13459_);
  and (_13512_, _13511_, _13510_);
  and (_13513_, _13482_, _13465_);
  or (_40860_, _13513_, _13512_);
  or (_13514_, _13473_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_13515_, _13514_, _13476_);
  or (_13516_, _13478_, _06852_);
  and (_13517_, _13516_, _13515_);
  and (_13518_, _13482_, _06891_);
  or (_40861_, _13518_, _13517_);
  nor (_13519_, _05004_, _04824_);
  nor (_13520_, _13519_, _05162_);
  and (_13521_, _04825_, _04565_);
  and (_13522_, _13521_, _13520_);
  or (_13523_, _13522_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_13524_, _06009_);
  nor (_13525_, _12246_, _13524_);
  nand (_13526_, _13525_, _12243_);
  and (_13527_, _13526_, _13523_);
  and (_13528_, _12227_, _04823_);
  and (_13529_, _13528_, _12226_);
  not (_13530_, _13522_);
  or (_13531_, _13530_, _13529_);
  and (_13532_, _13531_, _13527_);
  and (_13533_, _06009_, _05177_);
  and (_13534_, _13533_, _12232_);
  and (_13535_, _13534_, _12241_);
  or (_40865_, _13535_, _13532_);
  or (_13536_, _13522_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_13537_, _13536_, _13526_);
  and (_13538_, _12432_, _04823_);
  and (_13539_, _13538_, _12431_);
  or (_13540_, _13530_, _13539_);
  and (_13541_, _13540_, _13537_);
  and (_13542_, _13534_, _12440_);
  or (_40866_, _13542_, _13541_);
  or (_13543_, _13522_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_13544_, _13543_, _13526_);
  and (_13545_, _12639_, _04823_);
  and (_13546_, _13545_, _12636_);
  or (_13547_, _13530_, _13546_);
  and (_13548_, _13547_, _13544_);
  and (_13549_, _13534_, _12647_);
  or (_40868_, _13549_, _13548_);
  or (_13550_, _13522_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_13551_, _13550_, _13526_);
  and (_13552_, _12844_, _04823_);
  and (_13553_, _13552_, _12841_);
  or (_13554_, _13530_, _13553_);
  and (_13555_, _13554_, _13551_);
  and (_13556_, _13534_, _12852_);
  or (_40869_, _13556_, _13555_);
  or (_13557_, _13522_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_13558_, _13557_, _13526_);
  and (_13559_, _12049_, _04565_);
  nand (_13560_, _13559_, _12052_);
  or (_13561_, _13560_, _13054_);
  and (_13562_, _13561_, _13558_);
  and (_13563_, _13534_, _13062_);
  or (_40870_, _13563_, _13562_);
  or (_13564_, _13560_, _13256_);
  or (_13565_, _13522_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_13566_, _13565_, _13526_);
  and (_13567_, _13566_, _13564_);
  and (_13568_, _13534_, _13263_);
  or (_40871_, _13568_, _13567_);
  or (_13569_, _13522_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_13570_, _13569_, _13526_);
  and (_13571_, _13457_, _04823_);
  and (_13572_, _13571_, _13454_);
  or (_13573_, _13530_, _13572_);
  and (_13574_, _13573_, _13570_);
  and (_13575_, _13534_, _13465_);
  or (_40872_, _13575_, _13574_);
  or (_13576_, _13522_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_13577_, _13576_, _13526_);
  or (_13578_, _13560_, _06852_);
  and (_13579_, _13578_, _13577_);
  and (_13580_, _13534_, _06891_);
  or (_40874_, _13580_, _13579_);
  and (_13581_, _13520_, _04827_);
  or (_13582_, _13581_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_13583_, _12243_, _04569_);
  or (_13584_, _13583_, _12246_);
  and (_13585_, _13584_, _13582_);
  not (_13586_, _13581_);
  or (_13587_, _13586_, _13529_);
  and (_13588_, _13587_, _13585_);
  and (_13589_, _05177_, _04569_);
  and (_13590_, _13589_, _12232_);
  and (_13591_, _13590_, _12241_);
  or (_40878_, _13591_, _13588_);
  or (_13592_, _13581_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_13593_, _13592_, _13584_);
  or (_13594_, _13586_, _13539_);
  and (_13595_, _13594_, _13593_);
  and (_13596_, _13590_, _12440_);
  or (_40879_, _13596_, _13595_);
  or (_13597_, _13581_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_13598_, _13597_, _13584_);
  or (_13599_, _13586_, _13546_);
  and (_13600_, _13599_, _13598_);
  and (_13601_, _13590_, _12647_);
  or (_40880_, _13601_, _13600_);
  or (_13602_, _13581_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_13603_, _13602_, _13584_);
  or (_13604_, _13586_, _13553_);
  and (_13605_, _13604_, _13603_);
  and (_13606_, _13590_, _12852_);
  or (_40881_, _13606_, _13605_);
  or (_13607_, _13581_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_13608_, _13607_, _13584_);
  nand (_13609_, _12052_, _05187_);
  or (_13610_, _13609_, _13054_);
  and (_13611_, _13610_, _13608_);
  and (_13612_, _13590_, _13062_);
  or (_40882_, _13612_, _13611_);
  or (_13613_, _13581_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_13614_, _13613_, _13584_);
  and (_13615_, _13254_, _04823_);
  and (_13616_, _13615_, _13251_);
  or (_13617_, _13586_, _13616_);
  and (_13618_, _13617_, _13614_);
  and (_13619_, _13590_, _13263_);
  or (_40884_, _13619_, _13618_);
  or (_13620_, _13581_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_13621_, _13620_, _13584_);
  or (_13622_, _13586_, _13572_);
  and (_13623_, _13622_, _13621_);
  and (_13624_, _13590_, _13465_);
  or (_40885_, _13624_, _13623_);
  or (_13626_, _13581_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_13627_, _13626_, _13584_);
  or (_13628_, _13609_, _06852_);
  and (_13629_, _13628_, _13627_);
  and (_13630_, _13590_, _06891_);
  or (_40886_, _13630_, _13629_);
  and (_13631_, _12051_, _05004_);
  and (_13632_, _13631_, _12050_);
  not (_13633_, _13632_);
  or (_13635_, _13633_, _12229_);
  not (_13636_, _05172_);
  and (_13637_, _12231_, _13636_);
  and (_13638_, _13637_, _04570_);
  nor (_13639_, _13632_, \oc8051_golden_model_1.IRAM[4] [0]);
  nor (_13640_, _13639_, _13638_);
  and (_13641_, _13640_, _13635_);
  and (_13642_, _13638_, _12241_);
  or (_40890_, _13642_, _13641_);
  and (_13643_, _12244_, _13636_);
  nand (_13645_, _13643_, _04570_);
  nor (_13646_, _04824_, _04565_);
  nor (_13647_, _13646_, _04825_);
  and (_13648_, _05162_, _05004_);
  and (_13649_, _13648_, _13647_);
  or (_13650_, _13649_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_13651_, _13650_, _13645_);
  not (_13652_, _13649_);
  or (_13653_, _13652_, _13539_);
  and (_13654_, _13653_, _13651_);
  and (_13656_, _13638_, _12440_);
  or (_40891_, _13656_, _13654_);
  or (_13657_, _13649_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_13658_, _13657_, _13645_);
  or (_13659_, _13652_, _13546_);
  and (_13660_, _13659_, _13658_);
  and (_13661_, _13638_, _12647_);
  or (_40893_, _13661_, _13660_);
  or (_13662_, _13633_, _12846_);
  nor (_13663_, _13632_, \oc8051_golden_model_1.IRAM[4] [3]);
  nor (_13665_, _13663_, _13638_);
  and (_13666_, _13665_, _13662_);
  and (_13667_, _13638_, _12852_);
  or (_40894_, _13667_, _13666_);
  or (_13668_, _13649_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13669_, _13668_, _13645_);
  or (_13670_, _13633_, _13054_);
  and (_13671_, _13670_, _13669_);
  and (_13672_, _13638_, _13062_);
  or (_40895_, _13672_, _13671_);
  or (_13674_, _13649_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_13675_, _13674_, _13645_);
  or (_13676_, _13652_, _13616_);
  and (_13677_, _13676_, _13675_);
  and (_13678_, _13638_, _13263_);
  or (_40896_, _13678_, _13677_);
  or (_13679_, _13649_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13680_, _13679_, _13645_);
  or (_13681_, _13652_, _13572_);
  and (_13682_, _13681_, _13680_);
  and (_13684_, _13638_, _13465_);
  or (_40897_, _13684_, _13682_);
  or (_13685_, _13649_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13686_, _13685_, _13645_);
  or (_13687_, _13633_, _06852_);
  and (_13688_, _13687_, _13686_);
  and (_13689_, _13638_, _06891_);
  or (_40899_, _13689_, _13688_);
  and (_13690_, _13631_, _13472_);
  not (_13691_, _13690_);
  or (_13693_, _13691_, _12229_);
  and (_13694_, _13637_, _04887_);
  nor (_13695_, _13690_, \oc8051_golden_model_1.IRAM[5] [0]);
  nor (_13696_, _13695_, _13694_);
  and (_13697_, _13696_, _13693_);
  and (_13698_, _13694_, _12241_);
  or (_40902_, _13698_, _13697_);
  nand (_13699_, _13643_, _04887_);
  and (_13700_, _13646_, _04744_);
  and (_13701_, _13648_, _13700_);
  or (_13703_, _13701_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13704_, _13703_, _13699_);
  not (_13705_, _13701_);
  or (_13706_, _13705_, _13539_);
  and (_13707_, _13706_, _13704_);
  and (_13708_, _13694_, _12440_);
  or (_40904_, _13708_, _13707_);
  or (_13709_, _13701_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13710_, _13709_, _13699_);
  or (_13711_, _13705_, _13546_);
  and (_13713_, _13711_, _13710_);
  and (_13714_, _13694_, _12647_);
  or (_40905_, _13714_, _13713_);
  or (_13715_, _13691_, _12846_);
  nor (_13716_, _13690_, \oc8051_golden_model_1.IRAM[5] [3]);
  nor (_13717_, _13716_, _13694_);
  and (_13718_, _13717_, _13715_);
  and (_13719_, _13694_, _12852_);
  or (_40906_, _13719_, _13718_);
  or (_13720_, _13701_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13722_, _13720_, _13699_);
  or (_13723_, _13691_, _13054_);
  and (_13724_, _13723_, _13722_);
  and (_13725_, _13694_, _13062_);
  or (_40907_, _13725_, _13724_);
  or (_13726_, _13705_, _13616_);
  or (_13727_, _13701_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_13728_, _13727_, _13699_);
  and (_13729_, _13728_, _13726_);
  and (_13730_, _13694_, _13263_);
  or (_40908_, _13730_, _13729_);
  or (_13732_, _13701_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13733_, _13732_, _13699_);
  or (_13734_, _13705_, _13572_);
  and (_13735_, _13734_, _13733_);
  and (_13736_, _13694_, _13465_);
  or (_40910_, _13736_, _13735_);
  or (_13737_, _13701_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_13738_, _13737_, _13699_);
  or (_13739_, _13691_, _06852_);
  and (_13741_, _13739_, _13738_);
  and (_13742_, _13694_, _06891_);
  or (_40911_, _13742_, _13741_);
  and (_13743_, _13631_, _13559_);
  not (_13744_, _13743_);
  or (_13745_, _13744_, _12229_);
  and (_13746_, _13643_, _06009_);
  not (_13747_, _13746_);
  or (_13748_, _13743_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_13749_, _13748_, _13747_);
  and (_13751_, _13749_, _13745_);
  and (_13752_, _13746_, _12241_);
  or (_40914_, _13752_, _13751_);
  and (_13753_, _13648_, _13521_);
  or (_13754_, _13753_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_13755_, _13754_, _13747_);
  not (_13756_, _13753_);
  or (_13757_, _13756_, _13539_);
  and (_13758_, _13757_, _13755_);
  and (_13759_, _13746_, _12440_);
  or (_40916_, _13759_, _13758_);
  or (_13760_, _13753_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_13761_, _13760_, _13747_);
  or (_13762_, _13756_, _13546_);
  and (_13763_, _13762_, _13761_);
  and (_13764_, _13746_, _12647_);
  or (_40917_, _13764_, _13763_);
  or (_13765_, _13744_, _12846_);
  or (_13766_, _13743_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_13767_, _13766_, _13747_);
  and (_13768_, _13767_, _13765_);
  and (_13769_, _13746_, _12852_);
  or (_40918_, _13769_, _13768_);
  or (_13770_, _13753_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13771_, _13770_, _13747_);
  or (_13772_, _13744_, _13054_);
  and (_13773_, _13772_, _13771_);
  and (_13774_, _13746_, _13062_);
  or (_40919_, _13774_, _13773_);
  or (_13775_, _13753_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_13776_, _13775_, _13747_);
  or (_13777_, _13756_, _13616_);
  and (_13778_, _13777_, _13776_);
  and (_13779_, _13746_, _13263_);
  or (_40920_, _13779_, _13778_);
  or (_13780_, _13753_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13781_, _13780_, _13747_);
  or (_13782_, _13756_, _13572_);
  and (_13783_, _13782_, _13781_);
  and (_13784_, _13746_, _13465_);
  or (_40922_, _13784_, _13783_);
  or (_13785_, _13753_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13786_, _13785_, _13747_);
  or (_13787_, _13744_, _06852_);
  and (_13788_, _13787_, _13786_);
  and (_13789_, _13746_, _06891_);
  or (_40923_, _13789_, _13788_);
  and (_13790_, _13631_, _05187_);
  not (_13791_, _13790_);
  or (_13792_, _13791_, _12229_);
  and (_13793_, _13637_, _04569_);
  nor (_13794_, _13790_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_13795_, _13794_, _13793_);
  and (_13796_, _13795_, _13792_);
  and (_13797_, _13793_, _12241_);
  or (_40927_, _13797_, _13796_);
  nand (_13798_, _13643_, _04569_);
  and (_13799_, _13648_, _04827_);
  or (_13800_, _13799_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_13801_, _13800_, _13798_);
  not (_13802_, _13799_);
  or (_13803_, _13802_, _13539_);
  and (_13804_, _13803_, _13801_);
  and (_13805_, _13793_, _12440_);
  or (_40928_, _13805_, _13804_);
  or (_13806_, _13799_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_13807_, _13806_, _13798_);
  or (_13808_, _13802_, _13546_);
  and (_13809_, _13808_, _13807_);
  and (_13810_, _13793_, _12647_);
  or (_40929_, _13810_, _13809_);
  or (_13811_, _13791_, _12846_);
  nor (_13812_, _13790_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_13813_, _13812_, _13793_);
  and (_13814_, _13813_, _13811_);
  and (_13815_, _13793_, _12852_);
  or (_40930_, _13815_, _13814_);
  or (_13816_, _13799_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13817_, _13816_, _13798_);
  or (_13818_, _13791_, _13054_);
  and (_13819_, _13818_, _13817_);
  and (_13820_, _13793_, _13062_);
  or (_40931_, _13820_, _13819_);
  or (_13821_, _13799_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_13822_, _13821_, _13798_);
  or (_13823_, _13802_, _13616_);
  and (_13824_, _13823_, _13822_);
  and (_13825_, _13793_, _13263_);
  or (_40933_, _13825_, _13824_);
  or (_13826_, _13799_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13827_, _13826_, _13798_);
  or (_13828_, _13802_, _13572_);
  and (_13829_, _13828_, _13827_);
  and (_13830_, _13793_, _13465_);
  or (_40934_, _13830_, _13829_);
  or (_13831_, _13799_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13832_, _13831_, _13798_);
  or (_13833_, _13791_, _06852_);
  and (_13834_, _13833_, _13832_);
  and (_13835_, _13793_, _06891_);
  or (_40935_, _13835_, _13834_);
  and (_13836_, _05189_, _05161_);
  and (_13837_, _13836_, _12050_);
  or (_13838_, _13837_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_13839_, _05169_);
  and (_13840_, _05178_, _13839_);
  and (_13841_, _13840_, _04570_);
  not (_13842_, _13841_);
  and (_13843_, _13842_, _13838_);
  not (_13844_, _13837_);
  or (_13845_, _13844_, _12229_);
  and (_13846_, _13845_, _13843_);
  and (_13847_, _13841_, _12241_);
  or (_40939_, _13847_, _13846_);
  or (_13848_, _13837_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13849_, _13848_, _13842_);
  or (_13850_, _13844_, _12434_);
  and (_13851_, _13850_, _13849_);
  and (_13852_, _13841_, _12440_);
  or (_40940_, _13852_, _13851_);
  or (_13853_, _13837_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13854_, _13853_, _13842_);
  or (_13855_, _13844_, _12641_);
  and (_13856_, _13855_, _13854_);
  and (_13857_, _13841_, _12647_);
  or (_40942_, _13857_, _13856_);
  or (_13858_, _13844_, _12846_);
  or (_13859_, _13837_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13860_, _13859_, _13842_);
  and (_13861_, _13860_, _13858_);
  and (_13862_, _13841_, _12852_);
  or (_40943_, _13862_, _13861_);
  or (_13863_, _13837_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13864_, _13863_, _13842_);
  or (_13865_, _13844_, _13054_);
  and (_13866_, _13865_, _13864_);
  and (_13867_, _13841_, _13062_);
  or (_40944_, _13867_, _13866_);
  or (_13868_, _13837_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13869_, _13868_, _13842_);
  or (_13870_, _13844_, _13256_);
  and (_13871_, _13870_, _13869_);
  and (_13872_, _13841_, _13263_);
  or (_40945_, _13872_, _13871_);
  or (_13873_, _13837_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13874_, _13873_, _13842_);
  or (_13875_, _13844_, _13459_);
  and (_13876_, _13875_, _13874_);
  and (_13877_, _13841_, _13465_);
  or (_40946_, _13877_, _13876_);
  or (_13878_, _13837_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_13879_, _13878_, _13842_);
  or (_13880_, _13844_, _06852_);
  and (_13881_, _13880_, _13879_);
  and (_13882_, _13841_, _06891_);
  or (_40948_, _13882_, _13881_);
  and (_13883_, _13836_, _13472_);
  or (_13884_, _13883_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_13885_, _12245_, _04888_);
  and (_13886_, _13885_, _13884_);
  not (_13887_, _13883_);
  or (_13888_, _13887_, _12229_);
  and (_13889_, _13888_, _13886_);
  and (_13890_, _13840_, _04887_);
  and (_13891_, _13890_, _12241_);
  or (_40951_, _13891_, _13889_);
  or (_13892_, _13883_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13893_, _13892_, _13885_);
  or (_13894_, _13887_, _12434_);
  and (_13895_, _13894_, _13893_);
  and (_13896_, _13890_, _12440_);
  or (_40953_, _13896_, _13895_);
  or (_13897_, _13883_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13898_, _13897_, _13885_);
  or (_13899_, _13887_, _12641_);
  and (_13900_, _13899_, _13898_);
  and (_13901_, _13890_, _12647_);
  or (_40954_, _13901_, _13900_);
  or (_13902_, _13887_, _12846_);
  nor (_13903_, _13883_, \oc8051_golden_model_1.IRAM[9] [3]);
  nor (_13904_, _13903_, _13890_);
  and (_13905_, _13904_, _13902_);
  and (_13906_, _13890_, _12852_);
  or (_40955_, _13906_, _13905_);
  or (_13907_, _13883_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13908_, _13907_, _13885_);
  or (_13909_, _13887_, _13054_);
  and (_13910_, _13909_, _13908_);
  and (_13911_, _13890_, _13062_);
  or (_40956_, _13911_, _13910_);
  or (_13912_, _13883_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_13913_, _13912_, _13885_);
  or (_13914_, _13887_, _13256_);
  and (_13915_, _13914_, _13913_);
  and (_13916_, _13890_, _13263_);
  or (_40957_, _13916_, _13915_);
  or (_13917_, _13883_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13918_, _13917_, _13885_);
  or (_13919_, _13887_, _13459_);
  and (_13920_, _13919_, _13918_);
  and (_13921_, _13890_, _13465_);
  or (_40959_, _13921_, _13920_);
  or (_13922_, _13883_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13923_, _13922_, _13885_);
  or (_13924_, _13887_, _06852_);
  and (_13925_, _13924_, _13923_);
  and (_13926_, _13890_, _06891_);
  or (_40960_, _13926_, _13925_);
  and (_13927_, _13836_, _13559_);
  not (_13928_, _13927_);
  or (_13929_, _13928_, _12229_);
  or (_13930_, _13927_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13931_, _13840_, _06009_);
  not (_13932_, _13931_);
  and (_13933_, _13932_, _13930_);
  and (_13934_, _13933_, _13929_);
  and (_13935_, _13931_, _12241_);
  or (_40963_, _13935_, _13934_);
  or (_13936_, _13927_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13937_, _13936_, _13932_);
  or (_13938_, _13928_, _12434_);
  and (_13939_, _13938_, _13937_);
  and (_13940_, _13931_, _12440_);
  or (_40965_, _13940_, _13939_);
  or (_13941_, _13927_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13942_, _13941_, _13932_);
  or (_13943_, _13928_, _12641_);
  and (_13944_, _13943_, _13942_);
  and (_13945_, _13931_, _12647_);
  or (_40966_, _13945_, _13944_);
  or (_13946_, _13928_, _12846_);
  or (_13947_, _13927_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13948_, _13947_, _13932_);
  and (_13949_, _13948_, _13946_);
  and (_13950_, _13931_, _12852_);
  or (_40967_, _13950_, _13949_);
  or (_13951_, _13927_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13952_, _13951_, _13932_);
  or (_13953_, _13928_, _13054_);
  and (_13954_, _13953_, _13952_);
  and (_13955_, _13931_, _13062_);
  or (_40968_, _13955_, _13954_);
  or (_13956_, _13927_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13957_, _13956_, _13932_);
  or (_13958_, _13928_, _13256_);
  and (_13959_, _13958_, _13957_);
  and (_13960_, _13931_, _13263_);
  or (_40969_, _13960_, _13959_);
  or (_13961_, _13927_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13962_, _13961_, _13932_);
  or (_13963_, _13928_, _13459_);
  and (_13964_, _13963_, _13962_);
  and (_13965_, _13931_, _13465_);
  or (_40971_, _13965_, _13964_);
  or (_13966_, _13928_, _06852_);
  or (_13967_, _13927_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13968_, _13967_, _13932_);
  and (_13969_, _13968_, _13966_);
  and (_13970_, _13931_, _06891_);
  or (_40972_, _13970_, _13969_);
  and (_13971_, _13836_, _05187_);
  not (_13972_, _13971_);
  or (_13973_, _13972_, _12229_);
  or (_13974_, _13971_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13975_, _13840_, _04569_);
  not (_13976_, _13975_);
  and (_13977_, _13976_, _13974_);
  and (_13978_, _13977_, _13973_);
  and (_13979_, _13975_, _12241_);
  or (_40976_, _13979_, _13978_);
  or (_13980_, _13971_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13981_, _13980_, _13976_);
  or (_13982_, _13972_, _12434_);
  and (_13983_, _13982_, _13981_);
  and (_13984_, _13975_, _12440_);
  or (_40977_, _13984_, _13983_);
  or (_13985_, _13971_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13986_, _13985_, _13976_);
  or (_13987_, _13972_, _12641_);
  and (_13988_, _13987_, _13986_);
  and (_13989_, _13975_, _12647_);
  or (_40978_, _13989_, _13988_);
  or (_13990_, _13972_, _12846_);
  or (_13991_, _13971_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13992_, _13991_, _13976_);
  and (_13993_, _13992_, _13990_);
  and (_13994_, _13975_, _12852_);
  or (_40979_, _13994_, _13993_);
  or (_13995_, _13971_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13996_, _13995_, _13976_);
  or (_13997_, _13972_, _13054_);
  and (_13998_, _13997_, _13996_);
  and (_13999_, _13975_, _13062_);
  or (_40980_, _13999_, _13998_);
  or (_14000_, _13971_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_14001_, _14000_, _13976_);
  or (_14002_, _13972_, _13256_);
  and (_14003_, _14002_, _14001_);
  and (_14004_, _13975_, _13263_);
  or (_40982_, _14004_, _14003_);
  or (_14005_, _13971_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_14006_, _14005_, _13976_);
  or (_14007_, _13972_, _13459_);
  and (_14008_, _14007_, _14006_);
  and (_14009_, _13975_, _13465_);
  or (_40983_, _14009_, _14008_);
  or (_14010_, _13971_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_14011_, _14010_, _13976_);
  or (_14012_, _13972_, _06852_);
  and (_14013_, _14012_, _14011_);
  and (_14014_, _13975_, _06891_);
  or (_40984_, _14014_, _14013_);
  and (_14015_, _12050_, _05190_);
  not (_14016_, _14015_);
  or (_14017_, _14016_, _12229_);
  and (_14018_, _05179_, _04570_);
  not (_14019_, _14018_);
  or (_14020_, _14015_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_14021_, _14020_, _14019_);
  and (_14022_, _14021_, _14017_);
  and (_14023_, _14018_, _12241_);
  or (_40988_, _14023_, _14022_);
  and (_14024_, _13647_, _05164_);
  or (_14025_, _14024_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_14026_, _14025_, _14019_);
  not (_14027_, _14024_);
  or (_14028_, _14027_, _13539_);
  and (_14029_, _14028_, _14026_);
  and (_14030_, _14018_, _12440_);
  or (_40989_, _14030_, _14029_);
  or (_14031_, _14024_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_14032_, _14031_, _14019_);
  or (_14033_, _14027_, _13546_);
  and (_14034_, _14033_, _14032_);
  and (_14035_, _14018_, _12647_);
  or (_40990_, _14035_, _14034_);
  or (_14036_, _14016_, _12846_);
  or (_14037_, _14015_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_14038_, _14037_, _14019_);
  and (_14039_, _14038_, _14036_);
  and (_14040_, _14018_, _12852_);
  or (_40991_, _14040_, _14039_);
  or (_14041_, _14024_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_14042_, _14041_, _14019_);
  or (_14043_, _14016_, _13054_);
  and (_14044_, _14043_, _14042_);
  and (_14045_, _14018_, _13062_);
  or (_40993_, _14045_, _14044_);
  or (_14046_, _14024_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_14047_, _14046_, _14019_);
  or (_14048_, _14027_, _13616_);
  and (_14049_, _14048_, _14047_);
  and (_14050_, _14018_, _13263_);
  or (_40994_, _14050_, _14049_);
  or (_14051_, _14024_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_14052_, _14051_, _14019_);
  or (_14053_, _14027_, _13572_);
  and (_14054_, _14053_, _14052_);
  and (_14055_, _14018_, _13465_);
  or (_40995_, _14055_, _14054_);
  or (_14056_, _14024_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_14057_, _14056_, _14019_);
  or (_14058_, _14016_, _06852_);
  and (_14059_, _14058_, _14057_);
  and (_14060_, _14018_, _06891_);
  or (_40996_, _14060_, _14059_);
  and (_14061_, _13472_, _05190_);
  not (_14062_, _14061_);
  or (_14063_, _14062_, _12229_);
  and (_14064_, _05179_, _04887_);
  not (_14065_, _14064_);
  or (_14066_, _14061_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_14067_, _14066_, _14065_);
  and (_14068_, _14067_, _14063_);
  and (_14069_, _14064_, _12241_);
  or (_41000_, _14069_, _14068_);
  and (_14070_, _13700_, _05164_);
  or (_14071_, _14070_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_14072_, _14071_, _14065_);
  not (_14073_, _14070_);
  or (_14074_, _14073_, _13539_);
  and (_14075_, _14074_, _14072_);
  and (_14076_, _14064_, _12440_);
  or (_41001_, _14076_, _14075_);
  or (_14077_, _14070_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_14078_, _14077_, _14065_);
  or (_14079_, _14073_, _13546_);
  and (_14080_, _14079_, _14078_);
  and (_14081_, _14064_, _12647_);
  or (_41002_, _14081_, _14080_);
  or (_14082_, _14062_, _12846_);
  or (_14083_, _14061_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_14084_, _14083_, _14065_);
  and (_14085_, _14084_, _14082_);
  and (_14086_, _14064_, _12852_);
  or (_41004_, _14086_, _14085_);
  or (_14087_, _14070_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_14088_, _14087_, _14065_);
  or (_14089_, _14062_, _13054_);
  and (_14090_, _14089_, _14088_);
  and (_14091_, _14064_, _13062_);
  or (_41005_, _14091_, _14090_);
  or (_14092_, _14070_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_14093_, _14092_, _14065_);
  or (_14094_, _14073_, _13616_);
  and (_14095_, _14094_, _14093_);
  and (_14096_, _14064_, _13263_);
  or (_41006_, _14096_, _14095_);
  or (_14097_, _14070_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_14098_, _14097_, _14065_);
  or (_14099_, _14073_, _13572_);
  and (_14100_, _14099_, _14098_);
  and (_14101_, _14064_, _13465_);
  or (_41007_, _14101_, _14100_);
  or (_14102_, _14070_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_14103_, _14102_, _14065_);
  or (_14104_, _14062_, _06852_);
  and (_14105_, _14104_, _14103_);
  and (_14106_, _14064_, _06891_);
  or (_41008_, _14106_, _14105_);
  and (_14107_, _13559_, _05190_);
  not (_14108_, _14107_);
  or (_14109_, _14108_, _12229_);
  and (_14110_, _06009_, _05179_);
  not (_14111_, _14110_);
  or (_14112_, _14107_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_14113_, _14112_, _14111_);
  and (_14114_, _14113_, _14109_);
  and (_14115_, _14110_, _12241_);
  or (_41012_, _14115_, _14114_);
  and (_14116_, _13521_, _05164_);
  or (_14117_, _14116_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_14118_, _14117_, _14111_);
  not (_14119_, _14116_);
  or (_14120_, _14119_, _13539_);
  and (_14121_, _14120_, _14118_);
  and (_14122_, _14110_, _12440_);
  or (_41013_, _14122_, _14121_);
  or (_14123_, _14116_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_14124_, _14123_, _14111_);
  or (_14125_, _14119_, _13546_);
  and (_14126_, _14125_, _14124_);
  and (_14127_, _14110_, _12647_);
  or (_41014_, _14127_, _14126_);
  or (_14128_, _14108_, _12846_);
  or (_14129_, _14107_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_14130_, _14129_, _14111_);
  and (_14131_, _14130_, _14128_);
  and (_14132_, _14110_, _12852_);
  or (_41016_, _14132_, _14131_);
  or (_14133_, _14116_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_14134_, _14133_, _14111_);
  or (_14135_, _14108_, _13054_);
  and (_14136_, _14135_, _14134_);
  and (_14137_, _14110_, _13062_);
  or (_41017_, _14137_, _14136_);
  or (_14138_, _14116_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_14139_, _14138_, _14111_);
  or (_14140_, _14119_, _13616_);
  and (_14141_, _14140_, _14139_);
  and (_14142_, _14110_, _13263_);
  or (_41018_, _14142_, _14141_);
  or (_14143_, _14116_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_14144_, _14143_, _14111_);
  or (_14145_, _14119_, _13572_);
  and (_14146_, _14145_, _14144_);
  and (_14147_, _14110_, _13465_);
  or (_41019_, _14147_, _14146_);
  or (_14148_, _14116_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_14149_, _14148_, _14111_);
  or (_14150_, _14108_, _06852_);
  and (_14151_, _14150_, _14149_);
  and (_14152_, _14110_, _06891_);
  or (_41020_, _14152_, _14151_);
  or (_14153_, _12229_, _05192_);
  or (_14154_, _05191_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_14155_, _14154_, _05181_);
  and (_14156_, _14155_, _14153_);
  and (_14157_, _12241_, _05180_);
  or (_41024_, _14157_, _14156_);
  or (_14158_, _05165_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_14159_, _14158_, _05181_);
  not (_14160_, _05165_);
  or (_14161_, _13539_, _14160_);
  and (_14162_, _14161_, _14159_);
  and (_14163_, _12440_, _05180_);
  or (_41025_, _14163_, _14162_);
  or (_14164_, _05165_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_14165_, _14164_, _05181_);
  or (_14166_, _13546_, _14160_);
  and (_14167_, _14166_, _14165_);
  and (_14168_, _12647_, _05180_);
  or (_41026_, _14168_, _14167_);
  or (_14169_, _12846_, _05192_);
  or (_14170_, _05191_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_14171_, _14170_, _05181_);
  and (_14172_, _14171_, _14169_);
  and (_14173_, _12852_, _05180_);
  or (_41028_, _14173_, _14172_);
  or (_14174_, _05165_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_14175_, _14174_, _05181_);
  or (_14176_, _13054_, _05192_);
  and (_14177_, _14176_, _14175_);
  and (_14178_, _13062_, _05180_);
  or (_41029_, _14178_, _14177_);
  or (_14179_, _05165_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_14180_, _14179_, _05181_);
  or (_14181_, _13616_, _14160_);
  and (_14182_, _14181_, _14180_);
  and (_14183_, _13263_, _05180_);
  or (_41030_, _14183_, _14182_);
  or (_14184_, _05165_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_14185_, _14184_, _05181_);
  or (_14186_, _13572_, _14160_);
  and (_14187_, _14186_, _14185_);
  and (_14188_, _13465_, _05180_);
  or (_41031_, _14188_, _14187_);
  nor (_14189_, _43189_, _07480_);
  nor (_14190_, _05306_, _07480_);
  and (_14191_, _12183_, _05306_);
  or (_14192_, _14191_, _14190_);
  and (_14193_, _14192_, _03744_);
  nor (_14194_, _05722_, _06896_);
  or (_14195_, _14194_, _14190_);
  or (_14196_, _14195_, _04432_);
  and (_14197_, _05306_, \oc8051_golden_model_1.ACC [0]);
  or (_14198_, _14197_, _14190_);
  and (_14199_, _14198_, _04436_);
  nor (_14200_, _04436_, _07480_);
  or (_14201_, _14200_, _03534_);
  or (_14202_, _14201_, _14199_);
  and (_14203_, _14202_, _03470_);
  and (_14204_, _14203_, _14196_);
  and (_14205_, _12075_, _05929_);
  nor (_14206_, _05929_, _07480_);
  or (_14207_, _14206_, _14205_);
  and (_14208_, _14207_, _03469_);
  or (_14209_, _14208_, _14204_);
  and (_14210_, _14209_, _04457_);
  and (_14211_, _05306_, _04429_);
  or (_14212_, _14211_, _14190_);
  and (_14213_, _14212_, _03527_);
  or (_14214_, _14213_, _03530_);
  or (_14215_, _14214_, _14210_);
  or (_14216_, _14198_, _03531_);
  and (_14217_, _14216_, _03466_);
  and (_14218_, _14217_, _14215_);
  and (_14219_, _14190_, _03465_);
  or (_14220_, _14219_, _03458_);
  or (_14221_, _14220_, _14218_);
  or (_14222_, _14195_, _03459_);
  and (_14223_, _14222_, _14221_);
  or (_14224_, _14223_, _06933_);
  nor (_14225_, _07414_, _07412_);
  nor (_14226_, _14225_, _07415_);
  or (_14227_, _14226_, _07447_);
  and (_14228_, _14227_, _03453_);
  and (_14229_, _14228_, _14224_);
  nor (_14230_, _12106_, _07455_);
  or (_14231_, _14230_, _14206_);
  and (_14232_, _14231_, _03452_);
  or (_14233_, _14232_, _07454_);
  or (_14234_, _14233_, _14229_);
  or (_14235_, _14212_, _06903_);
  and (_14236_, _14235_, _04500_);
  and (_14237_, _14236_, _14234_);
  and (_14238_, _06617_, _05306_);
  or (_14239_, _14238_, _14190_);
  and (_14240_, _14239_, _04082_);
  or (_14241_, _14240_, _03224_);
  or (_14242_, _14241_, _14237_);
  nor (_14243_, _12164_, _06896_);
  or (_14244_, _14190_, _03521_);
  or (_14245_, _14244_, _14243_);
  and (_14246_, _14245_, _07474_);
  and (_14247_, _14246_, _14242_);
  nand (_14248_, _07827_, _03344_);
  or (_14249_, _07802_, _07791_);
  or (_14250_, _07827_, _14249_);
  and (_14251_, _14250_, _07468_);
  and (_14252_, _14251_, _14248_);
  or (_14253_, _14252_, _08905_);
  or (_14254_, _14253_, _14247_);
  and (_14255_, _12177_, _05306_);
  or (_14256_, _14190_, _04527_);
  or (_14257_, _14256_, _14255_);
  and (_14258_, _05306_, _06350_);
  or (_14259_, _14258_, _14190_);
  or (_14260_, _14259_, _04509_);
  and (_14261_, _14260_, _03745_);
  and (_14262_, _14261_, _14257_);
  and (_14263_, _14262_, _14254_);
  or (_14264_, _14263_, _14193_);
  and (_14265_, _14264_, _04523_);
  nand (_14266_, _14259_, _03611_);
  nor (_14267_, _14266_, _14194_);
  or (_14268_, _14267_, _14265_);
  and (_14269_, _14268_, _03734_);
  or (_14270_, _14190_, _05722_);
  and (_14271_, _14198_, _03733_);
  and (_14272_, _14271_, _14270_);
  or (_14273_, _14272_, _03618_);
  or (_14274_, _14273_, _14269_);
  nor (_14275_, _12057_, _06896_);
  or (_14276_, _14190_, _06453_);
  or (_14277_, _14276_, _14275_);
  and (_14278_, _14277_, _06458_);
  and (_14279_, _14278_, _14274_);
  nor (_14280_, _12181_, _06896_);
  or (_14281_, _14280_, _14190_);
  and (_14282_, _14281_, _03741_);
  or (_14283_, _14282_, _03767_);
  or (_14284_, _14283_, _14279_);
  or (_14285_, _14195_, _03948_);
  and (_14286_, _14285_, _03446_);
  and (_14287_, _14286_, _14284_);
  and (_14288_, _14190_, _03445_);
  or (_14289_, _14288_, _03473_);
  or (_14290_, _14289_, _14287_);
  or (_14291_, _14195_, _03474_);
  and (_14292_, _14291_, _43189_);
  and (_14293_, _14292_, _14290_);
  or (_14294_, _14293_, _14189_);
  and (_43732_, _14294_, _42003_);
  nor (_14295_, _43189_, _07475_);
  or (_14296_, _05306_, \oc8051_golden_model_1.B [1]);
  and (_14297_, _12265_, _05306_);
  not (_14298_, _14297_);
  and (_14299_, _14298_, _14296_);
  or (_14300_, _14299_, _04432_);
  nand (_14301_, _05306_, _03269_);
  and (_14302_, _14301_, _14296_);
  and (_14303_, _14302_, _04436_);
  nor (_14304_, _04436_, _07475_);
  or (_14305_, _14304_, _03534_);
  or (_14306_, _14305_, _14303_);
  and (_14307_, _14306_, _03470_);
  and (_14308_, _14307_, _14300_);
  and (_14309_, _12269_, _05929_);
  nor (_14310_, _05929_, _07475_);
  or (_14311_, _14310_, _03527_);
  or (_14312_, _14311_, _14309_);
  and (_14313_, _14312_, _03533_);
  or (_14314_, _14313_, _14308_);
  nor (_14315_, _05306_, _07475_);
  nor (_14316_, _06896_, _04635_);
  or (_14317_, _14316_, _14315_);
  or (_14318_, _14317_, _04457_);
  and (_14319_, _14318_, _14314_);
  or (_14320_, _14319_, _03530_);
  or (_14321_, _14302_, _03531_);
  and (_14322_, _14321_, _03466_);
  and (_14323_, _14322_, _14320_);
  and (_14324_, _12256_, _05929_);
  or (_14325_, _14324_, _14310_);
  and (_14326_, _14325_, _03465_);
  or (_14327_, _14326_, _14323_);
  and (_14328_, _14327_, _03459_);
  and (_14329_, _14309_, _12284_);
  or (_14330_, _14329_, _14310_);
  and (_14331_, _14330_, _03458_);
  or (_14332_, _14331_, _06933_);
  or (_14333_, _14332_, _14328_);
  or (_14334_, _07359_, _07358_);
  nand (_14335_, _14334_, _07416_);
  or (_14336_, _14334_, _07416_);
  and (_14337_, _14336_, _14335_);
  or (_14338_, _14337_, _07447_);
  and (_14339_, _14338_, _03453_);
  and (_14340_, _14339_, _14333_);
  nor (_14341_, _12301_, _07455_);
  or (_14342_, _14341_, _14310_);
  and (_14343_, _14342_, _03452_);
  or (_14344_, _14343_, _07454_);
  or (_14345_, _14344_, _14340_);
  or (_14346_, _14317_, _06903_);
  and (_14347_, _14346_, _14345_);
  or (_14348_, _14347_, _04082_);
  and (_14349_, _06572_, _05306_);
  or (_14350_, _14315_, _04500_);
  or (_14351_, _14350_, _14349_);
  and (_14352_, _14351_, _03521_);
  and (_14353_, _14352_, _14348_);
  nand (_14354_, _12360_, _05306_);
  and (_14355_, _14296_, _03224_);
  and (_14356_, _14355_, _14354_);
  or (_14357_, _14356_, _07468_);
  or (_14358_, _14357_, _14353_);
  nor (_14359_, _07803_, _07801_);
  or (_14360_, _14359_, _07804_);
  nor (_14361_, _14360_, _07827_);
  and (_14362_, _07827_, _07798_);
  or (_14363_, _14362_, _14361_);
  or (_14364_, _14363_, _07474_);
  and (_14365_, _14364_, _04509_);
  and (_14366_, _14365_, _14358_);
  nand (_14367_, _05306_, _04325_);
  and (_14368_, _14367_, _03624_);
  and (_14369_, _14368_, _14296_);
  or (_14370_, _14369_, _14366_);
  and (_14371_, _14370_, _04527_);
  or (_14372_, _12375_, _06896_);
  and (_14373_, _14296_, _03623_);
  and (_14374_, _14373_, _14372_);
  or (_14375_, _14374_, _14371_);
  and (_14376_, _14375_, _03745_);
  or (_14377_, _12381_, _06896_);
  and (_14378_, _14296_, _03744_);
  and (_14379_, _14378_, _14377_);
  or (_14380_, _14379_, _14376_);
  and (_14381_, _14380_, _04523_);
  or (_14382_, _12374_, _06896_);
  and (_14383_, _14296_, _03611_);
  and (_14384_, _14383_, _14382_);
  or (_14385_, _14384_, _14381_);
  and (_14386_, _14385_, _03734_);
  or (_14387_, _14315_, _05674_);
  and (_14388_, _14302_, _03733_);
  and (_14389_, _14388_, _14387_);
  or (_14390_, _14389_, _14386_);
  and (_14391_, _14390_, _03742_);
  or (_14392_, _14367_, _05674_);
  and (_14393_, _14296_, _03618_);
  and (_14394_, _14393_, _14392_);
  or (_14395_, _14301_, _05674_);
  and (_14396_, _14296_, _03741_);
  and (_14397_, _14396_, _14395_);
  or (_14398_, _14397_, _03767_);
  or (_14399_, _14398_, _14394_);
  or (_14400_, _14399_, _14391_);
  or (_14401_, _14299_, _03948_);
  and (_14402_, _14401_, _03446_);
  and (_14403_, _14402_, _14400_);
  and (_14404_, _14325_, _03445_);
  or (_14405_, _14404_, _03473_);
  or (_14406_, _14405_, _14403_);
  or (_14407_, _14315_, _03474_);
  or (_14408_, _14407_, _14297_);
  and (_14409_, _14408_, _43189_);
  and (_14410_, _14409_, _14406_);
  or (_14411_, _14410_, _14295_);
  and (_43733_, _14411_, _42003_);
  nor (_14412_, _43189_, _07528_);
  nor (_14413_, _05306_, _07528_);
  nor (_14414_, _06896_, _05073_);
  or (_14415_, _14414_, _14413_);
  or (_14416_, _14415_, _06903_);
  and (_14417_, _12462_, _05929_);
  and (_14418_, _14417_, _12491_);
  nor (_14419_, _05929_, _07528_);
  or (_14420_, _14419_, _03459_);
  or (_14421_, _14420_, _14418_);
  or (_14422_, _14415_, _04457_);
  nor (_14423_, _12467_, _06896_);
  or (_14424_, _14423_, _14413_);
  or (_14425_, _14424_, _04432_);
  and (_14426_, _05306_, \oc8051_golden_model_1.ACC [2]);
  or (_14427_, _14426_, _14413_);
  and (_14428_, _14427_, _04436_);
  nor (_14429_, _04436_, _07528_);
  or (_14430_, _14429_, _03534_);
  or (_14431_, _14430_, _14428_);
  and (_14432_, _14431_, _03470_);
  and (_14433_, _14432_, _14425_);
  or (_14434_, _14419_, _14417_);
  and (_14435_, _14434_, _03469_);
  or (_14436_, _14435_, _03527_);
  or (_14437_, _14436_, _14433_);
  and (_14438_, _14437_, _14422_);
  or (_14439_, _14438_, _03530_);
  or (_14440_, _14427_, _03531_);
  and (_14441_, _14440_, _03466_);
  and (_14442_, _14441_, _14439_);
  and (_14443_, _12460_, _05929_);
  or (_14444_, _14443_, _14419_);
  and (_14445_, _14444_, _03465_);
  or (_14446_, _14445_, _03458_);
  or (_14447_, _14446_, _14442_);
  and (_14448_, _14447_, _14421_);
  or (_14449_, _14448_, _06933_);
  nor (_14450_, _07418_, _07315_);
  nor (_14451_, _14450_, _07419_);
  or (_14452_, _14451_, _07447_);
  and (_14453_, _14452_, _03453_);
  and (_14454_, _14453_, _14449_);
  nor (_14455_, _12509_, _07455_);
  or (_14456_, _14455_, _14419_);
  and (_14457_, _14456_, _03452_);
  or (_14458_, _14457_, _07454_);
  or (_14459_, _14458_, _14454_);
  and (_14460_, _14459_, _14416_);
  or (_14461_, _14460_, _04082_);
  and (_14462_, _06710_, _05306_);
  or (_14463_, _14413_, _04500_);
  or (_14464_, _14463_, _14462_);
  and (_14465_, _14464_, _14461_);
  or (_14466_, _14465_, _03224_);
  nor (_14467_, _12568_, _06896_);
  or (_14468_, _14413_, _03521_);
  or (_14469_, _14468_, _14467_);
  and (_14470_, _14469_, _07474_);
  and (_14471_, _14470_, _14466_);
  nand (_14472_, _07827_, _07786_);
  nor (_14473_, _07804_, _07799_);
  not (_14474_, _14473_);
  and (_14475_, _14474_, _07789_);
  nor (_14476_, _14474_, _07789_);
  nor (_14477_, _14476_, _14475_);
  or (_14478_, _14477_, _07827_);
  and (_14479_, _14478_, _07468_);
  and (_14480_, _14479_, _14472_);
  or (_14481_, _14480_, _08905_);
  or (_14482_, _14481_, _14471_);
  and (_14483_, _12582_, _05306_);
  or (_14484_, _14413_, _04527_);
  or (_14485_, _14484_, _14483_);
  and (_14486_, _05306_, _06399_);
  or (_14487_, _14486_, _14413_);
  or (_14488_, _14487_, _04509_);
  and (_14489_, _14488_, _03745_);
  and (_14490_, _14489_, _14485_);
  and (_14491_, _14490_, _14482_);
  and (_14492_, _12588_, _05306_);
  or (_14493_, _14492_, _14413_);
  and (_14494_, _14493_, _03744_);
  or (_14495_, _14494_, _14491_);
  and (_14496_, _14495_, _04523_);
  or (_14497_, _14413_, _05772_);
  and (_14498_, _14487_, _03611_);
  and (_14499_, _14498_, _14497_);
  or (_14500_, _14499_, _14496_);
  and (_14501_, _14500_, _03734_);
  and (_14502_, _14427_, _03733_);
  and (_14503_, _14502_, _14497_);
  or (_14504_, _14503_, _03618_);
  or (_14505_, _14504_, _14501_);
  nor (_14506_, _12581_, _06896_);
  or (_14507_, _14413_, _06453_);
  or (_14508_, _14507_, _14506_);
  and (_14509_, _14508_, _06458_);
  and (_14510_, _14509_, _14505_);
  nor (_14511_, _12587_, _06896_);
  or (_14512_, _14511_, _14413_);
  and (_14513_, _14512_, _03741_);
  or (_14514_, _14513_, _03767_);
  or (_14515_, _14514_, _14510_);
  or (_14516_, _14424_, _03948_);
  and (_14517_, _14516_, _03446_);
  and (_14518_, _14517_, _14515_);
  and (_14519_, _14444_, _03445_);
  or (_14520_, _14519_, _03473_);
  or (_14521_, _14520_, _14518_);
  and (_14522_, _12638_, _05306_);
  or (_14523_, _14413_, _03474_);
  or (_14524_, _14523_, _14522_);
  and (_14525_, _14524_, _43189_);
  and (_14526_, _14525_, _14521_);
  or (_14527_, _14526_, _14412_);
  and (_43736_, _14527_, _42003_);
  nor (_14528_, _43189_, _07561_);
  nor (_14529_, _05306_, _07561_);
  nor (_14530_, _12773_, _06896_);
  or (_14531_, _14530_, _14529_);
  and (_14532_, _14531_, _03224_);
  nor (_14533_, _05929_, _07561_);
  and (_14534_, _12664_, _05929_);
  or (_14535_, _14534_, _14533_);
  or (_14536_, _14533_, _12691_);
  and (_14537_, _14536_, _14535_);
  or (_14538_, _14537_, _03459_);
  nor (_14539_, _12652_, _06896_);
  or (_14540_, _14539_, _14529_);
  or (_14541_, _14540_, _04432_);
  and (_14542_, _05306_, \oc8051_golden_model_1.ACC [3]);
  or (_14543_, _14542_, _14529_);
  and (_14544_, _14543_, _04436_);
  nor (_14545_, _04436_, _07561_);
  or (_14546_, _14545_, _03534_);
  or (_14547_, _14546_, _14544_);
  and (_14548_, _14547_, _03470_);
  and (_14549_, _14548_, _14541_);
  and (_14550_, _14535_, _03469_);
  or (_14551_, _14550_, _03527_);
  or (_14552_, _14551_, _14549_);
  nor (_14553_, _06896_, _04885_);
  or (_14554_, _14553_, _14529_);
  or (_14555_, _14554_, _04457_);
  and (_14556_, _14555_, _14552_);
  or (_14557_, _14556_, _03530_);
  or (_14558_, _14543_, _03531_);
  and (_14559_, _14558_, _03466_);
  and (_14560_, _14559_, _14557_);
  and (_14561_, _12662_, _05929_);
  or (_14562_, _14561_, _14533_);
  and (_14563_, _14562_, _03465_);
  or (_14564_, _14563_, _03458_);
  or (_14565_, _14564_, _14560_);
  and (_14566_, _14565_, _14538_);
  or (_14567_, _14566_, _06933_);
  nor (_14568_, _07421_, _07257_);
  nor (_14569_, _14568_, _07422_);
  or (_14570_, _14569_, _07447_);
  and (_14571_, _14570_, _03453_);
  and (_14572_, _14571_, _14567_);
  nor (_14573_, _12709_, _07455_);
  or (_14574_, _14573_, _14533_);
  and (_14575_, _14574_, _03452_);
  or (_14576_, _14575_, _07454_);
  or (_14577_, _14576_, _14572_);
  or (_14578_, _14554_, _06903_);
  and (_14579_, _14578_, _14577_);
  or (_14580_, _14579_, _04082_);
  and (_14581_, _06664_, _05306_);
  or (_14582_, _14529_, _04500_);
  or (_14583_, _14582_, _14581_);
  and (_14584_, _14583_, _03521_);
  and (_14585_, _14584_, _14580_);
  or (_14586_, _14585_, _14532_);
  and (_14587_, _14586_, _07474_);
  nand (_14588_, _07827_, _07777_);
  nor (_14589_, _14475_, _07788_);
  nor (_14590_, _14589_, _07780_);
  and (_14591_, _14589_, _07780_);
  or (_14592_, _14591_, _14590_);
  or (_14593_, _14592_, _07827_);
  and (_14594_, _14593_, _07468_);
  and (_14595_, _14594_, _14588_);
  or (_14596_, _14595_, _08905_);
  or (_14597_, _14596_, _14587_);
  and (_14598_, _12787_, _05306_);
  or (_14599_, _14529_, _04527_);
  or (_14600_, _14599_, _14598_);
  and (_14601_, _05306_, _06356_);
  or (_14602_, _14601_, _14529_);
  or (_14603_, _14602_, _04509_);
  and (_14604_, _14603_, _03745_);
  and (_14605_, _14604_, _14600_);
  and (_14606_, _14605_, _14597_);
  and (_14607_, _12793_, _05306_);
  or (_14608_, _14607_, _14529_);
  and (_14609_, _14608_, _03744_);
  or (_14610_, _14609_, _14606_);
  and (_14611_, _14610_, _04523_);
  or (_14612_, _14529_, _05625_);
  and (_14613_, _14602_, _03611_);
  and (_14614_, _14613_, _14612_);
  or (_14615_, _14614_, _14611_);
  and (_14616_, _14615_, _03734_);
  and (_14617_, _14543_, _03733_);
  and (_14618_, _14617_, _14612_);
  or (_14619_, _14618_, _03618_);
  or (_14620_, _14619_, _14616_);
  nor (_14621_, _12786_, _06896_);
  or (_14622_, _14529_, _06453_);
  or (_14623_, _14622_, _14621_);
  and (_14624_, _14623_, _06458_);
  and (_14625_, _14624_, _14620_);
  nor (_14626_, _12792_, _06896_);
  or (_14627_, _14626_, _14529_);
  and (_14628_, _14627_, _03741_);
  or (_14629_, _14628_, _03767_);
  or (_14630_, _14629_, _14625_);
  or (_14631_, _14540_, _03948_);
  and (_14632_, _14631_, _03446_);
  and (_14633_, _14632_, _14630_);
  and (_14634_, _14562_, _03445_);
  or (_14635_, _14634_, _03473_);
  or (_14636_, _14635_, _14633_);
  and (_14637_, _12843_, _05306_);
  or (_14638_, _14529_, _03474_);
  or (_14639_, _14638_, _14637_);
  and (_14640_, _14639_, _43189_);
  and (_14641_, _14640_, _14636_);
  or (_14642_, _14641_, _14528_);
  and (_43737_, _14642_, _42003_);
  nor (_14643_, _43189_, _07616_);
  nor (_14644_, _05306_, _07616_);
  nor (_14645_, _12972_, _06896_);
  or (_14646_, _14645_, _14644_);
  and (_14647_, _14646_, _03224_);
  nor (_14648_, _05929_, _07616_);
  and (_14649_, _12864_, _05929_);
  or (_14650_, _14649_, _14648_);
  and (_14651_, _14650_, _03465_);
  nor (_14652_, _12856_, _06896_);
  or (_14653_, _14652_, _14644_);
  and (_14654_, _14653_, _03534_);
  nor (_14655_, _04436_, _07616_);
  and (_14656_, _05306_, \oc8051_golden_model_1.ACC [4]);
  or (_14657_, _14656_, _14644_);
  and (_14658_, _14657_, _04436_);
  or (_14659_, _14658_, _14655_);
  and (_14660_, _14659_, _04432_);
  or (_14661_, _14660_, _03533_);
  or (_14662_, _14661_, _14654_);
  and (_14663_, _12866_, _05929_);
  or (_14664_, _14663_, _14648_);
  or (_14665_, _14664_, _03470_);
  nor (_14666_, _05831_, _06896_);
  or (_14667_, _14666_, _14644_);
  or (_14668_, _14667_, _04457_);
  and (_14669_, _14668_, _14665_);
  and (_14670_, _14669_, _14662_);
  or (_14671_, _14670_, _03530_);
  or (_14672_, _14657_, _03531_);
  and (_14673_, _14672_, _03466_);
  and (_14674_, _14673_, _14671_);
  or (_14675_, _14674_, _14651_);
  and (_14676_, _14675_, _03459_);
  or (_14677_, _14648_, _12894_);
  and (_14678_, _14677_, _03458_);
  and (_14679_, _14678_, _14664_);
  or (_14680_, _14679_, _06933_);
  or (_14681_, _14680_, _14676_);
  nor (_14682_, _07426_, _07424_);
  nor (_14683_, _14682_, _07427_);
  or (_14684_, _14683_, _07447_);
  and (_14685_, _14684_, _03453_);
  and (_14686_, _14685_, _14681_);
  nor (_14687_, _12912_, _07455_);
  or (_14688_, _14687_, _14648_);
  and (_14689_, _14688_, _03452_);
  or (_14690_, _14689_, _07454_);
  or (_14691_, _14690_, _14686_);
  or (_14692_, _14667_, _06903_);
  and (_14693_, _14692_, _14691_);
  or (_14694_, _14693_, _04082_);
  and (_14695_, _06802_, _05306_);
  or (_14696_, _14644_, _04500_);
  or (_14697_, _14696_, _14695_);
  and (_14698_, _14697_, _03521_);
  and (_14699_, _14698_, _14694_);
  or (_14700_, _14699_, _14647_);
  and (_14701_, _14700_, _07474_);
  nor (_14702_, _14589_, _07778_);
  or (_14703_, _14702_, _07779_);
  or (_14704_, _14703_, _07758_);
  nand (_14705_, _14703_, _07758_);
  nor (_14706_, _07827_, _07474_);
  and (_14707_, _14706_, _14705_);
  and (_14708_, _14707_, _14704_);
  and (_14709_, _07755_, _07468_);
  and (_14710_, _14709_, _07827_);
  or (_14711_, _14710_, _08905_);
  or (_14712_, _14711_, _14708_);
  or (_14713_, _14712_, _14701_);
  and (_14714_, _12986_, _05306_);
  or (_14715_, _14644_, _04527_);
  or (_14716_, _14715_, _14714_);
  and (_14717_, _06337_, _05306_);
  or (_14718_, _14717_, _14644_);
  or (_14719_, _14718_, _04509_);
  and (_14720_, _14719_, _03745_);
  and (_14721_, _14720_, _14716_);
  and (_14722_, _14721_, _14713_);
  and (_14723_, _12992_, _05306_);
  or (_14724_, _14723_, _14644_);
  and (_14725_, _14724_, _03744_);
  or (_14726_, _14725_, _14722_);
  and (_14727_, _14726_, _04523_);
  or (_14728_, _14644_, _05880_);
  and (_14729_, _14718_, _03611_);
  and (_14730_, _14729_, _14728_);
  or (_14731_, _14730_, _14727_);
  and (_14732_, _14731_, _03734_);
  and (_14733_, _14657_, _03733_);
  and (_14734_, _14733_, _14728_);
  or (_14735_, _14734_, _03618_);
  or (_14736_, _14735_, _14732_);
  nor (_14737_, _12985_, _06896_);
  or (_14738_, _14644_, _06453_);
  or (_14739_, _14738_, _14737_);
  and (_14740_, _14739_, _06458_);
  and (_14741_, _14740_, _14736_);
  nor (_14742_, _12991_, _06896_);
  or (_14743_, _14742_, _14644_);
  and (_14744_, _14743_, _03741_);
  or (_14745_, _14744_, _03767_);
  or (_14746_, _14745_, _14741_);
  or (_14747_, _14653_, _03948_);
  and (_14748_, _14747_, _03446_);
  and (_14749_, _14748_, _14746_);
  and (_14750_, _14650_, _03445_);
  or (_14751_, _14750_, _03473_);
  or (_14752_, _14751_, _14749_);
  and (_14753_, _13051_, _05306_);
  or (_14754_, _14644_, _03474_);
  or (_14755_, _14754_, _14753_);
  and (_14756_, _14755_, _43189_);
  and (_14757_, _14756_, _14752_);
  or (_14758_, _14757_, _14643_);
  and (_43738_, _14758_, _42003_);
  nor (_14759_, _43189_, _07607_);
  nor (_14760_, _05306_, _07607_);
  nor (_14761_, _13184_, _06896_);
  or (_14762_, _14761_, _14760_);
  and (_14763_, _14762_, _03224_);
  nor (_14764_, _05526_, _06896_);
  or (_14765_, _14764_, _14760_);
  or (_14766_, _14765_, _06903_);
  nor (_14767_, _05929_, _07607_);
  and (_14768_, _13078_, _05929_);
  or (_14769_, _14768_, _14767_);
  and (_14770_, _14769_, _03465_);
  nor (_14771_, _13070_, _06896_);
  or (_14772_, _14771_, _14760_);
  or (_14773_, _14772_, _04432_);
  and (_14774_, _05306_, \oc8051_golden_model_1.ACC [5]);
  or (_14775_, _14774_, _14760_);
  and (_14776_, _14775_, _04436_);
  nor (_14777_, _04436_, _07607_);
  or (_14778_, _14777_, _03534_);
  or (_14779_, _14778_, _14776_);
  and (_14780_, _14779_, _03470_);
  and (_14781_, _14780_, _14773_);
  and (_14782_, _13095_, _05929_);
  or (_14783_, _14782_, _14767_);
  and (_14784_, _14783_, _03469_);
  or (_14785_, _14784_, _03527_);
  or (_14786_, _14785_, _14781_);
  or (_14787_, _14765_, _04457_);
  and (_14788_, _14787_, _14786_);
  or (_14789_, _14788_, _03530_);
  or (_14790_, _14775_, _03531_);
  and (_14791_, _14790_, _03466_);
  and (_14792_, _14791_, _14789_);
  or (_14793_, _14792_, _14770_);
  and (_14794_, _14793_, _03459_);
  or (_14795_, _14767_, _13110_);
  and (_14796_, _14795_, _03458_);
  and (_14797_, _14796_, _14783_);
  or (_14798_, _14797_, _06933_);
  or (_14799_, _14798_, _14794_);
  nor (_14800_, _07429_, _07131_);
  nor (_14801_, _14800_, _07430_);
  or (_14802_, _14801_, _07447_);
  and (_14803_, _14802_, _03453_);
  and (_14804_, _14803_, _14799_);
  nor (_14805_, _13076_, _07455_);
  or (_14806_, _14805_, _14767_);
  and (_14807_, _14806_, _03452_);
  or (_14808_, _14807_, _07454_);
  or (_14809_, _14808_, _14804_);
  and (_14810_, _14809_, _14766_);
  or (_14811_, _14810_, _04082_);
  and (_14812_, _06757_, _05306_);
  or (_14813_, _14760_, _04500_);
  or (_14814_, _14813_, _14812_);
  and (_14815_, _14814_, _03521_);
  and (_14816_, _14815_, _14811_);
  or (_14817_, _14816_, _14763_);
  and (_14818_, _14817_, _07474_);
  not (_14819_, _07757_);
  and (_14820_, _14705_, _14819_);
  nor (_14821_, _14820_, _07768_);
  and (_14822_, _14820_, _07768_);
  or (_14823_, _14822_, _14821_);
  or (_14824_, _14823_, _07827_);
  nor (_14825_, _07765_, _07474_);
  or (_14826_, _14825_, _14706_);
  and (_14827_, _14826_, _14824_);
  or (_14828_, _14827_, _08905_);
  or (_14829_, _14828_, _14818_);
  and (_14830_, _13198_, _05306_);
  or (_14831_, _14760_, _04527_);
  or (_14832_, _14831_, _14830_);
  and (_14833_, _06295_, _05306_);
  or (_14834_, _14833_, _14760_);
  or (_14835_, _14834_, _04509_);
  and (_14836_, _14835_, _03745_);
  and (_14837_, _14836_, _14832_);
  and (_14838_, _14837_, _14829_);
  and (_14839_, _13204_, _05306_);
  or (_14840_, _14839_, _14760_);
  and (_14841_, _14840_, _03744_);
  or (_14842_, _14841_, _14838_);
  and (_14843_, _14842_, _04523_);
  or (_14844_, _14760_, _05576_);
  and (_14845_, _14834_, _03611_);
  and (_14846_, _14845_, _14844_);
  or (_14847_, _14846_, _14843_);
  and (_14848_, _14847_, _03734_);
  and (_14849_, _14775_, _03733_);
  and (_14850_, _14849_, _14844_);
  or (_14851_, _14850_, _03618_);
  or (_14852_, _14851_, _14848_);
  nor (_14853_, _13197_, _06896_);
  or (_14854_, _14760_, _06453_);
  or (_14855_, _14854_, _14853_);
  and (_14856_, _14855_, _06458_);
  and (_14857_, _14856_, _14852_);
  nor (_14858_, _13203_, _06896_);
  or (_14859_, _14858_, _14760_);
  and (_14860_, _14859_, _03741_);
  or (_14861_, _14860_, _03767_);
  or (_14862_, _14861_, _14857_);
  or (_14863_, _14772_, _03948_);
  and (_14864_, _14863_, _03446_);
  and (_14865_, _14864_, _14862_);
  and (_14866_, _14769_, _03445_);
  or (_14867_, _14866_, _03473_);
  or (_14868_, _14867_, _14865_);
  and (_14869_, _13253_, _05306_);
  or (_14870_, _14760_, _03474_);
  or (_14871_, _14870_, _14869_);
  and (_14872_, _14871_, _43189_);
  and (_14873_, _14872_, _14868_);
  or (_14874_, _14873_, _14759_);
  and (_43739_, _14874_, _42003_);
  nor (_14875_, _43189_, _07739_);
  nor (_14876_, _05306_, _07739_);
  nor (_14877_, _13387_, _06896_);
  or (_14878_, _14877_, _14876_);
  and (_14879_, _14878_, _03224_);
  nor (_14880_, _05417_, _06896_);
  or (_14881_, _14880_, _14876_);
  or (_14882_, _14881_, _06903_);
  nor (_14883_, _05929_, _07739_);
  and (_14884_, _13304_, _05929_);
  or (_14885_, _14884_, _14883_);
  and (_14886_, _14885_, _03465_);
  nor (_14887_, _13293_, _06896_);
  or (_14888_, _14887_, _14876_);
  or (_14889_, _14888_, _04432_);
  and (_14890_, _05306_, \oc8051_golden_model_1.ACC [6]);
  or (_14891_, _14890_, _14876_);
  and (_14892_, _14891_, _04436_);
  nor (_14893_, _04436_, _07739_);
  or (_14894_, _14893_, _03534_);
  or (_14895_, _14894_, _14892_);
  and (_14896_, _14895_, _03470_);
  and (_14897_, _14896_, _14889_);
  and (_14898_, _13280_, _05929_);
  or (_14899_, _14898_, _14883_);
  and (_14900_, _14899_, _03469_);
  or (_14901_, _14900_, _03527_);
  or (_14902_, _14901_, _14897_);
  or (_14903_, _14881_, _04457_);
  and (_14904_, _14903_, _14902_);
  or (_14905_, _14904_, _03530_);
  or (_14906_, _14891_, _03531_);
  and (_14907_, _14906_, _03466_);
  and (_14908_, _14907_, _14905_);
  or (_14909_, _14908_, _14886_);
  and (_14910_, _14909_, _03459_);
  or (_14911_, _14883_, _13311_);
  and (_14912_, _14911_, _03458_);
  and (_14913_, _14912_, _14899_);
  or (_14914_, _14913_, _06933_);
  or (_14915_, _14914_, _14910_);
  nor (_14916_, _07445_, _07432_);
  nor (_14917_, _14916_, _07446_);
  or (_14918_, _14917_, _07447_);
  and (_14919_, _14918_, _03453_);
  and (_14920_, _14919_, _14915_);
  nor (_14921_, _13329_, _07455_);
  or (_14922_, _14921_, _14883_);
  and (_14923_, _14922_, _03452_);
  or (_14924_, _14923_, _07454_);
  or (_14925_, _14924_, _14920_);
  and (_14926_, _14925_, _14882_);
  or (_14927_, _14926_, _04082_);
  and (_14928_, _06526_, _05306_);
  or (_14929_, _14876_, _04500_);
  or (_14930_, _14929_, _14928_);
  and (_14931_, _14930_, _03521_);
  and (_14932_, _14931_, _14927_);
  or (_14933_, _14932_, _14879_);
  and (_14934_, _14933_, _07474_);
  nor (_14935_, _14820_, _07766_);
  or (_14936_, _14935_, _07767_);
  nor (_14937_, _14936_, _07749_);
  and (_14938_, _14936_, _07749_);
  or (_14939_, _14938_, _14937_);
  or (_14940_, _14939_, _07827_);
  and (_14941_, _07745_, _07468_);
  or (_14942_, _14941_, _14706_);
  and (_14943_, _14942_, _14940_);
  or (_14944_, _14943_, _08905_);
  or (_14945_, _14944_, _14934_);
  and (_14946_, _13402_, _05306_);
  or (_14947_, _14876_, _04527_);
  or (_14948_, _14947_, _14946_);
  not (_14949_, _06262_);
  and (_14950_, _14949_, _05306_);
  or (_14951_, _14950_, _14876_);
  or (_14952_, _14951_, _04509_);
  and (_14953_, _14952_, _03745_);
  and (_14954_, _14953_, _14948_);
  and (_14955_, _14954_, _14945_);
  and (_14956_, _13407_, _05306_);
  or (_14957_, _14956_, _14876_);
  and (_14958_, _14957_, _03744_);
  or (_14959_, _14958_, _14955_);
  and (_14960_, _14959_, _04523_);
  or (_14961_, _14876_, _05469_);
  and (_14962_, _14951_, _03611_);
  and (_14963_, _14962_, _14961_);
  or (_14964_, _14963_, _14960_);
  and (_14965_, _14964_, _03734_);
  and (_14966_, _14891_, _03733_);
  and (_14967_, _14966_, _14961_);
  or (_14968_, _14967_, _03618_);
  or (_14969_, _14968_, _14965_);
  nor (_14970_, _13400_, _06896_);
  or (_14971_, _14876_, _06453_);
  or (_14972_, _14971_, _14970_);
  and (_14973_, _14972_, _06458_);
  and (_14974_, _14973_, _14969_);
  nor (_14975_, _13406_, _06896_);
  or (_14976_, _14975_, _14876_);
  and (_14977_, _14976_, _03741_);
  or (_14978_, _14977_, _03767_);
  or (_14979_, _14978_, _14974_);
  or (_14980_, _14888_, _03948_);
  and (_14981_, _14980_, _03446_);
  and (_14982_, _14981_, _14979_);
  and (_14983_, _14885_, _03445_);
  or (_14984_, _14983_, _03473_);
  or (_14985_, _14984_, _14982_);
  and (_14986_, _13456_, _05306_);
  or (_14987_, _14876_, _03474_);
  or (_14988_, _14987_, _14986_);
  and (_14989_, _14988_, _43189_);
  and (_14990_, _14989_, _14985_);
  or (_14991_, _14990_, _14875_);
  and (_43740_, _14991_, _42003_);
  nor (_14992_, _43189_, _03344_);
  nand (_14993_, _08815_, _06440_);
  nand (_14994_, _08415_, _03478_);
  and (_14995_, _14994_, _08786_);
  nand (_14996_, _08085_, _08595_);
  nand (_14997_, _08542_, _10159_);
  and (_14998_, _04462_, _03344_);
  nand (_14999_, _14998_, _07927_);
  or (_15000_, _08764_, _08510_);
  nor (_15001_, _05312_, _03344_);
  and (_15002_, _12177_, _05312_);
  nor (_15003_, _15002_, _15001_);
  nand (_15004_, _15003_, _03623_);
  or (_15005_, _12183_, _08486_);
  and (_15006_, _15005_, _07930_);
  nor (_15007_, _14998_, _07904_);
  and (_15008_, _08482_, _15007_);
  nand (_15009_, _03989_, _03262_);
  nor (_15010_, _12164_, _07936_);
  nor (_15011_, _15010_, _15001_);
  nor (_15012_, _15011_, _03521_);
  and (_15013_, _05312_, _04429_);
  nor (_15014_, _15013_, _15001_);
  nand (_15015_, _15014_, _07454_);
  nand (_15016_, _07988_, _07940_);
  or (_15017_, _08098_, _04429_);
  nor (_15018_, _04012_, _04007_);
  or (_15019_, _15018_, _06617_);
  nor (_15020_, _08380_, _08101_);
  or (_15021_, _08106_, _04429_);
  not (_15022_, _11680_);
  nor (_15023_, _08108_, _03344_);
  and (_15024_, _08108_, _03344_);
  or (_15025_, _15024_, _15023_);
  or (_15026_, _15025_, _15022_);
  and (_15027_, _15026_, _08101_);
  and (_15028_, _15027_, _15021_);
  or (_15029_, _15028_, _15020_);
  and (_15030_, _15029_, _11686_);
  or (_15031_, _15030_, _04012_);
  and (_15032_, _15031_, _04432_);
  and (_15033_, _15032_, _15019_);
  nor (_15034_, _05722_, _07936_);
  nor (_15035_, _15034_, _15001_);
  nor (_15036_, _15035_, _04432_);
  or (_15037_, _15036_, _03469_);
  or (_15038_, _15037_, _15033_);
  nor (_15039_, _05937_, _03344_);
  and (_15040_, _12075_, _05937_);
  nor (_15041_, _15040_, _15039_);
  nand (_15042_, _15041_, _03469_);
  and (_15043_, _15042_, _04457_);
  and (_15044_, _15043_, _15038_);
  nor (_15045_, _15014_, _04457_);
  or (_15046_, _15045_, _08099_);
  or (_15047_, _15046_, _15044_);
  and (_15048_, _15047_, _15017_);
  or (_15049_, _15048_, _04029_);
  or (_15050_, _06617_, _08160_);
  and (_15051_, _15050_, _03531_);
  and (_15052_, _15051_, _15049_);
  nor (_15053_, _08380_, _03531_);
  or (_15054_, _15053_, _08164_);
  or (_15055_, _15054_, _15052_);
  nand (_15056_, _08164_, _07545_);
  and (_15057_, _15056_, _15055_);
  or (_15058_, _15057_, _03465_);
  or (_15059_, _15001_, _03466_);
  and (_15060_, _15059_, _03459_);
  and (_15061_, _15060_, _15058_);
  nor (_15062_, _15035_, _03459_);
  or (_15063_, _15062_, _06933_);
  or (_15064_, _15063_, _15061_);
  not (_15065_, _07393_);
  nand (_15066_, _15065_, _06933_);
  and (_15067_, _15066_, _08191_);
  and (_15068_, _15067_, _15064_);
  nor (_15069_, _08241_, _03344_);
  nor (_15070_, _15069_, _08242_);
  nor (_15071_, _15070_, _08191_);
  or (_15072_, _15071_, _04066_);
  or (_15073_, _15072_, _15068_);
  nand (_15074_, _08085_, _04066_);
  and (_15075_, _15074_, _03599_);
  and (_15076_, _15075_, _15073_);
  nand (_15077_, _10306_, _07941_);
  and (_15078_, _15077_, _08267_);
  or (_15079_, _15078_, _15076_);
  and (_15080_, _15079_, _15016_);
  or (_15081_, _15080_, _03334_);
  nand (_15082_, _03989_, _03334_);
  and (_15083_, _15082_, _03453_);
  and (_15084_, _15083_, _15081_);
  nor (_15085_, _12106_, _08436_);
  nor (_15086_, _15085_, _15039_);
  nor (_15087_, _15086_, _03453_);
  or (_15088_, _15087_, _07454_);
  or (_15089_, _15088_, _15084_);
  and (_15090_, _15089_, _15015_);
  or (_15091_, _15090_, _04082_);
  and (_15092_, _06617_, _05312_);
  nor (_15093_, _15092_, _15001_);
  nand (_15094_, _15093_, _04082_);
  and (_15095_, _15094_, _03521_);
  and (_15096_, _15095_, _15091_);
  or (_15097_, _15096_, _15012_);
  and (_15098_, _15097_, _07474_);
  or (_15099_, _14706_, _03262_);
  or (_15100_, _15099_, _15098_);
  and (_15101_, _15100_, _15009_);
  or (_15102_, _15101_, _03624_);
  and (_15103_, _05312_, _06350_);
  nor (_15104_, _15103_, _15001_);
  nand (_15105_, _15104_, _03624_);
  and (_15106_, _15105_, _08462_);
  and (_15107_, _15106_, _15102_);
  nor (_15108_, _08462_, _03989_);
  or (_15109_, _15108_, _08469_);
  or (_15110_, _15109_, _15107_);
  or (_15111_, _08472_, _15007_);
  and (_15112_, _15111_, _08478_);
  and (_15113_, _15112_, _15110_);
  or (_15114_, _15113_, _15008_);
  and (_15115_, _15114_, _08487_);
  nor (_15116_, _06617_, \oc8051_golden_model_1.ACC [0]);
  nor (_15117_, _15116_, _08764_);
  and (_15118_, _15117_, _08481_);
  or (_15119_, _15118_, _03746_);
  or (_15120_, _15119_, _15115_);
  and (_15121_, _15120_, _15006_);
  and (_15122_, _10160_, _07929_);
  or (_15123_, _15122_, _03623_);
  or (_15124_, _15123_, _15121_);
  and (_15125_, _15124_, _15004_);
  or (_15126_, _15125_, _03744_);
  or (_15127_, _15001_, _03745_);
  and (_15128_, _15127_, _08506_);
  and (_15129_, _15128_, _15126_);
  and (_15130_, _08507_, _07904_);
  or (_15131_, _15130_, _04141_);
  or (_15132_, _15131_, _15129_);
  and (_15133_, _15132_, _15000_);
  or (_15134_, _15133_, _03735_);
  or (_15135_, _12182_, _08519_);
  and (_15136_, _15135_, _08518_);
  and (_15137_, _15136_, _15134_);
  and (_15138_, _08517_, _08831_);
  or (_15139_, _15138_, _15137_);
  and (_15140_, _15139_, _04523_);
  nor (_15141_, _15104_, _15034_);
  and (_15142_, _15141_, _03611_);
  or (_15143_, _15142_, _07927_);
  or (_15144_, _15143_, _15140_);
  and (_15145_, _15144_, _14999_);
  or (_15146_, _15145_, _08531_);
  nand (_15147_, _08531_, _14998_);
  and (_15148_, _15147_, _08533_);
  and (_15149_, _15148_, _15146_);
  nor (_15150_, _14998_, _08533_);
  or (_15151_, _15150_, _07923_);
  or (_15152_, _15151_, _15149_);
  nand (_15153_, _15116_, _07923_);
  and (_15154_, _15153_, _03740_);
  and (_15155_, _15154_, _15152_);
  not (_15156_, _11410_);
  nand (_15157_, _12181_, _08543_);
  and (_15158_, _15157_, _15156_);
  or (_15159_, _15158_, _15155_);
  and (_15160_, _15159_, _14997_);
  or (_15161_, _15160_, _03618_);
  nor (_15162_, _12057_, _07936_);
  nor (_15163_, _15162_, _15001_);
  nand (_15164_, _15163_, _03618_);
  and (_15165_, _15164_, _08564_);
  and (_15166_, _15165_, _15161_);
  nand (_15167_, _15070_, _08599_);
  and (_15168_, _15167_, _11940_);
  or (_15169_, _15168_, _15166_);
  and (_15170_, _15169_, _14996_);
  or (_15171_, _15170_, _03731_);
  nand (_15172_, _10306_, _03731_);
  and (_15173_, _15172_, _08709_);
  and (_15174_, _15173_, _15171_);
  nor (_15175_, _08709_, _07988_);
  or (_15176_, _15175_, _08707_);
  or (_15177_, _15176_, _15174_);
  and (_15178_, _08707_, _07982_);
  not (_15179_, _03188_);
  nor (_15180_, _10015_, _15179_);
  nor (_15181_, _15180_, _15178_);
  and (_15182_, _15181_, _15177_);
  and (_15183_, _15180_, _15007_);
  or (_15184_, _15183_, _04188_);
  or (_15185_, _15184_, _15182_);
  not (_15186_, _04188_);
  or (_15187_, _15007_, _15186_);
  and (_15188_, _15187_, _08742_);
  and (_15189_, _15188_, _15185_);
  and (_15190_, _15117_, _04184_);
  or (_15191_, _15190_, _03478_);
  or (_15192_, _15191_, _15189_);
  and (_15193_, _15192_, _14995_);
  and (_15194_, _08783_, _10160_);
  or (_15195_, _15194_, _08815_);
  or (_15196_, _15195_, _15193_);
  and (_15197_, _15196_, _14993_);
  or (_15198_, _15197_, _03767_);
  nand (_15199_, _15035_, _03767_);
  and (_15200_, _15199_, _08854_);
  and (_15201_, _15200_, _15198_);
  nor (_15202_, _08858_, _03344_);
  nor (_15203_, _15202_, _11998_);
  or (_15204_, _15203_, _15201_);
  nand (_15205_, _08858_, _03269_);
  and (_15206_, _15205_, _03446_);
  and (_15207_, _15206_, _15204_);
  and (_15208_, _15001_, _03445_);
  or (_15209_, _15208_, _03473_);
  or (_15210_, _15209_, _15207_);
  nand (_15211_, _15035_, _03473_);
  and (_15212_, _15211_, _08876_);
  and (_15213_, _15212_, _15210_);
  nor (_15214_, _08882_, _03344_);
  nor (_15215_, _15214_, _11392_);
  or (_15216_, _15215_, _15213_);
  nand (_15217_, _08882_, _03269_);
  and (_15218_, _15217_, _43189_);
  and (_15219_, _15218_, _15216_);
  or (_15220_, _15219_, _14992_);
  and (_43743_, _15220_, _42003_);
  nor (_15221_, _43189_, _03269_);
  nand (_15222_, _08815_, _03344_);
  nand (_15223_, _08542_, _07990_);
  not (_15224_, _11412_);
  nand (_15225_, _15224_, _07902_);
  or (_15226_, _12379_, _08519_);
  and (_15227_, _15226_, _08518_);
  nor (_15228_, _05312_, _03269_);
  and (_15229_, _15228_, _03744_);
  nand (_15230_, _04292_, _03262_);
  nor (_15231_, _07936_, _04635_);
  nor (_15232_, _15231_, _15228_);
  nand (_15233_, _15232_, _07454_);
  nand (_15234_, _07998_, _07940_);
  not (_15235_, _07993_);
  and (_15236_, _15235_, _04429_);
  nor (_15237_, _15236_, _07992_);
  and (_15238_, _15237_, _07903_);
  nor (_15239_, _15237_, _07903_);
  or (_15240_, _15239_, _15238_);
  or (_15241_, _15240_, _08191_);
  nor (_15242_, _05937_, _03269_);
  and (_15243_, _12269_, _05937_);
  and (_15244_, _15243_, _12284_);
  nor (_15245_, _15244_, _15242_);
  nor (_15246_, _15245_, _03459_);
  nand (_15247_, _08099_, _04635_);
  nor (_15248_, _08364_, _08101_);
  nor (_15249_, _08106_, _04635_);
  and (_15250_, _08108_, _03269_);
  nor (_15251_, _08108_, _03269_);
  or (_15252_, _15251_, _15250_);
  and (_15253_, _15252_, _08106_);
  or (_15254_, _15253_, _04007_);
  or (_15255_, _15254_, _15249_);
  and (_15256_, _15255_, _08101_);
  or (_15257_, _15256_, _15248_);
  and (_15258_, _15257_, _11686_);
  or (_15259_, _15258_, _04012_);
  or (_15260_, _15018_, _06572_);
  and (_15261_, _15260_, _15259_);
  or (_15262_, _15261_, _03534_);
  nor (_15263_, _05312_, \oc8051_golden_model_1.ACC [1]);
  and (_15264_, _12265_, _05312_);
  nor (_15265_, _15264_, _15263_);
  or (_15266_, _15265_, _04432_);
  and (_15267_, _15266_, _15262_);
  or (_15268_, _15267_, _08121_);
  nor (_15269_, _08128_, \oc8051_golden_model_1.PSW [6]);
  nor (_15270_, _15269_, \oc8051_golden_model_1.ACC [1]);
  and (_15271_, _15269_, \oc8051_golden_model_1.ACC [1]);
  nor (_15272_, _15271_, _15270_);
  nand (_15273_, _15272_, _08121_);
  and (_15274_, _15273_, _03532_);
  and (_15275_, _15274_, _15268_);
  nor (_15276_, _15243_, _15242_);
  nor (_15277_, _15276_, _03470_);
  nor (_15278_, _15232_, _04457_);
  or (_15279_, _15278_, _08099_);
  or (_15280_, _15279_, _15277_);
  or (_15281_, _15280_, _15275_);
  and (_15282_, _15281_, _15247_);
  or (_15283_, _15282_, _04029_);
  or (_15284_, _06572_, _08160_);
  and (_15285_, _15284_, _03531_);
  and (_15286_, _15285_, _15283_);
  nor (_15287_, _08364_, _03531_);
  or (_15288_, _15287_, _08164_);
  or (_15289_, _15288_, _15286_);
  nand (_15290_, _08164_, _07539_);
  and (_15291_, _15290_, _15289_);
  or (_15292_, _15291_, _03465_);
  and (_15293_, _12256_, _05937_);
  nor (_15294_, _15293_, _15242_);
  nand (_15295_, _15294_, _03465_);
  and (_15296_, _15295_, _03459_);
  and (_15297_, _15296_, _15292_);
  or (_15298_, _15297_, _15246_);
  and (_15299_, _15298_, _07447_);
  and (_15300_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_15301_, _15300_, _07794_);
  nor (_15302_, _15301_, _07394_);
  and (_15303_, _15302_, _06933_);
  nor (_15304_, _15303_, _08184_);
  nand (_15305_, _15304_, _08190_);
  or (_15306_, _15305_, _15299_);
  and (_15307_, _15306_, _15241_);
  or (_15308_, _15307_, _04066_);
  and (_15309_, _15235_, _06617_);
  nor (_15310_, _15309_, _07992_);
  and (_15311_, _15310_, _08763_);
  nor (_15312_, _15310_, _08763_);
  or (_15313_, _15312_, _15311_);
  or (_15314_, _15313_, _08024_);
  and (_15315_, _15314_, _03599_);
  and (_15316_, _15315_, _15308_);
  nand (_15317_, _10311_, _07941_);
  and (_15318_, _15317_, _08267_);
  or (_15319_, _15318_, _15316_);
  and (_15320_, _15319_, _15234_);
  or (_15321_, _15320_, _03334_);
  nand (_15322_, _04292_, _03334_);
  and (_15323_, _15322_, _03453_);
  and (_15324_, _15323_, _15321_);
  nor (_15325_, _12301_, _08436_);
  nor (_15326_, _15325_, _15242_);
  nor (_15327_, _15326_, _03453_);
  or (_15328_, _15327_, _07454_);
  or (_15329_, _15328_, _15324_);
  and (_15330_, _15329_, _15233_);
  or (_15331_, _15330_, _04082_);
  and (_15332_, _06572_, _05312_);
  nor (_15333_, _15332_, _15228_);
  nand (_15334_, _15333_, _04082_);
  and (_15335_, _15334_, _03521_);
  and (_15336_, _15335_, _15331_);
  nor (_15337_, _12360_, _07936_);
  nor (_15338_, _15337_, _15228_);
  nor (_15339_, _15338_, _03521_);
  or (_15340_, _15339_, _07468_);
  or (_15341_, _15340_, _15336_);
  or (_15342_, _07734_, _07474_);
  and (_15343_, _15342_, _15341_);
  or (_15344_, _15343_, _03262_);
  and (_15345_, _15344_, _15230_);
  or (_15346_, _15345_, _03624_);
  and (_15347_, _05312_, _04325_);
  nor (_15348_, _15347_, _15263_);
  or (_15349_, _15348_, _04509_);
  and (_15350_, _15349_, _08462_);
  and (_15351_, _15350_, _15346_);
  nor (_15352_, _08462_, _04292_);
  or (_15353_, _15352_, _08469_);
  or (_15354_, _15353_, _15351_);
  or (_15355_, _08472_, _07903_);
  and (_15356_, _15355_, _08475_);
  and (_15357_, _15356_, _15354_);
  or (_15358_, _08476_, _07903_);
  and (_15359_, _15358_, _08482_);
  or (_15360_, _15359_, _15357_);
  or (_15361_, _08477_, _07903_);
  and (_15362_, _15361_, _08487_);
  and (_15363_, _15362_, _15360_);
  and (_15364_, _08763_, _08481_);
  or (_15365_, _15364_, _03746_);
  or (_15366_, _15365_, _15363_);
  or (_15367_, _12381_, _08486_);
  and (_15368_, _15367_, _15366_);
  and (_15369_, _15368_, _07930_);
  and (_15370_, _07991_, _07929_);
  or (_15371_, _15370_, _03623_);
  or (_15372_, _15371_, _15369_);
  and (_15373_, _12375_, _05312_);
  nor (_15374_, _15373_, _15228_);
  nand (_15375_, _15374_, _03623_);
  and (_15376_, _15375_, _03745_);
  and (_15377_, _15376_, _15372_);
  or (_15378_, _15377_, _15229_);
  and (_15379_, _15378_, _08506_);
  and (_15380_, _08507_, _07901_);
  or (_15381_, _15380_, _15379_);
  and (_15382_, _15381_, _08510_);
  and (_15383_, _08761_, _04141_);
  or (_15384_, _15383_, _03735_);
  or (_15385_, _15384_, _15382_);
  and (_15386_, _15385_, _15227_);
  and (_15387_, _08517_, _07989_);
  or (_15388_, _15387_, _15386_);
  and (_15389_, _15388_, _04523_);
  and (_15390_, _12374_, _05312_);
  nor (_15391_, _15390_, _15228_);
  nor (_15392_, _15391_, _04523_);
  or (_15393_, _15392_, _15224_);
  or (_15394_, _15393_, _15389_);
  and (_15395_, _15394_, _15225_);
  or (_15396_, _15395_, _07923_);
  nand (_15397_, _08762_, _07923_);
  and (_15398_, _15397_, _03740_);
  and (_15399_, _15398_, _15396_);
  nand (_15400_, _12380_, _08543_);
  and (_15401_, _15400_, _15156_);
  or (_15402_, _15401_, _15399_);
  and (_15403_, _15402_, _15223_);
  or (_15404_, _15403_, _03618_);
  nor (_15405_, _12373_, _07936_);
  or (_15406_, _15405_, _15228_);
  or (_15407_, _15406_, _06453_);
  and (_15408_, _15407_, _08564_);
  and (_15409_, _15408_, _15404_);
  and (_15410_, _08576_, _08574_);
  nor (_15411_, _15410_, _08577_);
  or (_15412_, _15411_, _08595_);
  and (_15413_, _15412_, _11940_);
  or (_15414_, _15413_, _15409_);
  and (_15415_, _08608_, _08083_);
  nor (_15416_, _15415_, _08609_);
  or (_15417_, _15416_, _08599_);
  and (_15418_, _15417_, _15414_);
  or (_15419_, _15418_, _03731_);
  and (_15420_, _08688_, _08684_);
  nor (_15421_, _15420_, _08689_);
  or (_15422_, _15421_, _03732_);
  and (_15423_, _15422_, _08709_);
  and (_15424_, _15423_, _15419_);
  and (_15425_, _08718_, _08716_);
  nor (_15426_, _15425_, _08719_);
  and (_15427_, _15426_, _08627_);
  or (_15428_, _15427_, _08707_);
  or (_15429_, _15428_, _15424_);
  nand (_15430_, _08707_, _03344_);
  and (_15431_, _15430_, _07921_);
  and (_15432_, _15431_, _15429_);
  or (_15433_, _07904_, _07903_);
  nor (_15434_, _07921_, _07905_);
  and (_15435_, _15434_, _15433_);
  or (_15436_, _15435_, _04184_);
  or (_15437_, _15436_, _15432_);
  nor (_15438_, _08764_, _08763_);
  nor (_15439_, _15438_, _08765_);
  or (_15440_, _15439_, _08742_);
  and (_15441_, _15440_, _15437_);
  or (_15442_, _15441_, _03478_);
  and (_15443_, _08794_, _08413_);
  nor (_15444_, _15443_, _08795_);
  or (_15445_, _15444_, _03480_);
  and (_15446_, _15445_, _08786_);
  and (_15447_, _15446_, _15442_);
  nor (_15448_, _08831_, _07991_);
  nor (_15449_, _15448_, _08832_);
  and (_15450_, _15449_, _08783_);
  or (_15451_, _15450_, _08815_);
  or (_15452_, _15451_, _15447_);
  and (_15453_, _15452_, _15222_);
  or (_15454_, _15453_, _03767_);
  or (_15455_, _15265_, _03948_);
  and (_15456_, _15455_, _08854_);
  and (_15457_, _15456_, _15454_);
  nor (_15458_, _08883_, _08859_);
  nor (_15459_, _15458_, _08854_);
  or (_15460_, _15459_, _08858_);
  or (_15461_, _15460_, _15457_);
  nand (_15462_, _08858_, _07650_);
  and (_15463_, _15462_, _03446_);
  and (_15464_, _15463_, _15461_);
  nor (_15465_, _15294_, _03446_);
  or (_15466_, _15465_, _03473_);
  or (_15467_, _15466_, _15464_);
  nor (_15468_, _15264_, _15228_);
  nand (_15469_, _15468_, _03473_);
  and (_15470_, _15469_, _08876_);
  and (_15471_, _15470_, _15467_);
  nor (_15472_, _15458_, _08882_);
  nor (_15473_, _15472_, _11392_);
  or (_15474_, _15473_, _15471_);
  nand (_15475_, _08882_, _07650_);
  and (_15476_, _15475_, _43189_);
  and (_15477_, _15476_, _15474_);
  or (_15478_, _15477_, _15221_);
  and (_43744_, _15478_, _42003_);
  nor (_15479_, _43189_, _07650_);
  nand (_15480_, _08815_, _03269_);
  and (_15481_, _08720_, _07979_);
  nor (_15482_, _15481_, _08721_);
  or (_15483_, _15482_, _08709_);
  nand (_15484_, _08542_, _08828_);
  or (_15485_, _08757_, _08510_);
  nand (_15486_, _03944_, _03262_);
  nor (_15487_, _05312_, _07650_);
  nor (_15488_, _07936_, _05073_);
  nor (_15489_, _15488_, _15487_);
  nand (_15490_, _15489_, _07454_);
  nor (_15491_, _03989_, \oc8051_golden_model_1.ACC [0]);
  nor (_15492_, _15491_, _07991_);
  nor (_15493_, _15492_, _10130_);
  nor (_15494_, _08829_, _15493_);
  and (_15495_, _08829_, _15493_);
  nor (_15496_, _15495_, _15494_);
  not (_15497_, _10161_);
  or (_15498_, _15497_, _15496_);
  and (_15499_, _15498_, \oc8051_golden_model_1.PSW [7]);
  nor (_15500_, _15496_, \oc8051_golden_model_1.PSW [7]);
  or (_15501_, _15500_, _15499_);
  nand (_15502_, _15497_, _15496_);
  and (_15503_, _15502_, _15501_);
  nand (_15504_, _15503_, _07940_);
  nand (_15505_, _08099_, _05073_);
  nor (_15506_, _08350_, _08101_);
  nor (_15507_, _08106_, _05073_);
  and (_15508_, _08108_, _07650_);
  nor (_15509_, _08108_, _07650_);
  or (_15510_, _15509_, _15508_);
  and (_15511_, _15510_, _08106_);
  or (_15512_, _15511_, _04007_);
  or (_15513_, _15512_, _15507_);
  and (_15514_, _15513_, _08101_);
  or (_15515_, _15514_, _15506_);
  and (_15516_, _15515_, _11686_);
  or (_15517_, _15516_, _04012_);
  or (_15518_, _15018_, _06710_);
  and (_15519_, _15518_, _15517_);
  and (_15520_, _15519_, _04432_);
  nor (_15521_, _12467_, _07936_);
  nor (_15522_, _15521_, _15487_);
  nor (_15523_, _15522_, _04432_);
  or (_15524_, _15523_, _08121_);
  or (_15525_, _15524_, _15520_);
  nand (_15526_, _15269_, \oc8051_golden_model_1.ACC [2]);
  and (_15527_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_15528_, _15527_, _08127_);
  or (_15529_, _15528_, _15269_);
  and (_15530_, _15529_, _15526_);
  nand (_15531_, _15530_, _08121_);
  and (_15532_, _15531_, _03532_);
  and (_15533_, _15532_, _15525_);
  nor (_15534_, _05937_, _07650_);
  and (_15535_, _12462_, _05937_);
  nor (_15536_, _15535_, _15534_);
  nor (_15537_, _15536_, _03470_);
  nor (_15538_, _15489_, _04457_);
  or (_15539_, _15538_, _08099_);
  or (_15540_, _15539_, _15537_);
  or (_15541_, _15540_, _15533_);
  and (_15542_, _15541_, _15505_);
  or (_15543_, _15542_, _04029_);
  or (_15544_, _06710_, _08160_);
  and (_15545_, _15544_, _03531_);
  and (_15546_, _15545_, _15543_);
  nor (_15547_, _08350_, _03531_);
  or (_15548_, _15547_, _08164_);
  or (_15549_, _15548_, _15546_);
  nand (_15550_, _08164_, _07495_);
  and (_15551_, _15550_, _15549_);
  or (_15552_, _15551_, _03465_);
  and (_15553_, _12460_, _05937_);
  nor (_15554_, _15553_, _15534_);
  nand (_15555_, _15554_, _03465_);
  and (_15556_, _15555_, _03459_);
  and (_15557_, _15556_, _15552_);
  and (_15558_, _15535_, _12491_);
  nor (_15559_, _15558_, _15534_);
  nor (_15560_, _15559_, _03459_);
  or (_15561_, _15560_, _06933_);
  or (_15562_, _15561_, _15557_);
  nor (_15563_, _07396_, _07394_);
  nor (_15564_, _15563_, _07397_);
  or (_15565_, _15564_, _07447_);
  and (_15566_, _15565_, _08191_);
  and (_15567_, _15566_, _15562_);
  and (_15568_, _04635_, \oc8051_golden_model_1.ACC [1]);
  and (_15569_, _04429_, _03344_);
  nor (_15570_, _15569_, _07903_);
  nor (_15571_, _15570_, _15568_);
  nor (_15572_, _15571_, _07899_);
  and (_15573_, _15571_, _07899_);
  nor (_15574_, _15573_, _15572_);
  nor (_15575_, _15007_, _07903_);
  not (_15576_, _15575_);
  or (_15577_, _15576_, _15574_);
  and (_15578_, _15577_, \oc8051_golden_model_1.PSW [7]);
  nor (_15579_, _15574_, \oc8051_golden_model_1.PSW [7]);
  or (_15580_, _15579_, _15578_);
  nand (_15581_, _15576_, _15574_);
  and (_15582_, _15581_, _15580_);
  nor (_15583_, _15582_, _08191_);
  or (_15584_, _15583_, _15567_);
  or (_15585_, _15584_, _04066_);
  nor (_15586_, _06572_, _03269_);
  and (_15587_, _06617_, _03344_);
  nor (_15588_, _15587_, _08763_);
  nor (_15589_, _15588_, _15586_);
  nor (_15590_, _08759_, _15589_);
  and (_15591_, _08759_, _15589_);
  nor (_15592_, _15591_, _15590_);
  nor (_15593_, _15117_, _08763_);
  not (_15594_, _15593_);
  or (_15595_, _15594_, _15592_);
  and (_15596_, _15595_, \oc8051_golden_model_1.PSW [7]);
  nor (_15597_, _15592_, \oc8051_golden_model_1.PSW [7]);
  or (_15598_, _15597_, _15596_);
  nand (_15599_, _15594_, _15592_);
  and (_15600_, _15599_, _15598_);
  nand (_15601_, _15600_, _04066_);
  and (_15602_, _15601_, _03599_);
  and (_15603_, _15602_, _15585_);
  nor (_15604_, _08385_, _08383_);
  nor (_15605_, _15604_, _08386_);
  and (_15606_, _08416_, \oc8051_golden_model_1.PSW [7]);
  not (_15607_, _15606_);
  and (_15608_, _15607_, _15605_);
  or (_15609_, _15607_, _15605_);
  nand (_15610_, _15609_, _07941_);
  or (_15611_, _15610_, _15608_);
  and (_15612_, _15611_, _08267_);
  or (_15613_, _15612_, _15603_);
  and (_15614_, _15613_, _15504_);
  or (_15615_, _15614_, _03334_);
  nand (_15616_, _03944_, _03334_);
  and (_15617_, _15616_, _03453_);
  and (_15618_, _15617_, _15615_);
  nor (_15619_, _12509_, _08436_);
  nor (_15620_, _15619_, _15534_);
  nor (_15621_, _15620_, _03453_);
  or (_15622_, _15621_, _07454_);
  or (_15623_, _15622_, _15618_);
  and (_15624_, _15623_, _15490_);
  or (_15625_, _15624_, _04082_);
  and (_15626_, _06710_, _05312_);
  nor (_15627_, _15626_, _15487_);
  nand (_15628_, _15627_, _04082_);
  and (_15629_, _15628_, _03521_);
  and (_15630_, _15629_, _15625_);
  nor (_15631_, _12568_, _07936_);
  nor (_15632_, _15631_, _15487_);
  nor (_15633_, _15632_, _03521_);
  or (_15634_, _15633_, _07468_);
  or (_15635_, _15634_, _15630_);
  or (_15636_, _07670_, _07474_);
  and (_15637_, _15636_, _15635_);
  or (_15638_, _15637_, _03262_);
  and (_15639_, _15638_, _15486_);
  or (_15640_, _15639_, _03624_);
  and (_15641_, _05312_, _06399_);
  nor (_15642_, _15641_, _15487_);
  nand (_15643_, _15642_, _03624_);
  and (_15644_, _15643_, _08462_);
  and (_15645_, _15644_, _15640_);
  nor (_15646_, _08462_, _03944_);
  or (_15647_, _15646_, _08469_);
  or (_15648_, _15647_, _15645_);
  or (_15649_, _08472_, _07899_);
  and (_15650_, _03575_, _03171_);
  not (_15651_, _15650_);
  and (_15652_, _15651_, _08475_);
  and (_15653_, _15652_, _15649_);
  and (_15654_, _15653_, _15648_);
  nor (_15655_, _15652_, _07900_);
  or (_15656_, _15655_, _04132_);
  or (_15657_, _15656_, _15654_);
  not (_15658_, _04132_);
  or (_15659_, _07899_, _15658_);
  and (_15660_, _15659_, _08487_);
  and (_15661_, _15660_, _15657_);
  and (_15662_, _08759_, _08481_);
  or (_15663_, _15662_, _03746_);
  or (_15664_, _15663_, _15661_);
  or (_15665_, _12588_, _08486_);
  and (_15666_, _15665_, _07930_);
  and (_15667_, _15666_, _15664_);
  and (_15668_, _08829_, _07929_);
  or (_15669_, _15668_, _03623_);
  or (_15670_, _15669_, _15667_);
  and (_15671_, _12582_, _05312_);
  nor (_15672_, _15671_, _15487_);
  nand (_15673_, _15672_, _03623_);
  and (_15674_, _15673_, _03745_);
  and (_15675_, _15674_, _15670_);
  nor (_15676_, _06899_, _11900_);
  and (_15677_, _15487_, _03744_);
  or (_15678_, _15677_, _15676_);
  or (_15679_, _15678_, _15675_);
  or (_15680_, _05140_, _11900_);
  and (_15681_, _15680_, _04144_);
  not (_15682_, _07897_);
  nand (_15683_, _15676_, _15682_);
  and (_15684_, _15683_, _15681_);
  and (_15685_, _15684_, _15679_);
  nor (_15686_, _15681_, _15682_);
  or (_15687_, _15686_, _04141_);
  or (_15688_, _15687_, _15685_);
  and (_15689_, _15688_, _15485_);
  or (_15690_, _15689_, _03735_);
  or (_15691_, _12586_, _08519_);
  and (_15692_, _15691_, _08518_);
  and (_15694_, _15692_, _15690_);
  and (_15695_, _08517_, _08827_);
  or (_15696_, _15695_, _15694_);
  and (_15697_, _15696_, _04523_);
  or (_15698_, _05994_, _07926_);
  or (_15699_, _15642_, _12587_);
  or (_15700_, _15699_, _04523_);
  nand (_15701_, _15700_, _15698_);
  or (_15702_, _15701_, _15697_);
  and (_15703_, _03640_, _03177_);
  not (_15705_, _15703_);
  not (_15706_, _07898_);
  or (_15707_, _15698_, _15706_);
  and (_15708_, _15707_, _15705_);
  and (_15709_, _15708_, _15702_);
  nor (_15710_, _15705_, _07898_);
  or (_15711_, _15710_, _07923_);
  or (_15712_, _15711_, _15709_);
  nand (_15713_, _08758_, _07923_);
  and (_15714_, _15713_, _03740_);
  and (_15716_, _15714_, _15712_);
  nand (_15717_, _12587_, _08543_);
  and (_15718_, _15717_, _15156_);
  or (_15719_, _15718_, _15716_);
  and (_15720_, _15719_, _15484_);
  or (_15721_, _15720_, _03618_);
  nor (_15722_, _12581_, _07936_);
  nor (_15723_, _15722_, _15487_);
  nand (_15724_, _15723_, _03618_);
  and (_15725_, _15724_, _08564_);
  and (_15727_, _15725_, _15721_);
  not (_15728_, _08564_);
  and (_15729_, _08578_, _08233_);
  nor (_15730_, _15729_, _08579_);
  and (_15731_, _15730_, _15728_);
  or (_15732_, _15731_, _08595_);
  or (_15733_, _15732_, _15727_);
  and (_15734_, _08610_, _08065_);
  nor (_15735_, _15734_, _08611_);
  or (_15736_, _15735_, _08599_);
  and (_15738_, _15736_, _03732_);
  and (_15739_, _15738_, _15733_);
  and (_15740_, _08690_, _08678_);
  nor (_15741_, _15740_, _08691_);
  or (_15742_, _15741_, _08627_);
  and (_15743_, _15742_, _08629_);
  or (_15744_, _15743_, _15739_);
  and (_15745_, _15744_, _15483_);
  or (_15746_, _15745_, _08707_);
  nand (_15747_, _08707_, _03269_);
  and (_15749_, _15747_, _07921_);
  and (_15750_, _15749_, _15746_);
  and (_15751_, _07906_, _07900_);
  nor (_15752_, _15751_, _07907_);
  and (_15753_, _15752_, _07920_);
  or (_15754_, _15753_, _04184_);
  or (_15755_, _15754_, _15750_);
  and (_15756_, _08766_, _08760_);
  nor (_15757_, _15756_, _08767_);
  or (_15758_, _15757_, _08742_);
  and (_15760_, _15758_, _15755_);
  or (_15761_, _15760_, _03478_);
  and (_15762_, _08796_, _08385_);
  nor (_15763_, _15762_, _08797_);
  or (_15764_, _15763_, _03480_);
  and (_15765_, _15764_, _08786_);
  and (_15766_, _15765_, _15761_);
  and (_15767_, _08833_, _08830_);
  nor (_15768_, _15767_, _08834_);
  and (_15769_, _15768_, _08783_);
  or (_15771_, _15769_, _08815_);
  or (_15772_, _15771_, _15766_);
  and (_15773_, _15772_, _15480_);
  or (_15774_, _15773_, _03767_);
  nand (_15775_, _15522_, _03767_);
  and (_15776_, _15775_, _08854_);
  and (_15777_, _15776_, _15774_);
  and (_15778_, _08127_, _03344_);
  nor (_15779_, _08859_, _07650_);
  or (_15780_, _15779_, _15778_);
  nor (_15782_, _15780_, _08858_);
  nor (_15783_, _15782_, _11998_);
  or (_15784_, _15783_, _15777_);
  nand (_15785_, _08858_, _07644_);
  and (_15786_, _15785_, _03446_);
  and (_15787_, _15786_, _15784_);
  nor (_15788_, _15554_, _03446_);
  or (_15789_, _15788_, _03473_);
  or (_15790_, _15789_, _15787_);
  and (_15791_, _12638_, _05312_);
  nor (_15793_, _15791_, _15487_);
  nand (_15794_, _15793_, _03473_);
  and (_15795_, _15794_, _08876_);
  and (_15796_, _15795_, _15790_);
  and (_15797_, _08883_, \oc8051_golden_model_1.ACC [2]);
  nor (_15798_, _08883_, \oc8051_golden_model_1.ACC [2]);
  nor (_15799_, _15798_, _15797_);
  nor (_15800_, _15799_, _08882_);
  nor (_15801_, _15800_, _11392_);
  or (_15802_, _15801_, _15796_);
  nand (_15804_, _08882_, _07644_);
  and (_15805_, _15804_, _43189_);
  and (_15806_, _15805_, _15802_);
  or (_15807_, _15806_, _15479_);
  and (_43745_, _15807_, _42003_);
  nor (_15808_, _43189_, _07644_);
  nor (_15809_, _07896_, _07894_);
  nor (_15810_, _15809_, _07908_);
  and (_15811_, _15809_, _07908_);
  nor (_15812_, _15811_, _15810_);
  nand (_15814_, _15812_, _07920_);
  and (_15815_, _08580_, _08228_);
  nor (_15816_, _15815_, _08581_);
  and (_15817_, _15816_, _08566_);
  or (_15818_, _15817_, _08564_);
  and (_15819_, _08507_, _07894_);
  nor (_15820_, _05312_, _07644_);
  and (_15821_, _12787_, _05312_);
  nor (_15822_, _15821_, _15820_);
  nand (_15823_, _15822_, _03623_);
  nor (_15825_, _08753_, _08755_);
  or (_15826_, _15825_, _04130_);
  not (_15827_, _03171_);
  or (_15828_, _05994_, _15827_);
  and (_15829_, _15828_, _15651_);
  or (_15830_, _15829_, _15809_);
  nand (_15831_, _03440_, _03262_);
  nor (_15832_, _07936_, _04885_);
  nor (_15833_, _15832_, _15820_);
  nand (_15834_, _15833_, _07454_);
  and (_15836_, _03944_, \oc8051_golden_model_1.ACC [2]);
  nor (_15837_, _15494_, _15836_);
  nor (_15838_, _10127_, _15837_);
  and (_15839_, _10127_, _15837_);
  nor (_15840_, _15839_, _15838_);
  and (_15841_, _15840_, \oc8051_golden_model_1.PSW [7]);
  nor (_15842_, _15840_, \oc8051_golden_model_1.PSW [7]);
  nor (_15843_, _15842_, _15841_);
  and (_15844_, _15843_, _15499_);
  nor (_15845_, _15843_, _15499_);
  nor (_15847_, _15845_, _15844_);
  or (_15848_, _15847_, _07941_);
  and (_15849_, _05073_, \oc8051_golden_model_1.ACC [2]);
  nor (_15850_, _15572_, _15849_);
  nor (_15851_, _15850_, _15809_);
  and (_15852_, _15850_, _15809_);
  nor (_15853_, _15852_, _15851_);
  and (_15854_, _15853_, \oc8051_golden_model_1.PSW [7]);
  nor (_15855_, _15853_, \oc8051_golden_model_1.PSW [7]);
  nor (_15856_, _15855_, _15854_);
  and (_15858_, _15856_, _15578_);
  nor (_15859_, _15856_, _15578_);
  or (_15860_, _15859_, _15858_);
  nand (_15861_, _15860_, _08194_);
  nor (_15862_, _05937_, _07644_);
  and (_15863_, _12664_, _05937_);
  and (_15864_, _15863_, _12691_);
  nor (_15865_, _15864_, _15862_);
  nor (_15866_, _15865_, _03459_);
  nand (_15867_, _08099_, _04885_);
  or (_15868_, _15018_, _06664_);
  nor (_15869_, _08334_, _08101_);
  nor (_15870_, _08106_, _04885_);
  and (_15871_, _08108_, _07644_);
  nor (_15872_, _08108_, _07644_);
  or (_15873_, _15872_, _04007_);
  or (_15874_, _15873_, _15871_);
  and (_15875_, _15874_, _08106_);
  or (_15876_, _15875_, _15870_);
  and (_15877_, _15876_, _08101_);
  or (_15879_, _15877_, _15869_);
  and (_15880_, _15879_, _11686_);
  or (_15881_, _15880_, _04012_);
  and (_15882_, _15881_, _04432_);
  and (_15883_, _15882_, _15868_);
  nor (_15884_, _12652_, _07936_);
  nor (_15885_, _15884_, _15820_);
  nor (_15886_, _15885_, _04432_);
  or (_15887_, _15886_, _08121_);
  or (_15888_, _15887_, _15883_);
  not (_15890_, \oc8051_golden_model_1.PSW [6]);
  nor (_15891_, _08127_, _15890_);
  nor (_15892_, _15891_, \oc8051_golden_model_1.ACC [3]);
  nor (_15893_, _15892_, _08128_);
  not (_15894_, _15893_);
  nand (_15895_, _15894_, _08121_);
  and (_15896_, _15895_, _15888_);
  or (_15897_, _15896_, _03469_);
  nor (_15898_, _15863_, _15862_);
  nand (_15899_, _15898_, _03469_);
  and (_15901_, _15899_, _04457_);
  and (_15902_, _15901_, _15897_);
  nor (_15903_, _15833_, _04457_);
  or (_15904_, _15903_, _08099_);
  or (_15905_, _15904_, _15902_);
  and (_15906_, _15905_, _15867_);
  or (_15907_, _15906_, _04029_);
  or (_15908_, _06664_, _08160_);
  and (_15909_, _15908_, _03531_);
  and (_15910_, _15909_, _15907_);
  nor (_15912_, _08334_, _03531_);
  or (_15913_, _15912_, _08164_);
  or (_15914_, _15913_, _15910_);
  nand (_15915_, _08164_, _06440_);
  and (_15916_, _15915_, _15914_);
  or (_15917_, _15916_, _03465_);
  and (_15918_, _12662_, _05937_);
  nor (_15919_, _15918_, _15862_);
  nand (_15920_, _15919_, _03465_);
  and (_15921_, _15920_, _03459_);
  and (_15923_, _15921_, _15917_);
  or (_15924_, _15923_, _15866_);
  and (_15925_, _15924_, _07447_);
  nor (_15926_, _07399_, _07397_);
  nor (_15927_, _15926_, _07400_);
  nand (_15928_, _15927_, _06933_);
  nand (_15929_, _15928_, _08191_);
  or (_15930_, _15929_, _15925_);
  and (_15931_, _15930_, _15861_);
  or (_15932_, _15931_, _04066_);
  nor (_15934_, _06710_, _07650_);
  nor (_15935_, _15590_, _15934_);
  nor (_15936_, _15825_, _15935_);
  and (_15937_, _15825_, _15935_);
  nor (_15938_, _15937_, _15936_);
  and (_15939_, _15938_, \oc8051_golden_model_1.PSW [7]);
  nor (_15940_, _15938_, \oc8051_golden_model_1.PSW [7]);
  nor (_15941_, _15940_, _15939_);
  and (_15942_, _15941_, _15596_);
  nor (_15943_, _15941_, _15596_);
  nor (_15945_, _15943_, _15942_);
  or (_15946_, _15945_, _08024_);
  and (_15947_, _15946_, _03599_);
  and (_15948_, _15947_, _15932_);
  not (_15949_, _08411_);
  and (_15950_, _15949_, _08387_);
  nor (_15951_, _15949_, _08387_);
  nor (_15952_, _15951_, _15950_);
  and (_15953_, _15609_, _15952_);
  or (_15954_, _08418_, _07940_);
  or (_15956_, _15954_, _15953_);
  and (_15957_, _15956_, _08267_);
  or (_15958_, _15957_, _15948_);
  and (_15959_, _15958_, _15848_);
  or (_15960_, _15959_, _03334_);
  nand (_15961_, _03440_, _03334_);
  and (_15962_, _15961_, _03453_);
  and (_15963_, _15962_, _15960_);
  nor (_15964_, _12709_, _08436_);
  nor (_15965_, _15964_, _15862_);
  nor (_15967_, _15965_, _03453_);
  or (_15968_, _15967_, _07454_);
  or (_15969_, _15968_, _15963_);
  and (_15970_, _15969_, _15834_);
  or (_15971_, _15970_, _04082_);
  and (_15972_, _06664_, _05312_);
  nor (_15973_, _15972_, _15820_);
  nand (_15974_, _15973_, _04082_);
  and (_15975_, _15974_, _03521_);
  and (_15976_, _15975_, _15971_);
  nor (_15978_, _12773_, _07936_);
  nor (_15979_, _15978_, _15820_);
  nor (_15980_, _15979_, _03521_);
  or (_15981_, _15980_, _07468_);
  or (_15982_, _15981_, _15976_);
  or (_15983_, _07613_, _07474_);
  and (_15984_, _15983_, _15982_);
  or (_15985_, _15984_, _03262_);
  and (_15986_, _15985_, _15831_);
  or (_15987_, _15986_, _03624_);
  and (_15989_, _05312_, _06356_);
  nor (_15990_, _15989_, _15820_);
  nand (_15991_, _15990_, _03624_);
  and (_15992_, _15991_, _08462_);
  and (_15993_, _15992_, _15987_);
  or (_15994_, _08462_, _03440_);
  nand (_15995_, _15994_, _15829_);
  or (_15996_, _15995_, _15993_);
  and (_15997_, _15996_, _15830_);
  or (_15998_, _15997_, _04132_);
  and (_16000_, _03629_, _03171_);
  nor (_16001_, _15809_, _15658_);
  nor (_16002_, _16001_, _16000_);
  and (_16003_, _16002_, _15998_);
  and (_16004_, _15825_, _08481_);
  or (_16005_, _16004_, _04129_);
  or (_16006_, _16005_, _16003_);
  and (_16007_, _16006_, _15826_);
  or (_16008_, _16007_, _03746_);
  or (_16009_, _12793_, _08486_);
  and (_16011_, _16009_, _07930_);
  and (_16012_, _16011_, _16008_);
  and (_16013_, _10127_, _07929_);
  or (_16014_, _16013_, _03623_);
  or (_16015_, _16014_, _16012_);
  and (_16016_, _16015_, _15823_);
  or (_16017_, _16016_, _03744_);
  or (_16018_, _15820_, _03745_);
  and (_16019_, _16018_, _08506_);
  and (_16020_, _16019_, _16017_);
  or (_16022_, _16020_, _15819_);
  and (_16023_, _16022_, _08510_);
  and (_16024_, _08755_, _04141_);
  or (_16025_, _16024_, _03735_);
  or (_16026_, _16025_, _16023_);
  or (_16027_, _12791_, _08519_);
  and (_16028_, _16027_, _08518_);
  and (_16029_, _16028_, _16026_);
  and (_16030_, _08517_, _08825_);
  or (_16031_, _16030_, _16029_);
  and (_16033_, _16031_, _04523_);
  or (_16034_, _15990_, _12792_);
  nor (_16035_, _16034_, _04523_);
  or (_16036_, _16035_, _03902_);
  or (_16037_, _16036_, _16033_);
  nor (_16038_, _07896_, _03559_);
  or (_16039_, _16038_, _11412_);
  and (_16040_, _16039_, _16037_);
  and (_16041_, _03560_, _03177_);
  not (_16042_, _16041_);
  nor (_16044_, _16042_, _07896_);
  or (_16045_, _16044_, _07923_);
  or (_16046_, _16045_, _16040_);
  nand (_16047_, _08753_, _07923_);
  and (_16048_, _16047_, _03740_);
  and (_16049_, _16048_, _16046_);
  nand (_16050_, _12792_, _08543_);
  and (_16051_, _16050_, _15156_);
  or (_16052_, _16051_, _16049_);
  nand (_16053_, _08542_, _08826_);
  and (_16055_, _16053_, _06453_);
  and (_16056_, _16055_, _16052_);
  nor (_16057_, _12786_, _07936_);
  nor (_16058_, _16057_, _15820_);
  nor (_16059_, _16058_, _06453_);
  or (_16060_, _16059_, _08556_);
  or (_16061_, _16060_, _16056_);
  and (_16062_, _16061_, _15818_);
  and (_16063_, _15816_, _08565_);
  or (_16064_, _16063_, _08595_);
  or (_16066_, _16064_, _16062_);
  and (_16067_, _08612_, _08060_);
  nor (_16068_, _16067_, _08613_);
  or (_16069_, _16068_, _08599_);
  and (_16070_, _16069_, _03732_);
  and (_16071_, _16070_, _16066_);
  and (_16072_, _08692_, _08672_);
  nor (_16073_, _16072_, _08693_);
  or (_16074_, _16073_, _08627_);
  and (_16075_, _16074_, _08629_);
  or (_16077_, _16075_, _16071_);
  and (_16078_, _08722_, _07974_);
  nor (_16079_, _16078_, _08723_);
  or (_16080_, _16079_, _08709_);
  and (_16081_, _16080_, _08708_);
  and (_16082_, _16081_, _16077_);
  and (_16083_, _08707_, \oc8051_golden_model_1.ACC [2]);
  or (_16084_, _16083_, _07920_);
  or (_16085_, _16084_, _16082_);
  and (_16086_, _16085_, _15814_);
  or (_16088_, _16086_, _04184_);
  nor (_16089_, _08768_, _15825_);
  and (_16090_, _08768_, _15825_);
  nor (_16091_, _16090_, _16089_);
  nand (_16092_, _16091_, _04184_);
  and (_16093_, _16092_, _03480_);
  and (_16094_, _16093_, _16088_);
  nor (_16095_, _08798_, _08411_);
  and (_16096_, _08798_, _08411_);
  nor (_16097_, _16096_, _16095_);
  or (_16099_, _16097_, _08783_);
  and (_16100_, _16099_, _08785_);
  or (_16101_, _16100_, _16094_);
  nor (_16102_, _08835_, _10127_);
  and (_16103_, _08835_, _10127_);
  or (_16104_, _16103_, _16102_);
  or (_16105_, _16104_, _08786_);
  and (_16106_, _16105_, _08816_);
  and (_16107_, _16106_, _16101_);
  and (_16108_, _08815_, \oc8051_golden_model_1.ACC [2]);
  or (_16110_, _16108_, _03767_);
  or (_16111_, _16110_, _16107_);
  nand (_16112_, _15885_, _03767_);
  and (_16113_, _16112_, _08854_);
  and (_16114_, _16113_, _16111_);
  nor (_16115_, _15778_, _07644_);
  or (_16116_, _16115_, _08860_);
  and (_16117_, _16116_, _08853_);
  or (_16118_, _16117_, _08858_);
  or (_16119_, _16118_, _16114_);
  nand (_16121_, _08858_, _07545_);
  and (_16122_, _16121_, _03446_);
  and (_16123_, _16122_, _16119_);
  nor (_16124_, _15919_, _03446_);
  or (_16125_, _16124_, _03473_);
  or (_16126_, _16125_, _16123_);
  and (_16127_, _12843_, _05312_);
  nor (_16128_, _16127_, _15820_);
  nand (_16129_, _16128_, _03473_);
  and (_16130_, _16129_, _08876_);
  and (_16132_, _16130_, _16126_);
  or (_16133_, _15797_, \oc8051_golden_model_1.ACC [3]);
  and (_16134_, _16133_, _08884_);
  and (_16135_, _16134_, _08875_);
  or (_16136_, _16135_, _08882_);
  or (_16137_, _16136_, _16132_);
  nand (_16138_, _08882_, _07545_);
  and (_16139_, _16138_, _43189_);
  and (_16140_, _16139_, _16137_);
  or (_16141_, _16140_, _15808_);
  and (_43746_, _16141_, _42003_);
  nor (_16143_, _43189_, _07545_);
  nand (_16144_, _08815_, _07644_);
  and (_16145_, _08724_, _07968_);
  nor (_16146_, _16145_, _08725_);
  or (_16147_, _16146_, _08709_);
  nand (_16148_, _08542_, _08823_);
  and (_16149_, _03864_, _03177_);
  not (_16150_, _16149_);
  nor (_16151_, _07891_, _16150_);
  or (_16153_, _12990_, _08519_);
  and (_16154_, _16153_, _08518_);
  nor (_16155_, _05312_, _07545_);
  and (_16156_, _12986_, _05312_);
  nor (_16157_, _16156_, _16155_);
  nand (_16158_, _16157_, _03623_);
  nor (_16159_, _15650_, _04131_);
  or (_16160_, _16159_, _07892_);
  nor (_16161_, _06899_, _15827_);
  not (_16162_, _16161_);
  nor (_16164_, _08462_, _04257_);
  nand (_16165_, _04257_, _03262_);
  nor (_16166_, _05831_, _07936_);
  nor (_16167_, _16166_, _16155_);
  nand (_16168_, _16167_, _07454_);
  or (_16169_, _15858_, _15854_);
  nor (_16170_, _04885_, \oc8051_golden_model_1.ACC [3]);
  nand (_16171_, _04885_, \oc8051_golden_model_1.ACC [3]);
  and (_16172_, _15850_, _16171_);
  or (_16173_, _16172_, _16170_);
  nor (_16175_, _16173_, _07892_);
  and (_16176_, _16173_, _07892_);
  nor (_16177_, _16176_, _16175_);
  and (_16178_, _16177_, \oc8051_golden_model_1.PSW [7]);
  nor (_16179_, _16177_, \oc8051_golden_model_1.PSW [7]);
  nor (_16180_, _16179_, _16178_);
  and (_16181_, _16180_, _16169_);
  nor (_16182_, _16180_, _16169_);
  nor (_16183_, _16182_, _16181_);
  or (_16184_, _16183_, _08191_);
  nand (_16186_, _08099_, _05831_);
  nor (_16187_, _08320_, _08101_);
  or (_16188_, _06802_, _08103_);
  nor (_16189_, _08106_, _05831_);
  and (_16190_, _08108_, _07545_);
  nor (_16191_, _08108_, _07545_);
  or (_16192_, _16191_, _04007_);
  or (_16193_, _16192_, _16190_);
  and (_16194_, _16193_, _08106_);
  or (_16195_, _16194_, _16189_);
  and (_16197_, _16195_, _08101_);
  and (_16198_, _16197_, _16188_);
  or (_16199_, _16198_, _16187_);
  and (_16200_, _16199_, _08119_);
  nor (_16201_, _12856_, _07936_);
  nor (_16202_, _16201_, _16155_);
  nor (_16203_, _16202_, _04432_);
  or (_16204_, _16203_, _08121_);
  or (_16205_, _16204_, _16200_);
  nor (_16206_, _08128_, \oc8051_golden_model_1.ACC [4]);
  nor (_16208_, _16206_, _08134_);
  not (_16209_, _16208_);
  nand (_16210_, _16209_, _08121_);
  and (_16211_, _16210_, _03532_);
  and (_16212_, _16211_, _16205_);
  nor (_16213_, _05937_, _07545_);
  and (_16214_, _12866_, _05937_);
  nor (_16215_, _16214_, _16213_);
  nor (_16216_, _16215_, _03470_);
  nor (_16217_, _16167_, _04457_);
  or (_16219_, _16217_, _08099_);
  or (_16220_, _16219_, _16216_);
  or (_16221_, _16220_, _16212_);
  and (_16222_, _16221_, _16186_);
  or (_16223_, _16222_, _04029_);
  or (_16224_, _06802_, _08160_);
  and (_16225_, _16224_, _03531_);
  and (_16226_, _16225_, _16223_);
  nor (_16227_, _08320_, _03531_);
  or (_16228_, _16227_, _08164_);
  or (_16230_, _16228_, _16226_);
  nand (_16231_, _08164_, _03344_);
  and (_16232_, _16231_, _16230_);
  or (_16233_, _16232_, _03465_);
  and (_16234_, _12864_, _05937_);
  nor (_16235_, _16234_, _16213_);
  nand (_16236_, _16235_, _03465_);
  and (_16237_, _16236_, _03459_);
  and (_16238_, _16237_, _16233_);
  and (_16239_, _16214_, _12894_);
  nor (_16241_, _16239_, _16213_);
  nor (_16242_, _16241_, _03459_);
  or (_16243_, _16242_, _06933_);
  or (_16244_, _16243_, _16238_);
  nor (_16245_, _07402_, _07400_);
  nor (_16246_, _16245_, _07403_);
  or (_16247_, _16246_, _07447_);
  and (_16248_, _16247_, _16244_);
  or (_16249_, _16248_, _08194_);
  and (_16250_, _16249_, _08024_);
  and (_16252_, _16250_, _16184_);
  or (_16253_, _15942_, _15939_);
  and (_16254_, _06664_, _07644_);
  or (_16255_, _06664_, _07644_);
  and (_16256_, _16255_, _15935_);
  or (_16257_, _16256_, _16254_);
  nor (_16258_, _08752_, _16257_);
  and (_16259_, _08752_, _16257_);
  nor (_16260_, _16259_, _16258_);
  and (_16261_, _16260_, \oc8051_golden_model_1.PSW [7]);
  nor (_16263_, _16260_, \oc8051_golden_model_1.PSW [7]);
  nor (_16264_, _16263_, _16261_);
  and (_16265_, _16264_, _16253_);
  nor (_16266_, _16264_, _16253_);
  nor (_16267_, _16266_, _16265_);
  and (_16268_, _16267_, _04066_);
  or (_16269_, _16268_, _03594_);
  or (_16270_, _16269_, _16252_);
  and (_16271_, _08419_, _08410_);
  or (_16272_, _08420_, _03599_);
  or (_16274_, _16272_, _16271_);
  and (_16275_, _16274_, _07941_);
  and (_16276_, _16275_, _16270_);
  or (_16277_, _15844_, _15841_);
  nor (_16278_, _15837_, _10136_);
  nor (_16279_, _16278_, _10135_);
  nor (_16280_, _08824_, _16279_);
  and (_16281_, _08824_, _16279_);
  nor (_16282_, _16281_, _16280_);
  and (_16283_, _16282_, \oc8051_golden_model_1.PSW [7]);
  nor (_16285_, _16282_, \oc8051_golden_model_1.PSW [7]);
  nor (_16286_, _16285_, _16283_);
  and (_16287_, _16286_, _16277_);
  nor (_16288_, _16286_, _16277_);
  nor (_16289_, _16288_, _16287_);
  and (_16290_, _16289_, _07940_);
  or (_16291_, _16290_, _03334_);
  or (_16292_, _16291_, _16276_);
  nand (_16293_, _04257_, _03334_);
  and (_16294_, _16293_, _03453_);
  and (_16296_, _16294_, _16292_);
  nor (_16297_, _12912_, _08436_);
  nor (_16298_, _16297_, _16213_);
  nor (_16299_, _16298_, _03453_);
  or (_16300_, _16299_, _07454_);
  or (_16301_, _16300_, _16296_);
  and (_16302_, _16301_, _16168_);
  or (_16303_, _16302_, _04082_);
  and (_16304_, _06802_, _05312_);
  nor (_16305_, _16304_, _16155_);
  nand (_16307_, _16305_, _04082_);
  and (_16308_, _16307_, _03521_);
  and (_16309_, _16308_, _16303_);
  nor (_16310_, _12972_, _07936_);
  nor (_16311_, _16310_, _16155_);
  nor (_16312_, _16311_, _03521_);
  or (_16313_, _16312_, _07468_);
  or (_16314_, _16313_, _16309_);
  or (_16315_, _07558_, _07474_);
  and (_16316_, _16315_, _16314_);
  or (_16318_, _16316_, _03262_);
  and (_16319_, _16318_, _16165_);
  or (_16320_, _16319_, _03624_);
  and (_16321_, _06337_, _05312_);
  nor (_16322_, _16321_, _16155_);
  nand (_16323_, _16322_, _03624_);
  and (_16324_, _16323_, _08462_);
  and (_16325_, _16324_, _16320_);
  or (_16326_, _16325_, _16164_);
  and (_16327_, _16326_, _16162_);
  and (_16329_, _16161_, _07892_);
  or (_16330_, _16329_, _04131_);
  or (_16331_, _16330_, _15650_);
  or (_16332_, _16331_, _16327_);
  and (_16333_, _16332_, _16160_);
  or (_16334_, _16333_, _04132_);
  or (_16335_, _07892_, _15658_);
  and (_16336_, _16335_, _08487_);
  and (_16337_, _16336_, _16334_);
  and (_16338_, _08752_, _08481_);
  or (_16340_, _16338_, _03746_);
  or (_16341_, _16340_, _16337_);
  or (_16342_, _12992_, _08486_);
  and (_16343_, _16342_, _07930_);
  and (_16344_, _16343_, _16341_);
  and (_16345_, _08824_, _07929_);
  or (_16346_, _16345_, _03623_);
  or (_16347_, _16346_, _16344_);
  and (_16348_, _16347_, _16158_);
  or (_16349_, _16348_, _03744_);
  or (_16351_, _10015_, _11900_);
  or (_16352_, _16155_, _03745_);
  and (_16353_, _16352_, _16351_);
  and (_16354_, _16353_, _16349_);
  and (_16355_, _08507_, _07890_);
  or (_16356_, _16355_, _16354_);
  or (_16357_, _07890_, _04144_);
  and (_16358_, _16357_, _08510_);
  and (_16359_, _16358_, _16356_);
  and (_16360_, _08750_, _04141_);
  or (_16362_, _16360_, _03735_);
  or (_16363_, _16362_, _16359_);
  and (_16364_, _16363_, _16154_);
  and (_16365_, _08517_, _08822_);
  or (_16366_, _16365_, _16364_);
  and (_16367_, _16366_, _04523_);
  or (_16368_, _16322_, _12991_);
  nor (_16369_, _16368_, _04523_);
  or (_16370_, _16369_, _04334_);
  or (_16371_, _16370_, _16367_);
  nand (_16373_, _07891_, _04334_);
  and (_16374_, _16373_, _16150_);
  and (_16375_, _16374_, _16371_);
  or (_16376_, _16375_, _16151_);
  and (_16377_, _16376_, _16042_);
  nor (_16378_, _16042_, _07891_);
  or (_16379_, _16378_, _07923_);
  or (_16380_, _16379_, _16377_);
  nand (_16381_, _08751_, _07923_);
  and (_16382_, _16381_, _03740_);
  and (_16384_, _16382_, _16380_);
  nand (_16385_, _12991_, _08543_);
  and (_16386_, _16385_, _15156_);
  or (_16387_, _16386_, _16384_);
  and (_16388_, _16387_, _16148_);
  or (_16389_, _16388_, _03618_);
  nor (_16390_, _12985_, _07936_);
  nor (_16391_, _16390_, _16155_);
  nand (_16392_, _16391_, _03618_);
  and (_16393_, _16392_, _08564_);
  and (_16395_, _16393_, _16389_);
  and (_16396_, _08582_, _08220_);
  nor (_16397_, _16396_, _08583_);
  and (_16398_, _16397_, _15728_);
  or (_16399_, _16398_, _08595_);
  or (_16400_, _16399_, _16395_);
  and (_16401_, _08614_, _08051_);
  nor (_16402_, _16401_, _08615_);
  or (_16403_, _16402_, _08599_);
  and (_16404_, _16403_, _03732_);
  and (_16406_, _16404_, _16400_);
  and (_16407_, _08694_, _08666_);
  nor (_16408_, _16407_, _08695_);
  or (_16409_, _16408_, _08627_);
  and (_16410_, _16409_, _08629_);
  or (_16411_, _16410_, _16406_);
  and (_16412_, _16411_, _16147_);
  or (_16413_, _16412_, _08707_);
  nand (_16414_, _08707_, _07644_);
  and (_16415_, _16414_, _07921_);
  and (_16417_, _16415_, _16413_);
  and (_16418_, _07910_, _07893_);
  nor (_16419_, _16418_, _07911_);
  and (_16420_, _16419_, _07920_);
  or (_16421_, _16420_, _04184_);
  or (_16422_, _16421_, _16417_);
  nor (_16423_, _08770_, _08752_);
  nor (_16424_, _16423_, _08771_);
  or (_16425_, _16424_, _08742_);
  and (_16426_, _16425_, _16422_);
  or (_16428_, _16426_, _03478_);
  nor (_16429_, _08802_, _08790_);
  nor (_16430_, _16429_, _08803_);
  or (_16431_, _16430_, _03480_);
  and (_16432_, _16431_, _08786_);
  and (_16433_, _16432_, _16428_);
  nor (_16434_, _08837_, _08824_);
  nor (_16435_, _16434_, _08838_);
  and (_16436_, _16435_, _08783_);
  or (_16437_, _16436_, _08815_);
  or (_16439_, _16437_, _16433_);
  and (_16440_, _16439_, _16144_);
  or (_16441_, _16440_, _03767_);
  nand (_16442_, _16202_, _03767_);
  and (_16443_, _16442_, _08854_);
  and (_16444_, _16443_, _16441_);
  and (_16445_, _08860_, _07545_);
  nor (_16446_, _08860_, _07545_);
  nor (_16447_, _16446_, _16445_);
  not (_16448_, _16447_);
  and (_16450_, _16448_, _08853_);
  or (_16451_, _16450_, _08858_);
  or (_16452_, _16451_, _16444_);
  nand (_16453_, _08858_, _07539_);
  and (_16454_, _16453_, _03446_);
  and (_16455_, _16454_, _16452_);
  nor (_16456_, _16235_, _03446_);
  or (_16457_, _16456_, _03473_);
  or (_16458_, _16457_, _16455_);
  and (_16459_, _13051_, _05312_);
  nor (_16461_, _16459_, _16155_);
  nand (_16462_, _16461_, _03473_);
  and (_16463_, _16462_, _08876_);
  and (_16464_, _16463_, _16458_);
  and (_16465_, _08884_, _07545_);
  nor (_16466_, _16465_, _08885_);
  and (_16467_, _16466_, _08875_);
  or (_16468_, _16467_, _08882_);
  or (_16469_, _16468_, _16464_);
  nand (_16470_, _08882_, _07539_);
  and (_16472_, _16470_, _43189_);
  and (_16473_, _16472_, _16469_);
  or (_16474_, _16473_, _16143_);
  and (_43747_, _16474_, _42003_);
  nor (_16475_, _43189_, _07539_);
  and (_16476_, _07912_, _07889_);
  nor (_16477_, _16476_, _07913_);
  or (_16478_, _16477_, _07921_);
  and (_16479_, _08584_, _08215_);
  nor (_16480_, _16479_, _08585_);
  or (_16482_, _16480_, _08564_);
  or (_16483_, _13202_, _08519_);
  and (_16484_, _16483_, _08518_);
  or (_16485_, _15829_, _07888_);
  nand (_16486_, _03811_, _03262_);
  nor (_16487_, _05312_, _07539_);
  nor (_16488_, _05526_, _07936_);
  nor (_16489_, _16488_, _16487_);
  nand (_16490_, _16489_, _07454_);
  and (_16491_, _04257_, \oc8051_golden_model_1.ACC [4]);
  nor (_16493_, _16280_, _16491_);
  nor (_16494_, _10141_, _16493_);
  and (_16495_, _10141_, _16493_);
  nor (_16496_, _16495_, _16494_);
  and (_16497_, _16496_, \oc8051_golden_model_1.PSW [7]);
  nor (_16498_, _16496_, \oc8051_golden_model_1.PSW [7]);
  nor (_16499_, _16498_, _16497_);
  nor (_16500_, _16287_, _16283_);
  not (_16501_, _16500_);
  and (_16502_, _16501_, _16499_);
  nor (_16504_, _16501_, _16499_);
  nor (_16505_, _16504_, _16502_);
  or (_16506_, _16505_, _07941_);
  nor (_16507_, _06802_, _07545_);
  nor (_16508_, _16258_, _16507_);
  nor (_16509_, _08748_, _08746_);
  nor (_16510_, _16509_, _16508_);
  and (_16511_, _16509_, _16508_);
  nor (_16512_, _16511_, _16510_);
  and (_16513_, _16512_, \oc8051_golden_model_1.PSW [7]);
  nor (_16515_, _16512_, \oc8051_golden_model_1.PSW [7]);
  nor (_16516_, _16515_, _16513_);
  nor (_16517_, _16265_, _16261_);
  not (_16518_, _16517_);
  and (_16519_, _16518_, _16516_);
  nor (_16520_, _16518_, _16516_);
  nor (_16521_, _16520_, _16519_);
  and (_16522_, _16521_, _04066_);
  nor (_16523_, _05937_, _07539_);
  and (_16524_, _13095_, _05937_);
  and (_16526_, _16524_, _13110_);
  nor (_16527_, _16526_, _16523_);
  nor (_16528_, _16527_, _03459_);
  nand (_16529_, _08099_, _05526_);
  nor (_16530_, _08305_, _08101_);
  or (_16531_, _06757_, _08103_);
  nor (_16532_, _08106_, _05526_);
  and (_16533_, _08108_, _07539_);
  nor (_16534_, _08108_, _07539_);
  or (_16535_, _16534_, _16533_);
  and (_16537_, _16535_, _08106_);
  or (_16538_, _16537_, _04007_);
  or (_16539_, _16538_, _16532_);
  and (_16540_, _16539_, _08101_);
  and (_16541_, _16540_, _16531_);
  or (_16542_, _16541_, _16530_);
  and (_16543_, _16542_, _08119_);
  nor (_16544_, _13070_, _07936_);
  nor (_16545_, _16544_, _16487_);
  nor (_16546_, _16545_, _04432_);
  or (_16548_, _16546_, _08121_);
  or (_16549_, _16548_, _16543_);
  and (_16550_, _09991_, _08136_);
  nor (_16551_, _09991_, _08136_);
  nor (_16552_, _16551_, _16550_);
  nand (_16553_, _16552_, _08121_);
  and (_16554_, _16553_, _03532_);
  and (_16555_, _16554_, _16549_);
  nor (_16556_, _16524_, _16523_);
  nor (_16557_, _16556_, _03470_);
  nor (_16560_, _16489_, _04457_);
  or (_16561_, _16560_, _08099_);
  or (_16562_, _16561_, _16557_);
  or (_16563_, _16562_, _16555_);
  and (_16564_, _16563_, _16529_);
  or (_16565_, _16564_, _04029_);
  or (_16566_, _06757_, _08160_);
  and (_16567_, _16566_, _03531_);
  and (_16568_, _16567_, _16565_);
  nor (_16569_, _08305_, _03531_);
  or (_16571_, _16569_, _08164_);
  or (_16572_, _16571_, _16568_);
  nand (_16573_, _08164_, _03269_);
  and (_16574_, _16573_, _16572_);
  or (_16575_, _16574_, _03465_);
  and (_16576_, _13078_, _05937_);
  nor (_16577_, _16576_, _16523_);
  nand (_16578_, _16577_, _03465_);
  and (_16579_, _16578_, _03459_);
  and (_16580_, _16579_, _16575_);
  or (_16582_, _16580_, _16528_);
  and (_16583_, _16582_, _07447_);
  nor (_16584_, _07405_, _07403_);
  nor (_16585_, _16584_, _07406_);
  and (_16586_, _16585_, _06933_);
  or (_16587_, _16586_, _08194_);
  or (_16588_, _16587_, _16583_);
  and (_16589_, _05831_, \oc8051_golden_model_1.ACC [4]);
  nor (_16590_, _16175_, _16589_);
  nor (_16591_, _16590_, _07888_);
  and (_16593_, _16590_, _07888_);
  nor (_16594_, _16593_, _16591_);
  and (_16595_, _16594_, \oc8051_golden_model_1.PSW [7]);
  nor (_16596_, _16594_, \oc8051_golden_model_1.PSW [7]);
  nor (_16597_, _16596_, _16595_);
  nor (_16598_, _16181_, _16178_);
  not (_16599_, _16598_);
  and (_16600_, _16599_, _16597_);
  nor (_16601_, _16599_, _16597_);
  nor (_16602_, _16601_, _16600_);
  or (_16604_, _16602_, _08191_);
  and (_16605_, _16604_, _08024_);
  and (_16606_, _16605_, _16588_);
  or (_16607_, _16606_, _16522_);
  and (_16608_, _16607_, _03599_);
  and (_16609_, _08421_, _08408_);
  or (_16610_, _08422_, _07940_);
  or (_16611_, _16610_, _16609_);
  and (_16612_, _16611_, _08267_);
  or (_16613_, _16612_, _16608_);
  and (_16615_, _16613_, _16506_);
  or (_16616_, _16615_, _03334_);
  nand (_16617_, _03811_, _03334_);
  and (_16618_, _16617_, _03453_);
  and (_16619_, _16618_, _16616_);
  nor (_16620_, _13076_, _08436_);
  nor (_16621_, _16620_, _16523_);
  nor (_16622_, _16621_, _03453_);
  or (_16623_, _16622_, _07454_);
  or (_16624_, _16623_, _16619_);
  and (_16626_, _16624_, _16490_);
  or (_16627_, _16626_, _04082_);
  and (_16628_, _06757_, _05312_);
  nor (_16629_, _16628_, _16487_);
  nand (_16630_, _16629_, _04082_);
  and (_16631_, _16630_, _03521_);
  and (_16632_, _16631_, _16627_);
  nor (_16633_, _13184_, _07936_);
  nor (_16634_, _16633_, _16487_);
  nor (_16635_, _16634_, _03521_);
  or (_16637_, _16635_, _07468_);
  or (_16638_, _16637_, _16632_);
  or (_16639_, _07525_, _07474_);
  and (_16640_, _16639_, _16638_);
  or (_16641_, _16640_, _03262_);
  and (_16642_, _16641_, _16486_);
  or (_16643_, _16642_, _03624_);
  and (_16644_, _06295_, _05312_);
  nor (_16645_, _16644_, _16487_);
  nand (_16646_, _16645_, _03624_);
  and (_16648_, _16646_, _08462_);
  and (_16649_, _16648_, _16643_);
  or (_16650_, _08462_, _03811_);
  nand (_16651_, _16650_, _15829_);
  or (_16652_, _16651_, _16649_);
  and (_16653_, _16652_, _16485_);
  or (_16654_, _16653_, _04132_);
  or (_16655_, _07888_, _15658_);
  and (_16656_, _16655_, _08487_);
  and (_16657_, _16656_, _16654_);
  and (_16659_, _16509_, _08481_);
  or (_16660_, _16659_, _03746_);
  or (_16661_, _16660_, _16657_);
  or (_16662_, _13204_, _08486_);
  and (_16663_, _16662_, _16661_);
  and (_16664_, _16663_, _07930_);
  and (_16665_, _10141_, _07929_);
  or (_16666_, _16665_, _03623_);
  or (_16667_, _16666_, _16664_);
  and (_16668_, _13198_, _05312_);
  nor (_16670_, _16668_, _16487_);
  nand (_16671_, _16670_, _03623_);
  and (_16672_, _16671_, _03745_);
  and (_16673_, _16672_, _16667_);
  and (_16674_, _03572_, _03181_);
  and (_16675_, _16487_, _03744_);
  or (_16676_, _16675_, _16674_);
  or (_16677_, _16676_, _16673_);
  not (_16678_, _07886_);
  nand (_16679_, _16674_, _16678_);
  nor (_16681_, _03578_, _03566_);
  or (_16682_, _16681_, _11900_);
  and (_16683_, _15681_, _16682_);
  and (_16684_, _16683_, _16679_);
  and (_16685_, _16684_, _16677_);
  nor (_16686_, _16683_, _16678_);
  or (_16687_, _16686_, _16685_);
  and (_16688_, _16687_, _08510_);
  and (_16689_, _08748_, _04141_);
  or (_16690_, _16689_, _03735_);
  or (_16692_, _16690_, _16688_);
  and (_16693_, _16692_, _16484_);
  and (_16694_, _08517_, _08820_);
  or (_16695_, _16694_, _16693_);
  and (_16696_, _16695_, _04523_);
  or (_16697_, _16645_, _13203_);
  nor (_16698_, _16697_, _04523_);
  or (_16699_, _16698_, _07927_);
  or (_16700_, _16699_, _16696_);
  nor (_16701_, _15703_, _04155_);
  nand (_16703_, _07927_, _07887_);
  and (_16704_, _16703_, _16701_);
  and (_16705_, _16704_, _16700_);
  nor (_16706_, _16701_, _07887_);
  or (_16707_, _16706_, _07923_);
  or (_16708_, _16707_, _16705_);
  nand (_16709_, _08746_, _07923_);
  and (_16710_, _16709_, _03740_);
  and (_16711_, _16710_, _16708_);
  nand (_16712_, _13203_, _08543_);
  and (_16714_, _16712_, _15156_);
  or (_16715_, _16714_, _16711_);
  nand (_16716_, _08542_, _08821_);
  and (_16717_, _16716_, _06453_);
  and (_16718_, _16717_, _16715_);
  nor (_16719_, _13197_, _07936_);
  nor (_16720_, _16719_, _16487_);
  nor (_16721_, _16720_, _06453_);
  or (_16722_, _16721_, _15728_);
  or (_16723_, _16722_, _16718_);
  and (_16725_, _16723_, _16482_);
  or (_16726_, _16725_, _08595_);
  and (_16727_, _08616_, _08049_);
  nor (_16728_, _16727_, _08617_);
  or (_16729_, _16728_, _08599_);
  and (_16730_, _16729_, _03732_);
  and (_16731_, _16730_, _16726_);
  and (_16732_, _08696_, _08660_);
  nor (_16733_, _16732_, _08697_);
  or (_16734_, _16733_, _08627_);
  and (_16736_, _16734_, _08629_);
  or (_16737_, _16736_, _16731_);
  and (_16738_, _08726_, _07963_);
  nor (_16739_, _16738_, _08727_);
  or (_16740_, _16739_, _08709_);
  and (_16741_, _16740_, _08708_);
  and (_16742_, _16741_, _16737_);
  and (_16743_, _08707_, \oc8051_golden_model_1.ACC [4]);
  or (_16744_, _16743_, _07920_);
  or (_16745_, _16744_, _16742_);
  and (_16747_, _16745_, _16478_);
  or (_16748_, _16747_, _04184_);
  nor (_16749_, _08772_, _16509_);
  and (_16750_, _08772_, _16509_);
  or (_16751_, _16750_, _16749_);
  or (_16752_, _16751_, _08742_);
  and (_16753_, _16752_, _03480_);
  and (_16754_, _16753_, _16748_);
  and (_16755_, _08804_, _08404_);
  nor (_16756_, _16755_, _08805_);
  or (_16758_, _16756_, _08783_);
  and (_16759_, _16758_, _08785_);
  or (_16760_, _16759_, _16754_);
  not (_16761_, _10141_);
  nor (_16762_, _08839_, _16761_);
  and (_16763_, _08839_, _16761_);
  nor (_16764_, _16763_, _16762_);
  or (_16765_, _16764_, _08786_);
  and (_16766_, _16765_, _08816_);
  and (_16767_, _16766_, _16760_);
  and (_16769_, _08815_, \oc8051_golden_model_1.ACC [4]);
  or (_16770_, _16769_, _03767_);
  or (_16771_, _16770_, _16767_);
  nand (_16772_, _16545_, _03767_);
  and (_16773_, _16772_, _08854_);
  and (_16774_, _16773_, _16771_);
  nor (_16775_, _16445_, _07539_);
  or (_16776_, _16775_, _08861_);
  nor (_16777_, _16776_, _08858_);
  nor (_16778_, _16777_, _11998_);
  or (_16780_, _16778_, _16774_);
  nand (_16781_, _08858_, _07495_);
  and (_16782_, _16781_, _03446_);
  and (_16783_, _16782_, _16780_);
  nor (_16784_, _16577_, _03446_);
  or (_16785_, _16784_, _03473_);
  or (_16786_, _16785_, _16783_);
  and (_16787_, _13253_, _05312_);
  nor (_16788_, _16787_, _16487_);
  nand (_16789_, _16788_, _03473_);
  and (_16791_, _16789_, _08876_);
  and (_16792_, _16791_, _16786_);
  nor (_16793_, _08885_, \oc8051_golden_model_1.ACC [5]);
  nor (_16794_, _16793_, _08886_);
  and (_16795_, _16794_, _08875_);
  or (_16796_, _16795_, _08882_);
  or (_16797_, _16796_, _16792_);
  nand (_16798_, _08882_, _07495_);
  and (_16799_, _16798_, _43189_);
  and (_16800_, _16799_, _16797_);
  or (_16802_, _16800_, _16475_);
  and (_43748_, _16802_, _42003_);
  nor (_16803_, _43189_, _07495_);
  nand (_16804_, _08815_, _07539_);
  nand (_16805_, _08707_, _07539_);
  nand (_16806_, _08542_, _08818_);
  or (_16807_, _08743_, _08510_);
  nor (_16808_, _05312_, _07495_);
  and (_16809_, _13402_, _05312_);
  nor (_16810_, _16809_, _16808_);
  nand (_16812_, _16810_, _03623_);
  or (_16813_, _13407_, _08486_);
  and (_16814_, _16813_, _07930_);
  and (_16815_, _16161_, _07885_);
  nand (_16816_, _03511_, _03262_);
  nor (_16817_, _05417_, _07936_);
  nor (_16818_, _16817_, _16808_);
  nand (_16819_, _16818_, _07454_);
  and (_16820_, _08423_, _08403_);
  or (_16821_, _16820_, _08424_);
  or (_16823_, _16821_, _03599_);
  and (_16824_, _16823_, _07941_);
  nand (_16825_, _08099_, _05417_);
  nor (_16826_, _08287_, _08101_);
  or (_16827_, _06526_, _08103_);
  nor (_16828_, _08106_, _05417_);
  and (_16829_, _08108_, _07495_);
  nor (_16830_, _08108_, _07495_);
  or (_16831_, _16830_, _04007_);
  or (_16832_, _16831_, _16829_);
  and (_16834_, _16832_, _08106_);
  or (_16835_, _16834_, _16828_);
  and (_16836_, _16835_, _08101_);
  and (_16837_, _16836_, _16827_);
  or (_16838_, _16837_, _16826_);
  and (_16839_, _16838_, _08119_);
  nor (_16840_, _13293_, _07936_);
  nor (_16841_, _16840_, _16808_);
  nor (_16842_, _16841_, _04432_);
  or (_16843_, _16842_, _08121_);
  or (_16845_, _16843_, _16839_);
  not (_16846_, _08138_);
  nor (_16847_, _16551_, _16846_);
  and (_16848_, _09990_, _08139_);
  nor (_16849_, _16848_, _16847_);
  nand (_16850_, _16849_, _08121_);
  and (_16851_, _16850_, _03532_);
  and (_16852_, _16851_, _16845_);
  nor (_16853_, _05937_, _07495_);
  and (_16854_, _13280_, _05937_);
  nor (_16856_, _16854_, _16853_);
  nor (_16857_, _16856_, _03470_);
  nor (_16858_, _16818_, _04457_);
  or (_16859_, _16858_, _08099_);
  or (_16860_, _16859_, _16857_);
  or (_16861_, _16860_, _16852_);
  and (_16862_, _16861_, _16825_);
  or (_16863_, _16862_, _04029_);
  or (_16864_, _06526_, _08160_);
  and (_16865_, _16864_, _03531_);
  and (_16867_, _16865_, _16863_);
  nor (_16868_, _08287_, _03531_);
  or (_16869_, _16868_, _08164_);
  or (_16870_, _16869_, _16867_);
  nand (_16871_, _08164_, _07650_);
  and (_16872_, _16871_, _16870_);
  or (_16873_, _16872_, _03465_);
  and (_16874_, _13304_, _05937_);
  nor (_16875_, _16874_, _16853_);
  nand (_16876_, _16875_, _03465_);
  and (_16878_, _16876_, _03459_);
  and (_16879_, _16878_, _16873_);
  and (_16880_, _16854_, _13311_);
  nor (_16881_, _16880_, _16853_);
  nor (_16882_, _16881_, _03459_);
  or (_16883_, _16882_, _06933_);
  or (_16884_, _16883_, _16879_);
  nor (_16885_, _07408_, _07406_);
  nor (_16886_, _16885_, _07409_);
  or (_16887_, _16886_, _07447_);
  and (_16889_, _16887_, _08191_);
  and (_16890_, _16889_, _16884_);
  nand (_16891_, _05526_, \oc8051_golden_model_1.ACC [5]);
  nor (_16892_, _05526_, \oc8051_golden_model_1.ACC [5]);
  or (_16893_, _16590_, _16892_);
  and (_16894_, _16893_, _16891_);
  nor (_16895_, _16894_, _07885_);
  and (_16896_, _16894_, _07885_);
  nor (_16897_, _16896_, _16895_);
  nor (_16898_, _16600_, _16595_);
  and (_16900_, _16898_, \oc8051_golden_model_1.PSW [7]);
  or (_16901_, _16900_, _16897_);
  nand (_16902_, _16900_, _16897_);
  and (_16903_, _16902_, _16901_);
  and (_16904_, _16903_, _08194_);
  or (_16905_, _16904_, _04066_);
  or (_16906_, _16905_, _16890_);
  or (_16907_, _06757_, _07539_);
  and (_16908_, _06757_, _07539_);
  or (_16909_, _16508_, _16908_);
  and (_16911_, _16909_, _16907_);
  nor (_16912_, _16911_, _08745_);
  and (_16913_, _16911_, _08745_);
  nor (_16914_, _16913_, _16912_);
  nor (_16915_, _16519_, _16513_);
  and (_16916_, _16915_, \oc8051_golden_model_1.PSW [7]);
  nor (_16917_, _16916_, _16914_);
  and (_16918_, _16916_, _16914_);
  nor (_16919_, _16918_, _16917_);
  or (_16920_, _16919_, _08024_);
  and (_16922_, _16920_, _16906_);
  or (_16923_, _16922_, _03594_);
  and (_16924_, _16923_, _16824_);
  nor (_16925_, _16493_, _10147_);
  nor (_16926_, _16925_, _10146_);
  nor (_16927_, _16926_, _08819_);
  and (_16928_, _16926_, _08819_);
  nor (_16929_, _16928_, _16927_);
  nor (_16930_, _16502_, _16497_);
  and (_16931_, _16930_, \oc8051_golden_model_1.PSW [7]);
  or (_16933_, _16931_, _16929_);
  nand (_16934_, _16931_, _16929_);
  and (_16935_, _16934_, _16933_);
  and (_16936_, _16935_, _07940_);
  or (_16937_, _16936_, _03334_);
  or (_16938_, _16937_, _16924_);
  nand (_16939_, _03511_, _03334_);
  and (_16940_, _16939_, _03453_);
  and (_16941_, _16940_, _16938_);
  nor (_16942_, _13329_, _08436_);
  nor (_16944_, _16942_, _16853_);
  nor (_16945_, _16944_, _03453_);
  or (_16946_, _16945_, _07454_);
  or (_16947_, _16946_, _16941_);
  and (_16948_, _16947_, _16819_);
  or (_16949_, _16948_, _04082_);
  and (_16950_, _06526_, _05312_);
  nor (_16951_, _16950_, _16808_);
  nand (_16952_, _16951_, _04082_);
  and (_16953_, _16952_, _03521_);
  and (_16955_, _16953_, _16949_);
  nor (_16956_, _13387_, _07936_);
  nor (_16957_, _16956_, _16808_);
  nor (_16958_, _16957_, _03521_);
  or (_16959_, _16958_, _07468_);
  or (_16960_, _16959_, _16955_);
  not (_16961_, _07496_);
  and (_16962_, _07499_, _16961_);
  or (_16963_, _16962_, _07474_);
  and (_16964_, _16963_, _16960_);
  or (_16966_, _16964_, _03262_);
  and (_16967_, _16966_, _16816_);
  or (_16968_, _16967_, _03624_);
  and (_16969_, _14949_, _05312_);
  nor (_16970_, _16969_, _16808_);
  nand (_16971_, _16970_, _03624_);
  and (_16972_, _16971_, _08462_);
  and (_16973_, _16972_, _16968_);
  nor (_16974_, _08462_, _03511_);
  or (_16975_, _16974_, _16973_);
  and (_16977_, _16975_, _16162_);
  or (_16978_, _16977_, _16815_);
  and (_16979_, _16978_, _16159_);
  not (_16980_, _07885_);
  nor (_16981_, _16159_, _16980_);
  or (_16982_, _16981_, _04132_);
  or (_16983_, _16982_, _16979_);
  or (_16984_, _07885_, _15658_);
  and (_16985_, _16984_, _08487_);
  and (_16986_, _16985_, _16983_);
  and (_16988_, _08745_, _08481_);
  or (_16989_, _16988_, _03746_);
  or (_16990_, _16989_, _16986_);
  and (_16991_, _16990_, _16814_);
  and (_16992_, _08819_, _07929_);
  or (_16993_, _16992_, _03623_);
  or (_16994_, _16993_, _16991_);
  and (_16995_, _16994_, _16812_);
  or (_16996_, _16995_, _03744_);
  or (_16997_, _16808_, _03745_);
  and (_16999_, _16997_, _08506_);
  and (_17000_, _16999_, _16996_);
  and (_17001_, _08507_, _07883_);
  or (_17002_, _17001_, _04141_);
  or (_17003_, _17002_, _17000_);
  and (_17004_, _17003_, _16807_);
  or (_17005_, _17004_, _03735_);
  or (_17006_, _13276_, _08519_);
  and (_17007_, _17006_, _08518_);
  and (_17008_, _17007_, _17005_);
  and (_17010_, _08517_, _08817_);
  or (_17011_, _17010_, _17008_);
  and (_17012_, _17011_, _04523_);
  or (_17013_, _16970_, _13406_);
  nor (_17014_, _17013_, _04523_);
  or (_17015_, _17014_, _07927_);
  or (_17016_, _17015_, _17012_);
  nand (_17017_, _07927_, _07884_);
  and (_17018_, _17017_, _16701_);
  and (_17019_, _17018_, _17016_);
  nor (_17021_, _16701_, _07884_);
  or (_17022_, _17021_, _07923_);
  or (_17023_, _17022_, _17019_);
  nand (_17024_, _08744_, _07923_);
  and (_17025_, _17024_, _03740_);
  and (_17026_, _17025_, _17023_);
  nand (_17027_, _13406_, _08543_);
  and (_17028_, _17027_, _15156_);
  or (_17029_, _17028_, _17026_);
  and (_17030_, _17029_, _16806_);
  or (_17032_, _17030_, _03618_);
  nor (_17033_, _13400_, _07936_);
  nor (_17034_, _17033_, _16808_);
  nand (_17035_, _17034_, _03618_);
  and (_17036_, _17035_, _08564_);
  and (_17037_, _17036_, _17032_);
  and (_17038_, _08586_, _08568_);
  nor (_17039_, _17038_, _08587_);
  or (_17040_, _17039_, _08595_);
  and (_17041_, _17040_, _11940_);
  or (_17043_, _17041_, _17037_);
  and (_17044_, _08618_, _08601_);
  nor (_17045_, _17044_, _08619_);
  or (_17046_, _17045_, _08599_);
  and (_17047_, _17046_, _17043_);
  or (_17048_, _17047_, _03731_);
  and (_17049_, _08698_, _08654_);
  nor (_17050_, _17049_, _08699_);
  or (_17051_, _17050_, _03732_);
  and (_17052_, _17051_, _08709_);
  and (_17054_, _17052_, _17048_);
  and (_17055_, _08728_, _07957_);
  nor (_17056_, _17055_, _08729_);
  and (_17057_, _17056_, _08627_);
  or (_17058_, _17057_, _08707_);
  or (_17059_, _17058_, _17054_);
  and (_17060_, _17059_, _16805_);
  or (_17061_, _17060_, _07920_);
  nor (_17062_, _07914_, _07885_);
  nor (_17063_, _17062_, _07915_);
  or (_17065_, _17063_, _07921_);
  and (_17066_, _17065_, _08742_);
  and (_17067_, _17066_, _17061_);
  nor (_17068_, _08774_, _08745_);
  nor (_17069_, _17068_, _08775_);
  and (_17070_, _17069_, _04184_);
  or (_17071_, _17070_, _03478_);
  or (_17072_, _17071_, _17067_);
  and (_17073_, _08806_, _08290_);
  nor (_17074_, _17073_, _08807_);
  or (_17076_, _17074_, _03480_);
  and (_17077_, _17076_, _08786_);
  and (_17078_, _17077_, _17072_);
  nor (_17079_, _08841_, _08819_);
  nor (_17080_, _17079_, _08842_);
  and (_17081_, _17080_, _08783_);
  or (_17082_, _17081_, _08815_);
  or (_17083_, _17082_, _17078_);
  and (_17084_, _17083_, _16804_);
  or (_17085_, _17084_, _03767_);
  nand (_17087_, _16841_, _03767_);
  and (_17088_, _17087_, _08854_);
  and (_17089_, _17088_, _17085_);
  nor (_17090_, _08861_, _07495_);
  or (_17091_, _17090_, _08862_);
  and (_17092_, _17091_, _08853_);
  or (_17093_, _17092_, _08858_);
  or (_17094_, _17093_, _17089_);
  nand (_17095_, _08858_, _06440_);
  and (_17096_, _17095_, _03446_);
  and (_17098_, _17096_, _17094_);
  nor (_17099_, _16875_, _03446_);
  or (_17100_, _17099_, _03473_);
  or (_17101_, _17100_, _17098_);
  and (_17102_, _13456_, _05312_);
  nor (_17103_, _17102_, _16808_);
  nand (_17104_, _17103_, _03473_);
  and (_17105_, _17104_, _08876_);
  and (_17106_, _17105_, _17101_);
  nor (_17107_, _08886_, \oc8051_golden_model_1.ACC [6]);
  nor (_17109_, _17107_, _08887_);
  nor (_17110_, _17109_, _08882_);
  nor (_17111_, _17110_, _11392_);
  or (_17112_, _17111_, _17106_);
  nand (_17113_, _08882_, _06440_);
  and (_17114_, _17113_, _43189_);
  and (_17115_, _17114_, _17112_);
  or (_17116_, _17115_, _16803_);
  and (_43749_, _17116_, _42003_);
  not (_17117_, \oc8051_golden_model_1.DPL [0]);
  nor (_17119_, _43189_, _17117_);
  nor (_17120_, _05327_, _17117_);
  and (_17121_, _12183_, _05327_);
  or (_17122_, _17121_, _17120_);
  and (_17123_, _17122_, _03744_);
  and (_17124_, _08923_, _17117_);
  and (_17125_, _05327_, _04429_);
  or (_17126_, _17125_, _17120_);
  or (_17127_, _17126_, _04457_);
  nor (_17128_, _05722_, _08901_);
  or (_17130_, _17128_, _17120_);
  and (_17131_, _17130_, _03534_);
  nor (_17132_, _04436_, _17117_);
  and (_17133_, _05327_, \oc8051_golden_model_1.ACC [0]);
  or (_17134_, _17133_, _17120_);
  and (_17135_, _17134_, _04436_);
  or (_17136_, _17135_, _17132_);
  and (_17137_, _17136_, _04432_);
  or (_17138_, _17137_, _03527_);
  or (_17139_, _17138_, _17131_);
  and (_17141_, _17139_, _17127_);
  or (_17142_, _17141_, _03530_);
  or (_17143_, _17134_, _03531_);
  and (_17144_, _17143_, _08924_);
  and (_17145_, _17144_, _17142_);
  or (_17146_, _17145_, _17124_);
  and (_17147_, _17146_, _03622_);
  nor (_17148_, _04118_, _03622_);
  or (_17149_, _17148_, _07454_);
  or (_17150_, _17149_, _17147_);
  or (_17152_, _17126_, _06903_);
  and (_17153_, _17152_, _17150_);
  or (_17154_, _17153_, _04082_);
  and (_17155_, _06617_, _05327_);
  or (_17156_, _17120_, _04500_);
  or (_17157_, _17156_, _17155_);
  and (_17158_, _17157_, _03521_);
  and (_17159_, _17158_, _17154_);
  nor (_17160_, _12164_, _08901_);
  or (_17161_, _17160_, _17120_);
  and (_17163_, _17161_, _03224_);
  or (_17164_, _17163_, _17159_);
  or (_17165_, _17164_, _08905_);
  and (_17166_, _12177_, _05327_);
  or (_17167_, _17120_, _04527_);
  or (_17168_, _17167_, _17166_);
  and (_17169_, _05327_, _06350_);
  or (_17170_, _17169_, _17120_);
  or (_17171_, _17170_, _04509_);
  and (_17172_, _17171_, _03745_);
  and (_17174_, _17172_, _17168_);
  and (_17175_, _17174_, _17165_);
  or (_17176_, _17175_, _17123_);
  and (_17177_, _17176_, _04523_);
  nand (_17178_, _17170_, _03611_);
  nor (_17179_, _17178_, _17128_);
  or (_17180_, _17179_, _17177_);
  and (_17181_, _17180_, _03734_);
  or (_17182_, _17120_, _05722_);
  and (_17183_, _17134_, _03733_);
  and (_17185_, _17183_, _17182_);
  or (_17186_, _17185_, _03618_);
  or (_17187_, _17186_, _17181_);
  nor (_17188_, _12057_, _08901_);
  or (_17189_, _17120_, _06453_);
  or (_17190_, _17189_, _17188_);
  and (_17191_, _17190_, _06458_);
  and (_17192_, _17191_, _17187_);
  nor (_17193_, _12181_, _08901_);
  or (_17194_, _17193_, _17120_);
  and (_17196_, _17194_, _03741_);
  nor (_17197_, _03767_, _03473_);
  not (_17198_, _17197_);
  or (_17199_, _17198_, _17196_);
  or (_17200_, _17199_, _17192_);
  or (_17201_, _17197_, _17130_);
  and (_17202_, _17201_, _43189_);
  and (_17203_, _17202_, _17200_);
  or (_17204_, _17203_, _17119_);
  and (_43751_, _17204_, _42003_);
  not (_17206_, \oc8051_golden_model_1.DPL [1]);
  nor (_17207_, _43189_, _17206_);
  nor (_17208_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_17209_, _17208_, _08928_);
  and (_17210_, _17209_, _08923_);
  or (_17211_, _05327_, \oc8051_golden_model_1.DPL [1]);
  and (_17212_, _12265_, _05327_);
  not (_17213_, _17212_);
  and (_17214_, _17213_, _17211_);
  or (_17215_, _17214_, _04432_);
  nand (_17217_, _05327_, _03269_);
  and (_17218_, _17217_, _17211_);
  and (_17219_, _17218_, _04436_);
  nor (_17220_, _04436_, _17206_);
  or (_17221_, _17220_, _03534_);
  or (_17222_, _17221_, _17219_);
  and (_17223_, _17222_, _04457_);
  and (_17224_, _17223_, _17215_);
  nor (_17225_, _05327_, _17206_);
  nor (_17226_, _08901_, _04635_);
  or (_17228_, _17226_, _17225_);
  and (_17229_, _17228_, _03527_);
  or (_17230_, _17229_, _03530_);
  or (_17231_, _17230_, _17224_);
  or (_17232_, _17218_, _03531_);
  and (_17233_, _17232_, _08924_);
  and (_17234_, _17233_, _17231_);
  or (_17235_, _17234_, _17210_);
  and (_17236_, _17235_, _03622_);
  nor (_17237_, _04325_, _03622_);
  or (_17239_, _17237_, _07454_);
  or (_17240_, _17239_, _17236_);
  or (_17241_, _17228_, _06903_);
  and (_17242_, _17241_, _17240_);
  or (_17243_, _17242_, _04082_);
  and (_17244_, _06572_, _05327_);
  or (_17245_, _17225_, _04500_);
  or (_17246_, _17245_, _17244_);
  and (_17247_, _17246_, _03521_);
  and (_17248_, _17247_, _17243_);
  nor (_17250_, _12360_, _08901_);
  or (_17251_, _17250_, _17225_);
  and (_17252_, _17251_, _03224_);
  or (_17253_, _17252_, _17248_);
  and (_17254_, _17253_, _03625_);
  nand (_17255_, _05327_, _04325_);
  and (_17256_, _17211_, _03624_);
  and (_17257_, _17256_, _17255_);
  or (_17258_, _12375_, _08901_);
  and (_17259_, _17211_, _03623_);
  and (_17261_, _17259_, _17258_);
  or (_17262_, _17261_, _17257_);
  or (_17263_, _17262_, _17254_);
  and (_17264_, _17263_, _03745_);
  or (_17265_, _12381_, _08901_);
  and (_17266_, _17211_, _03744_);
  and (_17267_, _17266_, _17265_);
  or (_17268_, _17267_, _17264_);
  and (_17269_, _17268_, _04523_);
  or (_17270_, _12374_, _08901_);
  and (_17271_, _17211_, _03611_);
  and (_17272_, _17271_, _17270_);
  or (_17273_, _17272_, _17269_);
  and (_17274_, _17273_, _03734_);
  or (_17275_, _17225_, _05674_);
  and (_17276_, _17218_, _03733_);
  and (_17277_, _17276_, _17275_);
  or (_17278_, _17277_, _17274_);
  and (_17279_, _17278_, _03742_);
  or (_17280_, _17255_, _05674_);
  and (_17283_, _17211_, _03618_);
  and (_17284_, _17283_, _17280_);
  or (_17285_, _17217_, _05674_);
  and (_17286_, _17211_, _03741_);
  and (_17287_, _17286_, _17285_);
  or (_17288_, _17287_, _03767_);
  or (_17289_, _17288_, _17284_);
  or (_17290_, _17289_, _17279_);
  or (_17291_, _17214_, _03948_);
  and (_17292_, _17291_, _17290_);
  or (_17293_, _17292_, _03473_);
  or (_17294_, _17225_, _03474_);
  or (_17295_, _17294_, _17212_);
  and (_17296_, _17295_, _43189_);
  and (_17297_, _17296_, _17293_);
  or (_17298_, _17297_, _17207_);
  and (_43752_, _17298_, _42003_);
  not (_17299_, \oc8051_golden_model_1.DPL [2]);
  nor (_17300_, _43189_, _17299_);
  nor (_17301_, _05327_, _17299_);
  nor (_17304_, _12587_, _08901_);
  or (_17305_, _17304_, _17301_);
  and (_17306_, _17305_, _03741_);
  and (_17307_, _12588_, _05327_);
  or (_17308_, _17307_, _17301_);
  and (_17309_, _17308_, _03744_);
  nor (_17310_, _08901_, _05073_);
  or (_17311_, _17310_, _17301_);
  or (_17312_, _17311_, _06903_);
  nor (_17313_, _08928_, \oc8051_golden_model_1.DPL [2]);
  nor (_17315_, _17313_, _08929_);
  and (_17316_, _17315_, _08923_);
  nor (_17317_, _12467_, _08901_);
  or (_17318_, _17317_, _17301_);
  or (_17319_, _17318_, _04432_);
  and (_17320_, _05327_, \oc8051_golden_model_1.ACC [2]);
  or (_17321_, _17320_, _17301_);
  and (_17322_, _17321_, _04436_);
  nor (_17323_, _04436_, _17299_);
  or (_17324_, _17323_, _03534_);
  or (_17326_, _17324_, _17322_);
  and (_17327_, _17326_, _04457_);
  and (_17328_, _17327_, _17319_);
  and (_17329_, _17311_, _03527_);
  or (_17330_, _17329_, _03530_);
  or (_17331_, _17330_, _17328_);
  or (_17332_, _17321_, _03531_);
  and (_17333_, _17332_, _08924_);
  and (_17334_, _17333_, _17331_);
  or (_17335_, _17334_, _17316_);
  and (_17337_, _17335_, _03622_);
  nor (_17338_, _03855_, _03622_);
  or (_17339_, _17338_, _07454_);
  or (_17340_, _17339_, _17337_);
  and (_17341_, _17340_, _17312_);
  or (_17342_, _17341_, _04082_);
  and (_17343_, _06710_, _05327_);
  or (_17344_, _17301_, _04500_);
  or (_17345_, _17344_, _17343_);
  and (_17346_, _17345_, _03521_);
  and (_17348_, _17346_, _17342_);
  nor (_17349_, _12568_, _08901_);
  or (_17350_, _17349_, _17301_);
  and (_17351_, _17350_, _03224_);
  or (_17352_, _17351_, _17348_);
  or (_17353_, _17352_, _08905_);
  and (_17354_, _12582_, _05327_);
  or (_17355_, _17301_, _04527_);
  or (_17356_, _17355_, _17354_);
  and (_17357_, _05327_, _06399_);
  or (_17359_, _17357_, _17301_);
  or (_17360_, _17359_, _04509_);
  and (_17361_, _17360_, _03745_);
  and (_17362_, _17361_, _17356_);
  and (_17363_, _17362_, _17353_);
  or (_17364_, _17363_, _17309_);
  and (_17365_, _17364_, _04523_);
  or (_17366_, _17301_, _05772_);
  and (_17367_, _17359_, _03611_);
  and (_17368_, _17367_, _17366_);
  or (_17370_, _17368_, _17365_);
  and (_17371_, _17370_, _03734_);
  and (_17372_, _17321_, _03733_);
  and (_17373_, _17372_, _17366_);
  or (_17374_, _17373_, _03618_);
  or (_17375_, _17374_, _17371_);
  nor (_17376_, _12581_, _08901_);
  or (_17377_, _17301_, _06453_);
  or (_17378_, _17377_, _17376_);
  and (_17379_, _17378_, _06458_);
  and (_17381_, _17379_, _17375_);
  or (_17382_, _17381_, _17306_);
  and (_17383_, _17382_, _03948_);
  and (_17384_, _17318_, _03767_);
  or (_17385_, _17384_, _03473_);
  or (_17386_, _17385_, _17383_);
  and (_17387_, _12638_, _05327_);
  or (_17388_, _17301_, _03474_);
  or (_17389_, _17388_, _17387_);
  and (_17390_, _17389_, _43189_);
  and (_17392_, _17390_, _17386_);
  or (_17393_, _17392_, _17300_);
  and (_43753_, _17393_, _42003_);
  not (_17394_, \oc8051_golden_model_1.DPL [3]);
  nor (_17395_, _43189_, _17394_);
  nor (_17396_, _05327_, _17394_);
  nor (_17397_, _12792_, _08901_);
  or (_17398_, _17397_, _17396_);
  and (_17399_, _17398_, _03741_);
  and (_17400_, _12793_, _05327_);
  or (_17402_, _17400_, _17396_);
  and (_17403_, _17402_, _03744_);
  nor (_17404_, _08929_, \oc8051_golden_model_1.DPL [3]);
  nor (_17405_, _17404_, _08930_);
  and (_17406_, _17405_, _08923_);
  nor (_17407_, _12652_, _08901_);
  or (_17408_, _17407_, _17396_);
  or (_17409_, _17408_, _04432_);
  and (_17410_, _05327_, \oc8051_golden_model_1.ACC [3]);
  or (_17411_, _17410_, _17396_);
  and (_17413_, _17411_, _04436_);
  nor (_17414_, _04436_, _17394_);
  or (_17415_, _17414_, _03534_);
  or (_17416_, _17415_, _17413_);
  and (_17417_, _17416_, _04457_);
  and (_17418_, _17417_, _17409_);
  nor (_17419_, _08901_, _04885_);
  or (_17420_, _17419_, _17396_);
  and (_17421_, _17420_, _03527_);
  or (_17422_, _17421_, _03530_);
  or (_17424_, _17422_, _17418_);
  or (_17425_, _17411_, _03531_);
  and (_17426_, _17425_, _08924_);
  and (_17427_, _17426_, _17424_);
  or (_17428_, _17427_, _17406_);
  and (_17429_, _17428_, _03622_);
  nor (_17430_, _03725_, _03622_);
  or (_17431_, _17430_, _07454_);
  or (_17432_, _17431_, _17429_);
  or (_17433_, _17420_, _06903_);
  and (_17435_, _17433_, _17432_);
  or (_17436_, _17435_, _04082_);
  and (_17437_, _06664_, _05327_);
  or (_17438_, _17396_, _04500_);
  or (_17439_, _17438_, _17437_);
  and (_17440_, _17439_, _03521_);
  and (_17441_, _17440_, _17436_);
  nor (_17442_, _12773_, _08901_);
  or (_17443_, _17442_, _17396_);
  and (_17444_, _17443_, _03224_);
  or (_17446_, _17444_, _08905_);
  or (_17447_, _17446_, _17441_);
  and (_17448_, _12787_, _05327_);
  or (_17449_, _17396_, _04527_);
  or (_17450_, _17449_, _17448_);
  and (_17451_, _05327_, _06356_);
  or (_17452_, _17451_, _17396_);
  or (_17453_, _17452_, _04509_);
  and (_17454_, _17453_, _03745_);
  and (_17455_, _17454_, _17450_);
  and (_17457_, _17455_, _17447_);
  or (_17458_, _17457_, _17403_);
  and (_17459_, _17458_, _04523_);
  or (_17460_, _17396_, _05625_);
  and (_17461_, _17452_, _03611_);
  and (_17462_, _17461_, _17460_);
  or (_17463_, _17462_, _17459_);
  and (_17464_, _17463_, _03734_);
  and (_17465_, _17411_, _03733_);
  and (_17466_, _17465_, _17460_);
  or (_17468_, _17466_, _03618_);
  or (_17469_, _17468_, _17464_);
  nor (_17470_, _12786_, _08901_);
  or (_17471_, _17396_, _06453_);
  or (_17472_, _17471_, _17470_);
  and (_17473_, _17472_, _06458_);
  and (_17474_, _17473_, _17469_);
  or (_17475_, _17474_, _17399_);
  and (_17476_, _17475_, _03948_);
  and (_17477_, _17408_, _03767_);
  or (_17479_, _17477_, _03473_);
  or (_17480_, _17479_, _17476_);
  and (_17481_, _12843_, _05327_);
  or (_17482_, _17396_, _03474_);
  or (_17483_, _17482_, _17481_);
  and (_17484_, _17483_, _43189_);
  and (_17485_, _17484_, _17480_);
  or (_17486_, _17485_, _17395_);
  and (_43754_, _17486_, _42003_);
  not (_17487_, \oc8051_golden_model_1.DPL [4]);
  nor (_17489_, _43189_, _17487_);
  nor (_17490_, _05327_, _17487_);
  nor (_17491_, _12991_, _08901_);
  or (_17492_, _17491_, _17490_);
  and (_17493_, _17492_, _03741_);
  nor (_17494_, _05831_, _08901_);
  or (_17495_, _17494_, _17490_);
  or (_17496_, _17495_, _06903_);
  nor (_17497_, _12856_, _08901_);
  or (_17498_, _17497_, _17490_);
  or (_17500_, _17498_, _04432_);
  and (_17501_, _05327_, \oc8051_golden_model_1.ACC [4]);
  or (_17502_, _17501_, _17490_);
  and (_17503_, _17502_, _04436_);
  nor (_17504_, _04436_, _17487_);
  or (_17505_, _17504_, _03534_);
  or (_17506_, _17505_, _17503_);
  and (_17507_, _17506_, _04457_);
  and (_17508_, _17507_, _17500_);
  and (_17509_, _17495_, _03527_);
  or (_17511_, _17509_, _03530_);
  or (_17512_, _17511_, _17508_);
  or (_17513_, _17502_, _03531_);
  and (_17514_, _17513_, _08924_);
  and (_17515_, _17514_, _17512_);
  nor (_17516_, _08930_, \oc8051_golden_model_1.DPL [4]);
  nor (_17517_, _17516_, _08931_);
  and (_17518_, _17517_, _08923_);
  or (_17519_, _17518_, _17515_);
  and (_17520_, _17519_, _03622_);
  nor (_17522_, _06326_, _03622_);
  or (_17523_, _17522_, _07454_);
  or (_17524_, _17523_, _17520_);
  and (_17525_, _17524_, _17496_);
  or (_17526_, _17525_, _04082_);
  and (_17527_, _06802_, _05327_);
  or (_17528_, _17490_, _04500_);
  or (_17529_, _17528_, _17527_);
  and (_17530_, _17529_, _03521_);
  and (_17531_, _17530_, _17526_);
  nor (_17533_, _12972_, _08901_);
  or (_17534_, _17533_, _17490_);
  and (_17535_, _17534_, _03224_);
  or (_17536_, _17535_, _17531_);
  or (_17537_, _17536_, _08905_);
  and (_17538_, _12986_, _05327_);
  or (_17539_, _17490_, _04527_);
  or (_17540_, _17539_, _17538_);
  and (_17541_, _06337_, _05327_);
  or (_17542_, _17541_, _17490_);
  or (_17544_, _17542_, _04509_);
  and (_17545_, _17544_, _03745_);
  and (_17546_, _17545_, _17540_);
  and (_17547_, _17546_, _17537_);
  and (_17548_, _12992_, _05327_);
  or (_17549_, _17548_, _17490_);
  and (_17550_, _17549_, _03744_);
  or (_17551_, _17550_, _17547_);
  and (_17552_, _17551_, _04523_);
  or (_17553_, _17490_, _05880_);
  and (_17555_, _17542_, _03611_);
  and (_17556_, _17555_, _17553_);
  or (_17557_, _17556_, _17552_);
  and (_17558_, _17557_, _03734_);
  and (_17559_, _17502_, _03733_);
  and (_17560_, _17559_, _17553_);
  or (_17561_, _17560_, _03618_);
  or (_17562_, _17561_, _17558_);
  nor (_17563_, _12985_, _08901_);
  or (_17564_, _17490_, _06453_);
  or (_17566_, _17564_, _17563_);
  and (_17567_, _17566_, _06458_);
  and (_17568_, _17567_, _17562_);
  or (_17569_, _17568_, _17493_);
  and (_17570_, _17569_, _03948_);
  and (_17571_, _17498_, _03767_);
  or (_17572_, _17571_, _03473_);
  or (_17573_, _17572_, _17570_);
  and (_17574_, _13051_, _05327_);
  or (_17575_, _17490_, _03474_);
  or (_17577_, _17575_, _17574_);
  and (_17578_, _17577_, _43189_);
  and (_17579_, _17578_, _17573_);
  or (_17580_, _17579_, _17489_);
  and (_43757_, _17580_, _42003_);
  not (_17581_, \oc8051_golden_model_1.DPL [5]);
  nor (_17582_, _43189_, _17581_);
  nor (_17583_, _05327_, _17581_);
  nor (_17584_, _13203_, _08901_);
  or (_17585_, _17584_, _17583_);
  and (_17587_, _17585_, _03741_);
  nor (_17588_, _05526_, _08901_);
  or (_17589_, _17588_, _17583_);
  or (_17590_, _17589_, _06903_);
  nor (_17591_, _13070_, _08901_);
  or (_17592_, _17591_, _17583_);
  or (_17593_, _17592_, _04432_);
  and (_17594_, _05327_, \oc8051_golden_model_1.ACC [5]);
  or (_17595_, _17594_, _17583_);
  and (_17596_, _17595_, _04436_);
  nor (_17598_, _04436_, _17581_);
  or (_17599_, _17598_, _03534_);
  or (_17600_, _17599_, _17596_);
  and (_17601_, _17600_, _04457_);
  and (_17602_, _17601_, _17593_);
  and (_17603_, _17589_, _03527_);
  or (_17604_, _17603_, _03530_);
  or (_17605_, _17604_, _17602_);
  or (_17606_, _17595_, _03531_);
  and (_17607_, _17606_, _08924_);
  and (_17609_, _17607_, _17605_);
  nor (_17610_, _08931_, \oc8051_golden_model_1.DPL [5]);
  nor (_17611_, _17610_, _08932_);
  and (_17612_, _17611_, _08923_);
  or (_17613_, _17612_, _17609_);
  and (_17614_, _17613_, _03622_);
  nor (_17615_, _06294_, _03622_);
  or (_17616_, _17615_, _07454_);
  or (_17617_, _17616_, _17614_);
  and (_17618_, _17617_, _17590_);
  or (_17620_, _17618_, _04082_);
  and (_17621_, _06757_, _05327_);
  or (_17622_, _17583_, _04500_);
  or (_17623_, _17622_, _17621_);
  and (_17624_, _17623_, _03521_);
  and (_17625_, _17624_, _17620_);
  nor (_17626_, _13184_, _08901_);
  or (_17627_, _17626_, _17583_);
  and (_17628_, _17627_, _03224_);
  or (_17629_, _17628_, _17625_);
  or (_17631_, _17629_, _08905_);
  and (_17632_, _13198_, _05327_);
  or (_17633_, _17583_, _04527_);
  or (_17634_, _17633_, _17632_);
  and (_17635_, _06295_, _05327_);
  or (_17636_, _17635_, _17583_);
  or (_17637_, _17636_, _04509_);
  and (_17638_, _17637_, _03745_);
  and (_17639_, _17638_, _17634_);
  and (_17640_, _17639_, _17631_);
  and (_17642_, _13204_, _05327_);
  or (_17643_, _17642_, _17583_);
  and (_17644_, _17643_, _03744_);
  or (_17645_, _17644_, _17640_);
  and (_17646_, _17645_, _04523_);
  or (_17647_, _17583_, _05576_);
  and (_17648_, _17636_, _03611_);
  and (_17649_, _17648_, _17647_);
  or (_17650_, _17649_, _17646_);
  and (_17651_, _17650_, _03734_);
  and (_17653_, _17595_, _03733_);
  and (_17654_, _17653_, _17647_);
  or (_17655_, _17654_, _03618_);
  or (_17656_, _17655_, _17651_);
  nor (_17657_, _13197_, _08901_);
  or (_17658_, _17583_, _06453_);
  or (_17659_, _17658_, _17657_);
  and (_17660_, _17659_, _06458_);
  and (_17661_, _17660_, _17656_);
  or (_17662_, _17661_, _17587_);
  and (_17664_, _17662_, _03948_);
  and (_17665_, _17592_, _03767_);
  or (_17666_, _17665_, _03473_);
  or (_17667_, _17666_, _17664_);
  and (_17668_, _13253_, _05327_);
  or (_17669_, _17583_, _03474_);
  or (_17670_, _17669_, _17668_);
  and (_17671_, _17670_, _43189_);
  and (_17672_, _17671_, _17667_);
  or (_17673_, _17672_, _17582_);
  and (_43758_, _17673_, _42003_);
  not (_17675_, \oc8051_golden_model_1.DPL [6]);
  nor (_17676_, _43189_, _17675_);
  nor (_17677_, _05327_, _17675_);
  nor (_17678_, _13406_, _08901_);
  or (_17679_, _17678_, _17677_);
  and (_17680_, _17679_, _03741_);
  nor (_17681_, _05417_, _08901_);
  or (_17682_, _17681_, _17677_);
  or (_17683_, _17682_, _06903_);
  nor (_17685_, _13293_, _08901_);
  or (_17686_, _17685_, _17677_);
  or (_17687_, _17686_, _04432_);
  and (_17688_, _05327_, \oc8051_golden_model_1.ACC [6]);
  or (_17689_, _17688_, _17677_);
  and (_17690_, _17689_, _04436_);
  nor (_17691_, _04436_, _17675_);
  or (_17692_, _17691_, _03534_);
  or (_17693_, _17692_, _17690_);
  and (_17694_, _17693_, _04457_);
  and (_17696_, _17694_, _17687_);
  and (_17697_, _17682_, _03527_);
  or (_17698_, _17697_, _03530_);
  or (_17699_, _17698_, _17696_);
  or (_17700_, _17689_, _03531_);
  and (_17701_, _17700_, _08924_);
  and (_17702_, _17701_, _17699_);
  nor (_17703_, _08932_, \oc8051_golden_model_1.DPL [6]);
  nor (_17704_, _17703_, _08933_);
  and (_17705_, _17704_, _08923_);
  or (_17707_, _17705_, _17702_);
  and (_17708_, _17707_, _03622_);
  nor (_17709_, _06262_, _03622_);
  or (_17710_, _17709_, _07454_);
  or (_17711_, _17710_, _17708_);
  and (_17712_, _17711_, _17683_);
  or (_17713_, _17712_, _04082_);
  and (_17714_, _06526_, _05327_);
  or (_17715_, _17677_, _04500_);
  or (_17716_, _17715_, _17714_);
  and (_17718_, _17716_, _03521_);
  and (_17719_, _17718_, _17713_);
  nor (_17720_, _13387_, _08901_);
  or (_17721_, _17720_, _17677_);
  and (_17722_, _17721_, _03224_);
  or (_17723_, _17722_, _17719_);
  or (_17724_, _17723_, _08905_);
  and (_17725_, _13402_, _05327_);
  or (_17726_, _17677_, _04527_);
  or (_17727_, _17726_, _17725_);
  and (_17729_, _14949_, _05327_);
  or (_17730_, _17729_, _17677_);
  or (_17731_, _17730_, _04509_);
  and (_17732_, _17731_, _03745_);
  and (_17733_, _17732_, _17727_);
  and (_17734_, _17733_, _17724_);
  and (_17735_, _13407_, _05327_);
  or (_17736_, _17735_, _17677_);
  and (_17737_, _17736_, _03744_);
  or (_17738_, _17737_, _17734_);
  and (_17740_, _17738_, _04523_);
  or (_17741_, _17677_, _05469_);
  and (_17742_, _17730_, _03611_);
  and (_17743_, _17742_, _17741_);
  or (_17744_, _17743_, _17740_);
  and (_17745_, _17744_, _03734_);
  and (_17746_, _17689_, _03733_);
  and (_17747_, _17746_, _17741_);
  or (_17748_, _17747_, _03618_);
  or (_17749_, _17748_, _17745_);
  nor (_17751_, _13400_, _08901_);
  or (_17752_, _17677_, _06453_);
  or (_17753_, _17752_, _17751_);
  and (_17754_, _17753_, _06458_);
  and (_17755_, _17754_, _17749_);
  or (_17756_, _17755_, _17680_);
  and (_17757_, _17756_, _03948_);
  and (_17758_, _17686_, _03767_);
  or (_17759_, _17758_, _03473_);
  or (_17760_, _17759_, _17757_);
  and (_17762_, _13456_, _05327_);
  or (_17763_, _17677_, _03474_);
  or (_17764_, _17763_, _17762_);
  and (_17765_, _17764_, _43189_);
  and (_17766_, _17765_, _17760_);
  or (_17767_, _17766_, _17676_);
  and (_43759_, _17767_, _42003_);
  not (_17768_, \oc8051_golden_model_1.DPH [0]);
  nor (_17769_, _43189_, _17768_);
  nor (_17770_, _08935_, \oc8051_golden_model_1.DPH [0]);
  nor (_17772_, _17770_, _09028_);
  and (_17773_, _17772_, _08923_);
  nor (_17774_, _05320_, _17768_);
  nor (_17775_, _05722_, _09003_);
  or (_17776_, _17775_, _17774_);
  or (_17777_, _17776_, _04432_);
  and (_17778_, _05320_, \oc8051_golden_model_1.ACC [0]);
  or (_17779_, _17778_, _17774_);
  and (_17780_, _17779_, _04436_);
  nor (_17781_, _04436_, _17768_);
  or (_17783_, _17781_, _03534_);
  or (_17784_, _17783_, _17780_);
  and (_17785_, _17784_, _04457_);
  and (_17786_, _17785_, _17777_);
  and (_17787_, _05320_, _04429_);
  or (_17788_, _17787_, _17774_);
  and (_17789_, _17788_, _03527_);
  or (_17790_, _17789_, _03530_);
  or (_17791_, _17790_, _17786_);
  or (_17792_, _17779_, _03531_);
  and (_17794_, _17792_, _08924_);
  and (_17795_, _17794_, _17791_);
  or (_17796_, _17795_, _17773_);
  and (_17797_, _17796_, _03622_);
  nor (_17798_, _03989_, _03622_);
  or (_17799_, _17798_, _07454_);
  or (_17800_, _17799_, _17797_);
  or (_17801_, _17788_, _06903_);
  and (_17802_, _17801_, _17800_);
  or (_17803_, _17802_, _04082_);
  and (_17805_, _06617_, _05320_);
  or (_17806_, _17774_, _04500_);
  or (_17807_, _17806_, _17805_);
  and (_17808_, _17807_, _17803_);
  or (_17809_, _17808_, _03224_);
  nor (_17810_, _12164_, _09003_);
  or (_17811_, _17810_, _17774_);
  or (_17812_, _17811_, _03521_);
  and (_17813_, _17812_, _04509_);
  and (_17814_, _17813_, _17809_);
  and (_17816_, _05320_, _06350_);
  or (_17817_, _17816_, _17774_);
  and (_17818_, _17817_, _03624_);
  or (_17819_, _17818_, _03623_);
  or (_17820_, _17819_, _17814_);
  and (_17821_, _12177_, _05320_);
  or (_17822_, _17821_, _17774_);
  or (_17823_, _17822_, _04527_);
  and (_17824_, _17823_, _17820_);
  or (_17825_, _17824_, _03744_);
  and (_17827_, _12183_, _05320_);
  or (_17828_, _17827_, _17774_);
  or (_17829_, _17828_, _03745_);
  and (_17830_, _17829_, _04523_);
  and (_17831_, _17830_, _17825_);
  nand (_17832_, _17817_, _03611_);
  nor (_17833_, _17832_, _17775_);
  or (_17834_, _17833_, _17831_);
  and (_17835_, _17834_, _03734_);
  or (_17836_, _17774_, _05722_);
  and (_17838_, _17779_, _03733_);
  and (_17839_, _17838_, _17836_);
  or (_17840_, _17839_, _03618_);
  or (_17841_, _17840_, _17835_);
  nor (_17842_, _12057_, _09003_);
  or (_17843_, _17774_, _06453_);
  or (_17844_, _17843_, _17842_);
  and (_17845_, _17844_, _06458_);
  and (_17846_, _17845_, _17841_);
  nor (_17847_, _12181_, _09003_);
  or (_17849_, _17847_, _17774_);
  and (_17850_, _17849_, _03741_);
  or (_17851_, _17850_, _17198_);
  or (_17852_, _17851_, _17846_);
  or (_17853_, _17776_, _17197_);
  and (_17854_, _17853_, _43189_);
  and (_17855_, _17854_, _17852_);
  or (_17856_, _17855_, _17769_);
  and (_43761_, _17856_, _42003_);
  not (_17857_, \oc8051_golden_model_1.DPH [1]);
  nor (_17859_, _43189_, _17857_);
  or (_17860_, _05320_, \oc8051_golden_model_1.DPH [1]);
  and (_17861_, _12265_, _05320_);
  not (_17862_, _17861_);
  and (_17863_, _17862_, _17860_);
  or (_17864_, _17863_, _04432_);
  nand (_17865_, _05320_, _03269_);
  and (_17866_, _17865_, _17860_);
  and (_17867_, _17866_, _04436_);
  nor (_17868_, _04436_, _17857_);
  or (_17870_, _17868_, _03534_);
  or (_17871_, _17870_, _17867_);
  and (_17872_, _17871_, _04457_);
  and (_17873_, _17872_, _17864_);
  nor (_17874_, _05320_, _17857_);
  nor (_17875_, _09003_, _04635_);
  or (_17876_, _17875_, _17874_);
  and (_17877_, _17876_, _03527_);
  or (_17878_, _17877_, _03530_);
  or (_17879_, _17878_, _17873_);
  or (_17881_, _17866_, _03531_);
  and (_17882_, _17881_, _08924_);
  and (_17883_, _17882_, _17879_);
  nor (_17884_, _09028_, \oc8051_golden_model_1.DPH [1]);
  nor (_17885_, _17884_, _09029_);
  and (_17886_, _17885_, _08923_);
  or (_17887_, _17886_, _17883_);
  and (_17888_, _17887_, _03622_);
  nor (_17889_, _04292_, _03622_);
  or (_17890_, _17889_, _07454_);
  or (_17892_, _17890_, _17888_);
  or (_17893_, _17876_, _06903_);
  and (_17894_, _17893_, _17892_);
  or (_17895_, _17894_, _04082_);
  and (_17896_, _06572_, _05320_);
  or (_17897_, _17874_, _04500_);
  or (_17898_, _17897_, _17896_);
  and (_17899_, _17898_, _03521_);
  and (_17900_, _17899_, _17895_);
  nand (_17901_, _12360_, _05320_);
  and (_17903_, _17860_, _03224_);
  and (_17904_, _17903_, _17901_);
  or (_17905_, _17904_, _17900_);
  and (_17906_, _17905_, _03625_);
  or (_17907_, _12375_, _09003_);
  and (_17908_, _17907_, _03623_);
  nand (_17909_, _05320_, _04325_);
  and (_17910_, _17909_, _03624_);
  or (_17911_, _17910_, _17908_);
  and (_17912_, _17911_, _17860_);
  or (_17914_, _17912_, _17906_);
  and (_17915_, _17914_, _03745_);
  or (_17916_, _12381_, _09003_);
  and (_17917_, _17860_, _03744_);
  and (_17918_, _17917_, _17916_);
  or (_17919_, _17918_, _17915_);
  and (_17920_, _17919_, _04523_);
  or (_17921_, _12374_, _09003_);
  and (_17922_, _17860_, _03611_);
  and (_17923_, _17922_, _17921_);
  or (_17925_, _17923_, _17920_);
  and (_17926_, _17925_, _03734_);
  or (_17927_, _17874_, _05674_);
  and (_17928_, _17866_, _03733_);
  and (_17929_, _17928_, _17927_);
  or (_17930_, _17929_, _17926_);
  and (_17931_, _17930_, _03742_);
  or (_17932_, _17909_, _05674_);
  and (_17933_, _17860_, _03618_);
  and (_17934_, _17933_, _17932_);
  or (_17936_, _17865_, _05674_);
  and (_17937_, _17860_, _03741_);
  and (_17938_, _17937_, _17936_);
  or (_17939_, _17938_, _03767_);
  or (_17940_, _17939_, _17934_);
  or (_17941_, _17940_, _17931_);
  or (_17942_, _17863_, _03948_);
  and (_17943_, _17942_, _17941_);
  or (_17944_, _17943_, _03473_);
  or (_17945_, _17874_, _03474_);
  or (_17947_, _17945_, _17861_);
  and (_17948_, _17947_, _43189_);
  and (_17949_, _17948_, _17944_);
  or (_17950_, _17949_, _17859_);
  and (_43762_, _17950_, _42003_);
  not (_17951_, \oc8051_golden_model_1.DPH [2]);
  nor (_17952_, _43189_, _17951_);
  nor (_17953_, _05320_, _17951_);
  nor (_17954_, _12587_, _09003_);
  or (_17955_, _17954_, _17953_);
  and (_17957_, _17955_, _03741_);
  and (_17958_, _12588_, _05320_);
  or (_17959_, _17958_, _17953_);
  and (_17960_, _17959_, _03744_);
  nor (_17961_, _09003_, _05073_);
  or (_17962_, _17961_, _17953_);
  or (_17963_, _17962_, _06903_);
  nor (_17964_, _12467_, _09003_);
  or (_17965_, _17964_, _17953_);
  or (_17966_, _17965_, _04432_);
  and (_17968_, _05320_, \oc8051_golden_model_1.ACC [2]);
  or (_17969_, _17968_, _17953_);
  and (_17970_, _17969_, _04436_);
  nor (_17971_, _04436_, _17951_);
  or (_17972_, _17971_, _03534_);
  or (_17973_, _17972_, _17970_);
  and (_17974_, _17973_, _04457_);
  and (_17975_, _17974_, _17966_);
  and (_17976_, _17962_, _03527_);
  or (_17977_, _17976_, _03530_);
  or (_17979_, _17977_, _17975_);
  or (_17980_, _17969_, _03531_);
  and (_17981_, _17980_, _08924_);
  and (_17982_, _17981_, _17979_);
  or (_17983_, _09029_, \oc8051_golden_model_1.DPH [2]);
  nor (_17984_, _09030_, _08924_);
  and (_17985_, _17984_, _17983_);
  or (_17986_, _17985_, _17982_);
  and (_17987_, _17986_, _03622_);
  nor (_17988_, _03944_, _03622_);
  or (_17990_, _17988_, _07454_);
  or (_17991_, _17990_, _17987_);
  and (_17992_, _17991_, _17963_);
  or (_17993_, _17992_, _04082_);
  and (_17994_, _06710_, _05320_);
  or (_17995_, _17953_, _04500_);
  or (_17996_, _17995_, _17994_);
  and (_17997_, _17996_, _03521_);
  and (_17998_, _17997_, _17993_);
  nor (_17999_, _12568_, _09003_);
  or (_18001_, _17999_, _17953_);
  and (_18002_, _18001_, _03224_);
  or (_18003_, _18002_, _17998_);
  or (_18004_, _18003_, _08905_);
  and (_18005_, _12582_, _05320_);
  or (_18006_, _17953_, _04527_);
  or (_18007_, _18006_, _18005_);
  and (_18008_, _05320_, _06399_);
  or (_18009_, _18008_, _17953_);
  or (_18010_, _18009_, _04509_);
  and (_18012_, _18010_, _03745_);
  and (_18013_, _18012_, _18007_);
  and (_18014_, _18013_, _18004_);
  or (_18015_, _18014_, _17960_);
  and (_18016_, _18015_, _04523_);
  or (_18017_, _17953_, _05772_);
  and (_18018_, _18009_, _03611_);
  and (_18019_, _18018_, _18017_);
  or (_18020_, _18019_, _18016_);
  and (_18021_, _18020_, _03734_);
  and (_18023_, _17969_, _03733_);
  and (_18024_, _18023_, _18017_);
  or (_18025_, _18024_, _03618_);
  or (_18026_, _18025_, _18021_);
  nor (_18027_, _12581_, _09003_);
  or (_18028_, _17953_, _06453_);
  or (_18029_, _18028_, _18027_);
  and (_18030_, _18029_, _06458_);
  and (_18031_, _18030_, _18026_);
  or (_18032_, _18031_, _17957_);
  and (_18034_, _18032_, _03948_);
  and (_18035_, _17965_, _03767_);
  or (_18036_, _18035_, _03473_);
  or (_18037_, _18036_, _18034_);
  and (_18038_, _12638_, _05320_);
  or (_18039_, _17953_, _03474_);
  or (_18040_, _18039_, _18038_);
  and (_18041_, _18040_, _43189_);
  and (_18042_, _18041_, _18037_);
  or (_18043_, _18042_, _17952_);
  and (_43763_, _18043_, _42003_);
  not (_18045_, \oc8051_golden_model_1.DPH [3]);
  nor (_18046_, _43189_, _18045_);
  nor (_18047_, _05320_, _18045_);
  nor (_18048_, _12792_, _09003_);
  or (_18049_, _18048_, _18047_);
  and (_18050_, _18049_, _03741_);
  and (_18051_, _12793_, _05320_);
  or (_18052_, _18051_, _18047_);
  and (_18053_, _18052_, _03744_);
  nor (_18055_, _12652_, _09003_);
  or (_18056_, _18055_, _18047_);
  or (_18057_, _18056_, _04432_);
  and (_18058_, _05320_, \oc8051_golden_model_1.ACC [3]);
  or (_18059_, _18058_, _18047_);
  and (_18060_, _18059_, _04436_);
  nor (_18061_, _04436_, _18045_);
  or (_18062_, _18061_, _03534_);
  or (_18063_, _18062_, _18060_);
  and (_18064_, _18063_, _04457_);
  and (_18066_, _18064_, _18057_);
  nor (_18067_, _09003_, _04885_);
  or (_18068_, _18067_, _18047_);
  and (_18069_, _18068_, _03527_);
  or (_18070_, _18069_, _03530_);
  or (_18071_, _18070_, _18066_);
  or (_18072_, _18059_, _03531_);
  and (_18073_, _18072_, _08924_);
  and (_18074_, _18073_, _18071_);
  or (_18075_, _09030_, \oc8051_golden_model_1.DPH [3]);
  nor (_18077_, _09031_, _08924_);
  and (_18078_, _18077_, _18075_);
  or (_18079_, _18078_, _18074_);
  and (_18080_, _18079_, _03622_);
  nor (_18081_, _03622_, _03440_);
  or (_18082_, _18081_, _07454_);
  or (_18083_, _18082_, _18080_);
  or (_18084_, _18068_, _06903_);
  and (_18085_, _18084_, _18083_);
  or (_18086_, _18085_, _04082_);
  and (_18088_, _06664_, _05320_);
  or (_18089_, _18047_, _04500_);
  or (_18090_, _18089_, _18088_);
  and (_18091_, _18090_, _03521_);
  and (_18092_, _18091_, _18086_);
  nor (_18093_, _12773_, _09003_);
  or (_18094_, _18093_, _18047_);
  and (_18095_, _18094_, _03224_);
  or (_18096_, _18095_, _08905_);
  or (_18097_, _18096_, _18092_);
  and (_18099_, _12787_, _05320_);
  or (_18100_, _18047_, _04527_);
  or (_18101_, _18100_, _18099_);
  and (_18102_, _05320_, _06356_);
  or (_18103_, _18102_, _18047_);
  or (_18104_, _18103_, _04509_);
  and (_18105_, _18104_, _03745_);
  and (_18106_, _18105_, _18101_);
  and (_18107_, _18106_, _18097_);
  or (_18108_, _18107_, _18053_);
  and (_18110_, _18108_, _04523_);
  or (_18111_, _18047_, _05625_);
  and (_18112_, _18103_, _03611_);
  and (_18113_, _18112_, _18111_);
  or (_18114_, _18113_, _18110_);
  and (_18115_, _18114_, _03734_);
  and (_18116_, _18059_, _03733_);
  and (_18117_, _18116_, _18111_);
  or (_18118_, _18117_, _03618_);
  or (_18119_, _18118_, _18115_);
  nor (_18121_, _12786_, _09003_);
  or (_18122_, _18047_, _06453_);
  or (_18123_, _18122_, _18121_);
  and (_18124_, _18123_, _06458_);
  and (_18125_, _18124_, _18119_);
  or (_18126_, _18125_, _18050_);
  and (_18127_, _18126_, _03948_);
  and (_18128_, _18056_, _03767_);
  or (_18129_, _18128_, _03473_);
  or (_18130_, _18129_, _18127_);
  and (_18132_, _12843_, _05320_);
  or (_18133_, _18047_, _03474_);
  or (_18134_, _18133_, _18132_);
  and (_18135_, _18134_, _43189_);
  and (_18136_, _18135_, _18130_);
  or (_18137_, _18136_, _18046_);
  and (_43764_, _18137_, _42003_);
  not (_18138_, \oc8051_golden_model_1.DPH [4]);
  nor (_18139_, _43189_, _18138_);
  nor (_18140_, _05320_, _18138_);
  nor (_18142_, _12991_, _09003_);
  or (_18143_, _18142_, _18140_);
  and (_18144_, _18143_, _03741_);
  nor (_18145_, _05831_, _09003_);
  or (_18146_, _18145_, _18140_);
  or (_18147_, _18146_, _06903_);
  nor (_18148_, _12856_, _09003_);
  or (_18149_, _18148_, _18140_);
  or (_18150_, _18149_, _04432_);
  and (_18151_, _05320_, \oc8051_golden_model_1.ACC [4]);
  or (_18153_, _18151_, _18140_);
  and (_18154_, _18153_, _04436_);
  nor (_18155_, _04436_, _18138_);
  or (_18156_, _18155_, _03534_);
  or (_18157_, _18156_, _18154_);
  and (_18158_, _18157_, _04457_);
  and (_18159_, _18158_, _18150_);
  and (_18160_, _18146_, _03527_);
  or (_18161_, _18160_, _03530_);
  or (_18162_, _18161_, _18159_);
  or (_18164_, _18153_, _03531_);
  and (_18165_, _18164_, _08924_);
  and (_18166_, _18165_, _18162_);
  or (_18167_, _09031_, \oc8051_golden_model_1.DPH [4]);
  nor (_18168_, _09032_, _08924_);
  and (_18169_, _18168_, _18167_);
  or (_18170_, _18169_, _18166_);
  and (_18171_, _18170_, _03622_);
  nor (_18172_, _04257_, _03622_);
  or (_18173_, _18172_, _07454_);
  or (_18175_, _18173_, _18171_);
  and (_18176_, _18175_, _18147_);
  or (_18177_, _18176_, _04082_);
  and (_18178_, _06802_, _05320_);
  or (_18179_, _18140_, _04500_);
  or (_18180_, _18179_, _18178_);
  and (_18181_, _18180_, _03521_);
  and (_18182_, _18181_, _18177_);
  nor (_18183_, _12972_, _09003_);
  or (_18184_, _18183_, _18140_);
  and (_18186_, _18184_, _03224_);
  or (_18187_, _18186_, _18182_);
  or (_18188_, _18187_, _08905_);
  and (_18189_, _12986_, _05320_);
  or (_18190_, _18140_, _04527_);
  or (_18191_, _18190_, _18189_);
  and (_18192_, _06337_, _05320_);
  or (_18193_, _18192_, _18140_);
  or (_18194_, _18193_, _04509_);
  and (_18195_, _18194_, _03745_);
  and (_18197_, _18195_, _18191_);
  and (_18198_, _18197_, _18188_);
  and (_18199_, _12992_, _05320_);
  or (_18200_, _18199_, _18140_);
  and (_18201_, _18200_, _03744_);
  or (_18202_, _18201_, _18198_);
  and (_18203_, _18202_, _04523_);
  or (_18204_, _18140_, _05880_);
  and (_18205_, _18193_, _03611_);
  and (_18206_, _18205_, _18204_);
  or (_18208_, _18206_, _18203_);
  and (_18209_, _18208_, _03734_);
  and (_18210_, _18153_, _03733_);
  and (_18211_, _18210_, _18204_);
  or (_18212_, _18211_, _03618_);
  or (_18213_, _18212_, _18209_);
  nor (_18214_, _12985_, _09003_);
  or (_18215_, _18140_, _06453_);
  or (_18216_, _18215_, _18214_);
  and (_18217_, _18216_, _06458_);
  and (_18219_, _18217_, _18213_);
  or (_18220_, _18219_, _18144_);
  and (_18221_, _18220_, _03948_);
  and (_18222_, _18149_, _03767_);
  or (_18223_, _18222_, _03473_);
  or (_18224_, _18223_, _18221_);
  and (_18225_, _13051_, _05320_);
  or (_18226_, _18140_, _03474_);
  or (_18227_, _18226_, _18225_);
  and (_18228_, _18227_, _43189_);
  and (_18230_, _18228_, _18224_);
  or (_18231_, _18230_, _18139_);
  and (_43765_, _18231_, _42003_);
  not (_18232_, \oc8051_golden_model_1.DPH [5]);
  nor (_18233_, _43189_, _18232_);
  nor (_18234_, _05320_, _18232_);
  nor (_18235_, _13203_, _09003_);
  or (_18236_, _18235_, _18234_);
  and (_18237_, _18236_, _03741_);
  nor (_18238_, _05526_, _09003_);
  or (_18240_, _18238_, _18234_);
  or (_18241_, _18240_, _06903_);
  nor (_18242_, _13070_, _09003_);
  or (_18243_, _18242_, _18234_);
  or (_18244_, _18243_, _04432_);
  and (_18245_, _05320_, \oc8051_golden_model_1.ACC [5]);
  or (_18246_, _18245_, _18234_);
  and (_18247_, _18246_, _04436_);
  nor (_18248_, _04436_, _18232_);
  or (_18249_, _18248_, _03534_);
  or (_18251_, _18249_, _18247_);
  and (_18252_, _18251_, _04457_);
  and (_18253_, _18252_, _18244_);
  and (_18254_, _18240_, _03527_);
  or (_18255_, _18254_, _03530_);
  or (_18256_, _18255_, _18253_);
  or (_18257_, _18246_, _03531_);
  and (_18258_, _18257_, _08924_);
  and (_18259_, _18258_, _18256_);
  or (_18260_, _09032_, \oc8051_golden_model_1.DPH [5]);
  nor (_18262_, _09033_, _08924_);
  and (_18263_, _18262_, _18260_);
  or (_18264_, _18263_, _18259_);
  and (_18265_, _18264_, _03622_);
  nor (_18266_, _03811_, _03622_);
  or (_18267_, _18266_, _07454_);
  or (_18268_, _18267_, _18265_);
  and (_18269_, _18268_, _18241_);
  or (_18270_, _18269_, _04082_);
  and (_18271_, _06757_, _05320_);
  or (_18273_, _18234_, _04500_);
  or (_18274_, _18273_, _18271_);
  and (_18275_, _18274_, _03521_);
  and (_18276_, _18275_, _18270_);
  nor (_18277_, _13184_, _09003_);
  or (_18278_, _18277_, _18234_);
  and (_18279_, _18278_, _03224_);
  or (_18280_, _18279_, _18276_);
  or (_18281_, _18280_, _08905_);
  and (_18282_, _13198_, _05320_);
  or (_18284_, _18234_, _04527_);
  or (_18285_, _18284_, _18282_);
  and (_18286_, _06295_, _05320_);
  or (_18287_, _18286_, _18234_);
  or (_18288_, _18287_, _04509_);
  and (_18289_, _18288_, _03745_);
  and (_18290_, _18289_, _18285_);
  and (_18291_, _18290_, _18281_);
  and (_18292_, _13204_, _05320_);
  or (_18293_, _18292_, _18234_);
  and (_18295_, _18293_, _03744_);
  or (_18296_, _18295_, _18291_);
  and (_18297_, _18296_, _04523_);
  or (_18298_, _18234_, _05576_);
  and (_18299_, _18287_, _03611_);
  and (_18300_, _18299_, _18298_);
  or (_18301_, _18300_, _18297_);
  and (_18302_, _18301_, _03734_);
  and (_18303_, _18246_, _03733_);
  and (_18304_, _18303_, _18298_);
  or (_18306_, _18304_, _03618_);
  or (_18307_, _18306_, _18302_);
  nor (_18308_, _13197_, _09003_);
  or (_18309_, _18234_, _06453_);
  or (_18310_, _18309_, _18308_);
  and (_18311_, _18310_, _06458_);
  and (_18312_, _18311_, _18307_);
  or (_18313_, _18312_, _18237_);
  and (_18314_, _18313_, _03948_);
  and (_18315_, _18243_, _03767_);
  or (_18317_, _18315_, _03473_);
  or (_18318_, _18317_, _18314_);
  and (_18319_, _13253_, _05320_);
  or (_18320_, _18234_, _03474_);
  or (_18321_, _18320_, _18319_);
  and (_18322_, _18321_, _43189_);
  and (_18323_, _18322_, _18318_);
  or (_18324_, _18323_, _18233_);
  and (_43766_, _18324_, _42003_);
  not (_18325_, \oc8051_golden_model_1.DPH [6]);
  nor (_18327_, _43189_, _18325_);
  nor (_18328_, _05320_, _18325_);
  nor (_18329_, _13406_, _09003_);
  or (_18330_, _18329_, _18328_);
  and (_18331_, _18330_, _03741_);
  nor (_18332_, _05417_, _09003_);
  or (_18333_, _18332_, _18328_);
  or (_18334_, _18333_, _06903_);
  nor (_18335_, _13293_, _09003_);
  or (_18336_, _18335_, _18328_);
  or (_18338_, _18336_, _04432_);
  and (_18339_, _05320_, \oc8051_golden_model_1.ACC [6]);
  or (_18340_, _18339_, _18328_);
  and (_18341_, _18340_, _04436_);
  nor (_18342_, _04436_, _18325_);
  or (_18343_, _18342_, _03534_);
  or (_18344_, _18343_, _18341_);
  and (_18345_, _18344_, _04457_);
  and (_18346_, _18345_, _18338_);
  and (_18347_, _18333_, _03527_);
  or (_18349_, _18347_, _03530_);
  or (_18350_, _18349_, _18346_);
  or (_18351_, _18340_, _03531_);
  and (_18352_, _18351_, _08924_);
  and (_18353_, _18352_, _18350_);
  or (_18354_, _09033_, \oc8051_golden_model_1.DPH [6]);
  and (_18355_, _09034_, _08923_);
  and (_18356_, _18355_, _18354_);
  or (_18357_, _18356_, _18353_);
  and (_18358_, _18357_, _03622_);
  nor (_18360_, _03622_, _03511_);
  or (_18361_, _18360_, _07454_);
  or (_18362_, _18361_, _18358_);
  and (_18363_, _18362_, _18334_);
  or (_18364_, _18363_, _04082_);
  and (_18365_, _06526_, _05320_);
  or (_18366_, _18328_, _04500_);
  or (_18367_, _18366_, _18365_);
  and (_18368_, _18367_, _03521_);
  and (_18369_, _18368_, _18364_);
  nor (_18371_, _13387_, _09003_);
  or (_18372_, _18371_, _18328_);
  and (_18373_, _18372_, _03224_);
  or (_18374_, _18373_, _18369_);
  or (_18375_, _18374_, _08905_);
  and (_18376_, _13402_, _05320_);
  or (_18377_, _18328_, _04527_);
  or (_18378_, _18377_, _18376_);
  and (_18379_, _14949_, _05320_);
  or (_18380_, _18379_, _18328_);
  or (_18382_, _18380_, _04509_);
  and (_18383_, _18382_, _03745_);
  and (_18384_, _18383_, _18378_);
  and (_18385_, _18384_, _18375_);
  and (_18386_, _13407_, _05320_);
  or (_18387_, _18386_, _18328_);
  and (_18388_, _18387_, _03744_);
  or (_18389_, _18388_, _18385_);
  and (_18390_, _18389_, _04523_);
  or (_18391_, _18328_, _05469_);
  and (_18393_, _18380_, _03611_);
  and (_18394_, _18393_, _18391_);
  or (_18395_, _18394_, _18390_);
  and (_18396_, _18395_, _03734_);
  and (_18397_, _18340_, _03733_);
  and (_18398_, _18397_, _18391_);
  or (_18399_, _18398_, _03618_);
  or (_18400_, _18399_, _18396_);
  nor (_18401_, _13400_, _09003_);
  or (_18402_, _18328_, _06453_);
  or (_18404_, _18402_, _18401_);
  and (_18405_, _18404_, _06458_);
  and (_18406_, _18405_, _18400_);
  or (_18407_, _18406_, _18331_);
  and (_18408_, _18407_, _03948_);
  and (_18409_, _18336_, _03767_);
  or (_18410_, _18409_, _03473_);
  or (_18411_, _18410_, _18408_);
  and (_18412_, _13456_, _05320_);
  or (_18413_, _18328_, _03474_);
  or (_18415_, _18413_, _18412_);
  and (_18416_, _18415_, _43189_);
  and (_18417_, _18416_, _18411_);
  or (_18418_, _18417_, _18327_);
  and (_43767_, _18418_, _42003_);
  not (_18419_, \oc8051_golden_model_1.IE [0]);
  nor (_18420_, _05278_, _18419_);
  and (_18421_, _12183_, _05278_);
  nor (_18422_, _18421_, _18420_);
  nor (_18423_, _18422_, _03745_);
  and (_18425_, _05278_, _06350_);
  nor (_18426_, _18425_, _18420_);
  and (_18427_, _18426_, _03624_);
  and (_18428_, _05278_, _04429_);
  nor (_18429_, _18428_, _18420_);
  and (_18430_, _18429_, _07454_);
  and (_18431_, _05278_, \oc8051_golden_model_1.ACC [0]);
  nor (_18432_, _18431_, _18420_);
  nor (_18433_, _18432_, _04437_);
  nor (_18434_, _04436_, _18419_);
  or (_18436_, _18434_, _18433_);
  and (_18437_, _18436_, _04432_);
  nor (_18438_, _05722_, _09097_);
  nor (_18439_, _18438_, _18420_);
  nor (_18440_, _18439_, _04432_);
  or (_18441_, _18440_, _18437_);
  and (_18442_, _18441_, _03470_);
  nor (_18443_, _05944_, _18419_);
  and (_18444_, _12075_, _05944_);
  nor (_18445_, _18444_, _18443_);
  nor (_18447_, _18445_, _03470_);
  nor (_18448_, _18447_, _18442_);
  nor (_18449_, _18448_, _03527_);
  nor (_18450_, _18429_, _04457_);
  or (_18451_, _18450_, _18449_);
  and (_18452_, _18451_, _03531_);
  nor (_18453_, _18432_, _03531_);
  or (_18454_, _18453_, _18452_);
  and (_18455_, _18454_, _03466_);
  and (_18456_, _18420_, _03465_);
  or (_18458_, _18456_, _18455_);
  and (_18459_, _18458_, _03459_);
  nor (_18460_, _18439_, _03459_);
  or (_18461_, _18460_, _18459_);
  and (_18462_, _18461_, _03453_);
  nor (_18463_, _12106_, _09134_);
  nor (_18464_, _18463_, _18443_);
  nor (_18465_, _18464_, _03453_);
  or (_18466_, _18465_, _07454_);
  nor (_18467_, _18466_, _18462_);
  nor (_18469_, _18467_, _18430_);
  nor (_18470_, _18469_, _04082_);
  and (_18471_, _06617_, _05278_);
  nor (_18472_, _18420_, _04500_);
  not (_18473_, _18472_);
  nor (_18474_, _18473_, _18471_);
  or (_18475_, _18474_, _03224_);
  nor (_18476_, _18475_, _18470_);
  nor (_18477_, _12164_, _09097_);
  nor (_18478_, _18477_, _18420_);
  nor (_18480_, _18478_, _03521_);
  or (_18481_, _18480_, _03624_);
  nor (_18482_, _18481_, _18476_);
  nor (_18483_, _18482_, _18427_);
  or (_18484_, _18483_, _03623_);
  and (_18485_, _12177_, _05278_);
  or (_18486_, _18485_, _18420_);
  or (_18487_, _18486_, _04527_);
  and (_18488_, _18487_, _03745_);
  and (_18489_, _18488_, _18484_);
  nor (_18491_, _18489_, _18423_);
  nor (_18492_, _18491_, _03611_);
  or (_18493_, _18426_, _04523_);
  nor (_18494_, _18493_, _18438_);
  nor (_18495_, _18494_, _18492_);
  nor (_18496_, _18495_, _03733_);
  and (_18497_, _12182_, _05278_);
  or (_18498_, _18497_, _18420_);
  and (_18499_, _18498_, _03733_);
  or (_18500_, _18499_, _18496_);
  and (_18502_, _18500_, _06453_);
  nor (_18503_, _12057_, _09097_);
  nor (_18504_, _18503_, _18420_);
  nor (_18505_, _18504_, _06453_);
  or (_18506_, _18505_, _18502_);
  and (_18507_, _18506_, _06458_);
  nor (_18508_, _12181_, _09097_);
  nor (_18509_, _18508_, _18420_);
  nor (_18510_, _18509_, _06458_);
  or (_18511_, _18510_, _18507_);
  and (_18513_, _18511_, _03948_);
  nor (_18514_, _18439_, _03948_);
  or (_18515_, _18514_, _18513_);
  and (_18516_, _18515_, _03446_);
  and (_18517_, _18420_, _03445_);
  nor (_18518_, _18517_, _18516_);
  or (_18519_, _18518_, _03473_);
  or (_18520_, _18439_, _03474_);
  and (_18521_, _18520_, _18519_);
  nand (_18522_, _18521_, _43189_);
  or (_18524_, _43189_, \oc8051_golden_model_1.IE [0]);
  and (_18525_, _18524_, _42003_);
  and (_43769_, _18525_, _18522_);
  not (_18526_, _03742_);
  not (_18527_, \oc8051_golden_model_1.IE [1]);
  nor (_18528_, _05278_, _18527_);
  and (_18529_, _06572_, _05278_);
  or (_18530_, _18529_, _18528_);
  and (_18531_, _18530_, _04082_);
  nor (_18532_, _05278_, \oc8051_golden_model_1.IE [1]);
  and (_18534_, _05278_, _03269_);
  nor (_18535_, _18534_, _18532_);
  and (_18536_, _18535_, _04436_);
  nor (_18537_, _04436_, _18527_);
  or (_18538_, _18537_, _18536_);
  and (_18539_, _18538_, _04432_);
  and (_18540_, _12265_, _05278_);
  nor (_18541_, _18540_, _18532_);
  and (_18542_, _18541_, _03534_);
  or (_18543_, _18542_, _18539_);
  and (_18545_, _18543_, _03470_);
  and (_18546_, _12269_, _05944_);
  nor (_18547_, _05944_, _18527_);
  or (_18548_, _18547_, _03527_);
  or (_18549_, _18548_, _18546_);
  and (_18550_, _18549_, _03533_);
  nor (_18551_, _18550_, _18545_);
  nor (_18552_, _09097_, _04635_);
  nor (_18553_, _18552_, _18528_);
  and (_18554_, _18553_, _03527_);
  nor (_18556_, _18554_, _18551_);
  and (_18557_, _18556_, _03531_);
  and (_18558_, _18535_, _03530_);
  or (_18559_, _18558_, _18557_);
  and (_18560_, _18559_, _03466_);
  and (_18561_, _12256_, _05944_);
  nor (_18562_, _18561_, _18547_);
  nor (_18563_, _18562_, _03466_);
  or (_18564_, _18563_, _03458_);
  or (_18565_, _18564_, _18560_);
  and (_18567_, _18546_, _12284_);
  or (_18568_, _18547_, _03459_);
  or (_18569_, _18568_, _18567_);
  and (_18570_, _18569_, _18565_);
  and (_18571_, _18570_, _03453_);
  nor (_18572_, _12301_, _09134_);
  nor (_18573_, _18547_, _18572_);
  nor (_18574_, _18573_, _03453_);
  or (_18575_, _18574_, _07454_);
  nor (_18576_, _18575_, _18571_);
  and (_18578_, _18553_, _07454_);
  or (_18579_, _18578_, _04082_);
  nor (_18580_, _18579_, _18576_);
  or (_18581_, _18580_, _18531_);
  and (_18582_, _18581_, _03521_);
  nor (_18583_, _12360_, _09097_);
  nor (_18584_, _18583_, _18528_);
  nor (_18585_, _18584_, _03521_);
  nor (_18586_, _18585_, _18582_);
  nor (_18587_, _18586_, _08905_);
  not (_18589_, _18532_);
  nor (_18590_, _12375_, _09097_);
  nor (_18591_, _18590_, _04527_);
  and (_18592_, _05278_, _04325_);
  nor (_18593_, _18592_, _04509_);
  or (_18594_, _18593_, _18591_);
  and (_18595_, _18594_, _18589_);
  nor (_18596_, _18595_, _18587_);
  nor (_18597_, _18596_, _03744_);
  nor (_18598_, _12381_, _09097_);
  nor (_18600_, _18598_, _03745_);
  and (_18601_, _18600_, _18589_);
  nor (_18602_, _18601_, _18597_);
  nor (_18603_, _18602_, _03611_);
  nor (_18604_, _12374_, _09097_);
  nor (_18605_, _18604_, _04523_);
  and (_18606_, _18605_, _18589_);
  nor (_18607_, _18606_, _18603_);
  nor (_18608_, _18607_, _03733_);
  nor (_18609_, _18528_, _05674_);
  nor (_18611_, _18609_, _03734_);
  and (_18612_, _18611_, _18535_);
  nor (_18613_, _18612_, _18608_);
  or (_18614_, _18613_, _18526_);
  and (_18615_, _18592_, _05673_);
  nor (_18616_, _18615_, _06453_);
  and (_18617_, _18616_, _18589_);
  and (_18618_, _18534_, _05673_);
  or (_18619_, _18532_, _06458_);
  nor (_18620_, _18619_, _18618_);
  or (_18622_, _18620_, _03767_);
  nor (_18623_, _18622_, _18617_);
  and (_18624_, _18623_, _18614_);
  nor (_18625_, _18541_, _03948_);
  or (_18626_, _18625_, _03445_);
  nor (_18627_, _18626_, _18624_);
  nor (_18628_, _18562_, _03446_);
  or (_18629_, _18628_, _03473_);
  nor (_18630_, _18629_, _18627_);
  or (_18631_, _18528_, _03474_);
  nor (_18633_, _18631_, _18540_);
  nor (_18634_, _18633_, _18630_);
  or (_18635_, _18634_, _43193_);
  or (_18636_, _43189_, \oc8051_golden_model_1.IE [1]);
  and (_18637_, _18636_, _42003_);
  and (_43770_, _18637_, _18635_);
  not (_18638_, \oc8051_golden_model_1.IE [2]);
  nor (_18639_, _05278_, _18638_);
  and (_18640_, _05278_, _06399_);
  nor (_18641_, _18640_, _18639_);
  and (_18643_, _18641_, _03624_);
  nor (_18644_, _09097_, _05073_);
  nor (_18645_, _18644_, _18639_);
  and (_18646_, _18645_, _07454_);
  and (_18647_, _05278_, \oc8051_golden_model_1.ACC [2]);
  nor (_18648_, _18647_, _18639_);
  nor (_18649_, _18648_, _04437_);
  nor (_18650_, _04436_, _18638_);
  or (_18651_, _18650_, _18649_);
  and (_18652_, _18651_, _04432_);
  nor (_18654_, _12467_, _09097_);
  nor (_18655_, _18654_, _18639_);
  nor (_18656_, _18655_, _04432_);
  or (_18657_, _18656_, _18652_);
  and (_18658_, _18657_, _03470_);
  nor (_18659_, _05944_, _18638_);
  and (_18660_, _12462_, _05944_);
  nor (_18661_, _18660_, _18659_);
  nor (_18662_, _18661_, _03470_);
  or (_18663_, _18662_, _18658_);
  and (_18665_, _18663_, _04457_);
  nor (_18666_, _18645_, _04457_);
  or (_18667_, _18666_, _18665_);
  and (_18668_, _18667_, _03531_);
  nor (_18669_, _18648_, _03531_);
  or (_18670_, _18669_, _18668_);
  and (_18671_, _18670_, _03466_);
  and (_18672_, _12460_, _05944_);
  nor (_18673_, _18672_, _18659_);
  nor (_18674_, _18673_, _03466_);
  or (_18676_, _18674_, _03458_);
  or (_18677_, _18676_, _18671_);
  and (_18678_, _18660_, _12491_);
  or (_18679_, _18659_, _03459_);
  or (_18680_, _18679_, _18678_);
  and (_18681_, _18680_, _03453_);
  and (_18682_, _18681_, _18677_);
  nor (_18683_, _12509_, _09134_);
  nor (_18684_, _18683_, _18659_);
  nor (_18685_, _18684_, _03453_);
  nor (_18687_, _18685_, _07454_);
  not (_18688_, _18687_);
  nor (_18689_, _18688_, _18682_);
  nor (_18690_, _18689_, _18646_);
  nor (_18691_, _18690_, _04082_);
  and (_18692_, _06710_, _05278_);
  nor (_18693_, _18639_, _04500_);
  not (_18694_, _18693_);
  nor (_18695_, _18694_, _18692_);
  or (_18696_, _18695_, _03224_);
  nor (_18698_, _18696_, _18691_);
  nor (_18699_, _12568_, _09097_);
  nor (_18700_, _18639_, _18699_);
  nor (_18701_, _18700_, _03521_);
  or (_18702_, _18701_, _03624_);
  nor (_18703_, _18702_, _18698_);
  nor (_18704_, _18703_, _18643_);
  or (_18705_, _18704_, _03623_);
  and (_18706_, _12582_, _05278_);
  or (_18707_, _18706_, _18639_);
  or (_18709_, _18707_, _04527_);
  and (_18710_, _18709_, _03745_);
  and (_18711_, _18710_, _18705_);
  and (_18712_, _12588_, _05278_);
  nor (_18713_, _18712_, _18639_);
  nor (_18714_, _18713_, _03745_);
  nor (_18715_, _18714_, _18711_);
  nor (_18716_, _18715_, _03611_);
  nor (_18717_, _18639_, _05772_);
  not (_18718_, _18717_);
  nor (_18720_, _18641_, _04523_);
  and (_18721_, _18720_, _18718_);
  nor (_18722_, _18721_, _18716_);
  nor (_18723_, _18722_, _03733_);
  nor (_18724_, _18648_, _03734_);
  and (_18725_, _18724_, _18718_);
  or (_18726_, _18725_, _18723_);
  and (_18727_, _18726_, _06453_);
  nor (_18728_, _12581_, _09097_);
  nor (_18729_, _18728_, _18639_);
  nor (_18731_, _18729_, _06453_);
  or (_18732_, _18731_, _18727_);
  and (_18733_, _18732_, _06458_);
  nor (_18734_, _12587_, _09097_);
  nor (_18735_, _18734_, _18639_);
  nor (_18736_, _18735_, _06458_);
  or (_18737_, _18736_, _18733_);
  and (_18738_, _18737_, _03948_);
  nor (_18739_, _18655_, _03948_);
  or (_18740_, _18739_, _18738_);
  and (_18742_, _18740_, _03446_);
  nor (_18743_, _18673_, _03446_);
  or (_18744_, _18743_, _18742_);
  and (_18745_, _18744_, _03474_);
  and (_18746_, _12638_, _05278_);
  nor (_18747_, _18746_, _18639_);
  nor (_18748_, _18747_, _03474_);
  or (_18749_, _18748_, _18745_);
  or (_18750_, _18749_, _43193_);
  or (_18751_, _43189_, \oc8051_golden_model_1.IE [2]);
  and (_18753_, _18751_, _42003_);
  and (_43771_, _18753_, _18750_);
  not (_18754_, \oc8051_golden_model_1.IE [3]);
  nor (_18755_, _05278_, _18754_);
  and (_18756_, _05278_, _06356_);
  nor (_18757_, _18756_, _18755_);
  and (_18758_, _18757_, _03624_);
  nor (_18759_, _09097_, _04885_);
  nor (_18760_, _18759_, _18755_);
  and (_18761_, _18760_, _07454_);
  and (_18763_, _05278_, \oc8051_golden_model_1.ACC [3]);
  nor (_18764_, _18763_, _18755_);
  nor (_18765_, _18764_, _04437_);
  nor (_18766_, _04436_, _18754_);
  or (_18767_, _18766_, _18765_);
  and (_18768_, _18767_, _04432_);
  nor (_18769_, _12652_, _09097_);
  nor (_18770_, _18769_, _18755_);
  nor (_18771_, _18770_, _04432_);
  or (_18772_, _18771_, _18768_);
  and (_18774_, _18772_, _03470_);
  nor (_18775_, _05944_, _18754_);
  and (_18776_, _12664_, _05944_);
  nor (_18777_, _18776_, _18775_);
  nor (_18778_, _18777_, _03470_);
  or (_18779_, _18778_, _03527_);
  or (_18780_, _18779_, _18774_);
  nand (_18781_, _18760_, _03527_);
  and (_18782_, _18781_, _18780_);
  and (_18783_, _18782_, _03531_);
  nor (_18785_, _18764_, _03531_);
  or (_18786_, _18785_, _18783_);
  and (_18787_, _18786_, _03466_);
  and (_18788_, _12662_, _05944_);
  nor (_18789_, _18788_, _18775_);
  nor (_18790_, _18789_, _03466_);
  or (_18791_, _18790_, _03458_);
  or (_18792_, _18791_, _18787_);
  nor (_18793_, _18775_, _12691_);
  nor (_18794_, _18793_, _18777_);
  or (_18796_, _18794_, _03459_);
  and (_18797_, _18796_, _03453_);
  and (_18798_, _18797_, _18792_);
  nor (_18799_, _12709_, _09134_);
  nor (_18800_, _18799_, _18775_);
  nor (_18801_, _18800_, _03453_);
  nor (_18802_, _18801_, _07454_);
  not (_18803_, _18802_);
  nor (_18804_, _18803_, _18798_);
  nor (_18805_, _18804_, _18761_);
  nor (_18807_, _18805_, _04082_);
  and (_18808_, _06664_, _05278_);
  nor (_18809_, _18755_, _04500_);
  not (_18810_, _18809_);
  nor (_18811_, _18810_, _18808_);
  or (_18812_, _18811_, _03224_);
  nor (_18813_, _18812_, _18807_);
  nor (_18814_, _12773_, _09097_);
  nor (_18815_, _18755_, _18814_);
  nor (_18816_, _18815_, _03521_);
  or (_18818_, _18816_, _03624_);
  nor (_18819_, _18818_, _18813_);
  nor (_18820_, _18819_, _18758_);
  or (_18821_, _18820_, _03623_);
  and (_18822_, _12787_, _05278_);
  or (_18823_, _18822_, _18755_);
  or (_18824_, _18823_, _04527_);
  and (_18825_, _18824_, _03745_);
  and (_18826_, _18825_, _18821_);
  and (_18827_, _12793_, _05278_);
  nor (_18829_, _18827_, _18755_);
  nor (_18830_, _18829_, _03745_);
  nor (_18831_, _18830_, _18826_);
  nor (_18832_, _18831_, _03611_);
  nor (_18833_, _18755_, _05625_);
  not (_18834_, _18833_);
  nor (_18835_, _18757_, _04523_);
  and (_18836_, _18835_, _18834_);
  nor (_18837_, _18836_, _18832_);
  nor (_18838_, _18837_, _03733_);
  nor (_18840_, _18764_, _03734_);
  and (_18841_, _18840_, _18834_);
  nor (_18842_, _18841_, _03618_);
  not (_18843_, _18842_);
  nor (_18844_, _18843_, _18838_);
  nor (_18845_, _12786_, _09097_);
  or (_18846_, _18755_, _06453_);
  nor (_18847_, _18846_, _18845_);
  or (_18848_, _18847_, _03741_);
  nor (_18849_, _18848_, _18844_);
  nor (_18851_, _12792_, _09097_);
  nor (_18852_, _18851_, _18755_);
  nor (_18853_, _18852_, _06458_);
  or (_18854_, _18853_, _18849_);
  and (_18855_, _18854_, _03948_);
  nor (_18856_, _18770_, _03948_);
  or (_18857_, _18856_, _18855_);
  and (_18858_, _18857_, _03446_);
  nor (_18859_, _18789_, _03446_);
  or (_18860_, _18859_, _18858_);
  and (_18862_, _18860_, _03474_);
  and (_18863_, _12843_, _05278_);
  nor (_18864_, _18863_, _18755_);
  nor (_18865_, _18864_, _03474_);
  or (_18866_, _18865_, _18862_);
  or (_18867_, _18866_, _43193_);
  or (_18868_, _43189_, \oc8051_golden_model_1.IE [3]);
  and (_18869_, _18868_, _42003_);
  and (_43772_, _18869_, _18867_);
  not (_18870_, \oc8051_golden_model_1.IE [4]);
  nor (_18872_, _05278_, _18870_);
  nor (_18873_, _05831_, _09097_);
  nor (_18874_, _18873_, _18872_);
  and (_18875_, _18874_, _07454_);
  nor (_18876_, _05944_, _18870_);
  and (_18877_, _12864_, _05944_);
  nor (_18878_, _18877_, _18876_);
  nor (_18879_, _18878_, _03466_);
  and (_18880_, _05278_, \oc8051_golden_model_1.ACC [4]);
  nor (_18881_, _18880_, _18872_);
  nor (_18883_, _18881_, _04437_);
  nor (_18884_, _04436_, _18870_);
  or (_18885_, _18884_, _18883_);
  and (_18886_, _18885_, _04432_);
  nor (_18887_, _12856_, _09097_);
  nor (_18888_, _18887_, _18872_);
  nor (_18889_, _18888_, _04432_);
  or (_18890_, _18889_, _18886_);
  and (_18891_, _18890_, _03470_);
  and (_18892_, _12866_, _05944_);
  nor (_18894_, _18892_, _18876_);
  nor (_18895_, _18894_, _03470_);
  or (_18896_, _18895_, _03527_);
  or (_18897_, _18896_, _18891_);
  nand (_18898_, _18874_, _03527_);
  and (_18899_, _18898_, _18897_);
  and (_18900_, _18899_, _03531_);
  nor (_18901_, _18881_, _03531_);
  or (_18902_, _18901_, _18900_);
  and (_18903_, _18902_, _03466_);
  nor (_18905_, _18903_, _18879_);
  nor (_18906_, _18905_, _03458_);
  and (_18907_, _12895_, _05944_);
  nor (_18908_, _18907_, _18876_);
  nor (_18909_, _18908_, _03459_);
  nor (_18910_, _18909_, _18906_);
  nor (_18911_, _18910_, _03452_);
  nor (_18912_, _12912_, _09134_);
  nor (_18913_, _18912_, _18876_);
  nor (_18914_, _18913_, _03453_);
  nor (_18916_, _18914_, _07454_);
  not (_18917_, _18916_);
  nor (_18918_, _18917_, _18911_);
  nor (_18919_, _18918_, _18875_);
  nor (_18920_, _18919_, _04082_);
  and (_18921_, _06802_, _05278_);
  nor (_18922_, _18872_, _04500_);
  not (_18923_, _18922_);
  nor (_18924_, _18923_, _18921_);
  nor (_18925_, _18924_, _03224_);
  not (_18927_, _18925_);
  nor (_18928_, _18927_, _18920_);
  nor (_18929_, _12972_, _09097_);
  nor (_18930_, _18929_, _18872_);
  nor (_18931_, _18930_, _03521_);
  or (_18932_, _18931_, _08905_);
  or (_18933_, _18932_, _18928_);
  and (_18934_, _12986_, _05278_);
  or (_18935_, _18872_, _04527_);
  or (_18936_, _18935_, _18934_);
  and (_18938_, _06337_, _05278_);
  nor (_18939_, _18938_, _18872_);
  and (_18940_, _18939_, _03624_);
  nor (_18941_, _18940_, _03744_);
  and (_18942_, _18941_, _18936_);
  and (_18943_, _18942_, _18933_);
  and (_18944_, _12992_, _05278_);
  nor (_18945_, _18944_, _18872_);
  nor (_18946_, _18945_, _03745_);
  nor (_18947_, _18946_, _18943_);
  nor (_18949_, _18947_, _03611_);
  nor (_18950_, _18872_, _05880_);
  not (_18951_, _18950_);
  nor (_18952_, _18939_, _04523_);
  and (_18953_, _18952_, _18951_);
  nor (_18954_, _18953_, _18949_);
  nor (_18955_, _18954_, _03733_);
  nor (_18956_, _18881_, _03734_);
  and (_18957_, _18956_, _18951_);
  or (_18958_, _18957_, _18955_);
  and (_18960_, _18958_, _06453_);
  nor (_18961_, _12985_, _09097_);
  nor (_18962_, _18961_, _18872_);
  nor (_18963_, _18962_, _06453_);
  or (_18964_, _18963_, _18960_);
  and (_18965_, _18964_, _06458_);
  nor (_18966_, _12991_, _09097_);
  nor (_18967_, _18966_, _18872_);
  nor (_18968_, _18967_, _06458_);
  or (_18969_, _18968_, _18965_);
  and (_18971_, _18969_, _03948_);
  nor (_18972_, _18888_, _03948_);
  or (_18973_, _18972_, _18971_);
  and (_18974_, _18973_, _03446_);
  nor (_18975_, _18878_, _03446_);
  or (_18976_, _18975_, _18974_);
  and (_18977_, _18976_, _03474_);
  and (_18978_, _13051_, _05278_);
  nor (_18979_, _18978_, _18872_);
  nor (_18980_, _18979_, _03474_);
  or (_18982_, _18980_, _18977_);
  or (_18983_, _18982_, _43193_);
  or (_18984_, _43189_, \oc8051_golden_model_1.IE [4]);
  and (_18985_, _18984_, _42003_);
  and (_43773_, _18985_, _18983_);
  not (_18986_, \oc8051_golden_model_1.IE [5]);
  nor (_18987_, _05278_, _18986_);
  and (_18988_, _06757_, _05278_);
  or (_18989_, _18988_, _18987_);
  and (_18990_, _18989_, _04082_);
  and (_18992_, _05278_, \oc8051_golden_model_1.ACC [5]);
  nor (_18993_, _18992_, _18987_);
  nor (_18994_, _18993_, _04437_);
  nor (_18995_, _04436_, _18986_);
  or (_18996_, _18995_, _18994_);
  and (_18997_, _18996_, _04432_);
  nor (_18998_, _13070_, _09097_);
  nor (_18999_, _18998_, _18987_);
  nor (_19000_, _18999_, _04432_);
  or (_19001_, _19000_, _18997_);
  and (_19003_, _19001_, _03470_);
  nor (_19004_, _05944_, _18986_);
  and (_19005_, _13095_, _05944_);
  nor (_19006_, _19005_, _19004_);
  nor (_19007_, _19006_, _03470_);
  or (_19008_, _19007_, _03527_);
  or (_19009_, _19008_, _19003_);
  nor (_19010_, _05526_, _09097_);
  nor (_19011_, _19010_, _18987_);
  nand (_19012_, _19011_, _03527_);
  and (_19014_, _19012_, _19009_);
  and (_19015_, _19014_, _03531_);
  nor (_19016_, _18993_, _03531_);
  or (_19017_, _19016_, _19015_);
  and (_19018_, _19017_, _03466_);
  and (_19019_, _13078_, _05944_);
  nor (_19020_, _19019_, _19004_);
  nor (_19021_, _19020_, _03466_);
  or (_19022_, _19021_, _03458_);
  or (_19023_, _19022_, _19018_);
  nor (_19025_, _19004_, _13110_);
  nor (_19026_, _19025_, _19006_);
  or (_19027_, _19026_, _03459_);
  and (_19028_, _19027_, _03453_);
  and (_19029_, _19028_, _19023_);
  nor (_19030_, _13076_, _09134_);
  nor (_19031_, _19030_, _19004_);
  nor (_19032_, _19031_, _03453_);
  nor (_19033_, _19032_, _07454_);
  not (_19034_, _19033_);
  nor (_19036_, _19034_, _19029_);
  and (_19037_, _19011_, _07454_);
  or (_19038_, _19037_, _04082_);
  nor (_19039_, _19038_, _19036_);
  or (_19040_, _19039_, _18990_);
  and (_19041_, _19040_, _03521_);
  nor (_19042_, _13184_, _09097_);
  nor (_19043_, _19042_, _18987_);
  nor (_19044_, _19043_, _03521_);
  or (_19045_, _19044_, _08905_);
  or (_19047_, _19045_, _19041_);
  and (_19048_, _13198_, _05278_);
  or (_19049_, _18987_, _04527_);
  or (_19050_, _19049_, _19048_);
  and (_19051_, _06295_, _05278_);
  nor (_19052_, _19051_, _18987_);
  and (_19053_, _19052_, _03624_);
  nor (_19054_, _19053_, _03744_);
  and (_19055_, _19054_, _19050_);
  and (_19056_, _19055_, _19047_);
  and (_19058_, _13204_, _05278_);
  nor (_19059_, _19058_, _18987_);
  nor (_19060_, _19059_, _03745_);
  nor (_19061_, _19060_, _19056_);
  nor (_19062_, _19061_, _03611_);
  nor (_19063_, _18987_, _05576_);
  not (_19064_, _19063_);
  nor (_19065_, _19052_, _04523_);
  and (_19066_, _19065_, _19064_);
  nor (_19067_, _19066_, _19062_);
  nor (_19069_, _19067_, _03733_);
  nor (_19070_, _18993_, _03734_);
  and (_19071_, _19070_, _19064_);
  or (_19072_, _19071_, _19069_);
  and (_19073_, _19072_, _06453_);
  nor (_19074_, _13197_, _09097_);
  nor (_19075_, _19074_, _18987_);
  nor (_19076_, _19075_, _06453_);
  or (_19077_, _19076_, _19073_);
  and (_19078_, _19077_, _06458_);
  nor (_19080_, _13203_, _09097_);
  nor (_19081_, _19080_, _18987_);
  nor (_19082_, _19081_, _06458_);
  or (_19083_, _19082_, _19078_);
  and (_19084_, _19083_, _03948_);
  nor (_19085_, _18999_, _03948_);
  or (_19086_, _19085_, _19084_);
  and (_19087_, _19086_, _03446_);
  nor (_19088_, _19020_, _03446_);
  or (_19089_, _19088_, _19087_);
  and (_19091_, _19089_, _03474_);
  and (_19092_, _13253_, _05278_);
  nor (_19093_, _19092_, _18987_);
  nor (_19094_, _19093_, _03474_);
  or (_19095_, _19094_, _19091_);
  or (_19096_, _19095_, _43193_);
  or (_19097_, _43189_, \oc8051_golden_model_1.IE [5]);
  and (_19098_, _19097_, _42003_);
  and (_43774_, _19098_, _19096_);
  not (_19099_, \oc8051_golden_model_1.IE [6]);
  nor (_19101_, _05278_, _19099_);
  and (_19102_, _06526_, _05278_);
  or (_19103_, _19102_, _19101_);
  and (_19104_, _19103_, _04082_);
  and (_19105_, _05278_, \oc8051_golden_model_1.ACC [6]);
  nor (_19106_, _19105_, _19101_);
  nor (_19107_, _19106_, _04437_);
  nor (_19108_, _04436_, _19099_);
  or (_19109_, _19108_, _19107_);
  and (_19110_, _19109_, _04432_);
  nor (_19112_, _13293_, _09097_);
  nor (_19113_, _19112_, _19101_);
  nor (_19114_, _19113_, _04432_);
  or (_19115_, _19114_, _19110_);
  and (_19116_, _19115_, _03470_);
  nor (_19117_, _05944_, _19099_);
  and (_19118_, _13280_, _05944_);
  nor (_19119_, _19118_, _19117_);
  nor (_19120_, _19119_, _03470_);
  or (_19121_, _19120_, _03527_);
  or (_19123_, _19121_, _19116_);
  nor (_19124_, _05417_, _09097_);
  nor (_19125_, _19124_, _19101_);
  nand (_19126_, _19125_, _03527_);
  and (_19127_, _19126_, _19123_);
  and (_19128_, _19127_, _03531_);
  nor (_19129_, _19106_, _03531_);
  or (_19130_, _19129_, _19128_);
  and (_19131_, _19130_, _03466_);
  and (_19132_, _13304_, _05944_);
  nor (_19134_, _19132_, _19117_);
  nor (_19135_, _19134_, _03466_);
  or (_19136_, _19135_, _19131_);
  and (_19137_, _19136_, _03459_);
  nor (_19138_, _19117_, _13311_);
  nor (_19139_, _19138_, _19119_);
  and (_19140_, _19139_, _03458_);
  or (_19141_, _19140_, _19137_);
  and (_19142_, _19141_, _03453_);
  nor (_19143_, _13329_, _09134_);
  nor (_19145_, _19143_, _19117_);
  nor (_19146_, _19145_, _03453_);
  nor (_19147_, _19146_, _07454_);
  not (_19148_, _19147_);
  nor (_19149_, _19148_, _19142_);
  and (_19150_, _19125_, _07454_);
  or (_19151_, _19150_, _04082_);
  nor (_19152_, _19151_, _19149_);
  or (_19153_, _19152_, _19104_);
  and (_19154_, _19153_, _03521_);
  nor (_19156_, _13387_, _09097_);
  nor (_19157_, _19156_, _19101_);
  nor (_19158_, _19157_, _03521_);
  or (_19159_, _19158_, _08905_);
  or (_19160_, _19159_, _19154_);
  and (_19161_, _13402_, _05278_);
  or (_19162_, _19101_, _04527_);
  or (_19163_, _19162_, _19161_);
  and (_19164_, _14949_, _05278_);
  nor (_19165_, _19164_, _19101_);
  and (_19167_, _19165_, _03624_);
  nor (_19168_, _19167_, _03744_);
  and (_19169_, _19168_, _19163_);
  and (_19170_, _19169_, _19160_);
  and (_19171_, _13407_, _05278_);
  nor (_19172_, _19171_, _19101_);
  nor (_19173_, _19172_, _03745_);
  nor (_19174_, _19173_, _19170_);
  nor (_19175_, _19174_, _03611_);
  nor (_19176_, _19101_, _05469_);
  not (_19178_, _19176_);
  nor (_19179_, _19165_, _04523_);
  and (_19180_, _19179_, _19178_);
  nor (_19181_, _19180_, _19175_);
  nor (_19182_, _19181_, _03733_);
  nor (_19183_, _19106_, _03734_);
  and (_19184_, _19183_, _19178_);
  nor (_19185_, _19184_, _03618_);
  not (_19186_, _19185_);
  nor (_19187_, _19186_, _19182_);
  nor (_19189_, _13400_, _09097_);
  or (_19190_, _19101_, _06453_);
  nor (_19191_, _19190_, _19189_);
  or (_19192_, _19191_, _03741_);
  nor (_19193_, _19192_, _19187_);
  nor (_19194_, _13406_, _09097_);
  nor (_19195_, _19194_, _19101_);
  nor (_19196_, _19195_, _06458_);
  or (_19197_, _19196_, _19193_);
  and (_19198_, _19197_, _03948_);
  nor (_19200_, _19113_, _03948_);
  or (_19201_, _19200_, _19198_);
  and (_19202_, _19201_, _03446_);
  nor (_19203_, _19134_, _03446_);
  or (_19204_, _19203_, _19202_);
  and (_19205_, _19204_, _03474_);
  and (_19206_, _13456_, _05278_);
  nor (_19207_, _19206_, _19101_);
  nor (_19208_, _19207_, _03474_);
  or (_19209_, _19208_, _19205_);
  or (_19211_, _19209_, _43193_);
  or (_19212_, _43189_, \oc8051_golden_model_1.IE [6]);
  and (_19213_, _19212_, _42003_);
  and (_43775_, _19213_, _19211_);
  not (_19214_, \oc8051_golden_model_1.IP [0]);
  nor (_19215_, _05309_, _19214_);
  nor (_19216_, _05722_, _09204_);
  nor (_19217_, _19216_, _19215_);
  and (_19218_, _19217_, _03473_);
  and (_19219_, _12183_, _05309_);
  nor (_19221_, _19219_, _19215_);
  nor (_19222_, _19221_, _03745_);
  and (_19223_, _05309_, _06350_);
  nor (_19224_, _19223_, _19215_);
  and (_19225_, _19224_, _03624_);
  and (_19226_, _05309_, _04429_);
  nor (_19227_, _19226_, _19215_);
  and (_19228_, _19227_, _07454_);
  and (_19229_, _05309_, \oc8051_golden_model_1.ACC [0]);
  nor (_19230_, _19229_, _19215_);
  nor (_19232_, _19230_, _04437_);
  nor (_19233_, _04436_, _19214_);
  or (_19234_, _19233_, _19232_);
  and (_19235_, _19234_, _04432_);
  nor (_19236_, _19217_, _04432_);
  or (_19237_, _19236_, _19235_);
  and (_19238_, _19237_, _03470_);
  nor (_19239_, _05935_, _19214_);
  and (_19240_, _12075_, _05935_);
  nor (_19241_, _19240_, _19239_);
  nor (_19243_, _19241_, _03470_);
  nor (_19244_, _19243_, _19238_);
  nor (_19245_, _19244_, _03527_);
  nor (_19246_, _19227_, _04457_);
  or (_19247_, _19246_, _19245_);
  and (_19248_, _19247_, _03531_);
  nor (_19249_, _19230_, _03531_);
  or (_19250_, _19249_, _19248_);
  and (_19251_, _19250_, _03466_);
  and (_19252_, _19215_, _03465_);
  or (_19254_, _19252_, _19251_);
  and (_19255_, _19254_, _03459_);
  nor (_19256_, _19217_, _03459_);
  or (_19257_, _19256_, _19255_);
  and (_19258_, _19257_, _03453_);
  nor (_19259_, _12106_, _09241_);
  nor (_19260_, _19259_, _19239_);
  nor (_19261_, _19260_, _03453_);
  or (_19262_, _19261_, _07454_);
  nor (_19263_, _19262_, _19258_);
  nor (_19265_, _19263_, _19228_);
  nor (_19266_, _19265_, _04082_);
  and (_19267_, _06617_, _05309_);
  nor (_19268_, _19215_, _04500_);
  not (_19269_, _19268_);
  nor (_19270_, _19269_, _19267_);
  or (_19271_, _19270_, _03224_);
  nor (_19272_, _19271_, _19266_);
  nor (_19273_, _12164_, _09204_);
  nor (_19274_, _19273_, _19215_);
  nor (_19276_, _19274_, _03521_);
  or (_19277_, _19276_, _03624_);
  nor (_19278_, _19277_, _19272_);
  nor (_19279_, _19278_, _19225_);
  or (_19280_, _19279_, _03623_);
  and (_19281_, _12177_, _05309_);
  or (_19282_, _19281_, _19215_);
  or (_19283_, _19282_, _04527_);
  and (_19284_, _19283_, _03745_);
  and (_19285_, _19284_, _19280_);
  nor (_19287_, _19285_, _19222_);
  nor (_19288_, _19287_, _03611_);
  or (_19289_, _19224_, _04523_);
  nor (_19290_, _19289_, _19216_);
  nor (_19291_, _19290_, _19288_);
  nor (_19292_, _19291_, _03733_);
  and (_19293_, _12182_, _05309_);
  or (_19294_, _19293_, _19215_);
  and (_19295_, _19294_, _03733_);
  or (_19296_, _19295_, _19292_);
  and (_19298_, _19296_, _06453_);
  nor (_19299_, _12057_, _09204_);
  nor (_19300_, _19299_, _19215_);
  nor (_19301_, _19300_, _06453_);
  or (_19302_, _19301_, _19298_);
  and (_19303_, _19302_, _06458_);
  nor (_19304_, _12181_, _09204_);
  nor (_19305_, _19304_, _19215_);
  nor (_19306_, _19305_, _06458_);
  or (_19307_, _19306_, _19303_);
  and (_19309_, _19307_, _03948_);
  nor (_19310_, _19217_, _03948_);
  or (_19311_, _19310_, _19309_);
  and (_19312_, _19311_, _03446_);
  and (_19313_, _19215_, _03445_);
  nor (_19314_, _19313_, _03473_);
  not (_19315_, _19314_);
  nor (_19316_, _19315_, _19312_);
  nor (_19317_, _19316_, _19218_);
  or (_19318_, _19317_, _43193_);
  or (_19320_, _43189_, \oc8051_golden_model_1.IP [0]);
  and (_19321_, _19320_, _42003_);
  and (_43776_, _19321_, _19318_);
  not (_19322_, \oc8051_golden_model_1.IP [1]);
  nor (_19323_, _05309_, _19322_);
  and (_19324_, _06572_, _05309_);
  or (_19325_, _19324_, _19323_);
  and (_19326_, _19325_, _04082_);
  nor (_19327_, _05309_, \oc8051_golden_model_1.IP [1]);
  and (_19328_, _05309_, _03269_);
  nor (_19330_, _19328_, _19327_);
  and (_19331_, _19330_, _04436_);
  nor (_19332_, _04436_, _19322_);
  or (_19333_, _19332_, _19331_);
  and (_19334_, _19333_, _04432_);
  and (_19335_, _12265_, _05309_);
  nor (_19336_, _19335_, _19327_);
  and (_19337_, _19336_, _03534_);
  or (_19338_, _19337_, _19334_);
  and (_19339_, _19338_, _03470_);
  and (_19341_, _12269_, _05935_);
  nor (_19342_, _05935_, _19322_);
  or (_19343_, _19342_, _03527_);
  or (_19344_, _19343_, _19341_);
  and (_19345_, _19344_, _03533_);
  nor (_19346_, _19345_, _19339_);
  nor (_19347_, _09204_, _04635_);
  nor (_19348_, _19347_, _19323_);
  and (_19349_, _19348_, _03527_);
  nor (_19350_, _19349_, _19346_);
  and (_19352_, _19350_, _03531_);
  and (_19353_, _19330_, _03530_);
  or (_19354_, _19353_, _19352_);
  and (_19355_, _19354_, _03466_);
  and (_19356_, _12256_, _05935_);
  nor (_19357_, _19356_, _19342_);
  nor (_19358_, _19357_, _03466_);
  or (_19359_, _19358_, _19355_);
  and (_19360_, _19359_, _03459_);
  and (_19361_, _19341_, _12284_);
  or (_19363_, _19361_, _19342_);
  and (_19364_, _19363_, _03458_);
  or (_19365_, _19364_, _19360_);
  and (_19366_, _19365_, _03453_);
  nor (_19367_, _12301_, _09241_);
  nor (_19368_, _19342_, _19367_);
  nor (_19369_, _19368_, _03453_);
  or (_19370_, _19369_, _07454_);
  nor (_19371_, _19370_, _19366_);
  and (_19372_, _19348_, _07454_);
  or (_19374_, _19372_, _04082_);
  nor (_19375_, _19374_, _19371_);
  or (_19376_, _19375_, _19326_);
  and (_19377_, _19376_, _03521_);
  nor (_19378_, _12360_, _09204_);
  nor (_19379_, _19378_, _19323_);
  nor (_19380_, _19379_, _03521_);
  nor (_19381_, _19380_, _19377_);
  nor (_19382_, _19381_, _08905_);
  nor (_19383_, _12375_, _09204_);
  nor (_19385_, _19383_, _04527_);
  and (_19386_, _05309_, _04325_);
  nor (_19387_, _19386_, _04509_);
  nor (_19388_, _19387_, _19385_);
  nor (_19389_, _19388_, _19327_);
  nor (_19390_, _19389_, _19382_);
  nor (_19391_, _19390_, _03744_);
  not (_19392_, _19327_);
  nor (_19393_, _12381_, _09204_);
  nor (_19394_, _19393_, _03745_);
  and (_19396_, _19394_, _19392_);
  nor (_19397_, _19396_, _19391_);
  nor (_19398_, _19397_, _03611_);
  nor (_19399_, _12374_, _09204_);
  nor (_19400_, _19399_, _04523_);
  and (_19401_, _19400_, _19392_);
  nor (_19402_, _19401_, _19398_);
  nor (_19403_, _19402_, _03733_);
  nor (_19404_, _19323_, _05674_);
  nor (_19405_, _19404_, _03734_);
  and (_19407_, _19405_, _19330_);
  nor (_19408_, _19407_, _19403_);
  or (_19409_, _19408_, _18526_);
  and (_19410_, _19386_, _05673_);
  or (_19411_, _19327_, _06453_);
  or (_19412_, _19411_, _19410_);
  and (_19413_, _19328_, _05673_);
  or (_19414_, _19327_, _06458_);
  or (_19415_, _19414_, _19413_);
  and (_19416_, _19415_, _03948_);
  and (_19418_, _19416_, _19412_);
  and (_19419_, _19418_, _19409_);
  nor (_19420_, _19336_, _03948_);
  or (_19421_, _19420_, _03445_);
  nor (_19422_, _19421_, _19419_);
  nor (_19423_, _19357_, _03446_);
  or (_19424_, _19423_, _03473_);
  nor (_19425_, _19424_, _19422_);
  or (_19426_, _19323_, _03474_);
  nor (_19427_, _19426_, _19335_);
  nor (_19429_, _19427_, _19425_);
  or (_19430_, _19429_, _43193_);
  or (_19431_, _43189_, \oc8051_golden_model_1.IP [1]);
  and (_19432_, _19431_, _42003_);
  and (_43777_, _19432_, _19430_);
  not (_19433_, \oc8051_golden_model_1.IP [2]);
  nor (_19434_, _05309_, _19433_);
  and (_19435_, _05309_, _06399_);
  nor (_19436_, _19435_, _19434_);
  and (_19437_, _19436_, _03624_);
  nor (_19439_, _09204_, _05073_);
  nor (_19440_, _19439_, _19434_);
  and (_19441_, _19440_, _07454_);
  and (_19442_, _05309_, \oc8051_golden_model_1.ACC [2]);
  nor (_19443_, _19442_, _19434_);
  nor (_19444_, _19443_, _04437_);
  nor (_19445_, _04436_, _19433_);
  or (_19446_, _19445_, _19444_);
  and (_19447_, _19446_, _04432_);
  nor (_19448_, _12467_, _09204_);
  nor (_19450_, _19448_, _19434_);
  nor (_19451_, _19450_, _04432_);
  or (_19452_, _19451_, _19447_);
  and (_19453_, _19452_, _03470_);
  nor (_19454_, _05935_, _19433_);
  and (_19455_, _12462_, _05935_);
  nor (_19456_, _19455_, _19454_);
  nor (_19457_, _19456_, _03470_);
  or (_19458_, _19457_, _19453_);
  and (_19459_, _19458_, _04457_);
  nor (_19461_, _19440_, _04457_);
  or (_19462_, _19461_, _19459_);
  and (_19463_, _19462_, _03531_);
  nor (_19464_, _19443_, _03531_);
  or (_19465_, _19464_, _19463_);
  and (_19466_, _19465_, _03466_);
  and (_19467_, _12460_, _05935_);
  nor (_19468_, _19467_, _19454_);
  nor (_19469_, _19468_, _03466_);
  or (_19470_, _19469_, _03458_);
  or (_19472_, _19470_, _19466_);
  and (_19473_, _19455_, _12491_);
  or (_19474_, _19454_, _03459_);
  or (_19475_, _19474_, _19473_);
  and (_19476_, _19475_, _03453_);
  and (_19477_, _19476_, _19472_);
  nor (_19478_, _12509_, _09241_);
  nor (_19479_, _19478_, _19454_);
  nor (_19480_, _19479_, _03453_);
  nor (_19481_, _19480_, _07454_);
  not (_19483_, _19481_);
  nor (_19484_, _19483_, _19477_);
  nor (_19485_, _19484_, _19441_);
  nor (_19486_, _19485_, _04082_);
  and (_19487_, _06710_, _05309_);
  nor (_19488_, _19434_, _04500_);
  not (_19489_, _19488_);
  nor (_19490_, _19489_, _19487_);
  or (_19491_, _19490_, _03224_);
  nor (_19492_, _19491_, _19486_);
  nor (_19494_, _12568_, _09204_);
  nor (_19495_, _19434_, _19494_);
  nor (_19496_, _19495_, _03521_);
  or (_19497_, _19496_, _03624_);
  nor (_19498_, _19497_, _19492_);
  nor (_19499_, _19498_, _19437_);
  or (_19500_, _19499_, _03623_);
  and (_19501_, _12582_, _05309_);
  or (_19502_, _19501_, _19434_);
  or (_19503_, _19502_, _04527_);
  and (_19505_, _19503_, _03745_);
  and (_19506_, _19505_, _19500_);
  and (_19507_, _12588_, _05309_);
  nor (_19508_, _19507_, _19434_);
  nor (_19509_, _19508_, _03745_);
  nor (_19510_, _19509_, _19506_);
  nor (_19511_, _19510_, _03611_);
  nor (_19512_, _19434_, _05772_);
  not (_19513_, _19512_);
  nor (_19514_, _19436_, _04523_);
  and (_19516_, _19514_, _19513_);
  nor (_19517_, _19516_, _19511_);
  nor (_19518_, _19517_, _03733_);
  nor (_19519_, _19443_, _03734_);
  and (_19520_, _19519_, _19513_);
  nor (_19521_, _19520_, _03618_);
  not (_19522_, _19521_);
  nor (_19523_, _19522_, _19518_);
  nor (_19524_, _12581_, _09204_);
  or (_19525_, _19434_, _06453_);
  nor (_19527_, _19525_, _19524_);
  or (_19528_, _19527_, _03741_);
  nor (_19529_, _19528_, _19523_);
  nor (_19530_, _12587_, _09204_);
  nor (_19531_, _19530_, _19434_);
  nor (_19532_, _19531_, _06458_);
  or (_19533_, _19532_, _19529_);
  and (_19534_, _19533_, _03948_);
  nor (_19535_, _19450_, _03948_);
  or (_19536_, _19535_, _19534_);
  and (_19538_, _19536_, _03446_);
  nor (_19539_, _19468_, _03446_);
  or (_19540_, _19539_, _19538_);
  and (_19541_, _19540_, _03474_);
  and (_19542_, _12638_, _05309_);
  nor (_19543_, _19542_, _19434_);
  nor (_19544_, _19543_, _03474_);
  or (_19545_, _19544_, _19541_);
  or (_19546_, _19545_, _43193_);
  or (_19547_, _43189_, \oc8051_golden_model_1.IP [2]);
  and (_19549_, _19547_, _42003_);
  and (_43780_, _19549_, _19546_);
  not (_19550_, \oc8051_golden_model_1.IP [3]);
  nor (_19551_, _05309_, _19550_);
  and (_19552_, _05309_, _06356_);
  nor (_19553_, _19552_, _19551_);
  and (_19554_, _19553_, _03624_);
  nor (_19555_, _09204_, _04885_);
  nor (_19556_, _19555_, _19551_);
  and (_19557_, _19556_, _07454_);
  and (_19559_, _05309_, \oc8051_golden_model_1.ACC [3]);
  nor (_19560_, _19559_, _19551_);
  nor (_19561_, _19560_, _04437_);
  nor (_19562_, _04436_, _19550_);
  or (_19563_, _19562_, _19561_);
  and (_19564_, _19563_, _04432_);
  nor (_19565_, _12652_, _09204_);
  nor (_19566_, _19565_, _19551_);
  nor (_19567_, _19566_, _04432_);
  or (_19568_, _19567_, _19564_);
  and (_19570_, _19568_, _03470_);
  nor (_19571_, _05935_, _19550_);
  and (_19572_, _12664_, _05935_);
  nor (_19573_, _19572_, _19571_);
  nor (_19574_, _19573_, _03470_);
  or (_19575_, _19574_, _03527_);
  or (_19576_, _19575_, _19570_);
  nand (_19577_, _19556_, _03527_);
  and (_19578_, _19577_, _19576_);
  and (_19579_, _19578_, _03531_);
  nor (_19581_, _19560_, _03531_);
  or (_19582_, _19581_, _19579_);
  and (_19583_, _19582_, _03466_);
  and (_19584_, _12662_, _05935_);
  nor (_19585_, _19584_, _19571_);
  nor (_19586_, _19585_, _03466_);
  or (_19587_, _19586_, _19583_);
  and (_19588_, _19587_, _03459_);
  nor (_19589_, _19571_, _12691_);
  nor (_19590_, _19589_, _19573_);
  and (_19592_, _19590_, _03458_);
  or (_19593_, _19592_, _19588_);
  and (_19594_, _19593_, _03453_);
  nor (_19595_, _12709_, _09241_);
  nor (_19596_, _19595_, _19571_);
  nor (_19597_, _19596_, _03453_);
  nor (_19598_, _19597_, _07454_);
  not (_19599_, _19598_);
  nor (_19600_, _19599_, _19594_);
  nor (_19601_, _19600_, _19557_);
  nor (_19603_, _19601_, _04082_);
  and (_19604_, _06664_, _05309_);
  nor (_19605_, _19551_, _04500_);
  not (_19606_, _19605_);
  nor (_19607_, _19606_, _19604_);
  or (_19608_, _19607_, _03224_);
  nor (_19609_, _19608_, _19603_);
  nor (_19610_, _12773_, _09204_);
  nor (_19611_, _19551_, _19610_);
  nor (_19612_, _19611_, _03521_);
  or (_19614_, _19612_, _03624_);
  nor (_19615_, _19614_, _19609_);
  nor (_19616_, _19615_, _19554_);
  or (_19617_, _19616_, _03623_);
  and (_19618_, _12787_, _05309_);
  or (_19619_, _19618_, _19551_);
  or (_19620_, _19619_, _04527_);
  and (_19621_, _19620_, _03745_);
  and (_19622_, _19621_, _19617_);
  and (_19623_, _12793_, _05309_);
  nor (_19625_, _19623_, _19551_);
  nor (_19626_, _19625_, _03745_);
  nor (_19627_, _19626_, _19622_);
  nor (_19628_, _19627_, _03611_);
  nor (_19629_, _19551_, _05625_);
  not (_19630_, _19629_);
  nor (_19631_, _19553_, _04523_);
  and (_19632_, _19631_, _19630_);
  nor (_19633_, _19632_, _19628_);
  nor (_19634_, _19633_, _03733_);
  nor (_19636_, _19560_, _03734_);
  and (_19637_, _19636_, _19630_);
  nor (_19638_, _19637_, _03618_);
  not (_19639_, _19638_);
  nor (_19640_, _19639_, _19634_);
  nor (_19641_, _12786_, _09204_);
  or (_19642_, _19551_, _06453_);
  nor (_19643_, _19642_, _19641_);
  or (_19644_, _19643_, _03741_);
  nor (_19645_, _19644_, _19640_);
  nor (_19647_, _12792_, _09204_);
  nor (_19648_, _19647_, _19551_);
  nor (_19649_, _19648_, _06458_);
  or (_19650_, _19649_, _19645_);
  and (_19651_, _19650_, _03948_);
  nor (_19652_, _19566_, _03948_);
  or (_19653_, _19652_, _19651_);
  and (_19654_, _19653_, _03446_);
  nor (_19655_, _19585_, _03446_);
  or (_19656_, _19655_, _19654_);
  and (_19658_, _19656_, _03474_);
  and (_19659_, _12843_, _05309_);
  nor (_19660_, _19659_, _19551_);
  nor (_19661_, _19660_, _03474_);
  or (_19662_, _19661_, _19658_);
  or (_19663_, _19662_, _43193_);
  or (_19664_, _43189_, \oc8051_golden_model_1.IP [3]);
  and (_19665_, _19664_, _42003_);
  and (_43781_, _19665_, _19663_);
  not (_19666_, \oc8051_golden_model_1.IP [4]);
  nor (_19668_, _05309_, _19666_);
  nor (_19669_, _05831_, _09204_);
  nor (_19670_, _19669_, _19668_);
  and (_19671_, _19670_, _07454_);
  nor (_19672_, _05935_, _19666_);
  and (_19673_, _12864_, _05935_);
  nor (_19674_, _19673_, _19672_);
  nor (_19675_, _19674_, _03466_);
  and (_19676_, _05309_, \oc8051_golden_model_1.ACC [4]);
  nor (_19677_, _19676_, _19668_);
  nor (_19679_, _19677_, _04437_);
  nor (_19680_, _04436_, _19666_);
  or (_19681_, _19680_, _19679_);
  and (_19682_, _19681_, _04432_);
  nor (_19683_, _12856_, _09204_);
  nor (_19684_, _19683_, _19668_);
  nor (_19685_, _19684_, _04432_);
  or (_19686_, _19685_, _19682_);
  and (_19687_, _19686_, _03470_);
  and (_19688_, _12866_, _05935_);
  nor (_19690_, _19688_, _19672_);
  nor (_19691_, _19690_, _03470_);
  or (_19692_, _19691_, _03527_);
  or (_19693_, _19692_, _19687_);
  nand (_19694_, _19670_, _03527_);
  and (_19695_, _19694_, _19693_);
  and (_19696_, _19695_, _03531_);
  nor (_19697_, _19677_, _03531_);
  or (_19698_, _19697_, _19696_);
  and (_19699_, _19698_, _03466_);
  nor (_19701_, _19699_, _19675_);
  nor (_19702_, _19701_, _03458_);
  nor (_19703_, _19672_, _12894_);
  or (_19704_, _19690_, _03459_);
  nor (_19705_, _19704_, _19703_);
  nor (_19706_, _19705_, _19702_);
  nor (_19707_, _19706_, _03452_);
  nor (_19708_, _12912_, _09241_);
  nor (_19709_, _19708_, _19672_);
  nor (_19710_, _19709_, _03453_);
  nor (_19712_, _19710_, _07454_);
  not (_19713_, _19712_);
  nor (_19714_, _19713_, _19707_);
  nor (_19715_, _19714_, _19671_);
  nor (_19716_, _19715_, _04082_);
  and (_19717_, _06802_, _05309_);
  nor (_19718_, _19668_, _04500_);
  not (_19719_, _19718_);
  nor (_19720_, _19719_, _19717_);
  nor (_19721_, _19720_, _03224_);
  not (_19723_, _19721_);
  nor (_19724_, _19723_, _19716_);
  nor (_19725_, _12972_, _09204_);
  nor (_19726_, _19725_, _19668_);
  nor (_19727_, _19726_, _03521_);
  or (_19728_, _19727_, _08905_);
  or (_19729_, _19728_, _19724_);
  and (_19730_, _12986_, _05309_);
  or (_19731_, _19668_, _04527_);
  or (_19732_, _19731_, _19730_);
  and (_19734_, _06337_, _05309_);
  nor (_19735_, _19734_, _19668_);
  and (_19736_, _19735_, _03624_);
  nor (_19737_, _19736_, _03744_);
  and (_19738_, _19737_, _19732_);
  and (_19739_, _19738_, _19729_);
  and (_19740_, _12992_, _05309_);
  nor (_19741_, _19740_, _19668_);
  nor (_19742_, _19741_, _03745_);
  nor (_19743_, _19742_, _19739_);
  nor (_19745_, _19743_, _03611_);
  nor (_19746_, _19668_, _05880_);
  not (_19747_, _19746_);
  nor (_19748_, _19735_, _04523_);
  and (_19749_, _19748_, _19747_);
  nor (_19750_, _19749_, _19745_);
  nor (_19751_, _19750_, _03733_);
  nor (_19752_, _19677_, _03734_);
  and (_19753_, _19752_, _19747_);
  or (_19754_, _19753_, _19751_);
  and (_19756_, _19754_, _06453_);
  nor (_19757_, _12985_, _09204_);
  nor (_19758_, _19757_, _19668_);
  nor (_19759_, _19758_, _06453_);
  or (_19760_, _19759_, _19756_);
  and (_19761_, _19760_, _06458_);
  nor (_19762_, _12991_, _09204_);
  nor (_19763_, _19762_, _19668_);
  nor (_19764_, _19763_, _06458_);
  or (_19765_, _19764_, _19761_);
  and (_19767_, _19765_, _03948_);
  nor (_19768_, _19684_, _03948_);
  or (_19769_, _19768_, _19767_);
  and (_19770_, _19769_, _03446_);
  nor (_19771_, _19674_, _03446_);
  or (_19772_, _19771_, _19770_);
  and (_19773_, _19772_, _03474_);
  and (_19774_, _13051_, _05309_);
  nor (_19775_, _19774_, _19668_);
  nor (_19776_, _19775_, _03474_);
  or (_19778_, _19776_, _19773_);
  or (_19779_, _19778_, _43193_);
  or (_19780_, _43189_, \oc8051_golden_model_1.IP [4]);
  and (_19781_, _19780_, _42003_);
  and (_43782_, _19781_, _19779_);
  not (_19782_, \oc8051_golden_model_1.IP [5]);
  nor (_19783_, _05309_, _19782_);
  and (_19784_, _06757_, _05309_);
  or (_19785_, _19784_, _19783_);
  and (_19786_, _19785_, _04082_);
  and (_19788_, _05309_, \oc8051_golden_model_1.ACC [5]);
  nor (_19789_, _19788_, _19783_);
  nor (_19790_, _19789_, _04437_);
  nor (_19791_, _04436_, _19782_);
  or (_19792_, _19791_, _19790_);
  and (_19793_, _19792_, _04432_);
  nor (_19794_, _13070_, _09204_);
  nor (_19795_, _19794_, _19783_);
  nor (_19796_, _19795_, _04432_);
  or (_19797_, _19796_, _19793_);
  and (_19799_, _19797_, _03470_);
  nor (_19800_, _05935_, _19782_);
  and (_19801_, _13095_, _05935_);
  nor (_19802_, _19801_, _19800_);
  nor (_19803_, _19802_, _03470_);
  or (_19804_, _19803_, _03527_);
  or (_19805_, _19804_, _19799_);
  nor (_19806_, _05526_, _09204_);
  nor (_19807_, _19806_, _19783_);
  nand (_19808_, _19807_, _03527_);
  and (_19810_, _19808_, _19805_);
  and (_19811_, _19810_, _03531_);
  nor (_19812_, _19789_, _03531_);
  or (_19813_, _19812_, _19811_);
  and (_19814_, _19813_, _03466_);
  and (_19815_, _13078_, _05935_);
  nor (_19816_, _19815_, _19800_);
  nor (_19817_, _19816_, _03466_);
  or (_19818_, _19817_, _19814_);
  and (_19819_, _19818_, _03459_);
  nor (_19821_, _19800_, _13110_);
  nor (_19822_, _19821_, _19802_);
  and (_19823_, _19822_, _03458_);
  or (_19824_, _19823_, _19819_);
  and (_19825_, _19824_, _03453_);
  nor (_19826_, _13076_, _09241_);
  nor (_19827_, _19826_, _19800_);
  nor (_19828_, _19827_, _03453_);
  nor (_19829_, _19828_, _07454_);
  not (_19830_, _19829_);
  nor (_19832_, _19830_, _19825_);
  and (_19833_, _19807_, _07454_);
  or (_19834_, _19833_, _04082_);
  nor (_19835_, _19834_, _19832_);
  or (_19836_, _19835_, _19786_);
  and (_19837_, _19836_, _03521_);
  nor (_19838_, _13184_, _09204_);
  nor (_19839_, _19838_, _19783_);
  nor (_19840_, _19839_, _03521_);
  or (_19841_, _19840_, _08905_);
  or (_19843_, _19841_, _19837_);
  and (_19844_, _13198_, _05309_);
  or (_19845_, _19783_, _04527_);
  or (_19846_, _19845_, _19844_);
  and (_19847_, _06295_, _05309_);
  nor (_19848_, _19847_, _19783_);
  and (_19849_, _19848_, _03624_);
  nor (_19850_, _19849_, _03744_);
  and (_19851_, _19850_, _19846_);
  and (_19852_, _19851_, _19843_);
  and (_19854_, _13204_, _05309_);
  nor (_19855_, _19854_, _19783_);
  nor (_19856_, _19855_, _03745_);
  nor (_19857_, _19856_, _19852_);
  nor (_19858_, _19857_, _03611_);
  nor (_19859_, _19783_, _05576_);
  not (_19860_, _19859_);
  nor (_19861_, _19848_, _04523_);
  and (_19862_, _19861_, _19860_);
  nor (_19863_, _19862_, _19858_);
  nor (_19865_, _19863_, _03733_);
  nor (_19866_, _19789_, _03734_);
  and (_19867_, _19866_, _19860_);
  or (_19868_, _19867_, _19865_);
  and (_19869_, _19868_, _06453_);
  nor (_19870_, _13197_, _09204_);
  nor (_19871_, _19870_, _19783_);
  nor (_19872_, _19871_, _06453_);
  or (_19873_, _19872_, _19869_);
  and (_19874_, _19873_, _06458_);
  nor (_19876_, _13203_, _09204_);
  nor (_19877_, _19876_, _19783_);
  nor (_19878_, _19877_, _06458_);
  or (_19879_, _19878_, _19874_);
  and (_19880_, _19879_, _03948_);
  nor (_19881_, _19795_, _03948_);
  or (_19882_, _19881_, _19880_);
  and (_19883_, _19882_, _03446_);
  nor (_19884_, _19816_, _03446_);
  or (_19885_, _19884_, _19883_);
  and (_19887_, _19885_, _03474_);
  and (_19888_, _13253_, _05309_);
  nor (_19889_, _19888_, _19783_);
  nor (_19890_, _19889_, _03474_);
  or (_19891_, _19890_, _19887_);
  or (_19892_, _19891_, _43193_);
  or (_19893_, _43189_, \oc8051_golden_model_1.IP [5]);
  and (_19894_, _19893_, _42003_);
  and (_43783_, _19894_, _19892_);
  not (_19895_, \oc8051_golden_model_1.IP [6]);
  nor (_19897_, _05309_, _19895_);
  and (_19898_, _06526_, _05309_);
  or (_19899_, _19898_, _19897_);
  and (_19900_, _19899_, _04082_);
  and (_19901_, _05309_, \oc8051_golden_model_1.ACC [6]);
  nor (_19902_, _19901_, _19897_);
  nor (_19903_, _19902_, _04437_);
  nor (_19904_, _04436_, _19895_);
  or (_19905_, _19904_, _19903_);
  and (_19906_, _19905_, _04432_);
  nor (_19908_, _13293_, _09204_);
  nor (_19909_, _19908_, _19897_);
  nor (_19910_, _19909_, _04432_);
  or (_19911_, _19910_, _19906_);
  and (_19912_, _19911_, _03470_);
  nor (_19913_, _05935_, _19895_);
  and (_19914_, _13280_, _05935_);
  nor (_19915_, _19914_, _19913_);
  nor (_19916_, _19915_, _03470_);
  or (_19917_, _19916_, _03527_);
  or (_19919_, _19917_, _19912_);
  nor (_19920_, _05417_, _09204_);
  nor (_19921_, _19920_, _19897_);
  nand (_19922_, _19921_, _03527_);
  and (_19923_, _19922_, _19919_);
  and (_19924_, _19923_, _03531_);
  nor (_19925_, _19902_, _03531_);
  or (_19926_, _19925_, _19924_);
  and (_19927_, _19926_, _03466_);
  and (_19928_, _13304_, _05935_);
  nor (_19930_, _19928_, _19913_);
  nor (_19931_, _19930_, _03466_);
  or (_19932_, _19931_, _03458_);
  or (_19933_, _19932_, _19927_);
  nor (_19934_, _19913_, _13311_);
  nor (_19935_, _19934_, _19915_);
  or (_19936_, _19935_, _03459_);
  and (_19937_, _19936_, _03453_);
  and (_19938_, _19937_, _19933_);
  nor (_19939_, _13329_, _09241_);
  nor (_19941_, _19939_, _19913_);
  nor (_19942_, _19941_, _03453_);
  nor (_19943_, _19942_, _07454_);
  not (_19944_, _19943_);
  nor (_19945_, _19944_, _19938_);
  and (_19946_, _19921_, _07454_);
  or (_19947_, _19946_, _04082_);
  nor (_19948_, _19947_, _19945_);
  or (_19949_, _19948_, _19900_);
  and (_19950_, _19949_, _03521_);
  nor (_19952_, _13387_, _09204_);
  nor (_19953_, _19952_, _19897_);
  nor (_19954_, _19953_, _03521_);
  or (_19955_, _19954_, _08905_);
  or (_19956_, _19955_, _19950_);
  and (_19957_, _13402_, _05309_);
  or (_19958_, _19897_, _04527_);
  or (_19959_, _19958_, _19957_);
  and (_19960_, _14949_, _05309_);
  nor (_19961_, _19960_, _19897_);
  and (_19963_, _19961_, _03624_);
  nor (_19964_, _19963_, _03744_);
  and (_19965_, _19964_, _19959_);
  and (_19966_, _19965_, _19956_);
  and (_19967_, _13407_, _05309_);
  nor (_19968_, _19967_, _19897_);
  nor (_19969_, _19968_, _03745_);
  nor (_19970_, _19969_, _19966_);
  nor (_19971_, _19970_, _03611_);
  nor (_19972_, _19897_, _05469_);
  not (_19974_, _19972_);
  nor (_19975_, _19961_, _04523_);
  and (_19976_, _19975_, _19974_);
  nor (_19977_, _19976_, _19971_);
  nor (_19978_, _19977_, _03733_);
  nor (_19979_, _19902_, _03734_);
  and (_19980_, _19979_, _19974_);
  or (_19981_, _19980_, _19978_);
  and (_19982_, _19981_, _06453_);
  nor (_19983_, _13400_, _09204_);
  nor (_19985_, _19983_, _19897_);
  nor (_19986_, _19985_, _06453_);
  or (_19987_, _19986_, _19982_);
  and (_19988_, _19987_, _06458_);
  nor (_19989_, _13406_, _09204_);
  nor (_19990_, _19989_, _19897_);
  nor (_19991_, _19990_, _06458_);
  or (_19992_, _19991_, _19988_);
  and (_19993_, _19992_, _03948_);
  nor (_19994_, _19909_, _03948_);
  or (_19996_, _19994_, _19993_);
  and (_19997_, _19996_, _03446_);
  nor (_19998_, _19930_, _03446_);
  or (_19999_, _19998_, _19997_);
  and (_20000_, _19999_, _03474_);
  and (_20001_, _13456_, _05309_);
  nor (_20002_, _20001_, _19897_);
  nor (_20003_, _20002_, _03474_);
  or (_20004_, _20003_, _20000_);
  or (_20005_, _20004_, _43193_);
  or (_20007_, _43189_, \oc8051_golden_model_1.IP [6]);
  and (_20008_, _20007_, _42003_);
  and (_43784_, _20008_, _20005_);
  not (_20009_, \oc8051_golden_model_1.P0 [0]);
  nor (_20010_, _43189_, _20009_);
  or (_20011_, _20010_, rst);
  nor (_20012_, _05298_, _20009_);
  and (_20013_, _12183_, _05298_);
  or (_20014_, _20013_, _20012_);
  and (_20015_, _20014_, _03744_);
  and (_20017_, _05298_, _04429_);
  or (_20018_, _20017_, _20012_);
  or (_20019_, _20018_, _06903_);
  nor (_20020_, _05722_, _09311_);
  or (_20021_, _20020_, _20012_);
  or (_20022_, _20021_, _04432_);
  and (_20023_, _05298_, \oc8051_golden_model_1.ACC [0]);
  or (_20024_, _20023_, _20012_);
  and (_20025_, _20024_, _04436_);
  nor (_20026_, _04436_, _20009_);
  or (_20028_, _20026_, _03534_);
  or (_20029_, _20028_, _20025_);
  and (_20030_, _20029_, _03470_);
  and (_20031_, _20030_, _20022_);
  nor (_20032_, _05258_, _20009_);
  and (_20033_, _12075_, _05258_);
  or (_20034_, _20033_, _20032_);
  and (_20035_, _20034_, _03469_);
  or (_20036_, _20035_, _20031_);
  and (_20037_, _20036_, _04457_);
  and (_20039_, _20018_, _03527_);
  or (_20040_, _20039_, _03530_);
  or (_20041_, _20040_, _20037_);
  or (_20042_, _20024_, _03531_);
  and (_20043_, _20042_, _03466_);
  and (_20044_, _20043_, _20041_);
  and (_20045_, _20012_, _03465_);
  or (_20046_, _20045_, _03458_);
  or (_20047_, _20046_, _20044_);
  or (_20048_, _20021_, _03459_);
  and (_20050_, _20048_, _03453_);
  and (_20051_, _20050_, _20047_);
  or (_20052_, _12105_, _12063_);
  and (_20053_, _20052_, _05258_);
  or (_20054_, _20053_, _20032_);
  and (_20055_, _20054_, _03452_);
  or (_20056_, _20055_, _07454_);
  or (_20057_, _20056_, _20051_);
  and (_20058_, _20057_, _20019_);
  or (_20059_, _20058_, _04082_);
  and (_20061_, _06617_, _05298_);
  or (_20062_, _20012_, _04500_);
  or (_20063_, _20062_, _20061_);
  and (_20064_, _20063_, _03521_);
  and (_20065_, _20064_, _20059_);
  and (_20066_, _06329_, \oc8051_golden_model_1.P2 [0]);
  and (_20067_, _06334_, \oc8051_golden_model_1.P0 [0]);
  and (_20068_, _06340_, \oc8051_golden_model_1.P1 [0]);
  and (_20069_, _06344_, \oc8051_golden_model_1.P3 [0]);
  or (_20070_, _20069_, _20068_);
  or (_20072_, _20070_, _20067_);
  nor (_20073_, _20072_, _20066_);
  and (_20074_, _20073_, _12121_);
  and (_20075_, _20074_, _12145_);
  nand (_20076_, _20075_, _12161_);
  or (_20077_, _20076_, _12118_);
  and (_20078_, _20077_, _05298_);
  or (_20079_, _20078_, _20012_);
  and (_20080_, _20079_, _03224_);
  or (_20081_, _20080_, _20065_);
  or (_20083_, _20081_, _08905_);
  and (_20084_, _12177_, _05298_);
  or (_20085_, _20012_, _04527_);
  or (_20086_, _20085_, _20084_);
  and (_20087_, _05298_, _06350_);
  or (_20088_, _20087_, _20012_);
  or (_20089_, _20088_, _04509_);
  and (_20090_, _20089_, _03745_);
  and (_20091_, _20090_, _20086_);
  and (_20092_, _20091_, _20083_);
  or (_20094_, _20092_, _20015_);
  and (_20095_, _20094_, _04523_);
  nand (_20096_, _20088_, _03611_);
  nor (_20097_, _20096_, _20020_);
  or (_20098_, _20097_, _20095_);
  and (_20099_, _20098_, _03734_);
  or (_20100_, _20012_, _05722_);
  and (_20101_, _20024_, _03733_);
  and (_20102_, _20101_, _20100_);
  or (_20103_, _20102_, _03618_);
  or (_20105_, _20103_, _20099_);
  nor (_20106_, _12057_, _09311_);
  or (_20107_, _20012_, _06453_);
  or (_20108_, _20107_, _20106_);
  and (_20109_, _20108_, _06458_);
  and (_20110_, _20109_, _20105_);
  nor (_20111_, _12181_, _09311_);
  or (_20112_, _20111_, _20012_);
  and (_20113_, _20112_, _03741_);
  or (_20114_, _20113_, _03767_);
  or (_20116_, _20114_, _20110_);
  or (_20117_, _20021_, _03948_);
  and (_20118_, _20117_, _03446_);
  and (_20119_, _20118_, _20116_);
  and (_20120_, _20012_, _03445_);
  or (_20121_, _20120_, _03473_);
  or (_20122_, _20121_, _20119_);
  or (_20123_, _20021_, _03474_);
  and (_20124_, _20123_, _43189_);
  and (_20125_, _20124_, _20122_);
  or (_43787_, _20125_, _20011_);
  or (_20127_, _05298_, \oc8051_golden_model_1.P0 [1]);
  and (_20128_, _12265_, _05298_);
  not (_20129_, _20128_);
  and (_20130_, _20129_, _20127_);
  or (_20131_, _20130_, _04432_);
  nand (_20132_, _05298_, _03269_);
  and (_20133_, _20132_, _20127_);
  and (_20134_, _20133_, _04436_);
  and (_20135_, _04437_, \oc8051_golden_model_1.P0 [1]);
  or (_20137_, _20135_, _03534_);
  or (_20138_, _20137_, _20134_);
  and (_20139_, _20138_, _03470_);
  and (_20140_, _20139_, _20131_);
  and (_20141_, _12269_, _05258_);
  not (_20142_, _05258_);
  and (_20143_, _20142_, \oc8051_golden_model_1.P0 [1]);
  or (_20144_, _20143_, _03527_);
  or (_20145_, _20144_, _20141_);
  and (_20146_, _20145_, _03533_);
  or (_20148_, _20146_, _20140_);
  and (_20149_, _09311_, \oc8051_golden_model_1.P0 [1]);
  nor (_20150_, _09311_, _04635_);
  or (_20151_, _20150_, _20149_);
  or (_20152_, _20151_, _04457_);
  and (_20153_, _20152_, _20148_);
  or (_20154_, _20153_, _03530_);
  or (_20155_, _20133_, _03531_);
  and (_20156_, _20155_, _03466_);
  and (_20157_, _20156_, _20154_);
  and (_20159_, _12256_, _05258_);
  or (_20160_, _20159_, _20143_);
  and (_20161_, _20160_, _03465_);
  or (_20162_, _20161_, _03458_);
  or (_20163_, _20162_, _20157_);
  and (_20164_, _20141_, _12284_);
  or (_20165_, _20143_, _03459_);
  or (_20166_, _20165_, _20164_);
  and (_20167_, _20166_, _20163_);
  and (_20168_, _20167_, _03453_);
  or (_20170_, _12300_, _12256_);
  and (_20171_, _20170_, _05258_);
  or (_20172_, _20143_, _20171_);
  and (_20173_, _20172_, _03452_);
  or (_20174_, _20173_, _07454_);
  or (_20175_, _20174_, _20168_);
  or (_20176_, _20151_, _06903_);
  and (_20177_, _20176_, _20175_);
  or (_20178_, _20177_, _04082_);
  and (_20179_, _06572_, _05298_);
  or (_20181_, _20149_, _04500_);
  or (_20182_, _20181_, _20179_);
  and (_20183_, _20182_, _03521_);
  and (_20184_, _20183_, _20178_);
  and (_20185_, _06329_, \oc8051_golden_model_1.P2 [1]);
  and (_20186_, _06334_, \oc8051_golden_model_1.P0 [1]);
  and (_20187_, _06340_, \oc8051_golden_model_1.P1 [1]);
  and (_20188_, _06344_, \oc8051_golden_model_1.P3 [1]);
  or (_20189_, _20188_, _20187_);
  or (_20190_, _20189_, _20186_);
  nor (_20192_, _20190_, _20185_);
  and (_20193_, _20192_, _12326_);
  and (_20194_, _20193_, _12341_);
  nand (_20195_, _20194_, _12357_);
  or (_20196_, _20195_, _12314_);
  and (_20197_, _20196_, _05298_);
  or (_20198_, _20197_, _20149_);
  and (_20199_, _20198_, _03224_);
  or (_20200_, _20199_, _20184_);
  and (_20201_, _20200_, _03625_);
  or (_20203_, _12375_, _09311_);
  and (_20204_, _20203_, _03623_);
  nand (_20205_, _05298_, _04325_);
  and (_20206_, _20205_, _03624_);
  or (_20207_, _20206_, _20204_);
  and (_20208_, _20207_, _20127_);
  or (_20209_, _20208_, _20201_);
  and (_20210_, _20209_, _03745_);
  or (_20211_, _12381_, _09311_);
  and (_20212_, _20127_, _03744_);
  and (_20214_, _20212_, _20211_);
  or (_20215_, _20214_, _20210_);
  and (_20216_, _20215_, _04523_);
  or (_20217_, _12374_, _09311_);
  and (_20218_, _20127_, _03611_);
  and (_20219_, _20218_, _20217_);
  or (_20220_, _20219_, _20216_);
  and (_20221_, _20220_, _03734_);
  or (_20222_, _20149_, _05674_);
  and (_20223_, _20133_, _03733_);
  and (_20225_, _20223_, _20222_);
  or (_20226_, _20225_, _20221_);
  and (_20227_, _20226_, _03742_);
  or (_20228_, _20205_, _05674_);
  and (_20229_, _20127_, _03618_);
  and (_20230_, _20229_, _20228_);
  or (_20231_, _20132_, _05674_);
  and (_20232_, _20127_, _03741_);
  and (_20233_, _20232_, _20231_);
  or (_20234_, _20233_, _03767_);
  or (_20236_, _20234_, _20230_);
  or (_20237_, _20236_, _20227_);
  or (_20238_, _20130_, _03948_);
  and (_20239_, _20238_, _03446_);
  and (_20240_, _20239_, _20237_);
  and (_20241_, _20160_, _03445_);
  or (_20242_, _20241_, _03473_);
  or (_20243_, _20242_, _20240_);
  or (_20244_, _20149_, _03474_);
  or (_20245_, _20244_, _20128_);
  and (_20247_, _20245_, _43189_);
  and (_20248_, _20247_, _20243_);
  nor (_20249_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_20250_, _20249_, _05173_);
  or (_43788_, _20250_, _20248_);
  not (_20251_, \oc8051_golden_model_1.P0 [2]);
  nor (_20252_, _05298_, _20251_);
  nor (_20253_, _09311_, _05073_);
  or (_20254_, _20253_, _20252_);
  or (_20255_, _20254_, _06903_);
  and (_20257_, _20254_, _03527_);
  nor (_20258_, _05258_, _20251_);
  and (_20259_, _12462_, _05258_);
  or (_20260_, _20259_, _20258_);
  or (_20261_, _20260_, _03470_);
  nor (_20262_, _12467_, _09311_);
  or (_20263_, _20262_, _20252_);
  and (_20264_, _20263_, _03534_);
  nor (_20265_, _04436_, _20251_);
  and (_20266_, _05298_, \oc8051_golden_model_1.ACC [2]);
  or (_20268_, _20266_, _20252_);
  and (_20269_, _20268_, _04436_);
  or (_20270_, _20269_, _20265_);
  and (_20271_, _20270_, _04432_);
  or (_20272_, _20271_, _03469_);
  or (_20273_, _20272_, _20264_);
  and (_20274_, _20273_, _20261_);
  and (_20275_, _20274_, _04457_);
  or (_20276_, _20275_, _20257_);
  or (_20277_, _20276_, _03530_);
  or (_20279_, _20268_, _03531_);
  and (_20280_, _20279_, _03466_);
  and (_20281_, _20280_, _20277_);
  and (_20282_, _12460_, _05258_);
  or (_20283_, _20282_, _20258_);
  and (_20284_, _20283_, _03465_);
  or (_20285_, _20284_, _03458_);
  or (_20286_, _20285_, _20281_);
  or (_20287_, _20258_, _12491_);
  and (_20288_, _20287_, _20260_);
  or (_20290_, _20288_, _03459_);
  and (_20291_, _20290_, _03453_);
  and (_20292_, _20291_, _20286_);
  or (_20293_, _12508_, _12460_);
  and (_20294_, _20293_, _05258_);
  or (_20295_, _20294_, _20258_);
  and (_20296_, _20295_, _03452_);
  or (_20297_, _20296_, _07454_);
  or (_20298_, _20297_, _20292_);
  and (_20299_, _20298_, _20255_);
  or (_20301_, _20299_, _04082_);
  and (_20302_, _06710_, _05298_);
  or (_20303_, _20252_, _04500_);
  or (_20304_, _20303_, _20302_);
  and (_20305_, _20304_, _03521_);
  and (_20306_, _20305_, _20301_);
  and (_20307_, _06329_, \oc8051_golden_model_1.P2 [2]);
  and (_20308_, _06334_, \oc8051_golden_model_1.P0 [2]);
  and (_20309_, _06340_, \oc8051_golden_model_1.P1 [2]);
  and (_20310_, _06344_, \oc8051_golden_model_1.P3 [2]);
  or (_20312_, _20310_, _20309_);
  or (_20313_, _20312_, _20308_);
  nor (_20314_, _20313_, _20307_);
  and (_20315_, _20314_, _12534_);
  and (_20316_, _20315_, _12545_);
  nand (_20317_, _20316_, _12565_);
  or (_20318_, _20317_, _12522_);
  and (_20319_, _20318_, _05298_);
  or (_20320_, _20252_, _20319_);
  and (_20321_, _20320_, _03224_);
  or (_20323_, _20321_, _20306_);
  or (_20324_, _20323_, _08905_);
  and (_20325_, _12582_, _05298_);
  or (_20326_, _20252_, _04527_);
  or (_20327_, _20326_, _20325_);
  and (_20328_, _05298_, _06399_);
  or (_20329_, _20328_, _20252_);
  or (_20330_, _20329_, _04509_);
  and (_20331_, _20330_, _03745_);
  and (_20332_, _20331_, _20327_);
  and (_20334_, _20332_, _20324_);
  and (_20335_, _12588_, _05298_);
  or (_20336_, _20335_, _20252_);
  and (_20337_, _20336_, _03744_);
  or (_20338_, _20337_, _20334_);
  and (_20339_, _20338_, _04523_);
  or (_20340_, _20252_, _05772_);
  and (_20341_, _20329_, _03611_);
  and (_20342_, _20341_, _20340_);
  or (_20343_, _20342_, _20339_);
  and (_20345_, _20343_, _03734_);
  and (_20346_, _20268_, _03733_);
  and (_20347_, _20346_, _20340_);
  or (_20348_, _20347_, _03618_);
  or (_20349_, _20348_, _20345_);
  nor (_20350_, _12581_, _09311_);
  or (_20351_, _20252_, _06453_);
  or (_20352_, _20351_, _20350_);
  and (_20353_, _20352_, _06458_);
  and (_20354_, _20353_, _20349_);
  nor (_20356_, _12587_, _09311_);
  or (_20357_, _20356_, _20252_);
  and (_20358_, _20357_, _03741_);
  or (_20359_, _20358_, _03767_);
  or (_20360_, _20359_, _20354_);
  or (_20361_, _20263_, _03948_);
  and (_20362_, _20361_, _03446_);
  and (_20363_, _20362_, _20360_);
  and (_20364_, _20283_, _03445_);
  or (_20365_, _20364_, _03473_);
  or (_20367_, _20365_, _20363_);
  and (_20368_, _12638_, _05298_);
  or (_20369_, _20252_, _03474_);
  or (_20370_, _20369_, _20368_);
  and (_20371_, _20370_, _43189_);
  and (_20372_, _20371_, _20367_);
  nor (_20373_, _43189_, _20251_);
  or (_20374_, _20373_, rst);
  or (_43789_, _20374_, _20372_);
  not (_20375_, \oc8051_golden_model_1.P0 [3]);
  nor (_20377_, _43189_, _20375_);
  or (_20378_, _20377_, rst);
  nor (_20379_, _05298_, _20375_);
  nor (_20380_, _09311_, _04885_);
  or (_20381_, _20380_, _20379_);
  or (_20382_, _20381_, _06903_);
  nor (_20383_, _12652_, _09311_);
  or (_20384_, _20383_, _20379_);
  or (_20385_, _20384_, _04432_);
  and (_20386_, _05298_, \oc8051_golden_model_1.ACC [3]);
  or (_20388_, _20386_, _20379_);
  and (_20389_, _20388_, _04436_);
  nor (_20390_, _04436_, _20375_);
  or (_20391_, _20390_, _03534_);
  or (_20392_, _20391_, _20389_);
  and (_20393_, _20392_, _03470_);
  and (_20394_, _20393_, _20385_);
  nor (_20395_, _05258_, _20375_);
  and (_20396_, _12664_, _05258_);
  or (_20397_, _20396_, _20395_);
  and (_20399_, _20397_, _03469_);
  or (_20400_, _20399_, _03527_);
  or (_20401_, _20400_, _20394_);
  or (_20402_, _20381_, _04457_);
  and (_20403_, _20402_, _20401_);
  or (_20404_, _20403_, _03530_);
  or (_20405_, _20388_, _03531_);
  and (_20406_, _20405_, _03466_);
  and (_20407_, _20406_, _20404_);
  and (_20408_, _12662_, _05258_);
  or (_20410_, _20408_, _20395_);
  and (_20411_, _20410_, _03465_);
  or (_20412_, _20411_, _03458_);
  or (_20413_, _20412_, _20407_);
  or (_20414_, _20395_, _12691_);
  and (_20415_, _20414_, _20397_);
  or (_20416_, _20415_, _03459_);
  and (_20417_, _20416_, _03453_);
  and (_20418_, _20417_, _20413_);
  or (_20419_, _12662_, _12707_);
  and (_20421_, _20419_, _05258_);
  or (_20422_, _20421_, _20395_);
  and (_20423_, _20422_, _03452_);
  or (_20424_, _20423_, _07454_);
  or (_20425_, _20424_, _20418_);
  and (_20426_, _20425_, _20382_);
  or (_20427_, _20426_, _04082_);
  and (_20428_, _06664_, _05298_);
  or (_20429_, _20379_, _04500_);
  or (_20430_, _20429_, _20428_);
  and (_20432_, _20430_, _03521_);
  and (_20433_, _20432_, _20427_);
  and (_20434_, _06340_, \oc8051_golden_model_1.P1 [3]);
  and (_20435_, _06329_, \oc8051_golden_model_1.P2 [3]);
  and (_20436_, _06334_, \oc8051_golden_model_1.P0 [3]);
  or (_20437_, _20436_, _20435_);
  nor (_20438_, _20437_, _20434_);
  nand (_20439_, _20438_, _12735_);
  not (_20440_, _12765_);
  and (_20441_, _12757_, _20440_);
  nand (_20443_, _20441_, _12748_);
  or (_20444_, _12736_, _12738_);
  and (_20445_, _06344_, \oc8051_golden_model_1.P3 [3]);
  or (_20446_, _20445_, _12762_);
  or (_20447_, _20446_, _20444_);
  nor (_20448_, _12766_, _12763_);
  nand (_20449_, _20448_, _12760_);
  or (_20450_, _20449_, _20447_);
  or (_20451_, _20450_, _20443_);
  or (_20452_, _20451_, _20439_);
  or (_20454_, _20452_, _12722_);
  and (_20455_, _20454_, _05298_);
  or (_20456_, _20379_, _20455_);
  and (_20457_, _20456_, _03224_);
  or (_20458_, _20457_, _20433_);
  or (_20459_, _20458_, _08905_);
  and (_20460_, _12787_, _05298_);
  or (_20461_, _20379_, _04527_);
  or (_20462_, _20461_, _20460_);
  and (_20463_, _05298_, _06356_);
  or (_20465_, _20463_, _20379_);
  or (_20466_, _20465_, _04509_);
  and (_20467_, _20466_, _03745_);
  and (_20468_, _20467_, _20462_);
  and (_20469_, _20468_, _20459_);
  and (_20470_, _12793_, _05298_);
  or (_20471_, _20470_, _20379_);
  and (_20472_, _20471_, _03744_);
  or (_20473_, _20472_, _20469_);
  and (_20474_, _20473_, _04523_);
  or (_20476_, _20379_, _05625_);
  and (_20477_, _20465_, _03611_);
  and (_20478_, _20477_, _20476_);
  or (_20479_, _20478_, _20474_);
  and (_20480_, _20479_, _03734_);
  and (_20481_, _20388_, _03733_);
  and (_20482_, _20481_, _20476_);
  or (_20483_, _20482_, _03618_);
  or (_20484_, _20483_, _20480_);
  nor (_20485_, _12786_, _09311_);
  or (_20487_, _20379_, _06453_);
  or (_20488_, _20487_, _20485_);
  and (_20489_, _20488_, _06458_);
  and (_20490_, _20489_, _20484_);
  nor (_20491_, _12792_, _09311_);
  or (_20492_, _20491_, _20379_);
  and (_20493_, _20492_, _03741_);
  or (_20494_, _20493_, _03767_);
  or (_20495_, _20494_, _20490_);
  or (_20496_, _20384_, _03948_);
  and (_20498_, _20496_, _03446_);
  and (_20499_, _20498_, _20495_);
  and (_20500_, _20410_, _03445_);
  or (_20501_, _20500_, _03473_);
  or (_20502_, _20501_, _20499_);
  and (_20503_, _12843_, _05298_);
  or (_20504_, _20379_, _03474_);
  or (_20505_, _20504_, _20503_);
  and (_20506_, _20505_, _43189_);
  and (_20507_, _20506_, _20502_);
  or (_43790_, _20507_, _20378_);
  and (_20509_, _09311_, \oc8051_golden_model_1.P0 [4]);
  nor (_20510_, _05831_, _09311_);
  or (_20511_, _20510_, _20509_);
  or (_20512_, _20511_, _06903_);
  and (_20513_, _20142_, \oc8051_golden_model_1.P0 [4]);
  and (_20514_, _12864_, _05258_);
  or (_20515_, _20514_, _20513_);
  and (_20516_, _20515_, _03465_);
  nor (_20517_, _12856_, _09311_);
  or (_20519_, _20517_, _20509_);
  or (_20520_, _20519_, _04432_);
  and (_20521_, _05298_, \oc8051_golden_model_1.ACC [4]);
  or (_20522_, _20521_, _20509_);
  and (_20523_, _20522_, _04436_);
  and (_20524_, _04437_, \oc8051_golden_model_1.P0 [4]);
  or (_20525_, _20524_, _03534_);
  or (_20526_, _20525_, _20523_);
  and (_20527_, _20526_, _03470_);
  and (_20528_, _20527_, _20520_);
  and (_20529_, _12866_, _05258_);
  or (_20530_, _20529_, _20513_);
  and (_20531_, _20530_, _03469_);
  or (_20532_, _20531_, _03527_);
  or (_20533_, _20532_, _20528_);
  or (_20534_, _20511_, _04457_);
  and (_20535_, _20534_, _20533_);
  or (_20536_, _20535_, _03530_);
  or (_20537_, _20522_, _03531_);
  and (_20538_, _20537_, _03466_);
  and (_20540_, _20538_, _20536_);
  or (_20541_, _20540_, _20516_);
  and (_20542_, _20541_, _03459_);
  and (_20543_, _12895_, _05258_);
  or (_20544_, _20543_, _20513_);
  and (_20545_, _20544_, _03458_);
  or (_20546_, _20545_, _20542_);
  and (_20547_, _20546_, _03453_);
  or (_20548_, _12911_, _12864_);
  and (_20549_, _20548_, _05258_);
  or (_20551_, _20549_, _20513_);
  and (_20552_, _20551_, _03452_);
  or (_20553_, _20552_, _07454_);
  or (_20554_, _20553_, _20547_);
  and (_20555_, _20554_, _20512_);
  or (_20556_, _20555_, _04082_);
  and (_20557_, _06802_, _05298_);
  or (_20558_, _20509_, _04500_);
  or (_20559_, _20558_, _20557_);
  and (_20560_, _20559_, _03521_);
  and (_20562_, _20560_, _20556_);
  and (_20563_, _06329_, \oc8051_golden_model_1.P2 [4]);
  and (_20564_, _06334_, \oc8051_golden_model_1.P0 [4]);
  and (_20565_, _06340_, \oc8051_golden_model_1.P1 [4]);
  and (_20566_, _06344_, \oc8051_golden_model_1.P3 [4]);
  or (_20567_, _20566_, _20565_);
  or (_20568_, _20567_, _20564_);
  nor (_20569_, _20568_, _20563_);
  and (_20570_, _20569_, _12937_);
  and (_20571_, _20570_, _12952_);
  nand (_20572_, _20571_, _12969_);
  or (_20573_, _20572_, _12925_);
  and (_20574_, _20573_, _05298_);
  or (_20575_, _20574_, _20509_);
  and (_20576_, _20575_, _03224_);
  or (_20577_, _20576_, _08905_);
  or (_20578_, _20577_, _20562_);
  and (_20579_, _12986_, _05298_);
  or (_20580_, _20509_, _04527_);
  or (_20581_, _20580_, _20579_);
  and (_20583_, _06337_, _05298_);
  or (_20584_, _20583_, _20509_);
  or (_20585_, _20584_, _04509_);
  and (_20586_, _20585_, _03745_);
  and (_20587_, _20586_, _20581_);
  and (_20588_, _20587_, _20578_);
  and (_20589_, _12992_, _05298_);
  or (_20590_, _20589_, _20509_);
  and (_20591_, _20590_, _03744_);
  or (_20592_, _20591_, _20588_);
  and (_20594_, _20592_, _04523_);
  or (_20595_, _20509_, _05880_);
  and (_20596_, _20584_, _03611_);
  and (_20597_, _20596_, _20595_);
  or (_20598_, _20597_, _20594_);
  and (_20599_, _20598_, _03734_);
  and (_20600_, _20522_, _03733_);
  and (_20601_, _20600_, _20595_);
  or (_20602_, _20601_, _03618_);
  or (_20603_, _20602_, _20599_);
  nor (_20604_, _12985_, _09311_);
  or (_20605_, _20509_, _06453_);
  or (_20606_, _20605_, _20604_);
  and (_20607_, _20606_, _06458_);
  and (_20608_, _20607_, _20603_);
  nor (_20609_, _12991_, _09311_);
  or (_20610_, _20609_, _20509_);
  and (_20611_, _20610_, _03741_);
  or (_20612_, _20611_, _03767_);
  or (_20613_, _20612_, _20608_);
  or (_20615_, _20519_, _03948_);
  and (_20616_, _20615_, _03446_);
  and (_20617_, _20616_, _20613_);
  and (_20618_, _20515_, _03445_);
  or (_20619_, _20618_, _03473_);
  or (_20620_, _20619_, _20617_);
  and (_20621_, _13051_, _05298_);
  or (_20622_, _20509_, _03474_);
  or (_20623_, _20622_, _20621_);
  and (_20624_, _20623_, _43189_);
  and (_20626_, _20624_, _20620_);
  nor (_20627_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_20628_, _20627_, _05173_);
  or (_43791_, _20628_, _20626_);
  not (_20629_, \oc8051_golden_model_1.P0 [5]);
  nor (_20630_, _43189_, _20629_);
  or (_20631_, _20630_, rst);
  nor (_20632_, _05298_, _20629_);
  nor (_20633_, _13070_, _09311_);
  or (_20634_, _20633_, _20632_);
  or (_20635_, _20634_, _04432_);
  and (_20636_, _05298_, \oc8051_golden_model_1.ACC [5]);
  or (_20637_, _20636_, _20632_);
  and (_20638_, _20637_, _04436_);
  nor (_20639_, _04436_, _20629_);
  or (_20640_, _20639_, _03534_);
  or (_20641_, _20640_, _20638_);
  and (_20642_, _20641_, _03470_);
  and (_20643_, _20642_, _20635_);
  nor (_20644_, _05258_, _20629_);
  and (_20646_, _13095_, _05258_);
  or (_20647_, _20646_, _20644_);
  and (_20648_, _20647_, _03469_);
  or (_20649_, _20648_, _03527_);
  or (_20650_, _20649_, _20643_);
  nor (_20651_, _05526_, _09311_);
  or (_20652_, _20651_, _20632_);
  or (_20653_, _20652_, _04457_);
  and (_20654_, _20653_, _20650_);
  or (_20655_, _20654_, _03530_);
  or (_20657_, _20637_, _03531_);
  and (_20658_, _20657_, _03466_);
  and (_20659_, _20658_, _20655_);
  and (_20660_, _13078_, _05258_);
  or (_20661_, _20660_, _20644_);
  and (_20662_, _20661_, _03465_);
  or (_20663_, _20662_, _03458_);
  or (_20664_, _20663_, _20659_);
  or (_20665_, _20644_, _13110_);
  and (_20666_, _20665_, _20647_);
  or (_20667_, _20666_, _03459_);
  and (_20668_, _20667_, _03453_);
  and (_20669_, _20668_, _20664_);
  or (_20670_, _13078_, _13075_);
  and (_20671_, _20670_, _05258_);
  or (_20672_, _20671_, _20644_);
  and (_20673_, _20672_, _03452_);
  or (_20674_, _20673_, _07454_);
  or (_20675_, _20674_, _20669_);
  or (_20676_, _20652_, _06903_);
  and (_20678_, _20676_, _20675_);
  or (_20679_, _20678_, _04082_);
  and (_20680_, _06757_, _05298_);
  or (_20681_, _20632_, _04500_);
  or (_20682_, _20681_, _20680_);
  and (_20683_, _20682_, _03521_);
  and (_20684_, _20683_, _20679_);
  or (_20685_, _13147_, _13149_);
  and (_20686_, _06344_, \oc8051_golden_model_1.P3 [5]);
  or (_20687_, _20686_, _13173_);
  nor (_20689_, _20687_, _20685_);
  nand (_20690_, _20689_, _13146_);
  not (_20691_, _13176_);
  and (_20692_, _13168_, _20691_);
  nand (_20693_, _20692_, _13159_);
  nor (_20694_, _13177_, _13174_);
  nand (_20695_, _20694_, _13171_);
  and (_20696_, _06329_, \oc8051_golden_model_1.P2 [5]);
  and (_20697_, _06334_, \oc8051_golden_model_1.P0 [5]);
  and (_20698_, _06340_, \oc8051_golden_model_1.P1 [5]);
  or (_20699_, _20698_, _20697_);
  or (_20700_, _20699_, _20696_);
  or (_20701_, _20700_, _20695_);
  or (_20702_, _20701_, _20693_);
  or (_20703_, _20702_, _20690_);
  or (_20704_, _20703_, _13137_);
  and (_20705_, _20704_, _05298_);
  or (_20706_, _20705_, _20632_);
  and (_20707_, _20706_, _03224_);
  or (_20708_, _20707_, _08905_);
  or (_20710_, _20708_, _20684_);
  and (_20711_, _13198_, _05298_);
  or (_20712_, _20632_, _04527_);
  or (_20713_, _20712_, _20711_);
  and (_20714_, _06295_, _05298_);
  or (_20715_, _20714_, _20632_);
  or (_20716_, _20715_, _04509_);
  and (_20717_, _20716_, _03745_);
  and (_20718_, _20717_, _20713_);
  and (_20719_, _20718_, _20710_);
  and (_20721_, _13204_, _05298_);
  or (_20722_, _20721_, _20632_);
  and (_20723_, _20722_, _03744_);
  or (_20724_, _20723_, _20719_);
  and (_20725_, _20724_, _04523_);
  or (_20726_, _20632_, _05576_);
  and (_20727_, _20715_, _03611_);
  and (_20728_, _20727_, _20726_);
  or (_20729_, _20728_, _20725_);
  and (_20730_, _20729_, _03734_);
  and (_20731_, _20637_, _03733_);
  and (_20732_, _20731_, _20726_);
  or (_20733_, _20732_, _03618_);
  or (_20734_, _20733_, _20730_);
  nor (_20735_, _13197_, _09311_);
  or (_20736_, _20632_, _06453_);
  or (_20737_, _20736_, _20735_);
  and (_20738_, _20737_, _06458_);
  and (_20739_, _20738_, _20734_);
  nor (_20740_, _13203_, _09311_);
  or (_20742_, _20740_, _20632_);
  and (_20743_, _20742_, _03741_);
  or (_20744_, _20743_, _03767_);
  or (_20745_, _20744_, _20739_);
  or (_20746_, _20634_, _03948_);
  and (_20747_, _20746_, _03446_);
  and (_20748_, _20747_, _20745_);
  and (_20749_, _20661_, _03445_);
  or (_20750_, _20749_, _03473_);
  or (_20751_, _20750_, _20748_);
  and (_20753_, _13253_, _05298_);
  or (_20754_, _20632_, _03474_);
  or (_20755_, _20754_, _20753_);
  and (_20756_, _20755_, _43189_);
  and (_20757_, _20756_, _20751_);
  or (_43792_, _20757_, _20631_);
  and (_20758_, _09311_, \oc8051_golden_model_1.P0 [6]);
  nor (_20759_, _13293_, _09311_);
  or (_20760_, _20759_, _20758_);
  or (_20761_, _20760_, _04432_);
  and (_20762_, _05298_, \oc8051_golden_model_1.ACC [6]);
  or (_20763_, _20762_, _20758_);
  and (_20764_, _20763_, _04436_);
  and (_20765_, _04437_, \oc8051_golden_model_1.P0 [6]);
  or (_20766_, _20765_, _03534_);
  or (_20767_, _20766_, _20764_);
  and (_20768_, _20767_, _03470_);
  and (_20769_, _20768_, _20761_);
  and (_20770_, _20142_, \oc8051_golden_model_1.P0 [6]);
  and (_20771_, _13280_, _05258_);
  or (_20773_, _20771_, _20770_);
  and (_20774_, _20773_, _03469_);
  or (_20775_, _20774_, _03527_);
  or (_20776_, _20775_, _20769_);
  nor (_20777_, _05417_, _09311_);
  or (_20778_, _20777_, _20758_);
  or (_20779_, _20778_, _04457_);
  and (_20780_, _20779_, _20776_);
  or (_20781_, _20780_, _03530_);
  or (_20782_, _20763_, _03531_);
  and (_20784_, _20782_, _03466_);
  and (_20785_, _20784_, _20781_);
  and (_20786_, _13304_, _05258_);
  or (_20787_, _20786_, _20770_);
  and (_20788_, _20787_, _03465_);
  or (_20789_, _20788_, _03458_);
  or (_20790_, _20789_, _20785_);
  or (_20791_, _20770_, _13311_);
  and (_20792_, _20791_, _20773_);
  or (_20793_, _20792_, _03459_);
  and (_20794_, _20793_, _03453_);
  and (_20795_, _20794_, _20790_);
  or (_20796_, _13328_, _13304_);
  and (_20797_, _20796_, _05258_);
  or (_20798_, _20797_, _20770_);
  and (_20799_, _20798_, _03452_);
  or (_20800_, _20799_, _07454_);
  or (_20801_, _20800_, _20795_);
  or (_20802_, _20778_, _06903_);
  and (_20803_, _20802_, _20801_);
  or (_20805_, _20803_, _04082_);
  and (_20806_, _06526_, _05298_);
  or (_20807_, _20758_, _04500_);
  or (_20808_, _20807_, _20806_);
  and (_20809_, _20808_, _03521_);
  and (_20810_, _20809_, _20805_);
  and (_20811_, _06334_, \oc8051_golden_model_1.P0 [6]);
  and (_20812_, _06329_, \oc8051_golden_model_1.P2 [6]);
  and (_20813_, _06340_, \oc8051_golden_model_1.P1 [6]);
  and (_20814_, _06344_, \oc8051_golden_model_1.P3 [6]);
  or (_20816_, _20814_, _20813_);
  or (_20817_, _20816_, _20812_);
  nor (_20818_, _20817_, _20811_);
  and (_20819_, _20818_, _13348_);
  and (_20820_, _20819_, _13368_);
  nand (_20821_, _20820_, _13384_);
  or (_20822_, _20821_, _13341_);
  and (_20823_, _20822_, _05298_);
  or (_20824_, _20823_, _20758_);
  and (_20825_, _20824_, _03224_);
  or (_20826_, _20825_, _08905_);
  or (_20827_, _20826_, _20810_);
  and (_20828_, _13402_, _05298_);
  or (_20829_, _20758_, _04527_);
  or (_20830_, _20829_, _20828_);
  and (_20831_, _14949_, _05298_);
  or (_20832_, _20831_, _20758_);
  or (_20833_, _20832_, _04509_);
  and (_20834_, _20833_, _03745_);
  and (_20835_, _20834_, _20830_);
  and (_20837_, _20835_, _20827_);
  and (_20838_, _13407_, _05298_);
  or (_20839_, _20838_, _20758_);
  and (_20840_, _20839_, _03744_);
  or (_20841_, _20840_, _20837_);
  and (_20842_, _20841_, _04523_);
  or (_20843_, _20758_, _05469_);
  and (_20844_, _20832_, _03611_);
  and (_20845_, _20844_, _20843_);
  or (_20846_, _20845_, _20842_);
  and (_20848_, _20846_, _03734_);
  and (_20849_, _20763_, _03733_);
  and (_20850_, _20849_, _20843_);
  or (_20851_, _20850_, _03618_);
  or (_20852_, _20851_, _20848_);
  nor (_20853_, _13400_, _09311_);
  or (_20854_, _20758_, _06453_);
  or (_20855_, _20854_, _20853_);
  and (_20856_, _20855_, _06458_);
  and (_20857_, _20856_, _20852_);
  nor (_20858_, _13406_, _09311_);
  or (_20859_, _20858_, _20758_);
  and (_20860_, _20859_, _03741_);
  or (_20861_, _20860_, _03767_);
  or (_20862_, _20861_, _20857_);
  or (_20863_, _20760_, _03948_);
  and (_20864_, _20863_, _03446_);
  and (_20865_, _20864_, _20862_);
  and (_20866_, _20787_, _03445_);
  or (_20867_, _20866_, _03473_);
  or (_20869_, _20867_, _20865_);
  and (_20870_, _13456_, _05298_);
  or (_20871_, _20758_, _03474_);
  or (_20872_, _20871_, _20870_);
  and (_20873_, _20872_, _43189_);
  and (_20874_, _20873_, _20869_);
  nor (_20875_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_20876_, _20875_, _05173_);
  or (_43793_, _20876_, _20874_);
  nor (_20877_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_20879_, _20877_, _05173_);
  and (_20880_, _09427_, \oc8051_golden_model_1.P1 [0]);
  and (_20881_, _12183_, _05284_);
  or (_20882_, _20881_, _20880_);
  and (_20883_, _20882_, _03744_);
  and (_20884_, _05284_, _04429_);
  or (_20885_, _20884_, _20880_);
  or (_20886_, _20885_, _06903_);
  nor (_20887_, _05722_, _09427_);
  or (_20888_, _20887_, _20880_);
  or (_20889_, _20888_, _04432_);
  and (_20890_, _05284_, \oc8051_golden_model_1.ACC [0]);
  or (_20891_, _20890_, _20880_);
  and (_20892_, _20891_, _04436_);
  and (_20893_, _04437_, \oc8051_golden_model_1.P1 [0]);
  or (_20894_, _20893_, _03534_);
  or (_20895_, _20894_, _20892_);
  and (_20896_, _20895_, _03470_);
  and (_20897_, _20896_, _20889_);
  not (_20898_, _05951_);
  and (_20900_, _20898_, \oc8051_golden_model_1.P1 [0]);
  and (_20901_, _12075_, _05951_);
  or (_20902_, _20901_, _20900_);
  and (_20903_, _20902_, _03469_);
  or (_20904_, _20903_, _20897_);
  and (_20905_, _20904_, _04457_);
  and (_20906_, _20885_, _03527_);
  or (_20907_, _20906_, _03530_);
  or (_20908_, _20907_, _20905_);
  or (_20909_, _20891_, _03531_);
  and (_20911_, _20909_, _03466_);
  and (_20912_, _20911_, _20908_);
  and (_20913_, _20880_, _03465_);
  or (_20914_, _20913_, _03458_);
  or (_20915_, _20914_, _20912_);
  or (_20916_, _20888_, _03459_);
  and (_20917_, _20916_, _03453_);
  and (_20918_, _20917_, _20915_);
  and (_20919_, _20052_, _05951_);
  or (_20920_, _20919_, _20900_);
  and (_20921_, _20920_, _03452_);
  or (_20922_, _20921_, _07454_);
  or (_20923_, _20922_, _20918_);
  and (_20924_, _20923_, _20886_);
  or (_20925_, _20924_, _04082_);
  and (_20926_, _06617_, _05284_);
  or (_20927_, _20880_, _04500_);
  or (_20928_, _20927_, _20926_);
  and (_20929_, _20928_, _03521_);
  and (_20930_, _20929_, _20925_);
  and (_20932_, _20077_, _05284_);
  or (_20933_, _20932_, _20880_);
  and (_20934_, _20933_, _03224_);
  or (_20935_, _20934_, _20930_);
  or (_20936_, _20935_, _08905_);
  and (_20937_, _12177_, _05284_);
  or (_20938_, _20880_, _04527_);
  or (_20939_, _20938_, _20937_);
  and (_20940_, _05284_, _06350_);
  or (_20941_, _20940_, _20880_);
  or (_20943_, _20941_, _04509_);
  and (_20944_, _20943_, _03745_);
  and (_20945_, _20944_, _20939_);
  and (_20946_, _20945_, _20936_);
  or (_20947_, _20946_, _20883_);
  and (_20948_, _20947_, _04523_);
  nand (_20949_, _20941_, _03611_);
  nor (_20950_, _20949_, _20887_);
  or (_20951_, _20950_, _20948_);
  and (_20952_, _20951_, _03734_);
  or (_20954_, _20880_, _05722_);
  and (_20955_, _20891_, _03733_);
  and (_20956_, _20955_, _20954_);
  or (_20957_, _20956_, _03618_);
  or (_20958_, _20957_, _20952_);
  nor (_20959_, _12057_, _09427_);
  or (_20960_, _20880_, _06453_);
  or (_20961_, _20960_, _20959_);
  and (_20962_, _20961_, _06458_);
  and (_20963_, _20962_, _20958_);
  nor (_20964_, _12181_, _09427_);
  or (_20965_, _20964_, _20880_);
  and (_20966_, _20965_, _03741_);
  or (_20967_, _20966_, _03767_);
  or (_20968_, _20967_, _20963_);
  or (_20969_, _20888_, _03948_);
  and (_20970_, _20969_, _03446_);
  and (_20971_, _20970_, _20968_);
  and (_20972_, _20880_, _03445_);
  or (_20973_, _20972_, _03473_);
  or (_20975_, _20973_, _20971_);
  or (_20976_, _20888_, _03474_);
  and (_20977_, _20976_, _43189_);
  and (_20978_, _20977_, _20975_);
  or (_43794_, _20978_, _20879_);
  or (_20979_, _05284_, \oc8051_golden_model_1.P1 [1]);
  and (_20980_, _12265_, _05284_);
  not (_20981_, _20980_);
  and (_20982_, _20981_, _20979_);
  or (_20983_, _20982_, _04432_);
  nand (_20985_, _05284_, _03269_);
  and (_20986_, _20985_, _20979_);
  and (_20987_, _20986_, _04436_);
  and (_20988_, _04437_, \oc8051_golden_model_1.P1 [1]);
  or (_20989_, _20988_, _03534_);
  or (_20990_, _20989_, _20987_);
  and (_20991_, _20990_, _03470_);
  and (_20992_, _20991_, _20983_);
  and (_20993_, _12269_, _05951_);
  and (_20994_, _20898_, \oc8051_golden_model_1.P1 [1]);
  or (_20995_, _20994_, _03527_);
  or (_20996_, _20995_, _20993_);
  and (_20997_, _20996_, _03533_);
  or (_20998_, _20997_, _20992_);
  and (_20999_, _09427_, \oc8051_golden_model_1.P1 [1]);
  nor (_21000_, _09427_, _04635_);
  or (_21001_, _21000_, _20999_);
  or (_21002_, _21001_, _04457_);
  and (_21003_, _21002_, _20998_);
  or (_21004_, _21003_, _03530_);
  or (_21006_, _20986_, _03531_);
  and (_21007_, _21006_, _03466_);
  and (_21008_, _21007_, _21004_);
  and (_21009_, _12256_, _05951_);
  or (_21010_, _21009_, _20994_);
  and (_21011_, _21010_, _03465_);
  or (_21012_, _21011_, _03458_);
  or (_21013_, _21012_, _21008_);
  and (_21014_, _20993_, _12284_);
  or (_21015_, _20994_, _03459_);
  or (_21017_, _21015_, _21014_);
  and (_21018_, _21017_, _21013_);
  and (_21019_, _21018_, _03453_);
  and (_21020_, _20170_, _05951_);
  or (_21021_, _20994_, _21020_);
  and (_21022_, _21021_, _03452_);
  or (_21023_, _21022_, _07454_);
  or (_21024_, _21023_, _21019_);
  or (_21025_, _21001_, _06903_);
  and (_21026_, _21025_, _21024_);
  or (_21028_, _21026_, _04082_);
  and (_21029_, _06572_, _05284_);
  or (_21030_, _20999_, _04500_);
  or (_21031_, _21030_, _21029_);
  and (_21032_, _21031_, _03521_);
  and (_21033_, _21032_, _21028_);
  and (_21034_, _20196_, _05284_);
  or (_21035_, _21034_, _20999_);
  and (_21036_, _21035_, _03224_);
  or (_21037_, _21036_, _21033_);
  and (_21038_, _21037_, _03625_);
  or (_21039_, _12375_, _09427_);
  and (_21040_, _21039_, _03623_);
  nand (_21041_, _05284_, _04325_);
  and (_21042_, _21041_, _03624_);
  or (_21043_, _21042_, _21040_);
  and (_21044_, _21043_, _20979_);
  or (_21045_, _21044_, _21038_);
  and (_21046_, _21045_, _03745_);
  or (_21047_, _12381_, _09427_);
  and (_21049_, _20979_, _03744_);
  and (_21050_, _21049_, _21047_);
  or (_21051_, _21050_, _21046_);
  and (_21052_, _21051_, _04523_);
  or (_21053_, _12374_, _09427_);
  and (_21054_, _20979_, _03611_);
  and (_21055_, _21054_, _21053_);
  or (_21056_, _21055_, _21052_);
  and (_21057_, _21056_, _03734_);
  or (_21058_, _20999_, _05674_);
  and (_21060_, _20986_, _03733_);
  and (_21061_, _21060_, _21058_);
  or (_21062_, _21061_, _21057_);
  and (_21063_, _21062_, _03742_);
  or (_21064_, _21041_, _05674_);
  and (_21065_, _20979_, _03618_);
  and (_21066_, _21065_, _21064_);
  or (_21067_, _20985_, _05674_);
  and (_21068_, _20979_, _03741_);
  and (_21069_, _21068_, _21067_);
  or (_21070_, _21069_, _03767_);
  or (_21071_, _21070_, _21066_);
  or (_21072_, _21071_, _21063_);
  or (_21073_, _20982_, _03948_);
  and (_21074_, _21073_, _03446_);
  and (_21075_, _21074_, _21072_);
  and (_21076_, _21010_, _03445_);
  or (_21077_, _21076_, _03473_);
  or (_21078_, _21077_, _21075_);
  or (_21079_, _20999_, _03474_);
  or (_21081_, _21079_, _20980_);
  and (_21082_, _21081_, _43189_);
  and (_21083_, _21082_, _21078_);
  nor (_21084_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_21085_, _21084_, _05173_);
  or (_43795_, _21085_, _21083_);
  not (_21086_, \oc8051_golden_model_1.P1 [2]);
  nor (_21087_, _43189_, _21086_);
  or (_21088_, _21087_, rst);
  nor (_21089_, _05284_, _21086_);
  nor (_21091_, _09427_, _05073_);
  or (_21092_, _21091_, _21089_);
  or (_21093_, _21092_, _06903_);
  and (_21094_, _21092_, _03527_);
  nor (_21095_, _05951_, _21086_);
  and (_21096_, _12462_, _05951_);
  or (_21097_, _21096_, _21095_);
  or (_21098_, _21097_, _03470_);
  nor (_21099_, _12467_, _09427_);
  or (_21100_, _21099_, _21089_);
  and (_21102_, _21100_, _03534_);
  nor (_21103_, _04436_, _21086_);
  and (_21104_, _05284_, \oc8051_golden_model_1.ACC [2]);
  or (_21105_, _21104_, _21089_);
  and (_21106_, _21105_, _04436_);
  or (_21107_, _21106_, _21103_);
  and (_21108_, _21107_, _04432_);
  or (_21109_, _21108_, _03469_);
  or (_21110_, _21109_, _21102_);
  and (_21111_, _21110_, _21098_);
  and (_21113_, _21111_, _04457_);
  or (_21114_, _21113_, _21094_);
  or (_21115_, _21114_, _03530_);
  or (_21116_, _21105_, _03531_);
  and (_21117_, _21116_, _03466_);
  and (_21118_, _21117_, _21115_);
  and (_21119_, _12460_, _05951_);
  or (_21120_, _21119_, _21095_);
  and (_21121_, _21120_, _03465_);
  or (_21122_, _21121_, _03458_);
  or (_21124_, _21122_, _21118_);
  or (_21125_, _21095_, _12491_);
  and (_21126_, _21125_, _21097_);
  or (_21127_, _21126_, _03459_);
  and (_21128_, _21127_, _03453_);
  and (_21129_, _21128_, _21124_);
  and (_21130_, _20293_, _05951_);
  or (_21131_, _21130_, _21095_);
  and (_21132_, _21131_, _03452_);
  or (_21133_, _21132_, _07454_);
  or (_21135_, _21133_, _21129_);
  and (_21136_, _21135_, _21093_);
  or (_21137_, _21136_, _04082_);
  and (_21138_, _06710_, _05284_);
  or (_21139_, _21089_, _04500_);
  or (_21140_, _21139_, _21138_);
  and (_21141_, _21140_, _03521_);
  and (_21142_, _21141_, _21137_);
  and (_21143_, _20318_, _05284_);
  or (_21144_, _21089_, _21143_);
  and (_21146_, _21144_, _03224_);
  or (_21147_, _21146_, _21142_);
  or (_21148_, _21147_, _08905_);
  and (_21149_, _12582_, _05284_);
  or (_21150_, _21089_, _04527_);
  or (_21151_, _21150_, _21149_);
  and (_21152_, _05284_, _06399_);
  or (_21153_, _21152_, _21089_);
  or (_21154_, _21153_, _04509_);
  and (_21155_, _21154_, _03745_);
  and (_21157_, _21155_, _21151_);
  and (_21158_, _21157_, _21148_);
  and (_21159_, _12588_, _05284_);
  or (_21160_, _21159_, _21089_);
  and (_21161_, _21160_, _03744_);
  or (_21162_, _21161_, _21158_);
  and (_21163_, _21162_, _04523_);
  or (_21164_, _21089_, _05772_);
  and (_21165_, _21153_, _03611_);
  and (_21166_, _21165_, _21164_);
  or (_21168_, _21166_, _21163_);
  and (_21169_, _21168_, _03734_);
  and (_21170_, _21105_, _03733_);
  and (_21171_, _21170_, _21164_);
  or (_21172_, _21171_, _03618_);
  or (_21173_, _21172_, _21169_);
  nor (_21174_, _12581_, _09427_);
  or (_21175_, _21089_, _06453_);
  or (_21176_, _21175_, _21174_);
  and (_21177_, _21176_, _06458_);
  and (_21178_, _21177_, _21173_);
  nor (_21179_, _12587_, _09427_);
  or (_21180_, _21179_, _21089_);
  and (_21181_, _21180_, _03741_);
  or (_21182_, _21181_, _03767_);
  or (_21183_, _21182_, _21178_);
  or (_21184_, _21100_, _03948_);
  and (_21185_, _21184_, _03446_);
  and (_21186_, _21185_, _21183_);
  and (_21187_, _21120_, _03445_);
  or (_21188_, _21187_, _03473_);
  or (_21189_, _21188_, _21186_);
  and (_21190_, _12638_, _05284_);
  or (_21191_, _21089_, _03474_);
  or (_21192_, _21191_, _21190_);
  and (_21193_, _21192_, _43189_);
  and (_21194_, _21193_, _21189_);
  or (_43796_, _21194_, _21088_);
  and (_21195_, _09427_, \oc8051_golden_model_1.P1 [3]);
  nor (_21196_, _09427_, _04885_);
  or (_21198_, _21196_, _21195_);
  or (_21199_, _21198_, _06903_);
  nor (_21200_, _12652_, _09427_);
  or (_21201_, _21200_, _21195_);
  or (_21202_, _21201_, _04432_);
  and (_21203_, _05284_, \oc8051_golden_model_1.ACC [3]);
  or (_21204_, _21203_, _21195_);
  and (_21205_, _21204_, _04436_);
  and (_21206_, _04437_, \oc8051_golden_model_1.P1 [3]);
  or (_21207_, _21206_, _03534_);
  or (_21209_, _21207_, _21205_);
  and (_21210_, _21209_, _03470_);
  and (_21211_, _21210_, _21202_);
  and (_21212_, _20898_, \oc8051_golden_model_1.P1 [3]);
  and (_21213_, _12664_, _05951_);
  or (_21214_, _21213_, _21212_);
  and (_21215_, _21214_, _03469_);
  or (_21216_, _21215_, _03527_);
  or (_21217_, _21216_, _21211_);
  or (_21218_, _21198_, _04457_);
  and (_21220_, _21218_, _21217_);
  or (_21221_, _21220_, _03530_);
  or (_21222_, _21204_, _03531_);
  and (_21223_, _21222_, _03466_);
  and (_21224_, _21223_, _21221_);
  and (_21225_, _12662_, _05951_);
  or (_21226_, _21225_, _21212_);
  and (_21227_, _21226_, _03465_);
  or (_21228_, _21227_, _03458_);
  or (_21229_, _21228_, _21224_);
  or (_21231_, _21212_, _12691_);
  and (_21232_, _21231_, _21214_);
  or (_21233_, _21232_, _03459_);
  and (_21234_, _21233_, _03453_);
  and (_21235_, _21234_, _21229_);
  and (_21236_, _20419_, _05951_);
  or (_21237_, _21236_, _21212_);
  and (_21238_, _21237_, _03452_);
  or (_21239_, _21238_, _07454_);
  or (_21240_, _21239_, _21235_);
  and (_21242_, _21240_, _21199_);
  or (_21243_, _21242_, _04082_);
  and (_21244_, _06664_, _05284_);
  or (_21245_, _21195_, _04500_);
  or (_21246_, _21245_, _21244_);
  and (_21247_, _21246_, _03521_);
  and (_21248_, _21247_, _21243_);
  and (_21249_, _20454_, _05284_);
  or (_21250_, _21195_, _21249_);
  and (_21251_, _21250_, _03224_);
  or (_21253_, _21251_, _21248_);
  or (_21254_, _21253_, _08905_);
  and (_21255_, _12787_, _05284_);
  or (_21256_, _21195_, _04527_);
  or (_21257_, _21256_, _21255_);
  and (_21258_, _05284_, _06356_);
  or (_21259_, _21258_, _21195_);
  or (_21260_, _21259_, _04509_);
  and (_21261_, _21260_, _03745_);
  and (_21262_, _21261_, _21257_);
  and (_21264_, _21262_, _21254_);
  and (_21265_, _12793_, _05284_);
  or (_21266_, _21265_, _21195_);
  and (_21267_, _21266_, _03744_);
  or (_21268_, _21267_, _21264_);
  and (_21269_, _21268_, _04523_);
  or (_21270_, _21195_, _05625_);
  and (_21271_, _21259_, _03611_);
  and (_21272_, _21271_, _21270_);
  or (_21273_, _21272_, _21269_);
  and (_21275_, _21273_, _03734_);
  and (_21276_, _21204_, _03733_);
  and (_21277_, _21276_, _21270_);
  or (_21278_, _21277_, _03618_);
  or (_21279_, _21278_, _21275_);
  nor (_21280_, _12786_, _09427_);
  or (_21281_, _21195_, _06453_);
  or (_21282_, _21281_, _21280_);
  and (_21283_, _21282_, _06458_);
  and (_21284_, _21283_, _21279_);
  nor (_21286_, _12792_, _09427_);
  or (_21287_, _21286_, _21195_);
  and (_21288_, _21287_, _03741_);
  or (_21289_, _21288_, _03767_);
  or (_21290_, _21289_, _21284_);
  or (_21291_, _21201_, _03948_);
  and (_21292_, _21291_, _03446_);
  and (_21293_, _21292_, _21290_);
  and (_21294_, _21226_, _03445_);
  or (_21295_, _21294_, _03473_);
  or (_21297_, _21295_, _21293_);
  and (_21298_, _12843_, _05284_);
  or (_21299_, _21195_, _03474_);
  or (_21300_, _21299_, _21298_);
  and (_21301_, _21300_, _43189_);
  and (_21302_, _21301_, _21297_);
  nor (_21303_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_21304_, _21303_, _05173_);
  or (_43797_, _21304_, _21302_);
  nor (_21305_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_21307_, _21305_, _05173_);
  and (_21308_, _09427_, \oc8051_golden_model_1.P1 [4]);
  nor (_21309_, _05831_, _09427_);
  or (_21310_, _21309_, _21308_);
  or (_21311_, _21310_, _06903_);
  and (_21312_, _20898_, \oc8051_golden_model_1.P1 [4]);
  and (_21313_, _12864_, _05951_);
  or (_21314_, _21313_, _21312_);
  and (_21315_, _21314_, _03465_);
  nor (_21316_, _12856_, _09427_);
  or (_21318_, _21316_, _21308_);
  or (_21319_, _21318_, _04432_);
  and (_21320_, _05284_, \oc8051_golden_model_1.ACC [4]);
  or (_21321_, _21320_, _21308_);
  and (_21322_, _21321_, _04436_);
  and (_21323_, _04437_, \oc8051_golden_model_1.P1 [4]);
  or (_21324_, _21323_, _03534_);
  or (_21325_, _21324_, _21322_);
  and (_21326_, _21325_, _03470_);
  and (_21327_, _21326_, _21319_);
  and (_21329_, _12866_, _05951_);
  or (_21330_, _21329_, _21312_);
  and (_21331_, _21330_, _03469_);
  or (_21332_, _21331_, _03527_);
  or (_21333_, _21332_, _21327_);
  or (_21334_, _21310_, _04457_);
  and (_21335_, _21334_, _21333_);
  or (_21336_, _21335_, _03530_);
  or (_21337_, _21321_, _03531_);
  and (_21338_, _21337_, _03466_);
  and (_21340_, _21338_, _21336_);
  or (_21341_, _21340_, _21315_);
  and (_21342_, _21341_, _03459_);
  and (_21343_, _12895_, _05951_);
  or (_21344_, _21343_, _21312_);
  and (_21345_, _21344_, _03458_);
  or (_21346_, _21345_, _21342_);
  and (_21347_, _21346_, _03453_);
  and (_21348_, _20548_, _05951_);
  or (_21349_, _21348_, _21312_);
  and (_21351_, _21349_, _03452_);
  or (_21352_, _21351_, _07454_);
  or (_21353_, _21352_, _21347_);
  and (_21354_, _21353_, _21311_);
  or (_21355_, _21354_, _04082_);
  and (_21356_, _06802_, _05284_);
  or (_21357_, _21308_, _04500_);
  or (_21358_, _21357_, _21356_);
  and (_21359_, _21358_, _03521_);
  and (_21360_, _21359_, _21355_);
  and (_21362_, _20573_, _05284_);
  or (_21363_, _21362_, _21308_);
  and (_21364_, _21363_, _03224_);
  or (_21365_, _21364_, _08905_);
  or (_21366_, _21365_, _21360_);
  and (_21367_, _12986_, _05284_);
  or (_21368_, _21308_, _04527_);
  or (_21369_, _21368_, _21367_);
  and (_21370_, _06337_, _05284_);
  or (_21371_, _21370_, _21308_);
  or (_21373_, _21371_, _04509_);
  and (_21374_, _21373_, _03745_);
  and (_21375_, _21374_, _21369_);
  and (_21376_, _21375_, _21366_);
  and (_21377_, _12992_, _05284_);
  or (_21378_, _21377_, _21308_);
  and (_21379_, _21378_, _03744_);
  or (_21380_, _21379_, _21376_);
  and (_21381_, _21380_, _04523_);
  or (_21382_, _21308_, _05880_);
  and (_21384_, _21371_, _03611_);
  and (_21385_, _21384_, _21382_);
  or (_21386_, _21385_, _21381_);
  and (_21387_, _21386_, _03734_);
  and (_21388_, _21321_, _03733_);
  and (_21389_, _21388_, _21382_);
  or (_21390_, _21389_, _03618_);
  or (_21391_, _21390_, _21387_);
  nor (_21392_, _12985_, _09427_);
  or (_21393_, _21308_, _06453_);
  or (_21395_, _21393_, _21392_);
  and (_21396_, _21395_, _06458_);
  and (_21397_, _21396_, _21391_);
  nor (_21398_, _12991_, _09427_);
  or (_21399_, _21398_, _21308_);
  and (_21400_, _21399_, _03741_);
  or (_21401_, _21400_, _03767_);
  or (_21402_, _21401_, _21397_);
  or (_21403_, _21318_, _03948_);
  and (_21404_, _21403_, _03446_);
  and (_21406_, _21404_, _21402_);
  and (_21407_, _21314_, _03445_);
  or (_21408_, _21407_, _03473_);
  or (_21409_, _21408_, _21406_);
  and (_21410_, _13051_, _05284_);
  or (_21411_, _21308_, _03474_);
  or (_21412_, _21411_, _21410_);
  and (_21413_, _21412_, _43189_);
  and (_21414_, _21413_, _21409_);
  or (_43800_, _21414_, _21307_);
  and (_21416_, _09427_, \oc8051_golden_model_1.P1 [5]);
  nor (_21417_, _13070_, _09427_);
  or (_21418_, _21417_, _21416_);
  or (_21419_, _21418_, _04432_);
  and (_21420_, _05284_, \oc8051_golden_model_1.ACC [5]);
  or (_21421_, _21420_, _21416_);
  and (_21422_, _21421_, _04436_);
  and (_21423_, _04437_, \oc8051_golden_model_1.P1 [5]);
  or (_21424_, _21423_, _03534_);
  or (_21425_, _21424_, _21422_);
  and (_21427_, _21425_, _03470_);
  and (_21428_, _21427_, _21419_);
  and (_21429_, _20898_, \oc8051_golden_model_1.P1 [5]);
  and (_21430_, _13095_, _05951_);
  or (_21431_, _21430_, _21429_);
  and (_21432_, _21431_, _03469_);
  or (_21433_, _21432_, _03527_);
  or (_21434_, _21433_, _21428_);
  nor (_21435_, _05526_, _09427_);
  or (_21436_, _21435_, _21416_);
  or (_21438_, _21436_, _04457_);
  and (_21439_, _21438_, _21434_);
  or (_21440_, _21439_, _03530_);
  or (_21441_, _21421_, _03531_);
  and (_21442_, _21441_, _03466_);
  and (_21443_, _21442_, _21440_);
  and (_21444_, _13078_, _05951_);
  or (_21445_, _21444_, _21429_);
  and (_21446_, _21445_, _03465_);
  or (_21447_, _21446_, _03458_);
  or (_21449_, _21447_, _21443_);
  or (_21450_, _21429_, _13110_);
  and (_21451_, _21450_, _21431_);
  or (_21452_, _21451_, _03459_);
  and (_21453_, _21452_, _03453_);
  and (_21454_, _21453_, _21449_);
  and (_21455_, _20670_, _05951_);
  or (_21456_, _21455_, _21429_);
  and (_21457_, _21456_, _03452_);
  or (_21458_, _21457_, _07454_);
  or (_21460_, _21458_, _21454_);
  or (_21461_, _21436_, _06903_);
  and (_21462_, _21461_, _21460_);
  or (_21463_, _21462_, _04082_);
  and (_21464_, _06757_, _05284_);
  or (_21465_, _21416_, _04500_);
  or (_21466_, _21465_, _21464_);
  and (_21467_, _21466_, _03521_);
  and (_21468_, _21467_, _21463_);
  and (_21469_, _20704_, _05284_);
  or (_21471_, _21469_, _21416_);
  and (_21472_, _21471_, _03224_);
  or (_21473_, _21472_, _08905_);
  or (_21474_, _21473_, _21468_);
  and (_21475_, _13198_, _05284_);
  or (_21476_, _21416_, _04527_);
  or (_21477_, _21476_, _21475_);
  and (_21478_, _06295_, _05284_);
  or (_21479_, _21478_, _21416_);
  or (_21480_, _21479_, _04509_);
  and (_21482_, _21480_, _03745_);
  and (_21483_, _21482_, _21477_);
  and (_21484_, _21483_, _21474_);
  and (_21485_, _13204_, _05284_);
  or (_21486_, _21485_, _21416_);
  and (_21487_, _21486_, _03744_);
  or (_21488_, _21487_, _21484_);
  and (_21489_, _21488_, _04523_);
  or (_21490_, _21416_, _05576_);
  and (_21491_, _21479_, _03611_);
  and (_21494_, _21491_, _21490_);
  or (_21495_, _21494_, _21489_);
  and (_21496_, _21495_, _03734_);
  and (_21497_, _21421_, _03733_);
  and (_21498_, _21497_, _21490_);
  or (_21499_, _21498_, _03618_);
  or (_21500_, _21499_, _21496_);
  nor (_21501_, _13197_, _09427_);
  or (_21502_, _21416_, _06453_);
  or (_21503_, _21502_, _21501_);
  and (_21506_, _21503_, _06458_);
  and (_21507_, _21506_, _21500_);
  nor (_21508_, _13203_, _09427_);
  or (_21509_, _21508_, _21416_);
  and (_21510_, _21509_, _03741_);
  or (_21511_, _21510_, _03767_);
  or (_21512_, _21511_, _21507_);
  or (_21513_, _21418_, _03948_);
  and (_21514_, _21513_, _03446_);
  and (_21515_, _21514_, _21512_);
  and (_21518_, _21445_, _03445_);
  or (_21519_, _21518_, _03473_);
  or (_21520_, _21519_, _21515_);
  and (_21521_, _13253_, _05284_);
  or (_21522_, _21416_, _03474_);
  or (_21523_, _21522_, _21521_);
  and (_21524_, _21523_, _43189_);
  and (_21525_, _21524_, _21520_);
  nor (_21526_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_21527_, _21526_, _05173_);
  or (_43801_, _21527_, _21525_);
  and (_21530_, _09427_, \oc8051_golden_model_1.P1 [6]);
  nor (_21531_, _13293_, _09427_);
  or (_21532_, _21531_, _21530_);
  or (_21533_, _21532_, _04432_);
  and (_21534_, _05284_, \oc8051_golden_model_1.ACC [6]);
  or (_21535_, _21534_, _21530_);
  and (_21536_, _21535_, _04436_);
  and (_21537_, _04437_, \oc8051_golden_model_1.P1 [6]);
  or (_21538_, _21537_, _03534_);
  or (_21541_, _21538_, _21536_);
  and (_21542_, _21541_, _03470_);
  and (_21543_, _21542_, _21533_);
  and (_21544_, _20898_, \oc8051_golden_model_1.P1 [6]);
  and (_21545_, _13280_, _05951_);
  or (_21546_, _21545_, _21544_);
  and (_21547_, _21546_, _03469_);
  or (_21548_, _21547_, _03527_);
  or (_21549_, _21548_, _21543_);
  nor (_21550_, _05417_, _09427_);
  or (_21553_, _21550_, _21530_);
  or (_21554_, _21553_, _04457_);
  and (_21555_, _21554_, _21549_);
  or (_21556_, _21555_, _03530_);
  or (_21557_, _21535_, _03531_);
  and (_21558_, _21557_, _03466_);
  and (_21559_, _21558_, _21556_);
  and (_21560_, _13304_, _05951_);
  or (_21561_, _21560_, _21544_);
  and (_21562_, _21561_, _03465_);
  or (_21564_, _21562_, _03458_);
  or (_21565_, _21564_, _21559_);
  or (_21566_, _21544_, _13311_);
  and (_21567_, _21566_, _21546_);
  or (_21568_, _21567_, _03459_);
  and (_21569_, _21568_, _03453_);
  and (_21570_, _21569_, _21565_);
  and (_21571_, _20796_, _05951_);
  or (_21572_, _21571_, _21544_);
  and (_21573_, _21572_, _03452_);
  or (_21575_, _21573_, _07454_);
  or (_21576_, _21575_, _21570_);
  or (_21577_, _21553_, _06903_);
  and (_21578_, _21577_, _21576_);
  or (_21579_, _21578_, _04082_);
  and (_21580_, _06526_, _05284_);
  or (_21581_, _21530_, _04500_);
  or (_21582_, _21581_, _21580_);
  and (_21583_, _21582_, _03521_);
  and (_21584_, _21583_, _21579_);
  and (_21586_, _20822_, _05284_);
  or (_21587_, _21586_, _21530_);
  and (_21588_, _21587_, _03224_);
  or (_21589_, _21588_, _08905_);
  or (_21590_, _21589_, _21584_);
  and (_21591_, _13402_, _05284_);
  or (_21592_, _21530_, _04527_);
  or (_21593_, _21592_, _21591_);
  and (_21594_, _14949_, _05284_);
  or (_21595_, _21594_, _21530_);
  or (_21597_, _21595_, _04509_);
  and (_21598_, _21597_, _03745_);
  and (_21599_, _21598_, _21593_);
  and (_21600_, _21599_, _21590_);
  and (_21601_, _13407_, _05284_);
  or (_21602_, _21601_, _21530_);
  and (_21603_, _21602_, _03744_);
  or (_21604_, _21603_, _21600_);
  and (_21605_, _21604_, _04523_);
  or (_21606_, _21530_, _05469_);
  and (_21608_, _21595_, _03611_);
  and (_21609_, _21608_, _21606_);
  or (_21610_, _21609_, _21605_);
  and (_21611_, _21610_, _03734_);
  and (_21612_, _21535_, _03733_);
  and (_21613_, _21612_, _21606_);
  or (_21614_, _21613_, _03618_);
  or (_21615_, _21614_, _21611_);
  nor (_21616_, _13400_, _09427_);
  or (_21617_, _21530_, _06453_);
  or (_21619_, _21617_, _21616_);
  and (_21620_, _21619_, _06458_);
  and (_21621_, _21620_, _21615_);
  nor (_21622_, _13406_, _09427_);
  or (_21623_, _21622_, _21530_);
  and (_21624_, _21623_, _03741_);
  or (_21625_, _21624_, _03767_);
  or (_21626_, _21625_, _21621_);
  or (_21627_, _21532_, _03948_);
  and (_21628_, _21627_, _03446_);
  and (_21630_, _21628_, _21626_);
  and (_21631_, _21561_, _03445_);
  or (_21632_, _21631_, _03473_);
  or (_21633_, _21632_, _21630_);
  and (_21634_, _13456_, _05284_);
  or (_21635_, _21530_, _03474_);
  or (_21636_, _21635_, _21634_);
  and (_21637_, _21636_, _43189_);
  and (_21638_, _21637_, _21633_);
  nor (_21639_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_21641_, _21639_, _05173_);
  or (_43802_, _21641_, _21638_);
  and (_21642_, _09529_, \oc8051_golden_model_1.P2 [0]);
  and (_21643_, _12183_, _05289_);
  or (_21644_, _21643_, _21642_);
  and (_21645_, _21644_, _03744_);
  and (_21646_, _05289_, _04429_);
  or (_21647_, _21646_, _21642_);
  or (_21648_, _21647_, _06903_);
  nor (_21649_, _05722_, _09529_);
  or (_21651_, _21649_, _21642_);
  and (_21652_, _21651_, _03534_);
  and (_21653_, _04437_, \oc8051_golden_model_1.P2 [0]);
  and (_21654_, _05289_, \oc8051_golden_model_1.ACC [0]);
  or (_21655_, _21654_, _21642_);
  and (_21656_, _21655_, _04436_);
  or (_21657_, _21656_, _21653_);
  and (_21658_, _21657_, _04432_);
  or (_21659_, _21658_, _03469_);
  or (_21660_, _21659_, _21652_);
  and (_21662_, _12075_, _05948_);
  not (_21663_, _05948_);
  and (_21664_, _21663_, \oc8051_golden_model_1.P2 [0]);
  or (_21665_, _21664_, _03470_);
  or (_21666_, _21665_, _21662_);
  and (_21667_, _21666_, _04457_);
  and (_21668_, _21667_, _21660_);
  and (_21669_, _21647_, _03527_);
  or (_21670_, _21669_, _03530_);
  or (_21671_, _21670_, _21668_);
  or (_21673_, _21655_, _03531_);
  and (_21674_, _21673_, _03466_);
  and (_21675_, _21674_, _21671_);
  and (_21676_, _21642_, _03465_);
  or (_21677_, _21676_, _03458_);
  or (_21678_, _21677_, _21675_);
  or (_21679_, _21651_, _03459_);
  and (_21680_, _21679_, _03453_);
  and (_21681_, _21680_, _21678_);
  and (_21682_, _20052_, _05948_);
  or (_21684_, _21682_, _21664_);
  and (_21685_, _21684_, _03452_);
  or (_21686_, _21685_, _07454_);
  or (_21687_, _21686_, _21681_);
  and (_21688_, _21687_, _21648_);
  or (_21689_, _21688_, _04082_);
  and (_21690_, _06617_, _05289_);
  or (_21691_, _21642_, _04500_);
  or (_21692_, _21691_, _21690_);
  and (_21693_, _21692_, _03521_);
  and (_21695_, _21693_, _21689_);
  and (_21696_, _20077_, _05289_);
  or (_21697_, _21696_, _21642_);
  and (_21698_, _21697_, _03224_);
  or (_21699_, _21698_, _21695_);
  or (_21700_, _21699_, _08905_);
  and (_21701_, _12177_, _05289_);
  or (_21702_, _21642_, _04527_);
  or (_21703_, _21702_, _21701_);
  and (_21704_, _05289_, _06350_);
  or (_21706_, _21704_, _21642_);
  or (_21707_, _21706_, _04509_);
  and (_21708_, _21707_, _03745_);
  and (_21709_, _21708_, _21703_);
  and (_21710_, _21709_, _21700_);
  or (_21711_, _21710_, _21645_);
  and (_21712_, _21711_, _04523_);
  nand (_21713_, _21706_, _03611_);
  nor (_21714_, _21713_, _21649_);
  or (_21715_, _21714_, _21712_);
  and (_21717_, _21715_, _03734_);
  or (_21718_, _21642_, _05722_);
  and (_21719_, _21655_, _03733_);
  and (_21720_, _21719_, _21718_);
  or (_21721_, _21720_, _03618_);
  or (_21722_, _21721_, _21717_);
  nor (_21723_, _12057_, _09529_);
  or (_21724_, _21642_, _06453_);
  or (_21725_, _21724_, _21723_);
  and (_21726_, _21725_, _06458_);
  and (_21728_, _21726_, _21722_);
  nor (_21729_, _12181_, _09529_);
  or (_21730_, _21729_, _21642_);
  and (_21731_, _21730_, _03741_);
  or (_21732_, _21731_, _03767_);
  or (_21733_, _21732_, _21728_);
  or (_21734_, _21651_, _03948_);
  and (_21735_, _21734_, _03446_);
  and (_21736_, _21735_, _21733_);
  and (_21737_, _21642_, _03445_);
  or (_21739_, _21737_, _03473_);
  or (_21740_, _21739_, _21736_);
  or (_21741_, _21651_, _03474_);
  and (_21742_, _21741_, _43189_);
  and (_21743_, _21742_, _21740_);
  nor (_21744_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_21745_, _21744_, _05173_);
  or (_43805_, _21745_, _21743_);
  or (_21746_, _05289_, \oc8051_golden_model_1.P2 [1]);
  and (_21747_, _12265_, _05289_);
  not (_21749_, _21747_);
  and (_21750_, _21749_, _21746_);
  or (_21751_, _21750_, _04432_);
  nand (_21752_, _05289_, _03269_);
  and (_21753_, _21752_, _21746_);
  and (_21754_, _21753_, _04436_);
  and (_21755_, _04437_, \oc8051_golden_model_1.P2 [1]);
  or (_21756_, _21755_, _03534_);
  or (_21757_, _21756_, _21754_);
  and (_21758_, _21757_, _03470_);
  and (_21760_, _21758_, _21751_);
  and (_21761_, _12269_, _05948_);
  and (_21762_, _21663_, \oc8051_golden_model_1.P2 [1]);
  or (_21763_, _21762_, _03527_);
  or (_21764_, _21763_, _21761_);
  and (_21765_, _21764_, _03533_);
  or (_21766_, _21765_, _21760_);
  and (_21767_, _09529_, \oc8051_golden_model_1.P2 [1]);
  nor (_21768_, _09529_, _04635_);
  or (_21769_, _21768_, _21767_);
  or (_21771_, _21769_, _04457_);
  and (_21772_, _21771_, _21766_);
  or (_21773_, _21772_, _03530_);
  or (_21774_, _21753_, _03531_);
  and (_21775_, _21774_, _03466_);
  and (_21776_, _21775_, _21773_);
  and (_21777_, _12256_, _05948_);
  or (_21778_, _21777_, _21762_);
  and (_21779_, _21778_, _03465_);
  or (_21780_, _21779_, _03458_);
  or (_21782_, _21780_, _21776_);
  and (_21783_, _21761_, _12284_);
  or (_21784_, _21762_, _03459_);
  or (_21785_, _21784_, _21783_);
  and (_21786_, _21785_, _21782_);
  and (_21787_, _21786_, _03453_);
  and (_21788_, _20170_, _05948_);
  or (_21789_, _21762_, _21788_);
  and (_21790_, _21789_, _03452_);
  or (_21791_, _21790_, _07454_);
  or (_21793_, _21791_, _21787_);
  or (_21794_, _21769_, _06903_);
  and (_21795_, _21794_, _21793_);
  or (_21796_, _21795_, _04082_);
  and (_21797_, _06572_, _05289_);
  or (_21798_, _21767_, _04500_);
  or (_21799_, _21798_, _21797_);
  and (_21800_, _21799_, _03521_);
  and (_21801_, _21800_, _21796_);
  and (_21802_, _20196_, _05289_);
  or (_21804_, _21802_, _21767_);
  and (_21805_, _21804_, _03224_);
  or (_21806_, _21805_, _21801_);
  and (_21807_, _21806_, _03625_);
  or (_21808_, _12375_, _09529_);
  and (_21809_, _21808_, _03623_);
  nand (_21810_, _05289_, _04325_);
  and (_21811_, _21810_, _03624_);
  or (_21812_, _21811_, _21809_);
  and (_21813_, _21812_, _21746_);
  or (_21815_, _21813_, _21807_);
  and (_21816_, _21815_, _03745_);
  or (_21817_, _12381_, _09529_);
  and (_21818_, _21746_, _03744_);
  and (_21819_, _21818_, _21817_);
  or (_21820_, _21819_, _21816_);
  and (_21821_, _21820_, _04523_);
  or (_21822_, _12374_, _09529_);
  and (_21823_, _21746_, _03611_);
  and (_21824_, _21823_, _21822_);
  or (_21826_, _21824_, _21821_);
  and (_21827_, _21826_, _03734_);
  or (_21828_, _21767_, _05674_);
  and (_21829_, _21753_, _03733_);
  and (_21830_, _21829_, _21828_);
  or (_21831_, _21830_, _21827_);
  and (_21832_, _21831_, _03742_);
  or (_21833_, _21810_, _05674_);
  and (_21834_, _21746_, _03618_);
  and (_21835_, _21834_, _21833_);
  or (_21837_, _21752_, _05674_);
  and (_21838_, _21746_, _03741_);
  and (_21839_, _21838_, _21837_);
  or (_21840_, _21839_, _03767_);
  or (_21841_, _21840_, _21835_);
  or (_21842_, _21841_, _21832_);
  or (_21843_, _21750_, _03948_);
  and (_21844_, _21843_, _03446_);
  and (_21845_, _21844_, _21842_);
  and (_21846_, _21778_, _03445_);
  or (_21848_, _21846_, _03473_);
  or (_21849_, _21848_, _21845_);
  or (_21850_, _21767_, _03474_);
  or (_21851_, _21850_, _21747_);
  and (_21852_, _21851_, _43189_);
  and (_21853_, _21852_, _21849_);
  nor (_21854_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_21855_, _21854_, _05173_);
  or (_43806_, _21855_, _21853_);
  not (_21856_, \oc8051_golden_model_1.P2 [2]);
  nor (_21858_, _05289_, _21856_);
  nor (_21859_, _09529_, _05073_);
  or (_21860_, _21859_, _21858_);
  or (_21861_, _21860_, _06903_);
  and (_21862_, _21860_, _03527_);
  nor (_21863_, _05948_, _21856_);
  and (_21864_, _12462_, _05948_);
  or (_21865_, _21864_, _21863_);
  or (_21866_, _21865_, _03470_);
  nor (_21867_, _12467_, _09529_);
  or (_21869_, _21867_, _21858_);
  and (_21870_, _21869_, _03534_);
  nor (_21871_, _04436_, _21856_);
  and (_21872_, _05289_, \oc8051_golden_model_1.ACC [2]);
  or (_21873_, _21872_, _21858_);
  and (_21874_, _21873_, _04436_);
  or (_21875_, _21874_, _21871_);
  and (_21876_, _21875_, _04432_);
  or (_21877_, _21876_, _03469_);
  or (_21878_, _21877_, _21870_);
  and (_21880_, _21878_, _21866_);
  and (_21881_, _21880_, _04457_);
  or (_21882_, _21881_, _21862_);
  or (_21883_, _21882_, _03530_);
  or (_21884_, _21873_, _03531_);
  and (_21885_, _21884_, _03466_);
  and (_21886_, _21885_, _21883_);
  and (_21887_, _12460_, _05948_);
  or (_21888_, _21887_, _21863_);
  and (_21889_, _21888_, _03465_);
  or (_21891_, _21889_, _03458_);
  or (_21892_, _21891_, _21886_);
  or (_21893_, _21863_, _12491_);
  and (_21894_, _21893_, _21865_);
  or (_21895_, _21894_, _03459_);
  and (_21896_, _21895_, _03453_);
  and (_21897_, _21896_, _21892_);
  and (_21898_, _20293_, _05948_);
  or (_21899_, _21898_, _21863_);
  and (_21900_, _21899_, _03452_);
  or (_21902_, _21900_, _07454_);
  or (_21903_, _21902_, _21897_);
  and (_21904_, _21903_, _21861_);
  or (_21905_, _21904_, _04082_);
  and (_21906_, _06710_, _05289_);
  or (_21907_, _21858_, _04500_);
  or (_21908_, _21907_, _21906_);
  and (_21909_, _21908_, _03521_);
  and (_21910_, _21909_, _21905_);
  and (_21911_, _20318_, _05289_);
  or (_21913_, _21858_, _21911_);
  and (_21914_, _21913_, _03224_);
  or (_21915_, _21914_, _21910_);
  or (_21916_, _21915_, _08905_);
  and (_21917_, _12582_, _05289_);
  or (_21918_, _21858_, _04527_);
  or (_21919_, _21918_, _21917_);
  and (_21920_, _05289_, _06399_);
  or (_21921_, _21920_, _21858_);
  or (_21922_, _21921_, _04509_);
  and (_21924_, _21922_, _03745_);
  and (_21925_, _21924_, _21919_);
  and (_21926_, _21925_, _21916_);
  and (_21927_, _12588_, _05289_);
  or (_21928_, _21927_, _21858_);
  and (_21929_, _21928_, _03744_);
  or (_21930_, _21929_, _21926_);
  and (_21931_, _21930_, _04523_);
  or (_21932_, _21858_, _05772_);
  and (_21933_, _21921_, _03611_);
  and (_21935_, _21933_, _21932_);
  or (_21936_, _21935_, _21931_);
  and (_21937_, _21936_, _03734_);
  and (_21938_, _21873_, _03733_);
  and (_21939_, _21938_, _21932_);
  or (_21940_, _21939_, _03618_);
  or (_21941_, _21940_, _21937_);
  nor (_21942_, _12581_, _09529_);
  or (_21943_, _21858_, _06453_);
  or (_21944_, _21943_, _21942_);
  and (_21946_, _21944_, _06458_);
  and (_21947_, _21946_, _21941_);
  nor (_21948_, _12587_, _09529_);
  or (_21949_, _21948_, _21858_);
  and (_21950_, _21949_, _03741_);
  or (_21951_, _21950_, _03767_);
  or (_21952_, _21951_, _21947_);
  or (_21953_, _21869_, _03948_);
  and (_21954_, _21953_, _03446_);
  and (_21955_, _21954_, _21952_);
  and (_21957_, _21888_, _03445_);
  or (_21958_, _21957_, _03473_);
  or (_21959_, _21958_, _21955_);
  and (_21960_, _12638_, _05289_);
  or (_21961_, _21858_, _03474_);
  or (_21962_, _21961_, _21960_);
  and (_21963_, _21962_, _43189_);
  and (_21964_, _21963_, _21959_);
  nor (_21965_, _43189_, _21856_);
  or (_21966_, _21965_, rst);
  or (_43807_, _21966_, _21964_);
  and (_21968_, _09529_, \oc8051_golden_model_1.P2 [3]);
  nor (_21969_, _09529_, _04885_);
  or (_21970_, _21969_, _21968_);
  or (_21971_, _21970_, _06903_);
  nor (_21972_, _12652_, _09529_);
  or (_21973_, _21972_, _21968_);
  or (_21974_, _21973_, _04432_);
  and (_21975_, _05289_, \oc8051_golden_model_1.ACC [3]);
  or (_21976_, _21975_, _21968_);
  and (_21978_, _21976_, _04436_);
  and (_21979_, _04437_, \oc8051_golden_model_1.P2 [3]);
  or (_21980_, _21979_, _03534_);
  or (_21981_, _21980_, _21978_);
  and (_21982_, _21981_, _03470_);
  and (_21983_, _21982_, _21974_);
  and (_21984_, _21663_, \oc8051_golden_model_1.P2 [3]);
  and (_21985_, _12664_, _05948_);
  or (_21986_, _21985_, _21984_);
  and (_21987_, _21986_, _03469_);
  or (_21989_, _21987_, _03527_);
  or (_21990_, _21989_, _21983_);
  or (_21991_, _21970_, _04457_);
  and (_21992_, _21991_, _21990_);
  or (_21993_, _21992_, _03530_);
  or (_21994_, _21976_, _03531_);
  and (_21995_, _21994_, _03466_);
  and (_21996_, _21995_, _21993_);
  and (_21997_, _12662_, _05948_);
  or (_21998_, _21997_, _21984_);
  and (_22000_, _21998_, _03465_);
  or (_22001_, _22000_, _03458_);
  or (_22002_, _22001_, _21996_);
  or (_22003_, _21984_, _12691_);
  and (_22004_, _22003_, _21986_);
  or (_22005_, _22004_, _03459_);
  and (_22006_, _22005_, _03453_);
  and (_22007_, _22006_, _22002_);
  and (_22008_, _20419_, _05948_);
  or (_22009_, _22008_, _21984_);
  and (_22011_, _22009_, _03452_);
  or (_22012_, _22011_, _07454_);
  or (_22013_, _22012_, _22007_);
  and (_22014_, _22013_, _21971_);
  or (_22015_, _22014_, _04082_);
  and (_22016_, _06664_, _05289_);
  or (_22017_, _21968_, _04500_);
  or (_22018_, _22017_, _22016_);
  and (_22019_, _22018_, _03521_);
  and (_22020_, _22019_, _22015_);
  and (_22022_, _20454_, _05289_);
  or (_22023_, _21968_, _22022_);
  and (_22024_, _22023_, _03224_);
  or (_22025_, _22024_, _22020_);
  or (_22026_, _22025_, _08905_);
  and (_22027_, _12787_, _05289_);
  or (_22028_, _21968_, _04527_);
  or (_22029_, _22028_, _22027_);
  and (_22030_, _05289_, _06356_);
  or (_22031_, _22030_, _21968_);
  or (_22033_, _22031_, _04509_);
  and (_22034_, _22033_, _03745_);
  and (_22035_, _22034_, _22029_);
  and (_22036_, _22035_, _22026_);
  and (_22037_, _12793_, _05289_);
  or (_22038_, _22037_, _21968_);
  and (_22039_, _22038_, _03744_);
  or (_22040_, _22039_, _22036_);
  and (_22041_, _22040_, _04523_);
  or (_22042_, _21968_, _05625_);
  and (_22044_, _22031_, _03611_);
  and (_22045_, _22044_, _22042_);
  or (_22046_, _22045_, _22041_);
  and (_22047_, _22046_, _03734_);
  and (_22048_, _21976_, _03733_);
  and (_22049_, _22048_, _22042_);
  or (_22050_, _22049_, _03618_);
  or (_22051_, _22050_, _22047_);
  nor (_22052_, _12786_, _09529_);
  or (_22053_, _21968_, _06453_);
  or (_22054_, _22053_, _22052_);
  and (_22055_, _22054_, _06458_);
  and (_22056_, _22055_, _22051_);
  nor (_22057_, _12792_, _09529_);
  or (_22058_, _22057_, _21968_);
  and (_22059_, _22058_, _03741_);
  or (_22060_, _22059_, _03767_);
  or (_22061_, _22060_, _22056_);
  or (_22062_, _21973_, _03948_);
  and (_22063_, _22062_, _03446_);
  and (_22066_, _22063_, _22061_);
  and (_22067_, _21998_, _03445_);
  or (_22068_, _22067_, _03473_);
  or (_22069_, _22068_, _22066_);
  and (_22070_, _12843_, _05289_);
  or (_22071_, _21968_, _03474_);
  or (_22072_, _22071_, _22070_);
  and (_22073_, _22072_, _43189_);
  and (_22074_, _22073_, _22069_);
  nor (_22075_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_22077_, _22075_, _05173_);
  or (_43808_, _22077_, _22074_);
  nor (_22078_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_22079_, _22078_, _05173_);
  and (_22080_, _09529_, \oc8051_golden_model_1.P2 [4]);
  nor (_22081_, _05831_, _09529_);
  or (_22082_, _22081_, _22080_);
  or (_22083_, _22082_, _06903_);
  and (_22084_, _21663_, \oc8051_golden_model_1.P2 [4]);
  and (_22085_, _12864_, _05948_);
  or (_22087_, _22085_, _22084_);
  and (_22088_, _22087_, _03465_);
  nor (_22089_, _12856_, _09529_);
  or (_22090_, _22089_, _22080_);
  or (_22091_, _22090_, _04432_);
  and (_22092_, _05289_, \oc8051_golden_model_1.ACC [4]);
  or (_22093_, _22092_, _22080_);
  and (_22094_, _22093_, _04436_);
  and (_22095_, _04437_, \oc8051_golden_model_1.P2 [4]);
  or (_22096_, _22095_, _03534_);
  or (_22098_, _22096_, _22094_);
  and (_22099_, _22098_, _03470_);
  and (_22100_, _22099_, _22091_);
  and (_22101_, _12866_, _05948_);
  or (_22102_, _22101_, _22084_);
  and (_22103_, _22102_, _03469_);
  or (_22104_, _22103_, _03527_);
  or (_22105_, _22104_, _22100_);
  or (_22106_, _22082_, _04457_);
  and (_22107_, _22106_, _22105_);
  or (_22109_, _22107_, _03530_);
  or (_22110_, _22093_, _03531_);
  and (_22111_, _22110_, _03466_);
  and (_22112_, _22111_, _22109_);
  or (_22113_, _22112_, _22088_);
  and (_22114_, _22113_, _03459_);
  and (_22115_, _12895_, _05948_);
  or (_22116_, _22115_, _22084_);
  and (_22117_, _22116_, _03458_);
  or (_22118_, _22117_, _22114_);
  and (_22120_, _22118_, _03453_);
  and (_22121_, _20548_, _05948_);
  or (_22122_, _22121_, _22084_);
  and (_22123_, _22122_, _03452_);
  or (_22124_, _22123_, _07454_);
  or (_22125_, _22124_, _22120_);
  and (_22126_, _22125_, _22083_);
  or (_22127_, _22126_, _04082_);
  and (_22128_, _06802_, _05289_);
  or (_22129_, _22080_, _04500_);
  or (_22131_, _22129_, _22128_);
  and (_22132_, _22131_, _03521_);
  and (_22133_, _22132_, _22127_);
  and (_22134_, _20573_, _05289_);
  or (_22135_, _22134_, _22080_);
  and (_22136_, _22135_, _03224_);
  or (_22137_, _22136_, _08905_);
  or (_22138_, _22137_, _22133_);
  and (_22139_, _12986_, _05289_);
  or (_22140_, _22080_, _04527_);
  or (_22142_, _22140_, _22139_);
  and (_22143_, _06337_, _05289_);
  or (_22144_, _22143_, _22080_);
  or (_22145_, _22144_, _04509_);
  and (_22146_, _22145_, _03745_);
  and (_22147_, _22146_, _22142_);
  and (_22148_, _22147_, _22138_);
  and (_22149_, _12992_, _05289_);
  or (_22150_, _22149_, _22080_);
  and (_22151_, _22150_, _03744_);
  or (_22153_, _22151_, _22148_);
  and (_22154_, _22153_, _04523_);
  or (_22155_, _22080_, _05880_);
  and (_22156_, _22144_, _03611_);
  and (_22157_, _22156_, _22155_);
  or (_22158_, _22157_, _22154_);
  and (_22159_, _22158_, _03734_);
  and (_22160_, _22093_, _03733_);
  and (_22161_, _22160_, _22155_);
  or (_22162_, _22161_, _03618_);
  or (_22164_, _22162_, _22159_);
  nor (_22165_, _12985_, _09529_);
  or (_22166_, _22080_, _06453_);
  or (_22167_, _22166_, _22165_);
  and (_22168_, _22167_, _06458_);
  and (_22169_, _22168_, _22164_);
  nor (_22170_, _12991_, _09529_);
  or (_22171_, _22170_, _22080_);
  and (_22172_, _22171_, _03741_);
  or (_22173_, _22172_, _03767_);
  or (_22175_, _22173_, _22169_);
  or (_22176_, _22090_, _03948_);
  and (_22177_, _22176_, _03446_);
  and (_22178_, _22177_, _22175_);
  and (_22179_, _22087_, _03445_);
  or (_22180_, _22179_, _03473_);
  or (_22181_, _22180_, _22178_);
  and (_22182_, _13051_, _05289_);
  or (_22183_, _22080_, _03474_);
  or (_22184_, _22183_, _22182_);
  and (_22186_, _22184_, _43189_);
  and (_22187_, _22186_, _22181_);
  or (_43809_, _22187_, _22079_);
  and (_22188_, _09529_, \oc8051_golden_model_1.P2 [5]);
  nor (_22189_, _13070_, _09529_);
  or (_22190_, _22189_, _22188_);
  or (_22191_, _22190_, _04432_);
  and (_22192_, _05289_, \oc8051_golden_model_1.ACC [5]);
  or (_22193_, _22192_, _22188_);
  and (_22194_, _22193_, _04436_);
  and (_22196_, _04437_, \oc8051_golden_model_1.P2 [5]);
  or (_22197_, _22196_, _03534_);
  or (_22198_, _22197_, _22194_);
  and (_22199_, _22198_, _03470_);
  and (_22200_, _22199_, _22191_);
  and (_22201_, _21663_, \oc8051_golden_model_1.P2 [5]);
  and (_22202_, _13095_, _05948_);
  or (_22203_, _22202_, _22201_);
  and (_22204_, _22203_, _03469_);
  or (_22205_, _22204_, _03527_);
  or (_22207_, _22205_, _22200_);
  nor (_22208_, _05526_, _09529_);
  or (_22209_, _22208_, _22188_);
  or (_22210_, _22209_, _04457_);
  and (_22211_, _22210_, _22207_);
  or (_22212_, _22211_, _03530_);
  or (_22213_, _22193_, _03531_);
  and (_22214_, _22213_, _03466_);
  and (_22215_, _22214_, _22212_);
  and (_22216_, _13078_, _05948_);
  or (_22218_, _22216_, _22201_);
  and (_22219_, _22218_, _03465_);
  or (_22220_, _22219_, _03458_);
  or (_22221_, _22220_, _22215_);
  or (_22222_, _22201_, _13110_);
  and (_22223_, _22222_, _22203_);
  or (_22224_, _22223_, _03459_);
  and (_22225_, _22224_, _03453_);
  and (_22226_, _22225_, _22221_);
  and (_22227_, _20670_, _05948_);
  or (_22229_, _22227_, _22201_);
  and (_22230_, _22229_, _03452_);
  or (_22231_, _22230_, _07454_);
  or (_22232_, _22231_, _22226_);
  or (_22233_, _22209_, _06903_);
  and (_22234_, _22233_, _22232_);
  or (_22235_, _22234_, _04082_);
  and (_22236_, _06757_, _05289_);
  or (_22237_, _22188_, _04500_);
  or (_22238_, _22237_, _22236_);
  and (_22240_, _22238_, _03521_);
  and (_22241_, _22240_, _22235_);
  and (_22242_, _20704_, _05289_);
  or (_22243_, _22242_, _22188_);
  and (_22244_, _22243_, _03224_);
  or (_22245_, _22244_, _08905_);
  or (_22246_, _22245_, _22241_);
  and (_22247_, _13198_, _05289_);
  or (_22248_, _22188_, _04527_);
  or (_22249_, _22248_, _22247_);
  and (_22251_, _06295_, _05289_);
  or (_22252_, _22251_, _22188_);
  or (_22253_, _22252_, _04509_);
  and (_22254_, _22253_, _03745_);
  and (_22255_, _22254_, _22249_);
  and (_22256_, _22255_, _22246_);
  and (_22257_, _13204_, _05289_);
  or (_22258_, _22257_, _22188_);
  and (_22259_, _22258_, _03744_);
  or (_22260_, _22259_, _22256_);
  and (_22262_, _22260_, _04523_);
  or (_22263_, _22188_, _05576_);
  and (_22264_, _22252_, _03611_);
  and (_22265_, _22264_, _22263_);
  or (_22266_, _22265_, _22262_);
  and (_22267_, _22266_, _03734_);
  and (_22268_, _22193_, _03733_);
  and (_22269_, _22268_, _22263_);
  or (_22270_, _22269_, _03618_);
  or (_22271_, _22270_, _22267_);
  nor (_22273_, _13197_, _09529_);
  or (_22274_, _22188_, _06453_);
  or (_22275_, _22274_, _22273_);
  and (_22276_, _22275_, _06458_);
  and (_22277_, _22276_, _22271_);
  nor (_22278_, _13203_, _09529_);
  or (_22279_, _22278_, _22188_);
  and (_22280_, _22279_, _03741_);
  or (_22281_, _22280_, _03767_);
  or (_22282_, _22281_, _22277_);
  or (_22284_, _22190_, _03948_);
  and (_22285_, _22284_, _03446_);
  and (_22286_, _22285_, _22282_);
  and (_22287_, _22218_, _03445_);
  or (_22288_, _22287_, _03473_);
  or (_22289_, _22288_, _22286_);
  and (_22290_, _13253_, _05289_);
  or (_22291_, _22188_, _03474_);
  or (_22292_, _22291_, _22290_);
  and (_22293_, _22292_, _43189_);
  and (_22295_, _22293_, _22289_);
  nor (_22296_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_22297_, _22296_, _05173_);
  or (_43810_, _22297_, _22295_);
  nor (_22298_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_22299_, _22298_, _05173_);
  and (_22300_, _09529_, \oc8051_golden_model_1.P2 [6]);
  nor (_22301_, _13293_, _09529_);
  or (_22302_, _22301_, _22300_);
  or (_22303_, _22302_, _04432_);
  and (_22305_, _05289_, \oc8051_golden_model_1.ACC [6]);
  or (_22306_, _22305_, _22300_);
  and (_22307_, _22306_, _04436_);
  and (_22308_, _04437_, \oc8051_golden_model_1.P2 [6]);
  or (_22309_, _22308_, _03534_);
  or (_22310_, _22309_, _22307_);
  and (_22311_, _22310_, _03470_);
  and (_22312_, _22311_, _22303_);
  and (_22313_, _21663_, \oc8051_golden_model_1.P2 [6]);
  and (_22314_, _13280_, _05948_);
  or (_22316_, _22314_, _22313_);
  and (_22317_, _22316_, _03469_);
  or (_22318_, _22317_, _03527_);
  or (_22319_, _22318_, _22312_);
  nor (_22320_, _05417_, _09529_);
  or (_22321_, _22320_, _22300_);
  or (_22322_, _22321_, _04457_);
  and (_22323_, _22322_, _22319_);
  or (_22324_, _22323_, _03530_);
  or (_22325_, _22306_, _03531_);
  and (_22328_, _22325_, _03466_);
  and (_22329_, _22328_, _22324_);
  and (_22330_, _13304_, _05948_);
  or (_22331_, _22330_, _22313_);
  and (_22332_, _22331_, _03465_);
  or (_22333_, _22332_, _03458_);
  or (_22334_, _22333_, _22329_);
  or (_22335_, _22313_, _13311_);
  and (_22336_, _22335_, _22316_);
  or (_22337_, _22336_, _03459_);
  and (_22339_, _22337_, _03453_);
  and (_22340_, _22339_, _22334_);
  and (_22341_, _20796_, _05948_);
  or (_22342_, _22341_, _22313_);
  and (_22343_, _22342_, _03452_);
  or (_22344_, _22343_, _07454_);
  or (_22345_, _22344_, _22340_);
  or (_22346_, _22321_, _06903_);
  and (_22347_, _22346_, _22345_);
  or (_22348_, _22347_, _04082_);
  and (_22350_, _06526_, _05289_);
  or (_22351_, _22300_, _04500_);
  or (_22352_, _22351_, _22350_);
  and (_22353_, _22352_, _03521_);
  and (_22354_, _22353_, _22348_);
  and (_22355_, _20822_, _05289_);
  or (_22356_, _22355_, _22300_);
  and (_22357_, _22356_, _03224_);
  or (_22358_, _22357_, _08905_);
  or (_22359_, _22358_, _22354_);
  and (_22361_, _13402_, _05289_);
  or (_22362_, _22300_, _04527_);
  or (_22363_, _22362_, _22361_);
  and (_22364_, _14949_, _05289_);
  or (_22365_, _22364_, _22300_);
  or (_22366_, _22365_, _04509_);
  and (_22367_, _22366_, _03745_);
  and (_22368_, _22367_, _22363_);
  and (_22369_, _22368_, _22359_);
  and (_22370_, _13407_, _05289_);
  or (_22372_, _22370_, _22300_);
  and (_22373_, _22372_, _03744_);
  or (_22374_, _22373_, _22369_);
  and (_22375_, _22374_, _04523_);
  or (_22376_, _22300_, _05469_);
  and (_22377_, _22365_, _03611_);
  and (_22378_, _22377_, _22376_);
  or (_22379_, _22378_, _22375_);
  and (_22380_, _22379_, _03734_);
  and (_22381_, _22306_, _03733_);
  and (_22383_, _22381_, _22376_);
  or (_22384_, _22383_, _03618_);
  or (_22385_, _22384_, _22380_);
  nor (_22386_, _13400_, _09529_);
  or (_22387_, _22300_, _06453_);
  or (_22388_, _22387_, _22386_);
  and (_22389_, _22388_, _06458_);
  and (_22390_, _22389_, _22385_);
  nor (_22391_, _13406_, _09529_);
  or (_22392_, _22391_, _22300_);
  and (_22394_, _22392_, _03741_);
  or (_22395_, _22394_, _03767_);
  or (_22396_, _22395_, _22390_);
  or (_22397_, _22302_, _03948_);
  and (_22398_, _22397_, _03446_);
  and (_22399_, _22398_, _22396_);
  and (_22400_, _22331_, _03445_);
  or (_22401_, _22400_, _03473_);
  or (_22402_, _22401_, _22399_);
  and (_22403_, _13456_, _05289_);
  or (_22405_, _22300_, _03474_);
  or (_22406_, _22405_, _22403_);
  and (_22407_, _22406_, _43189_);
  and (_22408_, _22407_, _22402_);
  or (_43811_, _22408_, _22299_);
  and (_22409_, _09633_, \oc8051_golden_model_1.P3 [0]);
  and (_22410_, _12183_, _05293_);
  or (_22411_, _22410_, _22409_);
  and (_22412_, _22411_, _03744_);
  and (_22413_, _05293_, _04429_);
  or (_22415_, _22413_, _22409_);
  or (_22416_, _22415_, _06903_);
  nor (_22417_, _05722_, _09633_);
  or (_22418_, _22417_, _22409_);
  or (_22419_, _22418_, _04432_);
  and (_22420_, _05293_, \oc8051_golden_model_1.ACC [0]);
  or (_22421_, _22420_, _22409_);
  and (_22422_, _22421_, _04436_);
  and (_22423_, _04437_, \oc8051_golden_model_1.P3 [0]);
  or (_22424_, _22423_, _03534_);
  or (_22426_, _22424_, _22422_);
  and (_22427_, _22426_, _03470_);
  and (_22428_, _22427_, _22419_);
  not (_22429_, _05953_);
  and (_22430_, _22429_, \oc8051_golden_model_1.P3 [0]);
  and (_22431_, _12075_, _05953_);
  or (_22432_, _22431_, _22430_);
  and (_22433_, _22432_, _03469_);
  or (_22434_, _22433_, _22428_);
  and (_22435_, _22434_, _04457_);
  and (_22438_, _22415_, _03527_);
  or (_22439_, _22438_, _03530_);
  or (_22440_, _22439_, _22435_);
  or (_22441_, _22421_, _03531_);
  and (_22442_, _22441_, _03466_);
  and (_22443_, _22442_, _22440_);
  and (_22444_, _22409_, _03465_);
  or (_22445_, _22444_, _03458_);
  or (_22446_, _22445_, _22443_);
  or (_22447_, _22418_, _03459_);
  and (_22449_, _22447_, _03453_);
  and (_22450_, _22449_, _22446_);
  and (_22451_, _20052_, _05953_);
  or (_22452_, _22451_, _22430_);
  and (_22453_, _22452_, _03452_);
  or (_22454_, _22453_, _07454_);
  or (_22455_, _22454_, _22450_);
  and (_22456_, _22455_, _22416_);
  or (_22457_, _22456_, _04082_);
  and (_22458_, _06617_, _05293_);
  or (_22460_, _22409_, _04500_);
  or (_22461_, _22460_, _22458_);
  and (_22462_, _22461_, _03521_);
  and (_22463_, _22462_, _22457_);
  and (_22464_, _20077_, _05293_);
  or (_22465_, _22464_, _22409_);
  and (_22466_, _22465_, _03224_);
  or (_22467_, _22466_, _22463_);
  or (_22468_, _22467_, _08905_);
  and (_22469_, _12177_, _05293_);
  or (_22471_, _22409_, _04527_);
  or (_22472_, _22471_, _22469_);
  and (_22473_, _05293_, _06350_);
  or (_22474_, _22473_, _22409_);
  or (_22475_, _22474_, _04509_);
  and (_22476_, _22475_, _03745_);
  and (_22477_, _22476_, _22472_);
  and (_22478_, _22477_, _22468_);
  or (_22479_, _22478_, _22412_);
  and (_22480_, _22479_, _04523_);
  nand (_22482_, _22474_, _03611_);
  nor (_22483_, _22482_, _22417_);
  or (_22484_, _22483_, _22480_);
  and (_22485_, _22484_, _03734_);
  or (_22486_, _22409_, _05722_);
  and (_22487_, _22421_, _03733_);
  and (_22488_, _22487_, _22486_);
  or (_22489_, _22488_, _03618_);
  or (_22490_, _22489_, _22485_);
  nor (_22491_, _12057_, _09633_);
  or (_22493_, _22409_, _06453_);
  or (_22494_, _22493_, _22491_);
  and (_22495_, _22494_, _06458_);
  and (_22496_, _22495_, _22490_);
  nor (_22497_, _12181_, _09633_);
  or (_22498_, _22497_, _22409_);
  and (_22499_, _22498_, _03741_);
  or (_22500_, _22499_, _03767_);
  or (_22501_, _22500_, _22496_);
  or (_22502_, _22418_, _03948_);
  and (_22504_, _22502_, _03446_);
  and (_22505_, _22504_, _22501_);
  and (_22506_, _22409_, _03445_);
  or (_22507_, _22506_, _03473_);
  or (_22508_, _22507_, _22505_);
  or (_22509_, _22418_, _03474_);
  and (_22510_, _22509_, _43189_);
  and (_22511_, _22510_, _22508_);
  nor (_22512_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_22513_, _22512_, _05173_);
  or (_43812_, _22513_, _22511_);
  and (_22515_, _09633_, \oc8051_golden_model_1.P3 [1]);
  nor (_22516_, _09633_, _04635_);
  or (_22517_, _22516_, _22515_);
  and (_22518_, _22517_, _03527_);
  and (_22519_, _22429_, \oc8051_golden_model_1.P3 [1]);
  and (_22520_, _12269_, _05953_);
  or (_22521_, _22520_, _22519_);
  or (_22522_, _22521_, _03470_);
  or (_22523_, _05293_, \oc8051_golden_model_1.P3 [1]);
  and (_22525_, _12265_, _05293_);
  not (_22526_, _22525_);
  and (_22527_, _22526_, _22523_);
  and (_22528_, _22527_, _03534_);
  nand (_22529_, _05293_, _03269_);
  and (_22530_, _22529_, _22523_);
  and (_22531_, _22530_, _04436_);
  and (_22532_, _04437_, \oc8051_golden_model_1.P3 [1]);
  or (_22533_, _22532_, _22531_);
  and (_22534_, _22533_, _04432_);
  or (_22536_, _22534_, _03469_);
  or (_22537_, _22536_, _22528_);
  and (_22538_, _22537_, _22522_);
  and (_22539_, _22538_, _04457_);
  or (_22540_, _22539_, _22518_);
  or (_22541_, _22540_, _03530_);
  or (_22542_, _22530_, _03531_);
  and (_22543_, _22542_, _03466_);
  and (_22544_, _22543_, _22541_);
  and (_22545_, _12256_, _05953_);
  or (_22547_, _22545_, _22519_);
  and (_22548_, _22547_, _03465_);
  or (_22549_, _22548_, _03458_);
  or (_22550_, _22549_, _22544_);
  or (_22551_, _22519_, _12284_);
  and (_22552_, _22551_, _22521_);
  or (_22553_, _22552_, _03459_);
  and (_22554_, _22553_, _03453_);
  and (_22555_, _22554_, _22550_);
  and (_22556_, _20170_, _05953_);
  or (_22558_, _22556_, _22519_);
  and (_22559_, _22558_, _03452_);
  or (_22560_, _22559_, _07454_);
  or (_22561_, _22560_, _22555_);
  or (_22562_, _22517_, _06903_);
  and (_22563_, _22562_, _22561_);
  or (_22564_, _22563_, _04082_);
  and (_22565_, _06572_, _05293_);
  or (_22566_, _22515_, _04500_);
  or (_22567_, _22566_, _22565_);
  and (_22569_, _22567_, _03521_);
  and (_22570_, _22569_, _22564_);
  and (_22571_, _20196_, _05293_);
  or (_22572_, _22571_, _22515_);
  and (_22573_, _22572_, _03224_);
  or (_22574_, _22573_, _22570_);
  and (_22575_, _22574_, _03625_);
  or (_22576_, _12375_, _09633_);
  and (_22577_, _22576_, _03623_);
  nand (_22578_, _05293_, _04325_);
  and (_22580_, _22578_, _03624_);
  or (_22581_, _22580_, _22577_);
  and (_22582_, _22581_, _22523_);
  or (_22583_, _22582_, _22575_);
  and (_22584_, _22583_, _03745_);
  or (_22585_, _12381_, _09633_);
  and (_22586_, _22523_, _03744_);
  and (_22587_, _22586_, _22585_);
  or (_22588_, _22587_, _22584_);
  and (_22589_, _22588_, _04523_);
  or (_22591_, _12374_, _09633_);
  and (_22592_, _22523_, _03611_);
  and (_22593_, _22592_, _22591_);
  or (_22594_, _22593_, _22589_);
  and (_22595_, _22594_, _03734_);
  or (_22596_, _22515_, _05674_);
  and (_22597_, _22530_, _03733_);
  and (_22598_, _22597_, _22596_);
  or (_22599_, _22598_, _22595_);
  and (_22600_, _22599_, _03742_);
  or (_22602_, _22578_, _05674_);
  and (_22603_, _22523_, _03618_);
  and (_22604_, _22603_, _22602_);
  or (_22605_, _22529_, _05674_);
  and (_22606_, _22523_, _03741_);
  and (_22607_, _22606_, _22605_);
  or (_22608_, _22607_, _03767_);
  or (_22609_, _22608_, _22604_);
  or (_22610_, _22609_, _22600_);
  or (_22611_, _22527_, _03948_);
  and (_22613_, _22611_, _03446_);
  and (_22614_, _22613_, _22610_);
  and (_22615_, _22547_, _03445_);
  or (_22616_, _22615_, _03473_);
  or (_22617_, _22616_, _22614_);
  or (_22618_, _22515_, _03474_);
  or (_22619_, _22618_, _22525_);
  and (_22620_, _22619_, _43189_);
  and (_22621_, _22620_, _22617_);
  nor (_22622_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_22624_, _22622_, _05173_);
  or (_43813_, _22624_, _22621_);
  not (_22625_, \oc8051_golden_model_1.P3 [2]);
  nor (_22626_, _05293_, _22625_);
  nor (_22627_, _09633_, _05073_);
  or (_22628_, _22627_, _22626_);
  or (_22629_, _22628_, _06903_);
  or (_22630_, _22628_, _04457_);
  nor (_22631_, _12467_, _09633_);
  or (_22632_, _22631_, _22626_);
  or (_22634_, _22632_, _04432_);
  and (_22635_, _05293_, \oc8051_golden_model_1.ACC [2]);
  or (_22636_, _22635_, _22626_);
  and (_22637_, _22636_, _04436_);
  nor (_22638_, _04436_, _22625_);
  or (_22639_, _22638_, _03534_);
  or (_22640_, _22639_, _22637_);
  and (_22641_, _22640_, _03470_);
  and (_22642_, _22641_, _22634_);
  nor (_22643_, _05953_, _22625_);
  and (_22645_, _12462_, _05953_);
  or (_22646_, _22645_, _22643_);
  and (_22647_, _22646_, _03469_);
  or (_22648_, _22647_, _03527_);
  or (_22649_, _22648_, _22642_);
  and (_22650_, _22649_, _22630_);
  or (_22651_, _22650_, _03530_);
  or (_22652_, _22636_, _03531_);
  and (_22653_, _22652_, _03466_);
  and (_22654_, _22653_, _22651_);
  and (_22656_, _12460_, _05953_);
  or (_22657_, _22656_, _22643_);
  and (_22658_, _22657_, _03465_);
  or (_22659_, _22658_, _03458_);
  or (_22660_, _22659_, _22654_);
  and (_22661_, _22645_, _12491_);
  or (_22662_, _22643_, _03459_);
  or (_22663_, _22662_, _22661_);
  and (_22664_, _22663_, _03453_);
  and (_22665_, _22664_, _22660_);
  and (_22667_, _20293_, _05953_);
  or (_22668_, _22667_, _22643_);
  and (_22669_, _22668_, _03452_);
  or (_22670_, _22669_, _07454_);
  or (_22671_, _22670_, _22665_);
  and (_22672_, _22671_, _22629_);
  or (_22673_, _22672_, _04082_);
  and (_22674_, _06710_, _05293_);
  or (_22675_, _22626_, _04500_);
  or (_22676_, _22675_, _22674_);
  and (_22678_, _22676_, _03521_);
  and (_22679_, _22678_, _22673_);
  and (_22680_, _20318_, _05293_);
  or (_22681_, _22626_, _22680_);
  and (_22682_, _22681_, _03224_);
  or (_22683_, _22682_, _22679_);
  or (_22684_, _22683_, _08905_);
  and (_22685_, _12582_, _05293_);
  or (_22686_, _22626_, _04527_);
  or (_22687_, _22686_, _22685_);
  and (_22689_, _05293_, _06399_);
  or (_22690_, _22689_, _22626_);
  or (_22691_, _22690_, _04509_);
  and (_22692_, _22691_, _03745_);
  and (_22693_, _22692_, _22687_);
  and (_22694_, _22693_, _22684_);
  and (_22695_, _12588_, _05293_);
  or (_22696_, _22695_, _22626_);
  and (_22697_, _22696_, _03744_);
  or (_22698_, _22697_, _22694_);
  and (_22700_, _22698_, _04523_);
  or (_22701_, _22626_, _05772_);
  and (_22702_, _22690_, _03611_);
  and (_22703_, _22702_, _22701_);
  or (_22704_, _22703_, _22700_);
  and (_22705_, _22704_, _03734_);
  and (_22706_, _22636_, _03733_);
  and (_22707_, _22706_, _22701_);
  or (_22708_, _22707_, _03618_);
  or (_22709_, _22708_, _22705_);
  nor (_22711_, _12581_, _09633_);
  or (_22712_, _22626_, _06453_);
  or (_22713_, _22712_, _22711_);
  and (_22714_, _22713_, _06458_);
  and (_22715_, _22714_, _22709_);
  nor (_22716_, _12587_, _09633_);
  or (_22717_, _22716_, _22626_);
  and (_22718_, _22717_, _03741_);
  or (_22719_, _22718_, _03767_);
  or (_22720_, _22719_, _22715_);
  or (_22722_, _22632_, _03948_);
  and (_22723_, _22722_, _03446_);
  and (_22724_, _22723_, _22720_);
  and (_22725_, _22657_, _03445_);
  or (_22726_, _22725_, _03473_);
  or (_22727_, _22726_, _22724_);
  and (_22728_, _12638_, _05293_);
  or (_22729_, _22626_, _03474_);
  or (_22730_, _22729_, _22728_);
  and (_22731_, _22730_, _43189_);
  and (_22733_, _22731_, _22727_);
  nor (_22734_, _43189_, _22625_);
  or (_22735_, _22734_, rst);
  or (_43814_, _22735_, _22733_);
  and (_22736_, _09633_, \oc8051_golden_model_1.P3 [3]);
  nor (_22737_, _09633_, _04885_);
  or (_22738_, _22737_, _22736_);
  or (_22739_, _22738_, _06903_);
  nor (_22740_, _12652_, _09633_);
  or (_22741_, _22740_, _22736_);
  or (_22743_, _22741_, _04432_);
  and (_22744_, _05293_, \oc8051_golden_model_1.ACC [3]);
  or (_22745_, _22744_, _22736_);
  and (_22746_, _22745_, _04436_);
  and (_22747_, _04437_, \oc8051_golden_model_1.P3 [3]);
  or (_22748_, _22747_, _03534_);
  or (_22749_, _22748_, _22746_);
  and (_22750_, _22749_, _03470_);
  and (_22751_, _22750_, _22743_);
  and (_22752_, _22429_, \oc8051_golden_model_1.P3 [3]);
  and (_22754_, _12664_, _05953_);
  or (_22755_, _22754_, _22752_);
  and (_22756_, _22755_, _03469_);
  or (_22757_, _22756_, _03527_);
  or (_22758_, _22757_, _22751_);
  or (_22759_, _22738_, _04457_);
  and (_22760_, _22759_, _22758_);
  or (_22761_, _22760_, _03530_);
  or (_22762_, _22745_, _03531_);
  and (_22763_, _22762_, _03466_);
  and (_22765_, _22763_, _22761_);
  and (_22766_, _12662_, _05953_);
  or (_22767_, _22766_, _22752_);
  and (_22768_, _22767_, _03465_);
  or (_22769_, _22768_, _03458_);
  or (_22770_, _22769_, _22765_);
  or (_22771_, _22752_, _12691_);
  and (_22772_, _22771_, _22755_);
  or (_22773_, _22772_, _03459_);
  and (_22774_, _22773_, _03453_);
  and (_22776_, _22774_, _22770_);
  and (_22777_, _20419_, _05953_);
  or (_22778_, _22777_, _22752_);
  and (_22779_, _22778_, _03452_);
  or (_22780_, _22779_, _07454_);
  or (_22781_, _22780_, _22776_);
  and (_22782_, _22781_, _22739_);
  or (_22783_, _22782_, _04082_);
  and (_22784_, _06664_, _05293_);
  or (_22785_, _22736_, _04500_);
  or (_22787_, _22785_, _22784_);
  and (_22788_, _22787_, _03521_);
  and (_22789_, _22788_, _22783_);
  and (_22790_, _20454_, _05293_);
  or (_22791_, _22736_, _22790_);
  and (_22792_, _22791_, _03224_);
  or (_22793_, _22792_, _22789_);
  or (_22794_, _22793_, _08905_);
  and (_22795_, _12787_, _05293_);
  or (_22796_, _22736_, _04527_);
  or (_22798_, _22796_, _22795_);
  and (_22799_, _05293_, _06356_);
  or (_22800_, _22799_, _22736_);
  or (_22801_, _22800_, _04509_);
  and (_22802_, _22801_, _03745_);
  and (_22803_, _22802_, _22798_);
  and (_22804_, _22803_, _22794_);
  and (_22805_, _12793_, _05293_);
  or (_22806_, _22805_, _22736_);
  and (_22807_, _22806_, _03744_);
  or (_22809_, _22807_, _22804_);
  and (_22810_, _22809_, _04523_);
  or (_22811_, _22736_, _05625_);
  and (_22812_, _22800_, _03611_);
  and (_22813_, _22812_, _22811_);
  or (_22814_, _22813_, _22810_);
  and (_22815_, _22814_, _03734_);
  and (_22816_, _22745_, _03733_);
  and (_22817_, _22816_, _22811_);
  or (_22818_, _22817_, _03618_);
  or (_22820_, _22818_, _22815_);
  nor (_22821_, _12786_, _09633_);
  or (_22822_, _22736_, _06453_);
  or (_22823_, _22822_, _22821_);
  and (_22824_, _22823_, _06458_);
  and (_22825_, _22824_, _22820_);
  nor (_22826_, _12792_, _09633_);
  or (_22827_, _22826_, _22736_);
  and (_22828_, _22827_, _03741_);
  or (_22829_, _22828_, _03767_);
  or (_22831_, _22829_, _22825_);
  or (_22832_, _22741_, _03948_);
  and (_22833_, _22832_, _03446_);
  and (_22834_, _22833_, _22831_);
  and (_22835_, _22767_, _03445_);
  or (_22836_, _22835_, _03473_);
  or (_22837_, _22836_, _22834_);
  and (_22838_, _12843_, _05293_);
  or (_22839_, _22736_, _03474_);
  or (_22840_, _22839_, _22838_);
  and (_22842_, _22840_, _43189_);
  and (_22843_, _22842_, _22837_);
  nor (_22844_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_22845_, _22844_, _05173_);
  or (_43815_, _22845_, _22843_);
  and (_22846_, _09633_, \oc8051_golden_model_1.P3 [4]);
  nor (_22847_, _05831_, _09633_);
  or (_22848_, _22847_, _22846_);
  or (_22849_, _22848_, _06903_);
  and (_22850_, _22429_, \oc8051_golden_model_1.P3 [4]);
  and (_22852_, _12864_, _05953_);
  or (_22853_, _22852_, _22850_);
  and (_22854_, _22853_, _03465_);
  nor (_22855_, _12856_, _09633_);
  or (_22856_, _22855_, _22846_);
  or (_22857_, _22856_, _04432_);
  and (_22858_, _05293_, \oc8051_golden_model_1.ACC [4]);
  or (_22859_, _22858_, _22846_);
  and (_22860_, _22859_, _04436_);
  and (_22861_, _04437_, \oc8051_golden_model_1.P3 [4]);
  or (_22863_, _22861_, _03534_);
  or (_22864_, _22863_, _22860_);
  and (_22865_, _22864_, _03470_);
  and (_22866_, _22865_, _22857_);
  and (_22867_, _12866_, _05953_);
  or (_22868_, _22867_, _22850_);
  and (_22869_, _22868_, _03469_);
  or (_22870_, _22869_, _03527_);
  or (_22871_, _22870_, _22866_);
  or (_22872_, _22848_, _04457_);
  and (_22874_, _22872_, _22871_);
  or (_22875_, _22874_, _03530_);
  or (_22876_, _22859_, _03531_);
  and (_22877_, _22876_, _03466_);
  and (_22878_, _22877_, _22875_);
  or (_22879_, _22878_, _22854_);
  and (_22880_, _22879_, _03459_);
  or (_22881_, _22850_, _12894_);
  and (_22882_, _22881_, _03458_);
  and (_22883_, _22882_, _22868_);
  or (_22885_, _22883_, _22880_);
  and (_22886_, _22885_, _03453_);
  and (_22887_, _20548_, _05953_);
  or (_22888_, _22887_, _22850_);
  and (_22889_, _22888_, _03452_);
  or (_22890_, _22889_, _07454_);
  or (_22891_, _22890_, _22886_);
  and (_22892_, _22891_, _22849_);
  or (_22893_, _22892_, _04082_);
  and (_22894_, _06802_, _05293_);
  or (_22896_, _22846_, _04500_);
  or (_22897_, _22896_, _22894_);
  and (_22898_, _22897_, _03521_);
  and (_22899_, _22898_, _22893_);
  and (_22900_, _20573_, _05293_);
  or (_22901_, _22900_, _22846_);
  and (_22902_, _22901_, _03224_);
  or (_22903_, _22902_, _08905_);
  or (_22904_, _22903_, _22899_);
  and (_22905_, _12986_, _05293_);
  or (_22907_, _22846_, _04527_);
  or (_22908_, _22907_, _22905_);
  and (_22909_, _06337_, _05293_);
  or (_22910_, _22909_, _22846_);
  or (_22911_, _22910_, _04509_);
  and (_22912_, _22911_, _03745_);
  and (_22913_, _22912_, _22908_);
  and (_22914_, _22913_, _22904_);
  and (_22915_, _12992_, _05293_);
  or (_22916_, _22915_, _22846_);
  and (_22918_, _22916_, _03744_);
  or (_22919_, _22918_, _22914_);
  and (_22920_, _22919_, _04523_);
  or (_22921_, _22846_, _05880_);
  and (_22922_, _22910_, _03611_);
  and (_22923_, _22922_, _22921_);
  or (_22924_, _22923_, _22920_);
  and (_22925_, _22924_, _03734_);
  and (_22926_, _22859_, _03733_);
  and (_22927_, _22926_, _22921_);
  or (_22929_, _22927_, _03618_);
  or (_22930_, _22929_, _22925_);
  nor (_22931_, _12985_, _09633_);
  or (_22932_, _22846_, _06453_);
  or (_22933_, _22932_, _22931_);
  and (_22934_, _22933_, _06458_);
  and (_22935_, _22934_, _22930_);
  nor (_22936_, _12991_, _09633_);
  or (_22937_, _22936_, _22846_);
  and (_22938_, _22937_, _03741_);
  or (_22940_, _22938_, _03767_);
  or (_22941_, _22940_, _22935_);
  or (_22942_, _22856_, _03948_);
  and (_22943_, _22942_, _03446_);
  and (_22944_, _22943_, _22941_);
  and (_22945_, _22853_, _03445_);
  or (_22946_, _22945_, _03473_);
  or (_22947_, _22946_, _22944_);
  and (_22948_, _13051_, _05293_);
  or (_22949_, _22846_, _03474_);
  or (_22951_, _22949_, _22948_);
  and (_22952_, _22951_, _43189_);
  and (_22953_, _22952_, _22947_);
  nor (_22954_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_22955_, _22954_, _05173_);
  or (_43816_, _22955_, _22953_);
  nor (_22956_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_22957_, _22956_, _05173_);
  and (_22958_, _09633_, \oc8051_golden_model_1.P3 [5]);
  nor (_22959_, _13070_, _09633_);
  or (_22961_, _22959_, _22958_);
  or (_22962_, _22961_, _04432_);
  and (_22963_, _05293_, \oc8051_golden_model_1.ACC [5]);
  or (_22964_, _22963_, _22958_);
  and (_22965_, _22964_, _04436_);
  and (_22966_, _04437_, \oc8051_golden_model_1.P3 [5]);
  or (_22967_, _22966_, _03534_);
  or (_22968_, _22967_, _22965_);
  and (_22969_, _22968_, _03470_);
  and (_22970_, _22969_, _22962_);
  and (_22972_, _22429_, \oc8051_golden_model_1.P3 [5]);
  and (_22973_, _13095_, _05953_);
  or (_22974_, _22973_, _22972_);
  and (_22975_, _22974_, _03469_);
  or (_22976_, _22975_, _03527_);
  or (_22977_, _22976_, _22970_);
  nor (_22978_, _05526_, _09633_);
  or (_22979_, _22978_, _22958_);
  or (_22980_, _22979_, _04457_);
  and (_22981_, _22980_, _22977_);
  or (_22983_, _22981_, _03530_);
  or (_22984_, _22964_, _03531_);
  and (_22985_, _22984_, _03466_);
  and (_22986_, _22985_, _22983_);
  and (_22987_, _13078_, _05953_);
  or (_22988_, _22987_, _22972_);
  and (_22989_, _22988_, _03465_);
  or (_22990_, _22989_, _03458_);
  or (_22991_, _22990_, _22986_);
  or (_22992_, _22972_, _13110_);
  and (_22993_, _22992_, _22974_);
  or (_22994_, _22993_, _03459_);
  and (_22995_, _22994_, _03453_);
  and (_22996_, _22995_, _22991_);
  and (_22997_, _20670_, _05953_);
  or (_22998_, _22997_, _22972_);
  and (_22999_, _22998_, _03452_);
  or (_23000_, _22999_, _07454_);
  or (_23001_, _23000_, _22996_);
  or (_23002_, _22979_, _06903_);
  and (_23005_, _23002_, _23001_);
  or (_23006_, _23005_, _04082_);
  and (_23007_, _06757_, _05293_);
  or (_23008_, _22958_, _04500_);
  or (_23009_, _23008_, _23007_);
  and (_23010_, _23009_, _03521_);
  and (_23011_, _23010_, _23006_);
  and (_23012_, _20704_, _05293_);
  or (_23013_, _23012_, _22958_);
  and (_23014_, _23013_, _03224_);
  or (_23016_, _23014_, _08905_);
  or (_23017_, _23016_, _23011_);
  and (_23018_, _13198_, _05293_);
  or (_23019_, _22958_, _04527_);
  or (_23020_, _23019_, _23018_);
  and (_23021_, _06295_, _05293_);
  or (_23022_, _23021_, _22958_);
  or (_23023_, _23022_, _04509_);
  and (_23024_, _23023_, _03745_);
  and (_23025_, _23024_, _23020_);
  and (_23026_, _23025_, _23017_);
  and (_23027_, _13204_, _05293_);
  or (_23028_, _23027_, _22958_);
  and (_23029_, _23028_, _03744_);
  or (_23030_, _23029_, _23026_);
  and (_23031_, _23030_, _04523_);
  or (_23032_, _22958_, _05576_);
  and (_23033_, _23022_, _03611_);
  and (_23034_, _23033_, _23032_);
  or (_23035_, _23034_, _23031_);
  and (_23038_, _23035_, _03734_);
  and (_23039_, _22964_, _03733_);
  and (_23040_, _23039_, _23032_);
  or (_23041_, _23040_, _03618_);
  or (_23042_, _23041_, _23038_);
  nor (_23043_, _13197_, _09633_);
  or (_23044_, _22958_, _06453_);
  or (_23045_, _23044_, _23043_);
  and (_23046_, _23045_, _06458_);
  and (_23047_, _23046_, _23042_);
  nor (_23049_, _13203_, _09633_);
  or (_23050_, _23049_, _22958_);
  and (_23051_, _23050_, _03741_);
  or (_23052_, _23051_, _03767_);
  or (_23053_, _23052_, _23047_);
  or (_23054_, _22961_, _03948_);
  and (_23055_, _23054_, _03446_);
  and (_23056_, _23055_, _23053_);
  and (_23057_, _22988_, _03445_);
  or (_23058_, _23057_, _03473_);
  or (_23059_, _23058_, _23056_);
  and (_23060_, _13253_, _05293_);
  or (_23061_, _22958_, _03474_);
  or (_23062_, _23061_, _23060_);
  and (_23063_, _23062_, _43189_);
  and (_23064_, _23063_, _23059_);
  or (_43817_, _23064_, _22957_);
  and (_23065_, _09633_, \oc8051_golden_model_1.P3 [6]);
  nor (_23066_, _13293_, _09633_);
  or (_23067_, _23066_, _23065_);
  or (_23070_, _23067_, _04432_);
  and (_23071_, _05293_, \oc8051_golden_model_1.ACC [6]);
  or (_23072_, _23071_, _23065_);
  and (_23073_, _23072_, _04436_);
  and (_23074_, _04437_, \oc8051_golden_model_1.P3 [6]);
  or (_23075_, _23074_, _03534_);
  or (_23076_, _23075_, _23073_);
  and (_23077_, _23076_, _03470_);
  and (_23078_, _23077_, _23070_);
  and (_23079_, _22429_, \oc8051_golden_model_1.P3 [6]);
  and (_23081_, _13280_, _05953_);
  or (_23082_, _23081_, _23079_);
  and (_23083_, _23082_, _03469_);
  or (_23084_, _23083_, _03527_);
  or (_23085_, _23084_, _23078_);
  nor (_23086_, _05417_, _09633_);
  or (_23087_, _23086_, _23065_);
  or (_23088_, _23087_, _04457_);
  and (_23089_, _23088_, _23085_);
  or (_23090_, _23089_, _03530_);
  or (_23091_, _23072_, _03531_);
  and (_23092_, _23091_, _03466_);
  and (_23093_, _23092_, _23090_);
  and (_23094_, _13304_, _05953_);
  or (_23095_, _23094_, _23079_);
  and (_23096_, _23095_, _03465_);
  or (_23097_, _23096_, _03458_);
  or (_23098_, _23097_, _23093_);
  or (_23099_, _23079_, _13311_);
  and (_23100_, _23099_, _23082_);
  or (_23103_, _23100_, _03459_);
  and (_23104_, _23103_, _03453_);
  and (_23105_, _23104_, _23098_);
  and (_23106_, _20796_, _05953_);
  or (_23107_, _23106_, _23079_);
  and (_23108_, _23107_, _03452_);
  or (_23109_, _23108_, _07454_);
  or (_23110_, _23109_, _23105_);
  or (_23111_, _23087_, _06903_);
  and (_23112_, _23111_, _23110_);
  or (_23114_, _23112_, _04082_);
  and (_23115_, _06526_, _05293_);
  or (_23116_, _23065_, _04500_);
  or (_23117_, _23116_, _23115_);
  and (_23118_, _23117_, _03521_);
  and (_23119_, _23118_, _23114_);
  and (_23120_, _20822_, _05293_);
  or (_23121_, _23120_, _23065_);
  and (_23122_, _23121_, _03224_);
  or (_23123_, _23122_, _08905_);
  or (_23124_, _23123_, _23119_);
  and (_23125_, _13402_, _05293_);
  or (_23126_, _23065_, _04527_);
  or (_23127_, _23126_, _23125_);
  and (_23128_, _14949_, _05293_);
  or (_23129_, _23128_, _23065_);
  or (_23130_, _23129_, _04509_);
  and (_23131_, _23130_, _03745_);
  and (_23132_, _23131_, _23127_);
  and (_23133_, _23132_, _23124_);
  and (_23136_, _13407_, _05293_);
  or (_23137_, _23136_, _23065_);
  and (_23138_, _23137_, _03744_);
  or (_23139_, _23138_, _23133_);
  and (_23140_, _23139_, _04523_);
  or (_23141_, _23065_, _05469_);
  and (_23142_, _23129_, _03611_);
  and (_23143_, _23142_, _23141_);
  or (_23144_, _23143_, _23140_);
  and (_23145_, _23144_, _03734_);
  and (_23147_, _23072_, _03733_);
  and (_23148_, _23147_, _23141_);
  or (_23149_, _23148_, _03618_);
  or (_23150_, _23149_, _23145_);
  nor (_23151_, _13400_, _09633_);
  or (_23152_, _23065_, _06453_);
  or (_23153_, _23152_, _23151_);
  and (_23154_, _23153_, _06458_);
  and (_23155_, _23154_, _23150_);
  nor (_23156_, _13406_, _09633_);
  or (_23157_, _23156_, _23065_);
  and (_23158_, _23157_, _03741_);
  or (_23159_, _23158_, _03767_);
  or (_23160_, _23159_, _23155_);
  or (_23161_, _23067_, _03948_);
  and (_23162_, _23161_, _03446_);
  and (_23163_, _23162_, _23160_);
  and (_23164_, _23095_, _03445_);
  or (_23165_, _23164_, _03473_);
  or (_23166_, _23165_, _23163_);
  and (_23169_, _13456_, _05293_);
  or (_23170_, _23065_, _03474_);
  or (_23171_, _23170_, _23169_);
  and (_23172_, _23171_, _43189_);
  and (_23173_, _23172_, _23166_);
  nor (_23174_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_23175_, _23174_, _05173_);
  or (_43820_, _23175_, _23173_);
  not (_23176_, \oc8051_golden_model_1.PSW [0]);
  nor (_23177_, _43189_, _23176_);
  nor (_23179_, _07591_, _07590_);
  nor (_23180_, _23179_, _07495_);
  and (_23181_, _23179_, _07495_);
  nor (_23182_, _23181_, _23180_);
  nor (_23183_, _07511_, _07510_);
  nor (_23184_, _23183_, _15458_);
  and (_23185_, _23183_, _15458_);
  nor (_23186_, _23185_, _23184_);
  and (_23187_, _23186_, _23182_);
  nor (_23188_, _23186_, _23182_);
  nor (_23189_, _23188_, _23187_);
  nor (_23190_, _23189_, _06440_);
  and (_23191_, _23189_, _06440_);
  nor (_23192_, _23191_, _23190_);
  not (_23193_, _11989_);
  and (_23194_, _03188_, _03442_);
  nor (_23195_, _23194_, _23193_);
  or (_23196_, _23195_, _23192_);
  and (_23197_, _11815_, _05915_);
  or (_23198_, _23197_, _23192_);
  and (_23201_, _15232_, _15014_);
  nor (_23202_, _15232_, _15014_);
  nor (_23203_, _23202_, _23201_);
  and (_23204_, _23203_, _15489_);
  nor (_23205_, _23203_, _15489_);
  or (_23206_, _23205_, _23204_);
  and (_23207_, _23206_, _15833_);
  nor (_23208_, _23206_, _15833_);
  or (_23209_, _23208_, _23207_);
  not (_23210_, _16818_);
  nor (_23212_, _16489_, _16167_);
  and (_23213_, _16489_, _16167_);
  nor (_23214_, _23213_, _23212_);
  nor (_23215_, _23214_, _23210_);
  and (_23216_, _23214_, _23210_);
  nor (_23217_, _23216_, _23215_);
  nor (_23218_, _23217_, _23209_);
  and (_23219_, _23217_, _23209_);
  nor (_23220_, _23219_, _23218_);
  and (_23221_, _23220_, _07938_);
  nor (_23223_, _23220_, _07938_);
  or (_23224_, _23223_, _23221_);
  and (_23225_, _23224_, _07454_);
  or (_23226_, _23225_, _04082_);
  nor (_23227_, _15240_, _15070_);
  and (_23228_, _15240_, _15070_);
  nor (_23229_, _23228_, _23227_);
  or (_23230_, _23229_, _15860_);
  nand (_23231_, _23229_, _15860_);
  and (_23232_, _23231_, _23230_);
  or (_23234_, _23232_, _15582_);
  nand (_23235_, _23232_, _15582_);
  and (_23236_, _23235_, _23234_);
  nor (_23237_, _23236_, _16183_);
  and (_23238_, _23236_, _16183_);
  nor (_23239_, _23238_, _23237_);
  or (_23240_, _23239_, _16602_);
  nand (_23241_, _23239_, _16602_);
  and (_23242_, _23241_, _23240_);
  and (_23243_, _23242_, _16903_);
  nor (_23245_, _23242_, _16903_);
  nor (_23246_, _23245_, _23243_);
  nor (_23247_, _23246_, _08260_);
  and (_23248_, _23246_, _08260_);
  or (_23249_, _23248_, _23247_);
  or (_23250_, _23249_, _08191_);
  nor (_23251_, _15294_, _15001_);
  and (_23252_, _15294_, _15001_);
  nor (_23253_, _23252_, _23251_);
  not (_23254_, _15919_);
  and (_23256_, _23254_, _15554_);
  nor (_23257_, _23254_, _15554_);
  nor (_23258_, _23257_, _23256_);
  and (_23259_, _23258_, _23253_);
  nor (_23260_, _23258_, _23253_);
  or (_23261_, _23260_, _23259_);
  nor (_23262_, _16577_, _16235_);
  and (_23263_, _16577_, _16235_);
  nor (_23264_, _23263_, _23262_);
  and (_23265_, _23264_, _16875_);
  nor (_23267_, _23264_, _16875_);
  nor (_23268_, _23267_, _23265_);
  and (_23269_, _23268_, _23261_);
  nor (_23270_, _23268_, _23261_);
  or (_23271_, _23270_, _23269_);
  or (_23272_, _23271_, _08172_);
  nand (_23273_, _23271_, _08172_);
  and (_23274_, _23273_, _23272_);
  and (_23275_, _23274_, _03465_);
  nor (_23276_, _08334_, _08287_);
  and (_23278_, _08334_, _08287_);
  nor (_23279_, _23278_, _23276_);
  nor (_23280_, _23279_, _08632_);
  and (_23281_, _23279_, _08632_);
  nor (_23282_, _23281_, _23280_);
  nor (_23283_, _08380_, _08634_);
  and (_23284_, _08380_, _08634_);
  nor (_23285_, _23284_, _23283_);
  and (_23286_, _08364_, _08305_);
  nor (_23287_, _08364_, _08305_);
  or (_23289_, _23287_, _23286_);
  and (_23290_, _23289_, _23285_);
  nor (_23291_, _23289_, _23285_);
  or (_23292_, _23291_, _23290_);
  nor (_23293_, _23292_, _23282_);
  and (_23294_, _23292_, _23282_);
  nor (_23295_, _23294_, _23293_);
  nor (_23296_, _23295_, _10288_);
  and (_23297_, _23295_, _10288_);
  or (_23298_, _23297_, _23296_);
  and (_23300_, _23298_, _03536_);
  nor (_23301_, _06840_, _06711_);
  not (_23302_, _23301_);
  nand (_23303_, _23302_, _12411_);
  or (_23304_, _23302_, _12411_);
  and (_23305_, _23304_, _23303_);
  nor (_23306_, _06842_, _06803_);
  nand (_23307_, _23306_, _06527_);
  or (_23308_, _23306_, _06527_);
  and (_23309_, _23308_, _23307_);
  and (_23311_, _23309_, _23305_);
  nor (_23312_, _23309_, _23305_);
  or (_23313_, _23312_, _23311_);
  nor (_23314_, _23313_, _06114_);
  and (_23315_, _23313_, _06114_);
  or (_23316_, _23315_, _23314_);
  or (_23317_, _23316_, _08103_);
  and (_23318_, _05897_, _05526_);
  nor (_23319_, _05897_, _05526_);
  nor (_23320_, _23319_, _23318_);
  nor (_23322_, _05985_, _05891_);
  not (_23323_, _23322_);
  nor (_23324_, _12251_, _05889_);
  and (_23325_, _12251_, _05889_);
  nor (_23326_, _23325_, _23324_);
  and (_23327_, _23326_, _23323_);
  nor (_23328_, _23326_, _23323_);
  nor (_23329_, _23328_, _23327_);
  or (_23330_, _23329_, _23320_);
  nand (_23331_, _23329_, _23320_);
  and (_23333_, _23331_, _23330_);
  and (_23334_, _23333_, _08105_);
  and (_23335_, _11683_, _10754_);
  or (_23336_, _23335_, _23192_);
  nand (_23337_, _23335_, _23176_);
  and (_23338_, _23337_, _23336_);
  or (_23339_, _23338_, _04007_);
  and (_23340_, _23339_, _08106_);
  or (_23341_, _23340_, _23334_);
  and (_23342_, _23341_, _08101_);
  and (_23344_, _23342_, _23317_);
  or (_23345_, _23344_, _23300_);
  and (_23346_, _05997_, _03209_);
  and (_23347_, _23346_, _11686_);
  and (_23348_, _23347_, _23345_);
  not (_23349_, _23192_);
  nor (_23350_, _23346_, _23349_);
  or (_23351_, _23350_, _04012_);
  or (_23352_, _23351_, _23348_);
  nor (_23353_, _23183_, \oc8051_golden_model_1.ACC [6]);
  and (_23355_, _23183_, \oc8051_golden_model_1.ACC [6]);
  nor (_23356_, _23355_, _23353_);
  nor (_23357_, _23356_, \oc8051_golden_model_1.ACC [7]);
  and (_23358_, _23356_, \oc8051_golden_model_1.ACC [7]);
  nor (_23359_, _23358_, _23357_);
  and (_23360_, _23359_, _23305_);
  nor (_23361_, _23359_, _23305_);
  or (_23362_, _23361_, _23360_);
  or (_23363_, _23362_, _06008_);
  and (_23364_, _23363_, _04432_);
  and (_23366_, _23364_, _23352_);
  not (_23367_, _16841_);
  not (_23368_, _15035_);
  nor (_23369_, _15265_, _23368_);
  and (_23370_, _15265_, _23368_);
  nor (_23371_, _23370_, _23369_);
  and (_23372_, _23371_, _15522_);
  nor (_23373_, _23371_, _15522_);
  nor (_23374_, _23373_, _23372_);
  and (_23375_, _23374_, _16545_);
  nor (_23377_, _23374_, _16545_);
  or (_23378_, _23377_, _23375_);
  nor (_23379_, _16202_, _15885_);
  and (_23380_, _16202_, _15885_);
  nor (_23381_, _23380_, _23379_);
  and (_23382_, _23381_, _23378_);
  nor (_23383_, _23381_, _23378_);
  nor (_23384_, _23383_, _23382_);
  nor (_23385_, _23384_, _23367_);
  and (_23386_, _23384_, _23367_);
  or (_23388_, _23386_, _23385_);
  and (_23389_, _23388_, _08123_);
  nor (_23390_, _23388_, _08123_);
  or (_23391_, _23390_, _23389_);
  and (_23392_, _23391_, _03534_);
  or (_23393_, _23392_, _08121_);
  or (_23394_, _23393_, _23366_);
  and (_23395_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_23396_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_23397_, _23396_, _23395_);
  and (_23398_, _23397_, _15271_);
  nor (_23399_, _23397_, _15271_);
  nor (_23400_, _23399_, _23398_);
  and (_23401_, _16209_, _15893_);
  and (_23402_, _16208_, _15894_);
  nor (_23403_, _23402_, _23401_);
  nor (_23404_, _23403_, _23400_);
  and (_23405_, _23403_, _23400_);
  or (_23406_, _23405_, _23404_);
  nor (_23407_, _23406_, _16552_);
  and (_23409_, _23406_, _16552_);
  or (_23410_, _23409_, _23407_);
  nor (_23411_, _16849_, _08146_);
  and (_23412_, _16849_, _08146_);
  nor (_23413_, _23412_, _23411_);
  nor (_23414_, _23413_, _23410_);
  and (_23415_, _23413_, _23410_);
  nor (_23416_, _23415_, _23414_);
  nand (_23417_, _23416_, _08121_);
  and (_23418_, _23417_, _23394_);
  or (_23420_, _23418_, _09994_);
  nand (_23421_, _23349_, _09994_);
  and (_23422_, _23421_, _03470_);
  and (_23423_, _23422_, _23420_);
  and (_23424_, _15276_, _15041_);
  nor (_23425_, _15276_, _15041_);
  or (_23426_, _23425_, _23424_);
  nor (_23427_, _15898_, _15536_);
  and (_23428_, _15898_, _15536_);
  nor (_23429_, _23428_, _23427_);
  nor (_23430_, _23429_, _23426_);
  and (_23431_, _23429_, _23426_);
  nor (_23432_, _23431_, _23430_);
  not (_23433_, _16856_);
  nor (_23434_, _16556_, _16215_);
  and (_23435_, _16556_, _16215_);
  nor (_23436_, _23435_, _23434_);
  nor (_23437_, _23436_, _23433_);
  and (_23438_, _23436_, _23433_);
  nor (_23439_, _23438_, _23437_);
  nor (_23440_, _23439_, _23432_);
  and (_23441_, _23439_, _23432_);
  or (_23442_, _23441_, _23440_);
  and (_23443_, _23442_, _08152_);
  nor (_23444_, _23442_, _08152_);
  or (_23445_, _23444_, _23443_);
  and (_23446_, _23445_, _03469_);
  or (_23447_, _23446_, _23423_);
  and (_23448_, _23447_, _03202_);
  nor (_23449_, _23349_, _03202_);
  or (_23450_, _23449_, _23448_);
  or (_23451_, _23450_, _03527_);
  or (_23452_, _23224_, _04457_);
  and (_23453_, _23452_, _08098_);
  and (_23454_, _23453_, _23451_);
  or (_23455_, _23333_, _04029_);
  and (_23456_, _23455_, _11716_);
  or (_23457_, _23456_, _23454_);
  or (_23458_, _23316_, _08160_);
  and (_23459_, _23458_, _03531_);
  and (_23460_, _23459_, _23457_);
  and (_23461_, _23298_, _03530_);
  or (_23462_, _23461_, _11724_);
  or (_23463_, _23462_, _23460_);
  or (_23464_, _23192_, _11723_);
  and (_23465_, _23464_, _03466_);
  and (_23466_, _23465_, _23463_);
  or (_23467_, _23466_, _23275_);
  nand (_23468_, _03572_, _03457_);
  and (_23469_, _23468_, _03639_);
  nor (_23470_, _03641_, _03547_);
  and (_23471_, _23470_, _10112_);
  and (_23472_, _23471_, _11728_);
  and (_23473_, _23472_, _23469_);
  and (_23474_, _23473_, _23467_);
  nor (_23475_, _23473_, _23349_);
  or (_23476_, _23475_, _10124_);
  or (_23477_, _23476_, _23474_);
  or (_23478_, _23192_, _10123_);
  and (_23479_, _23478_, _03459_);
  and (_23481_, _23479_, _23477_);
  nor (_23482_, _15865_, _23368_);
  and (_23483_, _15865_, _23368_);
  nor (_23484_, _23483_, _23482_);
  nor (_23485_, _23484_, _16241_);
  and (_23486_, _23484_, _16241_);
  or (_23487_, _23486_, _23485_);
  not (_23488_, _15559_);
  and (_23489_, _23488_, _15245_);
  nor (_23490_, _23488_, _15245_);
  nor (_23492_, _23490_, _23489_);
  nor (_23493_, _23492_, _16527_);
  and (_23494_, _23492_, _16527_);
  nor (_23495_, _23494_, _23493_);
  and (_23496_, _23495_, _23487_);
  nor (_23497_, _23495_, _23487_);
  nor (_23498_, _23497_, _23496_);
  not (_23499_, _16881_);
  and (_23500_, _23499_, _08177_);
  nor (_23501_, _23499_, _08177_);
  nor (_23502_, _23501_, _23500_);
  or (_23503_, _23502_, _23498_);
  nand (_23504_, _23502_, _23498_);
  and (_23505_, _23504_, _03458_);
  and (_23506_, _23505_, _23503_);
  or (_23507_, _23506_, _23481_);
  nor (_23508_, _03522_, _04755_);
  and (_23509_, _23508_, _03582_);
  and (_23510_, _23509_, _23507_);
  and (_23511_, _03629_, _03558_);
  or (_23513_, _11421_, _23511_);
  or (_23514_, _04054_, _03562_);
  nor (_23515_, _23514_, _23513_);
  or (_23516_, _23509_, _23349_);
  nand (_23517_, _23516_, _23515_);
  or (_23518_, _23517_, _23510_);
  or (_23519_, _23515_, _23192_);
  and (_23520_, _23519_, _07447_);
  nand (_23521_, _23520_, _23518_);
  and (_23522_, _11777_, _08924_);
  nor (_23524_, _15301_, _07393_);
  nor (_23525_, _15302_, _15065_);
  nor (_23526_, _23525_, _23524_);
  nor (_23527_, _23526_, _15564_);
  and (_23528_, _23526_, _15564_);
  nor (_23529_, _23528_, _23527_);
  nor (_23530_, _23529_, _15927_);
  and (_23531_, _23529_, _15927_);
  or (_23532_, _23531_, _23530_);
  not (_23533_, _23532_);
  nor (_23535_, _23533_, _16246_);
  and (_23536_, _23533_, _16246_);
  nor (_23537_, _23536_, _23535_);
  nor (_23538_, _23537_, _16585_);
  and (_23539_, _23537_, _16585_);
  or (_23540_, _23539_, _23538_);
  and (_23541_, _23540_, _16886_);
  nor (_23542_, _23540_, _16886_);
  nor (_23543_, _23542_, _23541_);
  nor (_23544_, _23543_, _08182_);
  and (_23546_, _23543_, _08182_);
  or (_23547_, _23546_, _07447_);
  or (_23548_, _23547_, _23544_);
  and (_23549_, _23548_, _23522_);
  and (_23550_, _23549_, _23521_);
  nor (_23551_, _23522_, _23192_);
  or (_23552_, _23551_, _03586_);
  nor (_23553_, _23552_, _23550_);
  nand (_23554_, _23192_, _03586_);
  nand (_23555_, _23554_, _08191_);
  or (_23557_, _23555_, _23553_);
  and (_23558_, _23557_, _23250_);
  or (_23559_, _23558_, _04066_);
  not (_23560_, _08085_);
  and (_23561_, _15313_, _23560_);
  or (_23562_, _23561_, _08086_);
  nor (_23563_, _23562_, _15600_);
  and (_23564_, _23562_, _15600_);
  or (_23565_, _23564_, _23563_);
  nor (_23566_, _23565_, _15945_);
  and (_23567_, _23565_, _15945_);
  nor (_23568_, _23567_, _23566_);
  nor (_23569_, _23568_, _16267_);
  and (_23570_, _23568_, _16267_);
  nor (_23571_, _23570_, _23569_);
  nor (_23572_, _23571_, _16521_);
  and (_23573_, _23571_, _16521_);
  or (_23574_, _23573_, _23572_);
  nor (_23575_, _23574_, _16919_);
  and (_23576_, _23574_, _16919_);
  nor (_23578_, _23576_, _23575_);
  or (_23579_, _23578_, _08096_);
  and (_23580_, _08095_, _04066_);
  nand (_23581_, _23580_, _23578_);
  and (_23582_, _23581_, _03599_);
  and (_23583_, _23582_, _23579_);
  and (_23584_, _23583_, _23559_);
  not (_23585_, _16820_);
  not (_23586_, _08408_);
  not (_23587_, _16271_);
  not (_23589_, _15952_);
  or (_23590_, _10311_, _10306_);
  and (_23591_, _23590_, _10312_);
  nor (_23592_, _23591_, _15608_);
  and (_23593_, _23591_, _15608_);
  nor (_23594_, _23593_, _23592_);
  and (_23595_, _23594_, _23589_);
  nor (_23596_, _23594_, _23589_);
  nor (_23597_, _23596_, _23595_);
  and (_23598_, _23597_, _23587_);
  nor (_23600_, _23597_, _23587_);
  nor (_23601_, _23600_, _23598_);
  and (_23602_, _23601_, _23586_);
  nor (_23603_, _23601_, _23586_);
  nor (_23604_, _23603_, _23602_);
  nor (_23605_, _23604_, _23585_);
  and (_23606_, _23604_, _23585_);
  nor (_23607_, _23606_, _23605_);
  and (_23608_, _23607_, _08401_);
  nor (_23609_, _23607_, _08401_);
  or (_23611_, _23609_, _07940_);
  or (_23612_, _23611_, _23608_);
  and (_23613_, _23612_, _08267_);
  or (_23614_, _23613_, _23584_);
  not (_23615_, _16289_);
  or (_23616_, _07998_, _07988_);
  and (_23617_, _23616_, _07999_);
  nand (_23618_, _23617_, _15503_);
  or (_23619_, _23617_, _15503_);
  and (_23620_, _23619_, _23618_);
  nor (_23622_, _23620_, _15847_);
  and (_23623_, _23620_, _15847_);
  or (_23624_, _23623_, _23622_);
  and (_23625_, _23624_, _23615_);
  nor (_23626_, _23624_, _23615_);
  nor (_23627_, _23626_, _23625_);
  or (_23628_, _23627_, _16505_);
  nand (_23629_, _23627_, _16505_);
  and (_23630_, _23629_, _23628_);
  nor (_23631_, _23630_, _16935_);
  and (_23632_, _23630_, _16935_);
  nor (_23633_, _23632_, _23631_);
  nor (_23634_, _23633_, _08022_);
  and (_23635_, _23633_, _08022_);
  or (_23636_, _23635_, _23634_);
  or (_23637_, _23636_, _07941_);
  and (_23638_, _23637_, _23614_);
  or (_23639_, _23638_, _03334_);
  nor (_23640_, _05255_, _03512_);
  nor (_23641_, _05276_, _05268_);
  nor (_23643_, _05337_, _05282_);
  nor (_23644_, _05325_, _05264_);
  and (_23645_, _23644_, _23643_);
  nor (_23646_, _23644_, _23643_);
  nor (_23647_, _23646_, _23645_);
  and (_23648_, _23647_, _23641_);
  nor (_23649_, _23647_, _23641_);
  nor (_23650_, _23649_, _23648_);
  nor (_23651_, _23650_, _23640_);
  and (_23652_, _23650_, _23640_);
  or (_23654_, _23652_, _23651_);
  or (_23655_, _23654_, _03233_);
  and (_23656_, _23655_, _03453_);
  and (_23657_, _23656_, _23639_);
  nor (_23658_, _03621_, _03219_);
  not (_23659_, _23658_);
  not (_23660_, _15965_);
  and (_23661_, _23660_, _15620_);
  nor (_23662_, _23660_, _15620_);
  nor (_23663_, _23662_, _23661_);
  nor (_23665_, _16621_, _16298_);
  and (_23666_, _16621_, _16298_);
  nor (_23667_, _23666_, _23665_);
  nor (_23668_, _23667_, _23663_);
  and (_23669_, _23667_, _23663_);
  nor (_23670_, _23669_, _23668_);
  and (_23671_, _15326_, _15086_);
  nor (_23672_, _15326_, _15086_);
  nor (_23673_, _23672_, _23671_);
  and (_23674_, _16944_, _08438_);
  nor (_23676_, _16944_, _08438_);
  nor (_23677_, _23676_, _23674_);
  not (_23678_, _23677_);
  and (_23679_, _23678_, _23673_);
  nor (_23680_, _23678_, _23673_);
  nor (_23681_, _23680_, _23679_);
  or (_23682_, _23681_, _23670_);
  nand (_23683_, _23681_, _23670_);
  and (_23684_, _23683_, _23682_);
  and (_23685_, _23684_, _03452_);
  or (_23687_, _23685_, _23659_);
  or (_23688_, _23687_, _23657_);
  or (_23689_, _23658_, _23192_);
  and (_23690_, _23689_, _06903_);
  and (_23691_, _23690_, _23688_);
  or (_23692_, _23691_, _23226_);
  not (_23693_, _16629_);
  and (_23694_, _23693_, _16305_);
  nor (_23695_, _23693_, _16305_);
  nor (_23696_, _23695_, _23694_);
  not (_23697_, _23696_);
  and (_23698_, _15333_, _15093_);
  nor (_23699_, _15333_, _15093_);
  nor (_23700_, _23699_, _23698_);
  and (_23701_, _23700_, _15627_);
  nor (_23702_, _23700_, _15627_);
  or (_23703_, _23702_, _23701_);
  nand (_23704_, _23703_, _15973_);
  or (_23705_, _23703_, _15973_);
  and (_23706_, _23705_, _23704_);
  nor (_23708_, _23706_, _23697_);
  and (_23709_, _23706_, _23697_);
  nor (_23710_, _23709_, _23708_);
  and (_23711_, _23710_, _16951_);
  nor (_23712_, _23710_, _16951_);
  or (_23713_, _23712_, _23711_);
  and (_23714_, _23713_, _08445_);
  nor (_23715_, _23713_, _08445_);
  or (_23716_, _23715_, _04500_);
  or (_23717_, _23716_, _23714_);
  and (_23719_, _23717_, _03521_);
  and (_23720_, _23719_, _23692_);
  and (_23721_, _15338_, _15011_);
  nor (_23722_, _15338_, _15011_);
  nor (_23723_, _23722_, _23721_);
  not (_23724_, _23723_);
  not (_23725_, _15979_);
  and (_23726_, _23725_, _15632_);
  nor (_23727_, _23725_, _15632_);
  nor (_23728_, _23727_, _23726_);
  and (_23730_, _23728_, _23724_);
  nor (_23731_, _23728_, _23724_);
  or (_23732_, _23731_, _23730_);
  nor (_23733_, _16957_, _16634_);
  and (_23734_, _16957_, _16634_);
  nor (_23735_, _23734_, _23733_);
  not (_23736_, _16311_);
  and (_23737_, _23736_, _08450_);
  nor (_23738_, _23736_, _08450_);
  nor (_23739_, _23738_, _23737_);
  nor (_23741_, _23739_, _23735_);
  and (_23742_, _23739_, _23735_);
  nor (_23743_, _23742_, _23741_);
  nand (_23744_, _23743_, _23732_);
  or (_23745_, _23743_, _23732_);
  and (_23746_, _23745_, _03224_);
  and (_23747_, _23746_, _23744_);
  or (_23748_, _23747_, _23720_);
  and (_23749_, _23748_, _07474_);
  and (_23750_, _07525_, _16962_);
  nor (_23752_, _07525_, _16962_);
  nor (_23753_, _23752_, _23750_);
  not (_23754_, _23753_);
  nor (_23755_, _07613_, _07562_);
  and (_23756_, _07613_, _07562_);
  nor (_23757_, _23756_, _23755_);
  not (_23758_, _23757_);
  and (_23759_, _23758_, _07670_);
  nor (_23760_, _23758_, _07670_);
  nor (_23761_, _23760_, _23759_);
  and (_23762_, _23761_, _23754_);
  nor (_23763_, _23761_, _23754_);
  nor (_23764_, _23763_, _23762_);
  nand (_23765_, _23764_, _08454_);
  or (_23766_, _23764_, _08454_);
  and (_23767_, _23766_, _23765_);
  nor (_23768_, _23767_, _07734_);
  and (_23769_, _23767_, _07734_);
  nor (_23770_, _23769_, _23768_);
  nor (_23771_, _23770_, _07827_);
  and (_23773_, _23770_, _07827_);
  or (_23774_, _23773_, _23771_);
  and (_23775_, _23774_, _07468_);
  or (_23776_, _23775_, _23749_);
  and (_23777_, _23776_, _03263_);
  nand (_23778_, _23654_, _03262_);
  nand (_23779_, _23778_, _23197_);
  or (_23780_, _23779_, _23777_);
  and (_23781_, _23780_, _23198_);
  or (_23782_, _23781_, _05913_);
  nand (_23784_, _23349_, _05913_);
  and (_23785_, _23784_, _04509_);
  and (_23786_, _23785_, _23782_);
  nor (_23787_, _15348_, _15104_);
  and (_23788_, _15348_, _15104_);
  or (_23789_, _23788_, _23787_);
  nor (_23790_, _15990_, _15642_);
  and (_23791_, _15990_, _15642_);
  nor (_23792_, _23791_, _23790_);
  nor (_23793_, _23792_, _23789_);
  and (_23795_, _23792_, _23789_);
  or (_23796_, _23795_, _23793_);
  nor (_23797_, _16645_, _16322_);
  and (_23798_, _16645_, _16322_);
  nor (_23799_, _23798_, _23797_);
  and (_23800_, _23799_, _16970_);
  nor (_23801_, _23799_, _16970_);
  nor (_23802_, _23801_, _23800_);
  and (_23803_, _23802_, _23796_);
  nor (_23804_, _23802_, _23796_);
  or (_23806_, _23804_, _23803_);
  or (_23807_, _23806_, _08464_);
  nand (_23808_, _23806_, _08464_);
  and (_23809_, _23808_, _03624_);
  and (_23810_, _23809_, _23807_);
  or (_23811_, _23810_, _23786_);
  and (_23812_, _23811_, _08462_);
  nand (_23813_, _23654_, _08461_);
  not (_23814_, _11828_);
  and (_23815_, _11864_, _23814_);
  nand (_23817_, _23815_, _23813_);
  or (_23818_, _23817_, _23812_);
  not (_23819_, _11868_);
  or (_23820_, _23815_, _23192_);
  and (_23821_, _23820_, _23819_);
  and (_23822_, _23821_, _23818_);
  nand (_23823_, _23192_, _11868_);
  nand (_23824_, _23823_, _11415_);
  or (_23825_, _23824_, _23822_);
  and (_23826_, _15809_, _07899_);
  nor (_23827_, _15809_, _07899_);
  nor (_23828_, _23827_, _23826_);
  and (_23829_, _15007_, _07903_);
  nor (_23830_, _23829_, _15575_);
  nor (_23831_, _23830_, _23828_);
  and (_23832_, _23830_, _23828_);
  nor (_23833_, _23832_, _23831_);
  and (_23834_, _07892_, _07888_);
  nor (_23835_, _07892_, _07888_);
  nor (_23836_, _23835_, _23834_);
  nor (_23838_, _23836_, _23833_);
  and (_23839_, _23836_, _23833_);
  nor (_23840_, _23839_, _23838_);
  and (_23841_, _23840_, _16980_);
  nor (_23842_, _23840_, _16980_);
  nor (_23843_, _23842_, _23841_);
  nor (_23844_, _23843_, _07882_);
  and (_23845_, _23843_, _07882_);
  or (_23846_, _23845_, _23844_);
  or (_23847_, _23846_, _11415_);
  and (_23849_, _23847_, _23825_);
  or (_23850_, _23849_, _08481_);
  nor (_23851_, _15825_, _08759_);
  and (_23852_, _15825_, _08759_);
  nor (_23853_, _23852_, _23851_);
  and (_23854_, _15117_, _08763_);
  nor (_23855_, _23854_, _15593_);
  nor (_23856_, _23855_, _23853_);
  and (_23857_, _23855_, _23853_);
  nor (_23858_, _23857_, _23856_);
  nor (_23860_, _16509_, _08752_);
  and (_23861_, _16509_, _08752_);
  nor (_23862_, _23861_, _23860_);
  nor (_23863_, _23862_, _23858_);
  and (_23864_, _23862_, _23858_);
  nor (_23865_, _23864_, _23863_);
  or (_23866_, _23865_, _08745_);
  nand (_23867_, _23865_, _08745_);
  and (_23868_, _23867_, _23866_);
  nand (_23869_, _23868_, _08489_);
  or (_23871_, _23868_, _08489_);
  and (_23872_, _23871_, _23869_);
  or (_23873_, _23872_, _08487_);
  and (_23874_, _23873_, _08486_);
  and (_23875_, _23874_, _23850_);
  nor (_23876_, _12793_, _12588_);
  and (_23877_, _12793_, _12588_);
  nor (_23878_, _23877_, _23876_);
  nor (_23879_, _12381_, _12183_);
  and (_23880_, _12381_, _12183_);
  nor (_23882_, _23880_, _23879_);
  not (_23883_, _23882_);
  and (_23884_, _23883_, _23878_);
  nor (_23885_, _23883_, _23878_);
  nor (_23886_, _23885_, _23884_);
  or (_23887_, _23886_, _12992_);
  nand (_23888_, _23886_, _12992_);
  and (_23889_, _23888_, _23887_);
  or (_23890_, _23889_, _13204_);
  nand (_23891_, _23889_, _13204_);
  and (_23893_, _23891_, _23890_);
  not (_23894_, _13407_);
  and (_23895_, _23894_, _06443_);
  nor (_23896_, _23894_, _06443_);
  nor (_23897_, _23896_, _23895_);
  or (_23898_, _23897_, _23893_);
  nand (_23899_, _23897_, _23893_);
  and (_23900_, _23899_, _03746_);
  and (_23901_, _23900_, _23898_);
  or (_23902_, _23901_, _07929_);
  or (_23904_, _23902_, _23875_);
  and (_23905_, _10127_, _08829_);
  nor (_23906_, _23905_, _10128_);
  and (_23907_, _10160_, _07991_);
  nor (_23908_, _23907_, _10161_);
  nor (_23909_, _16761_, _08824_);
  and (_23910_, _16761_, _08824_);
  or (_23911_, _23910_, _23909_);
  nand (_23912_, _23911_, _23908_);
  or (_23913_, _23911_, _23908_);
  and (_23914_, _23913_, _23912_);
  or (_23915_, _23914_, _23906_);
  nand (_23916_, _23914_, _23906_);
  and (_23917_, _23916_, _23915_);
  and (_23918_, _08819_, _07933_);
  nor (_23919_, _10143_, _23918_);
  not (_23920_, _23919_);
  nor (_23921_, _23920_, _23917_);
  and (_23922_, _23920_, _23917_);
  or (_23923_, _23922_, _23921_);
  or (_23925_, _23923_, _07930_);
  and (_23926_, _23925_, _04527_);
  and (_23927_, _23926_, _23904_);
  and (_23928_, _15374_, _15003_);
  nor (_23929_, _15374_, _15003_);
  nor (_23930_, _23929_, _23928_);
  not (_23931_, _23930_);
  not (_23932_, _15822_);
  and (_23933_, _23932_, _15672_);
  nor (_23934_, _23932_, _15672_);
  nor (_23936_, _23934_, _23933_);
  and (_23937_, _23936_, _23931_);
  nor (_23938_, _23936_, _23931_);
  or (_23939_, _23938_, _23937_);
  nor (_23940_, _16810_, _16670_);
  and (_23941_, _16810_, _16670_);
  nor (_23942_, _23941_, _23940_);
  not (_23943_, _16157_);
  and (_23944_, _23943_, _08501_);
  nor (_23945_, _23943_, _08501_);
  nor (_23947_, _23945_, _23944_);
  nor (_23948_, _23947_, _23942_);
  and (_23949_, _23947_, _23942_);
  nor (_23950_, _23949_, _23948_);
  or (_23951_, _23950_, _23939_);
  nand (_23952_, _23950_, _23939_);
  and (_23953_, _23952_, _03623_);
  and (_23954_, _23953_, _23951_);
  or (_23955_, _23954_, _23927_);
  and (_23956_, _23955_, _03745_);
  nor (_23958_, _11889_, _03172_);
  nand (_23959_, _23192_, _03744_);
  or (_23960_, _23959_, _05312_);
  nand (_23961_, _23960_, _23958_);
  or (_23962_, _23961_, _23956_);
  or (_23963_, _23958_, _23192_);
  and (_23964_, _23963_, _08506_);
  and (_23965_, _23964_, _23962_);
  or (_23966_, _07904_, _07901_);
  nand (_23967_, _07904_, _07901_);
  and (_23969_, _23967_, _23966_);
  and (_23970_, _15682_, _07894_);
  and (_23971_, _07897_, _07895_);
  nor (_23972_, _23971_, _23970_);
  not (_23973_, _23972_);
  and (_23974_, _23973_, _23969_);
  nor (_23975_, _23973_, _23969_);
  nor (_23976_, _23975_, _23974_);
  nor (_23977_, _07890_, _07883_);
  and (_23978_, _07890_, _07883_);
  nor (_23979_, _23978_, _23977_);
  nor (_23980_, _23979_, _16678_);
  and (_23981_, _23979_, _16678_);
  nor (_23982_, _23981_, _23980_);
  not (_23983_, _23982_);
  nor (_23984_, _23983_, _23976_);
  and (_23985_, _23983_, _23976_);
  nor (_23986_, _23985_, _23984_);
  or (_23987_, _23986_, _07881_);
  nand (_23988_, _23986_, _07881_);
  and (_23990_, _23988_, _08507_);
  and (_23991_, _23990_, _23987_);
  or (_23992_, _23991_, _04141_);
  or (_23993_, _23992_, _23965_);
  or (_23994_, _08764_, _08761_);
  nand (_23995_, _08764_, _08761_);
  and (_23996_, _23995_, _23994_);
  nor (_23997_, _08756_, _08757_);
  and (_23998_, _08756_, _08757_);
  nor (_23999_, _23998_, _23997_);
  not (_24001_, _23999_);
  and (_24002_, _24001_, _23996_);
  nor (_24003_, _24001_, _23996_);
  nor (_24004_, _24003_, _24002_);
  nor (_24005_, _08750_, _08743_);
  and (_24006_, _08750_, _08743_);
  nor (_24007_, _24006_, _24005_);
  nor (_24008_, _24007_, _08749_);
  and (_24009_, _24007_, _08749_);
  nor (_24010_, _24009_, _24008_);
  nor (_24012_, _24010_, _24004_);
  and (_24013_, _24010_, _24004_);
  nor (_24014_, _24013_, _24012_);
  and (_24015_, _24014_, _08488_);
  nor (_24016_, _24014_, _08488_);
  or (_24017_, _24016_, _08510_);
  or (_24018_, _24017_, _24015_);
  and (_24019_, _24018_, _08519_);
  and (_24020_, _24019_, _23993_);
  nor (_24021_, _12379_, _12182_);
  and (_24023_, _12379_, _12182_);
  nor (_24024_, _24023_, _24021_);
  not (_24025_, _12791_);
  and (_24026_, _24025_, _12586_);
  nor (_24027_, _24025_, _12586_);
  nor (_24028_, _24027_, _24026_);
  and (_24029_, _24028_, _24024_);
  nor (_24030_, _24028_, _24024_);
  nor (_24031_, _24030_, _24029_);
  not (_24032_, _13276_);
  nor (_24034_, _13202_, _12990_);
  and (_24035_, _13202_, _12990_);
  nor (_24036_, _24035_, _24034_);
  nor (_24037_, _24036_, _24032_);
  and (_24038_, _24036_, _24032_);
  nor (_24039_, _24038_, _24037_);
  and (_24040_, _24039_, _24031_);
  nor (_24041_, _24039_, _24031_);
  or (_24042_, _24041_, _24040_);
  nor (_24043_, _24042_, _06441_);
  and (_24045_, _24042_, _06441_);
  or (_24046_, _24045_, _24043_);
  and (_24047_, _24046_, _03735_);
  or (_24048_, _24047_, _08517_);
  or (_24049_, _24048_, _24020_);
  or (_24050_, _08831_, _07989_);
  nand (_24051_, _08831_, _07989_);
  and (_24052_, _24051_, _24050_);
  not (_24053_, _08825_);
  and (_24054_, _24053_, _08827_);
  nor (_24056_, _24053_, _08827_);
  nor (_24057_, _24056_, _24054_);
  and (_24058_, _24057_, _24052_);
  nor (_24059_, _24057_, _24052_);
  nor (_24060_, _24059_, _24058_);
  or (_24061_, _24060_, _08822_);
  nand (_24062_, _24060_, _08822_);
  and (_24063_, _24062_, _24061_);
  or (_24064_, _24063_, _08820_);
  nand (_24065_, _24063_, _08820_);
  and (_24067_, _24065_, _24064_);
  or (_24068_, _24067_, _08817_);
  nand (_24069_, _24067_, _08817_);
  and (_24070_, _24069_, _24068_);
  and (_24071_, _24070_, _07931_);
  nor (_24072_, _24070_, _07931_);
  or (_24073_, _24072_, _24071_);
  or (_24074_, _24073_, _08518_);
  and (_24075_, _24074_, _04523_);
  and (_24076_, _24075_, _24049_);
  not (_24078_, _11915_);
  and (_24079_, _24078_, _10828_);
  nor (_24080_, _15699_, _15141_);
  and (_24081_, _15699_, _15141_);
  nor (_24082_, _24081_, _24080_);
  nor (_24083_, _17013_, _16368_);
  and (_24084_, _17013_, _16368_);
  nor (_24085_, _24084_, _24083_);
  and (_24086_, _24085_, _24082_);
  nor (_24087_, _24085_, _24082_);
  nor (_24089_, _24087_, _24086_);
  nor (_24090_, _16034_, _15391_);
  and (_24091_, _16034_, _15391_);
  nor (_24092_, _24091_, _24090_);
  nor (_24093_, _16697_, _08526_);
  and (_24094_, _16697_, _08526_);
  nor (_24095_, _24094_, _24093_);
  and (_24096_, _24095_, _24092_);
  nor (_24097_, _24095_, _24092_);
  nor (_24098_, _24097_, _24096_);
  not (_24100_, _24098_);
  nand (_24101_, _24100_, _24089_);
  or (_24102_, _24100_, _24089_);
  and (_24103_, _24102_, _03611_);
  nand (_24104_, _24103_, _24101_);
  nand (_24105_, _24104_, _24079_);
  or (_24106_, _24105_, _24076_);
  or (_24107_, _23192_, _24079_);
  and (_24108_, _24107_, _11412_);
  and (_24109_, _24108_, _24106_);
  nor (_24111_, _14998_, _07902_);
  and (_24112_, _14998_, _07902_);
  nor (_24113_, _24112_, _24111_);
  and (_24114_, _24113_, _07898_);
  nor (_24115_, _24113_, _07898_);
  or (_24116_, _24115_, _24114_);
  and (_24117_, _24116_, _07896_);
  nor (_24118_, _24116_, _07896_);
  or (_24119_, _24118_, _24117_);
  not (_24120_, _07887_);
  nor (_24122_, _07891_, _07884_);
  and (_24123_, _07891_, _07884_);
  nor (_24124_, _24123_, _24122_);
  nor (_24125_, _24124_, _24120_);
  and (_24126_, _24124_, _24120_);
  nor (_24127_, _24126_, _24125_);
  not (_24128_, _24127_);
  nor (_24129_, _24128_, _24119_);
  and (_24130_, _24128_, _24119_);
  or (_24131_, _24130_, _24129_);
  and (_24133_, _24131_, _07880_);
  nor (_24134_, _24131_, _07880_);
  or (_24135_, _24134_, _24133_);
  and (_24136_, _24135_, _15224_);
  or (_24137_, _24136_, _07923_);
  or (_24138_, _24137_, _24109_);
  nor (_24139_, _15116_, _08762_);
  and (_24140_, _15116_, _08762_);
  nor (_24141_, _24140_, _24139_);
  not (_24142_, _24141_);
  nor (_24144_, _08754_, _08758_);
  and (_24145_, _08754_, _08758_);
  nor (_24146_, _24145_, _24144_);
  nor (_24147_, _24146_, _24142_);
  and (_24148_, _24146_, _24142_);
  nor (_24149_, _24148_, _24147_);
  nor (_24150_, _08751_, _08744_);
  and (_24151_, _08751_, _08744_);
  nor (_24152_, _24151_, _24150_);
  nor (_24153_, _24152_, _08747_);
  and (_24155_, _24152_, _08747_);
  nor (_24156_, _24155_, _24153_);
  nor (_24157_, _24156_, _24149_);
  and (_24158_, _24156_, _24149_);
  nor (_24159_, _24158_, _24157_);
  nor (_24160_, _24159_, _07924_);
  and (_24161_, _24159_, _07924_);
  or (_24162_, _24161_, _24160_);
  or (_24163_, _24162_, _11411_);
  and (_24164_, _24163_, _03740_);
  and (_24166_, _24164_, _24138_);
  nor (_24167_, _12380_, _12181_);
  and (_24168_, _12380_, _12181_);
  nor (_24169_, _24168_, _24167_);
  and (_24170_, _24169_, _12587_);
  nor (_24171_, _24169_, _12587_);
  or (_24172_, _24171_, _24170_);
  nand (_24173_, _24172_, _12792_);
  or (_24174_, _24172_, _12792_);
  and (_24175_, _24174_, _24173_);
  nor (_24177_, _13203_, _12991_);
  and (_24178_, _13203_, _12991_);
  nor (_24179_, _24178_, _24177_);
  nor (_24180_, _24179_, _13406_);
  and (_24181_, _24179_, _13406_);
  nor (_24182_, _24181_, _24180_);
  not (_24183_, _24182_);
  nor (_24184_, _24183_, _24175_);
  and (_24185_, _24183_, _24175_);
  nor (_24186_, _24185_, _24184_);
  or (_24189_, _24186_, _06442_);
  nand (_24190_, _24186_, _06442_);
  and (_24191_, _24190_, _03739_);
  and (_24192_, _24191_, _24189_);
  or (_24193_, _24192_, _08542_);
  or (_24194_, _24193_, _24166_);
  nor (_24195_, _10159_, _07990_);
  and (_24196_, _10159_, _07990_);
  nor (_24197_, _24196_, _24195_);
  not (_24198_, _08826_);
  and (_24201_, _24198_, _08828_);
  nor (_24202_, _24198_, _08828_);
  nor (_24203_, _24202_, _24201_);
  and (_24204_, _24203_, _24197_);
  nor (_24205_, _24203_, _24197_);
  nor (_24206_, _24205_, _24204_);
  not (_24207_, _08823_);
  nor (_24208_, _08821_, _08818_);
  and (_24209_, _08821_, _08818_);
  nor (_24210_, _24209_, _24208_);
  nor (_24213_, _24210_, _24207_);
  and (_24214_, _24210_, _24207_);
  nor (_24215_, _24214_, _24213_);
  and (_24216_, _24215_, _24206_);
  nor (_24217_, _24215_, _24206_);
  or (_24218_, _24217_, _24216_);
  and (_24219_, _24218_, _07932_);
  nor (_24220_, _24218_, _07932_);
  or (_24221_, _24220_, _24219_);
  or (_24222_, _24221_, _08543_);
  and (_24225_, _24222_, _06453_);
  and (_24226_, _24225_, _24194_);
  and (_24227_, _11942_, _11932_);
  nor (_24228_, _15406_, _15163_);
  and (_24229_, _15406_, _15163_);
  or (_24230_, _24229_, _24228_);
  nor (_24231_, _16058_, _15723_);
  and (_24232_, _16058_, _15723_);
  nor (_24233_, _24232_, _24231_);
  nor (_24234_, _24233_, _24230_);
  and (_24237_, _24233_, _24230_);
  nor (_24238_, _24237_, _24234_);
  nor (_24239_, _17034_, _16720_);
  and (_24240_, _17034_, _16720_);
  nor (_24241_, _24240_, _24239_);
  not (_24242_, _16391_);
  and (_24243_, _24242_, _08551_);
  nor (_24244_, _24242_, _08551_);
  nor (_24245_, _24244_, _24243_);
  nor (_24246_, _24245_, _24241_);
  and (_24249_, _24245_, _24241_);
  nor (_24250_, _24249_, _24246_);
  not (_24251_, _24250_);
  nand (_24252_, _24251_, _24238_);
  or (_24253_, _24251_, _24238_);
  and (_24254_, _24253_, _03618_);
  nand (_24255_, _24254_, _24252_);
  nand (_24256_, _24255_, _24227_);
  or (_24257_, _24256_, _24226_);
  or (_24258_, _23192_, _24227_);
  and (_24261_, _24258_, _08564_);
  and (_24262_, _24261_, _24257_);
  nor (_24263_, _15411_, _15070_);
  and (_24264_, _15411_, _15070_);
  or (_24265_, _24264_, _24263_);
  nor (_24266_, _24265_, _15730_);
  and (_24267_, _24265_, _15730_);
  nor (_24268_, _24267_, _24266_);
  nor (_24269_, _24268_, _15816_);
  and (_24270_, _24268_, _15816_);
  or (_24272_, _24270_, _24269_);
  nor (_24273_, _24272_, _16397_);
  and (_24274_, _24272_, _16397_);
  or (_24275_, _24274_, _24273_);
  nor (_24276_, _24275_, _16480_);
  and (_24277_, _24275_, _16480_);
  or (_24278_, _24277_, _24276_);
  and (_24279_, _24278_, _17039_);
  nor (_24280_, _24278_, _17039_);
  or (_24281_, _24280_, _24279_);
  nand (_24283_, _24281_, _08591_);
  or (_24284_, _24281_, _08591_);
  and (_24285_, _24284_, _24283_);
  and (_24286_, _24285_, _15728_);
  or (_24287_, _24286_, _08595_);
  or (_24288_, _24287_, _24262_);
  nor (_24289_, _08085_, _08083_);
  nor (_24290_, _15416_, _23560_);
  nor (_24291_, _24290_, _24289_);
  nor (_24292_, _24291_, _15735_);
  and (_24294_, _24291_, _15735_);
  nor (_24295_, _24294_, _24292_);
  nor (_24296_, _24295_, _16068_);
  and (_24297_, _24295_, _16068_);
  or (_24298_, _24297_, _24296_);
  nor (_24299_, _24298_, _16402_);
  and (_24300_, _24298_, _16402_);
  or (_24301_, _24300_, _24299_);
  and (_24302_, _24301_, _16728_);
  nor (_24303_, _24301_, _16728_);
  or (_24305_, _24303_, _24302_);
  and (_24306_, _24305_, _17045_);
  nor (_24307_, _24305_, _17045_);
  nor (_24308_, _24307_, _24306_);
  nor (_24309_, _24308_, _08623_);
  and (_24310_, _24308_, _08623_);
  or (_24311_, _24310_, _24309_);
  or (_24312_, _24311_, _08599_);
  and (_24313_, _24312_, _03732_);
  and (_24314_, _24313_, _24288_);
  and (_24316_, _15421_, _10306_);
  nor (_24317_, _15421_, _10306_);
  nor (_24318_, _24317_, _24316_);
  nor (_24319_, _24318_, _15741_);
  and (_24320_, _24318_, _15741_);
  nor (_24321_, _24320_, _24319_);
  nor (_24322_, _24321_, _16073_);
  and (_24323_, _24321_, _16073_);
  or (_24324_, _24323_, _24322_);
  nor (_24325_, _24324_, _16408_);
  and (_24327_, _24324_, _16408_);
  or (_24328_, _24327_, _24325_);
  nor (_24329_, _24328_, _16733_);
  and (_24330_, _24328_, _16733_);
  or (_24331_, _24330_, _24329_);
  and (_24332_, _24331_, _17050_);
  nor (_24333_, _24331_, _17050_);
  or (_24334_, _24333_, _24332_);
  nor (_24335_, _24334_, _08703_);
  and (_24336_, _24334_, _08703_);
  or (_24338_, _24336_, _24335_);
  and (_24339_, _24338_, _03731_);
  or (_24340_, _24339_, _08627_);
  or (_24341_, _24340_, _24314_);
  and (_24342_, _15426_, _07988_);
  nor (_24343_, _15426_, _07988_);
  nor (_24344_, _24343_, _24342_);
  nor (_24345_, _24344_, _15482_);
  and (_24346_, _24344_, _15482_);
  nor (_24347_, _24346_, _24345_);
  nor (_24349_, _24347_, _16079_);
  and (_24350_, _24347_, _16079_);
  nor (_24351_, _24350_, _24349_);
  nor (_24352_, _24351_, _16146_);
  and (_24353_, _24351_, _16146_);
  or (_24354_, _24353_, _24352_);
  nor (_24355_, _24354_, _16739_);
  and (_24356_, _24354_, _16739_);
  or (_24357_, _24356_, _24355_);
  and (_24358_, _24357_, _17056_);
  nor (_24360_, _24357_, _17056_);
  nor (_24361_, _24360_, _24358_);
  nor (_24362_, _24361_, _08733_);
  and (_24363_, _24361_, _08733_);
  or (_24364_, _24363_, _24362_);
  or (_24365_, _24364_, _08709_);
  and (_24366_, _24365_, _08708_);
  and (_24367_, _24366_, _24341_);
  nor (_24368_, _07993_, _07992_);
  nor (_24369_, _15528_, \oc8051_golden_model_1.ACC [3]);
  and (_24371_, _15528_, \oc8051_golden_model_1.ACC [3]);
  nor (_24372_, _24371_, _24369_);
  and (_24373_, _24372_, _23356_);
  nor (_24374_, _24372_, _23356_);
  nor (_24375_, _24374_, _24373_);
  not (_24376_, _24375_);
  nand (_24377_, _24376_, _24368_);
  or (_24378_, _24376_, _24368_);
  and (_24379_, _24378_, _24377_);
  nand (_24380_, _24379_, _08707_);
  and (_24382_, _10848_, _03814_);
  nand (_24383_, _24382_, _24380_);
  or (_24384_, _24383_, _24367_);
  or (_24385_, _24382_, _23192_);
  and (_24386_, _24385_, _07921_);
  and (_24387_, _24386_, _24384_);
  not (_24388_, _14998_);
  and (_24389_, _24388_, _07903_);
  nor (_24390_, _24388_, _07903_);
  nor (_24391_, _24390_, _24389_);
  and (_24393_, _24391_, _15752_);
  nor (_24394_, _24391_, _15752_);
  nor (_24395_, _24394_, _24393_);
  and (_24396_, _24395_, _15812_);
  nor (_24397_, _24395_, _15812_);
  nor (_24398_, _24397_, _24396_);
  and (_24399_, _24398_, _16419_);
  nor (_24400_, _24398_, _16419_);
  nor (_24401_, _24400_, _24399_);
  nor (_24402_, _24401_, _16477_);
  and (_24404_, _24401_, _16477_);
  or (_24405_, _24404_, _24402_);
  and (_24406_, _24405_, _17063_);
  nor (_24407_, _24405_, _17063_);
  or (_24408_, _24407_, _24406_);
  nor (_24409_, _24408_, _07919_);
  and (_24410_, _24408_, _07919_);
  or (_24411_, _24410_, _24409_);
  and (_24412_, _24411_, _07920_);
  or (_24413_, _24412_, _04184_);
  or (_24415_, _24413_, _24387_);
  not (_24416_, _15116_);
  and (_24417_, _24416_, _08763_);
  nor (_24418_, _24416_, _08763_);
  nor (_24419_, _24418_, _24417_);
  and (_24420_, _24419_, _15757_);
  nor (_24421_, _24419_, _15757_);
  nor (_24422_, _24421_, _24420_);
  and (_24423_, _24422_, _16091_);
  nor (_24424_, _24422_, _16091_);
  nor (_24426_, _24424_, _24423_);
  and (_24427_, _24426_, _16424_);
  nor (_24428_, _24426_, _16424_);
  nor (_24429_, _24428_, _24427_);
  and (_24430_, _24429_, _16751_);
  nor (_24431_, _24429_, _16751_);
  nor (_24432_, _24431_, _24430_);
  and (_24433_, _24432_, _17069_);
  nor (_24434_, _24432_, _17069_);
  nor (_24435_, _24434_, _24433_);
  nor (_24437_, _24435_, _08779_);
  and (_24438_, _24435_, _08779_);
  or (_24439_, _24438_, _24437_);
  or (_24440_, _24439_, _08742_);
  and (_24441_, _24440_, _08784_);
  and (_24442_, _24441_, _24415_);
  not (_24443_, _08811_);
  not (_24444_, _16756_);
  not (_24445_, _15763_);
  nor (_24446_, _15444_, _08415_);
  and (_24448_, _15444_, _08415_);
  or (_24449_, _24448_, _24446_);
  and (_24450_, _24449_, _24445_);
  nor (_24451_, _24449_, _24445_);
  nor (_24452_, _24451_, _24450_);
  and (_24453_, _24452_, _16097_);
  nor (_24454_, _24452_, _16097_);
  nor (_24455_, _24454_, _24453_);
  nor (_24456_, _24455_, _16430_);
  and (_24457_, _24455_, _16430_);
  or (_24459_, _24457_, _24456_);
  and (_24460_, _24459_, _24444_);
  nor (_24461_, _24459_, _24444_);
  nor (_24462_, _24461_, _24460_);
  nor (_24463_, _24462_, _17074_);
  and (_24464_, _24462_, _17074_);
  nor (_24465_, _24464_, _24463_);
  nor (_24466_, _24465_, _24443_);
  and (_24467_, _24465_, _24443_);
  or (_24468_, _24467_, _24466_);
  and (_24470_, _24468_, _03478_);
  not (_24471_, _10159_);
  and (_24472_, _24471_, _07991_);
  nor (_24473_, _24471_, _07991_);
  nor (_24474_, _24473_, _24472_);
  and (_24475_, _24474_, _15768_);
  nor (_24476_, _24474_, _15768_);
  nor (_24477_, _24476_, _24475_);
  and (_24478_, _24477_, _16104_);
  nor (_24479_, _24477_, _16104_);
  nor (_24481_, _24479_, _24478_);
  nor (_24482_, _24481_, _16435_);
  and (_24483_, _24481_, _16435_);
  or (_24484_, _24483_, _24482_);
  nor (_24485_, _24484_, _16764_);
  and (_24486_, _24484_, _16764_);
  nor (_24487_, _24486_, _24485_);
  nor (_24488_, _24487_, _17080_);
  and (_24489_, _24487_, _17080_);
  nor (_24490_, _24489_, _24488_);
  and (_24492_, _24490_, _08846_);
  nor (_24493_, _24490_, _08846_);
  or (_24494_, _24493_, _24492_);
  nand (_24495_, _24494_, _08783_);
  nand (_24496_, _24495_, _23195_);
  or (_24497_, _24496_, _24470_);
  or (_24498_, _24497_, _24442_);
  and (_24499_, _24498_, _23196_);
  nor (_24500_, _05912_, _05139_);
  or (_24501_, _24500_, _24499_);
  nand (_24503_, _24500_, _23349_);
  and (_24504_, _24503_, _03948_);
  and (_24505_, _24504_, _24501_);
  and (_24506_, _23391_, _03767_);
  or (_24507_, _24506_, _08853_);
  or (_24508_, _24507_, _24505_);
  not (_24509_, _08859_);
  and (_24510_, _15528_, _24509_);
  and (_24511_, _24510_, \oc8051_golden_model_1.ACC [3]);
  nor (_24512_, _24510_, \oc8051_golden_model_1.ACC [3]);
  nor (_24514_, _24512_, _24511_);
  and (_24515_, _24514_, _16448_);
  nor (_24516_, _24514_, _16448_);
  nor (_24517_, _24516_, _24515_);
  and (_24518_, _16775_, _07495_);
  nor (_24519_, _16775_, _07495_);
  nor (_24520_, _24519_, _24518_);
  nor (_24521_, _24520_, _24517_);
  and (_24522_, _24520_, _24517_);
  or (_24523_, _24522_, _24521_);
  nor (_24525_, _24523_, _08865_);
  and (_24526_, _24523_, _08865_);
  nor (_24527_, _24526_, _24525_);
  and (_24528_, _24527_, _08853_);
  nor (_24529_, _24528_, _08858_);
  and (_24530_, _24529_, _24508_);
  and (_24531_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_24532_, _24531_, _08142_);
  or (_24533_, _24532_, _24375_);
  nand (_24534_, _24532_, _24375_);
  and (_24536_, _24534_, _24533_);
  nand (_24537_, _24536_, _08858_);
  nand (_24538_, _24537_, _04553_);
  or (_24539_, _24538_, _24530_);
  or (_24540_, _23192_, _04553_);
  and (_24541_, _24540_, _03446_);
  and (_24542_, _24541_, _24539_);
  not (_24543_, _04795_);
  and (_24544_, _24543_, _04790_);
  nand (_24545_, _23274_, _03445_);
  nand (_24547_, _24545_, _24544_);
  or (_24548_, _24547_, _24542_);
  nor (_24549_, _04734_, _04215_);
  or (_24550_, _23192_, _24544_);
  and (_24551_, _24550_, _24549_);
  and (_24552_, _24551_, _24548_);
  nor (_24553_, _23349_, _24549_);
  or (_24554_, _24553_, _03473_);
  or (_24555_, _24554_, _24552_);
  nor (_24556_, _15468_, _15035_);
  and (_24558_, _15468_, _15035_);
  nor (_24559_, _24558_, _24556_);
  nor (_24560_, _24559_, _15793_);
  and (_24561_, _24559_, _15793_);
  nor (_24562_, _24561_, _24560_);
  and (_24563_, _24562_, _16788_);
  nor (_24564_, _24562_, _16788_);
  or (_24565_, _24564_, _24563_);
  not (_24566_, _16128_);
  nor (_24567_, _16461_, _24566_);
  and (_24569_, _16461_, _24566_);
  nor (_24570_, _24569_, _24567_);
  and (_24571_, _24570_, _24565_);
  nor (_24572_, _24570_, _24565_);
  nor (_24573_, _24572_, _24571_);
  not (_24574_, _17103_);
  nand (_24575_, _24574_, _08878_);
  or (_24576_, _24574_, _08878_);
  and (_24577_, _24576_, _24575_);
  and (_24578_, _24577_, _24573_);
  nor (_24580_, _24577_, _24573_);
  or (_24581_, _24580_, _03474_);
  or (_24582_, _24581_, _24578_);
  and (_24583_, _24582_, _08876_);
  and (_24584_, _24583_, _24555_);
  not (_24585_, _08883_);
  and (_24586_, _15528_, _24585_);
  and (_24587_, _24586_, _07644_);
  nor (_24588_, _24586_, _07644_);
  nor (_24589_, _24588_, _24587_);
  nor (_24591_, _24589_, _16466_);
  and (_24592_, _24589_, _16466_);
  or (_24593_, _24592_, _24591_);
  and (_24594_, _24593_, _17109_);
  nor (_24595_, _24593_, _17109_);
  nor (_24596_, _24595_, _24594_);
  nor (_24597_, _16794_, _08890_);
  and (_24598_, _16794_, _08890_);
  nor (_24599_, _24598_, _24597_);
  nor (_24600_, _24599_, _24596_);
  and (_24602_, _24599_, _24596_);
  or (_24603_, _24602_, _24600_);
  nand (_24604_, _24603_, _08875_);
  nor (_24605_, _03615_, _03194_);
  nor (_24606_, _12031_, _08882_);
  and (_24607_, _24606_, _24605_);
  nand (_24608_, _24607_, _24604_);
  or (_24609_, _24608_, _24584_);
  or (_24610_, _24607_, _23192_);
  and (_24611_, _24610_, _43189_);
  and (_24613_, _24611_, _24609_);
  or (_24614_, _24613_, _23177_);
  and (_43821_, _24614_, _42003_);
  or (_24615_, _05303_, \oc8051_golden_model_1.PSW [1]);
  and (_24616_, _12265_, _05303_);
  not (_24617_, _24616_);
  and (_24618_, _24617_, _24615_);
  or (_24619_, _24618_, _04432_);
  nand (_24620_, _05303_, _03269_);
  and (_24621_, _24620_, _24615_);
  and (_24624_, _24621_, _04436_);
  not (_24625_, \oc8051_golden_model_1.PSW [1]);
  nor (_24626_, _04436_, _24625_);
  or (_24627_, _24626_, _03534_);
  or (_24628_, _24627_, _24624_);
  and (_24629_, _24628_, _03470_);
  and (_24630_, _24629_, _24619_);
  and (_24631_, _12269_, _05932_);
  nor (_24632_, _05932_, _24625_);
  or (_24633_, _24632_, _03527_);
  or (_24635_, _24633_, _24631_);
  and (_24636_, _24635_, _03533_);
  or (_24637_, _24636_, _24630_);
  nor (_24638_, _05303_, _24625_);
  nor (_24639_, _09753_, _04635_);
  or (_24640_, _24639_, _24638_);
  or (_24641_, _24640_, _04457_);
  and (_24642_, _24641_, _24637_);
  or (_24643_, _24642_, _03530_);
  or (_24644_, _24621_, _03531_);
  and (_24646_, _24644_, _03466_);
  and (_24647_, _24646_, _24643_);
  and (_24648_, _12256_, _05932_);
  or (_24649_, _24648_, _24632_);
  and (_24650_, _24649_, _03465_);
  or (_24651_, _24650_, _03458_);
  or (_24652_, _24651_, _24647_);
  and (_24653_, _24631_, _12284_);
  or (_24654_, _24632_, _03459_);
  or (_24655_, _24654_, _24653_);
  and (_24657_, _24655_, _24652_);
  and (_24658_, _24657_, _03453_);
  not (_24659_, _05932_);
  nor (_24660_, _12301_, _24659_);
  or (_24661_, _24632_, _24660_);
  and (_24662_, _24661_, _03452_);
  or (_24663_, _24662_, _07454_);
  or (_24664_, _24663_, _24658_);
  or (_24665_, _24640_, _06903_);
  and (_24666_, _24665_, _24664_);
  or (_24668_, _24666_, _04082_);
  and (_24669_, _06572_, _05303_);
  or (_24670_, _24638_, _04500_);
  or (_24671_, _24670_, _24669_);
  and (_24672_, _24671_, _03521_);
  and (_24673_, _24672_, _24668_);
  nor (_24674_, _12360_, _09753_);
  or (_24675_, _24674_, _24638_);
  and (_24676_, _24675_, _03224_);
  or (_24677_, _24676_, _24673_);
  and (_24679_, _24677_, _03625_);
  or (_24680_, _12375_, _09753_);
  and (_24681_, _24680_, _03623_);
  nand (_24682_, _05303_, _04325_);
  and (_24683_, _24682_, _03624_);
  or (_24684_, _24683_, _24681_);
  and (_24685_, _24684_, _24615_);
  or (_24686_, _24685_, _24679_);
  and (_24687_, _24686_, _03745_);
  or (_24688_, _12381_, _09753_);
  and (_24690_, _24615_, _03744_);
  and (_24691_, _24690_, _24688_);
  or (_24692_, _24691_, _24687_);
  and (_24693_, _24692_, _04523_);
  or (_24694_, _12374_, _09753_);
  and (_24695_, _24615_, _03611_);
  and (_24696_, _24695_, _24694_);
  or (_24697_, _24696_, _24693_);
  and (_24698_, _24697_, _03734_);
  or (_24699_, _24638_, _05674_);
  and (_24701_, _24621_, _03733_);
  and (_24702_, _24701_, _24699_);
  or (_24703_, _24702_, _24698_);
  and (_24704_, _24703_, _03742_);
  or (_24705_, _24682_, _05674_);
  and (_24706_, _24615_, _03618_);
  and (_24707_, _24706_, _24705_);
  or (_24708_, _24620_, _05674_);
  and (_24709_, _24615_, _03741_);
  and (_24710_, _24709_, _24708_);
  or (_24712_, _24710_, _03767_);
  or (_24713_, _24712_, _24707_);
  or (_24714_, _24713_, _24704_);
  or (_24715_, _24618_, _03948_);
  and (_24716_, _24715_, _03446_);
  and (_24717_, _24716_, _24714_);
  and (_24718_, _24649_, _03445_);
  or (_24719_, _24718_, _03473_);
  or (_24720_, _24719_, _24717_);
  or (_24721_, _24638_, _03474_);
  or (_24723_, _24721_, _24616_);
  and (_24724_, _24723_, _24720_);
  or (_24725_, _24724_, _43193_);
  or (_24726_, _43189_, \oc8051_golden_model_1.PSW [1]);
  and (_24727_, _24726_, _42003_);
  and (_43822_, _24727_, _24725_);
  not (_24728_, \oc8051_golden_model_1.PSW [2]);
  nor (_24729_, _05303_, _24728_);
  nor (_24730_, _12568_, _09753_);
  or (_24731_, _24730_, _24729_);
  and (_24733_, _24731_, _03224_);
  nor (_24734_, _09753_, _05073_);
  or (_24735_, _24734_, _24729_);
  or (_24736_, _24735_, _06903_);
  and (_24737_, _09744_, _08488_);
  nor (_24738_, _08026_, \oc8051_golden_model_1.ACC [7]);
  nor (_24739_, _24738_, _24737_);
  and (_24740_, _24739_, _09766_);
  nor (_24741_, _24739_, _09766_);
  or (_24742_, _24741_, _24740_);
  and (_24744_, _24742_, _08095_);
  nor (_24745_, _24742_, _08095_);
  or (_24746_, _24745_, _24744_);
  or (_24747_, _24746_, _08024_);
  and (_24748_, _24735_, _03527_);
  nor (_24749_, _05932_, _24728_);
  and (_24750_, _12462_, _05932_);
  or (_24751_, _24750_, _24749_);
  or (_24752_, _24751_, _03470_);
  nor (_24753_, _12467_, _09753_);
  or (_24755_, _24753_, _24729_);
  and (_24756_, _24755_, _03534_);
  nor (_24757_, _04436_, _24728_);
  and (_24758_, _05303_, \oc8051_golden_model_1.ACC [2]);
  or (_24759_, _24758_, _24729_);
  and (_24760_, _24759_, _04436_);
  or (_24761_, _24760_, _24757_);
  and (_24762_, _24761_, _04432_);
  or (_24763_, _24762_, _03469_);
  or (_24764_, _24763_, _24756_);
  and (_24766_, _24764_, _24752_);
  and (_24767_, _24766_, _04457_);
  or (_24768_, _24767_, _24748_);
  or (_24769_, _24768_, _03530_);
  or (_24770_, _24759_, _03531_);
  and (_24771_, _24770_, _03466_);
  and (_24772_, _24771_, _24769_);
  and (_24773_, _12460_, _05932_);
  or (_24774_, _24773_, _24749_);
  and (_24775_, _24774_, _03465_);
  or (_24777_, _24775_, _24772_);
  and (_24778_, _24777_, _03459_);
  or (_24779_, _24749_, _12491_);
  and (_24780_, _24779_, _03458_);
  and (_24781_, _24780_, _24751_);
  or (_24782_, _24781_, _24778_);
  and (_24783_, _24782_, _07447_);
  or (_24784_, _14226_, _07449_);
  or (_24785_, _24784_, _14337_);
  or (_24786_, _24785_, _14451_);
  or (_24788_, _24786_, _14569_);
  or (_24789_, _24788_, _14683_);
  nor (_24790_, _24789_, _14801_);
  nand (_24791_, _24790_, _14916_);
  and (_24792_, _24791_, _06933_);
  or (_24793_, _24792_, _08194_);
  or (_24794_, _24793_, _24783_);
  nor (_24795_, _08198_, \oc8051_golden_model_1.ACC [7]);
  and (_24796_, _08198_, \oc8051_golden_model_1.ACC [7]);
  nor (_24797_, _24796_, _24795_);
  and (_24799_, _24797_, _10278_);
  nor (_24800_, _24797_, _10278_);
  or (_24801_, _24800_, _24799_);
  and (_24802_, _24801_, _08260_);
  nor (_24803_, _24801_, _08260_);
  or (_24804_, _24803_, _24802_);
  or (_24805_, _24804_, _08191_);
  and (_24806_, _24805_, _24794_);
  or (_24807_, _24806_, _04066_);
  and (_24808_, _24807_, _03599_);
  and (_24810_, _24808_, _24747_);
  nor (_24811_, _10319_, _08652_);
  or (_24812_, _24811_, _08653_);
  not (_24813_, _08644_);
  and (_24814_, _10323_, _24813_);
  nor (_24815_, _10323_, _24813_);
  nor (_24816_, _24815_, _24814_);
  nand (_24817_, _24816_, _24812_);
  or (_24818_, _24816_, _24812_);
  and (_24819_, _24818_, _03594_);
  and (_24821_, _24819_, _24817_);
  or (_24822_, _24821_, _07940_);
  or (_24823_, _24822_, _24810_);
  not (_24824_, _07947_);
  and (_24825_, _08019_, _24824_);
  nor (_24826_, _24825_, _10336_);
  and (_24827_, _24825_, _10336_);
  or (_24828_, _24827_, _07941_);
  or (_24829_, _24828_, _24826_);
  and (_24830_, _24829_, _03453_);
  and (_24832_, _24830_, _24823_);
  nor (_24833_, _12509_, _24659_);
  or (_24834_, _24833_, _24749_);
  and (_24835_, _24834_, _03452_);
  or (_24836_, _24835_, _07454_);
  or (_24837_, _24836_, _24832_);
  and (_24838_, _24837_, _24736_);
  or (_24839_, _24838_, _04082_);
  and (_24840_, _06710_, _05303_);
  or (_24841_, _24729_, _04500_);
  or (_24843_, _24841_, _24840_);
  and (_24844_, _24843_, _03521_);
  and (_24845_, _24844_, _24839_);
  or (_24846_, _24845_, _24733_);
  and (_24847_, _24846_, _07474_);
  nor (_24848_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_24849_, _24848_, _07493_);
  nand (_24850_, _24849_, _07468_);
  nand (_24851_, _24850_, _03625_);
  or (_24852_, _24851_, _24847_);
  and (_24854_, _12582_, _05303_);
  or (_24855_, _24729_, _04527_);
  or (_24856_, _24855_, _24854_);
  and (_24857_, _05303_, _06399_);
  or (_24858_, _24857_, _24729_);
  or (_24859_, _24858_, _04509_);
  and (_24860_, _24859_, _03745_);
  and (_24861_, _24860_, _24856_);
  and (_24862_, _24861_, _24852_);
  and (_24863_, _12588_, _05303_);
  or (_24865_, _24863_, _24729_);
  and (_24866_, _24865_, _03744_);
  or (_24867_, _24866_, _24862_);
  and (_24868_, _24867_, _04523_);
  or (_24869_, _24729_, _05772_);
  and (_24870_, _24858_, _03611_);
  and (_24871_, _24870_, _24869_);
  or (_24872_, _24871_, _24868_);
  and (_24873_, _24872_, _03734_);
  and (_24874_, _24759_, _03733_);
  and (_24876_, _24874_, _24869_);
  or (_24877_, _24876_, _03618_);
  or (_24878_, _24877_, _24873_);
  nor (_24879_, _12581_, _09753_);
  or (_24880_, _24729_, _06453_);
  or (_24881_, _24880_, _24879_);
  and (_24882_, _24881_, _06458_);
  and (_24883_, _24882_, _24878_);
  nor (_24884_, _12587_, _09753_);
  or (_24885_, _24884_, _24729_);
  and (_24887_, _24885_, _03741_);
  or (_24888_, _24887_, _08556_);
  or (_24889_, _24888_, _24883_);
  and (_24890_, _24797_, _10393_);
  nor (_24891_, _24890_, _24796_);
  and (_24892_, _24891_, _08591_);
  and (_24893_, _24796_, _08588_);
  or (_24894_, _24893_, _24892_);
  and (_24895_, _24894_, _08566_);
  or (_24896_, _24895_, _08564_);
  and (_24898_, _24896_, _24889_);
  and (_24899_, _24894_, _08565_);
  or (_24900_, _24899_, _08595_);
  or (_24901_, _24900_, _24898_);
  and (_24902_, _24737_, _08620_);
  and (_24903_, _24739_, _09742_);
  nor (_24904_, _24903_, _24737_);
  and (_24905_, _24904_, _08623_);
  or (_24906_, _24905_, _24902_);
  or (_24907_, _24906_, _08599_);
  and (_24909_, _24907_, _03732_);
  and (_24910_, _24909_, _24901_);
  nor (_24911_, _08642_, _10429_);
  nor (_24912_, _08643_, \oc8051_golden_model_1.ACC [7]);
  nor (_24913_, _24912_, _10404_);
  nor (_24914_, _24913_, _24911_);
  nand (_24915_, _24914_, _08703_);
  nand (_24916_, _24911_, _08700_);
  and (_24917_, _24916_, _24915_);
  nor (_24918_, _24917_, _03732_);
  or (_24920_, _24918_, _08627_);
  or (_24921_, _24920_, _24910_);
  and (_24922_, _07946_, \oc8051_golden_model_1.ACC [7]);
  and (_24923_, _24922_, _08730_);
  nor (_24924_, _07949_, _07946_);
  or (_24925_, _24924_, _08709_);
  or (_24926_, _24925_, _08731_);
  and (_24927_, _24926_, _08734_);
  or (_24928_, _24927_, _24923_);
  and (_24929_, _24928_, _07921_);
  and (_24931_, _24929_, _24921_);
  or (_24932_, _07916_, _07880_);
  or (_24933_, _10416_, _07915_);
  and (_24934_, _24933_, _07920_);
  and (_24935_, _24934_, _24932_);
  or (_24936_, _24935_, _24931_);
  and (_24937_, _24936_, _08742_);
  nand (_24938_, _08776_, _10422_);
  and (_24939_, _24938_, _10424_);
  or (_24940_, _24939_, _24937_);
  and (_24942_, _24940_, _08784_);
  or (_24943_, _08808_, _08268_);
  and (_24944_, _24943_, _10431_);
  nand (_24945_, _08843_, _09731_);
  and (_24946_, _24945_, _09733_);
  or (_24947_, _24946_, _03767_);
  or (_24948_, _24947_, _24944_);
  or (_24949_, _24948_, _24942_);
  or (_24950_, _24755_, _03948_);
  and (_24951_, _24950_, _03446_);
  and (_24953_, _24951_, _24949_);
  and (_24954_, _24774_, _03445_);
  or (_24955_, _24954_, _03473_);
  or (_24956_, _24955_, _24953_);
  and (_24957_, _12638_, _05303_);
  or (_24958_, _24729_, _03474_);
  or (_24959_, _24958_, _24957_);
  and (_24960_, _24959_, _24956_);
  or (_24961_, _24960_, _43193_);
  or (_24962_, _43189_, \oc8051_golden_model_1.PSW [2]);
  and (_24964_, _24962_, _42003_);
  and (_43825_, _24964_, _24961_);
  not (_24965_, \oc8051_golden_model_1.PSW [3]);
  nor (_24966_, _05303_, _24965_);
  and (_24967_, _05303_, _06356_);
  nor (_24968_, _24967_, _24966_);
  and (_24969_, _24968_, _03624_);
  nor (_24970_, _09753_, _04885_);
  nor (_24971_, _24970_, _24966_);
  and (_24972_, _24971_, _07454_);
  and (_24974_, _05303_, \oc8051_golden_model_1.ACC [3]);
  nor (_24975_, _24974_, _24966_);
  nor (_24976_, _24975_, _04437_);
  nor (_24977_, _04436_, _24965_);
  or (_24978_, _24977_, _24976_);
  and (_24979_, _24978_, _04432_);
  nor (_24980_, _12652_, _09753_);
  nor (_24981_, _24980_, _24966_);
  nor (_24982_, _24981_, _04432_);
  or (_24983_, _24982_, _24979_);
  and (_24985_, _24983_, _03470_);
  nor (_24986_, _05932_, _24965_);
  and (_24987_, _12664_, _05932_);
  nor (_24988_, _24987_, _24986_);
  nor (_24989_, _24988_, _03470_);
  or (_24990_, _24989_, _03527_);
  or (_24991_, _24990_, _24985_);
  nand (_24992_, _24971_, _03527_);
  and (_24993_, _24992_, _24991_);
  and (_24994_, _24993_, _03531_);
  nor (_24996_, _24975_, _03531_);
  or (_24997_, _24996_, _24994_);
  and (_24998_, _24997_, _03466_);
  and (_24999_, _12662_, _05932_);
  nor (_25000_, _24999_, _24986_);
  nor (_25001_, _25000_, _03466_);
  or (_25002_, _25001_, _03458_);
  or (_25003_, _25002_, _24998_);
  nor (_25004_, _24986_, _12691_);
  nor (_25005_, _25004_, _24988_);
  or (_25007_, _25005_, _03459_);
  and (_25008_, _25007_, _03453_);
  and (_25009_, _25008_, _25003_);
  nor (_25010_, _12709_, _24659_);
  nor (_25011_, _25010_, _24986_);
  nor (_25012_, _25011_, _03453_);
  nor (_25013_, _25012_, _07454_);
  not (_25014_, _25013_);
  nor (_25015_, _25014_, _25009_);
  nor (_25016_, _25015_, _24972_);
  nor (_25018_, _25016_, _04082_);
  and (_25019_, _06664_, _05303_);
  nor (_25020_, _24966_, _04500_);
  not (_25021_, _25020_);
  nor (_25022_, _25021_, _25019_);
  or (_25023_, _25022_, _03224_);
  nor (_25024_, _25023_, _25018_);
  nor (_25025_, _12773_, _09753_);
  nor (_25026_, _24966_, _25025_);
  nor (_25027_, _25026_, _03521_);
  or (_25029_, _25027_, _03624_);
  nor (_25030_, _25029_, _25024_);
  nor (_25031_, _25030_, _24969_);
  or (_25032_, _25031_, _03623_);
  and (_25033_, _12787_, _05303_);
  or (_25034_, _25033_, _24966_);
  or (_25035_, _25034_, _04527_);
  and (_25036_, _25035_, _03745_);
  and (_25037_, _25036_, _25032_);
  and (_25038_, _12793_, _05303_);
  nor (_25040_, _25038_, _24966_);
  nor (_25041_, _25040_, _03745_);
  nor (_25042_, _25041_, _25037_);
  nor (_25043_, _25042_, _03611_);
  nor (_25044_, _24966_, _05625_);
  not (_25045_, _25044_);
  nor (_25046_, _24968_, _04523_);
  and (_25047_, _25046_, _25045_);
  nor (_25048_, _25047_, _25043_);
  nor (_25049_, _25048_, _03733_);
  nor (_25051_, _24975_, _03734_);
  and (_25052_, _25051_, _25045_);
  nor (_25053_, _25052_, _03618_);
  not (_25054_, _25053_);
  nor (_25055_, _25054_, _25049_);
  nor (_25056_, _12786_, _09753_);
  or (_25057_, _24966_, _06453_);
  nor (_25058_, _25057_, _25056_);
  or (_25059_, _25058_, _03741_);
  nor (_25060_, _25059_, _25055_);
  nor (_25062_, _12792_, _09753_);
  nor (_25063_, _25062_, _24966_);
  nor (_25064_, _25063_, _06458_);
  or (_25065_, _25064_, _25060_);
  and (_25066_, _25065_, _03948_);
  nor (_25067_, _24981_, _03948_);
  or (_25068_, _25067_, _25066_);
  and (_25069_, _25068_, _03446_);
  nor (_25070_, _25000_, _03446_);
  or (_25071_, _25070_, _25069_);
  and (_25073_, _25071_, _03474_);
  and (_25074_, _12843_, _05303_);
  nor (_25075_, _25074_, _24966_);
  nor (_25076_, _25075_, _03474_);
  or (_25077_, _25076_, _25073_);
  or (_25078_, _25077_, _43193_);
  or (_25079_, _43189_, \oc8051_golden_model_1.PSW [3]);
  and (_25080_, _25079_, _42003_);
  and (_43826_, _25080_, _25078_);
  not (_25081_, \oc8051_golden_model_1.PSW [4]);
  nor (_25083_, _05303_, _25081_);
  nor (_25084_, _05831_, _09753_);
  nor (_25085_, _25084_, _25083_);
  and (_25086_, _25085_, _07454_);
  nor (_25087_, _05932_, _25081_);
  and (_25088_, _12864_, _05932_);
  nor (_25089_, _25088_, _25087_);
  nor (_25090_, _25089_, _03466_);
  and (_25091_, _05303_, \oc8051_golden_model_1.ACC [4]);
  nor (_25092_, _25091_, _25083_);
  nor (_25094_, _25092_, _04437_);
  nor (_25095_, _04436_, _25081_);
  or (_25096_, _25095_, _25094_);
  and (_25097_, _25096_, _04432_);
  nor (_25098_, _12856_, _09753_);
  nor (_25099_, _25098_, _25083_);
  nor (_25100_, _25099_, _04432_);
  or (_25101_, _25100_, _25097_);
  and (_25102_, _25101_, _03470_);
  and (_25103_, _12866_, _05932_);
  nor (_25104_, _25103_, _25087_);
  nor (_25105_, _25104_, _03470_);
  or (_25106_, _25105_, _03527_);
  or (_25107_, _25106_, _25102_);
  nand (_25108_, _25085_, _03527_);
  and (_25109_, _25108_, _25107_);
  and (_25110_, _25109_, _03531_);
  nor (_25111_, _25092_, _03531_);
  or (_25112_, _25111_, _25110_);
  and (_25113_, _25112_, _03466_);
  nor (_25116_, _25113_, _25090_);
  nor (_25117_, _25116_, _03458_);
  nor (_25118_, _25087_, _12894_);
  or (_25119_, _25104_, _03459_);
  nor (_25120_, _25119_, _25118_);
  nor (_25121_, _25120_, _25117_);
  nor (_25122_, _25121_, _03452_);
  nor (_25123_, _12912_, _24659_);
  nor (_25124_, _25123_, _25087_);
  nor (_25125_, _25124_, _03453_);
  nor (_25127_, _25125_, _07454_);
  not (_25128_, _25127_);
  nor (_25129_, _25128_, _25122_);
  nor (_25130_, _25129_, _25086_);
  nor (_25131_, _25130_, _04082_);
  and (_25132_, _06802_, _05303_);
  nor (_25133_, _25083_, _04500_);
  not (_25134_, _25133_);
  nor (_25135_, _25134_, _25132_);
  nor (_25136_, _25135_, _03224_);
  not (_25138_, _25136_);
  nor (_25139_, _25138_, _25131_);
  nor (_25140_, _12972_, _09753_);
  nor (_25141_, _25140_, _25083_);
  nor (_25142_, _25141_, _03521_);
  or (_25143_, _25142_, _08905_);
  or (_25144_, _25143_, _25139_);
  and (_25145_, _12986_, _05303_);
  or (_25146_, _25083_, _04527_);
  or (_25147_, _25146_, _25145_);
  and (_25148_, _06337_, _05303_);
  nor (_25149_, _25148_, _25083_);
  and (_25150_, _25149_, _03624_);
  nor (_25151_, _25150_, _03744_);
  and (_25152_, _25151_, _25147_);
  and (_25153_, _25152_, _25144_);
  and (_25154_, _12992_, _05303_);
  nor (_25155_, _25154_, _25083_);
  nor (_25156_, _25155_, _03745_);
  nor (_25157_, _25156_, _25153_);
  nor (_25160_, _25157_, _03611_);
  nor (_25161_, _25083_, _05880_);
  not (_25162_, _25161_);
  nor (_25163_, _25149_, _04523_);
  and (_25164_, _25163_, _25162_);
  nor (_25165_, _25164_, _25160_);
  nor (_25166_, _25165_, _03733_);
  nor (_25167_, _25092_, _03734_);
  and (_25168_, _25167_, _25162_);
  nor (_25169_, _25168_, _03618_);
  not (_25171_, _25169_);
  nor (_25172_, _25171_, _25166_);
  nor (_25173_, _12985_, _09753_);
  or (_25174_, _25083_, _06453_);
  nor (_25175_, _25174_, _25173_);
  or (_25176_, _25175_, _03741_);
  nor (_25177_, _25176_, _25172_);
  nor (_25178_, _12991_, _09753_);
  nor (_25179_, _25178_, _25083_);
  nor (_25180_, _25179_, _06458_);
  or (_25181_, _25180_, _25177_);
  and (_25182_, _25181_, _03948_);
  nor (_25183_, _25099_, _03948_);
  or (_25184_, _25183_, _25182_);
  and (_25185_, _25184_, _03446_);
  nor (_25186_, _25089_, _03446_);
  or (_25187_, _25186_, _25185_);
  and (_25188_, _25187_, _03474_);
  and (_25189_, _13051_, _05303_);
  nor (_25190_, _25189_, _25083_);
  nor (_25193_, _25190_, _03474_);
  or (_25194_, _25193_, _25188_);
  or (_25195_, _25194_, _43193_);
  or (_25196_, _43189_, \oc8051_golden_model_1.PSW [4]);
  and (_25197_, _25196_, _42003_);
  and (_43827_, _25197_, _25195_);
  not (_25198_, \oc8051_golden_model_1.PSW [5]);
  nor (_25199_, _05303_, _25198_);
  and (_25200_, _06757_, _05303_);
  or (_25201_, _25200_, _25199_);
  and (_25203_, _25201_, _04082_);
  and (_25204_, _05303_, \oc8051_golden_model_1.ACC [5]);
  nor (_25205_, _25204_, _25199_);
  nor (_25206_, _25205_, _04437_);
  nor (_25207_, _04436_, _25198_);
  or (_25208_, _25207_, _25206_);
  and (_25209_, _25208_, _04432_);
  nor (_25210_, _13070_, _09753_);
  nor (_25211_, _25210_, _25199_);
  nor (_25212_, _25211_, _04432_);
  or (_25214_, _25212_, _25209_);
  and (_25215_, _25214_, _03470_);
  nor (_25216_, _05932_, _25198_);
  and (_25217_, _13095_, _05932_);
  nor (_25218_, _25217_, _25216_);
  nor (_25219_, _25218_, _03470_);
  or (_25220_, _25219_, _03527_);
  or (_25221_, _25220_, _25215_);
  nor (_25222_, _05526_, _09753_);
  nor (_25223_, _25222_, _25199_);
  nand (_25225_, _25223_, _03527_);
  and (_25226_, _25225_, _25221_);
  and (_25227_, _25226_, _03531_);
  nor (_25228_, _25205_, _03531_);
  or (_25229_, _25228_, _25227_);
  and (_25230_, _25229_, _03466_);
  and (_25231_, _13078_, _05932_);
  nor (_25232_, _25231_, _25216_);
  nor (_25233_, _25232_, _03466_);
  or (_25234_, _25233_, _25230_);
  and (_25235_, _25234_, _03459_);
  nor (_25236_, _25216_, _13110_);
  nor (_25237_, _25236_, _25218_);
  and (_25238_, _25237_, _03458_);
  or (_25239_, _25238_, _25235_);
  and (_25240_, _25239_, _03453_);
  nor (_25241_, _13076_, _24659_);
  nor (_25242_, _25241_, _25216_);
  nor (_25243_, _25242_, _03453_);
  nor (_25244_, _25243_, _07454_);
  not (_25247_, _25244_);
  nor (_25248_, _25247_, _25240_);
  and (_25249_, _25223_, _07454_);
  or (_25250_, _25249_, _04082_);
  nor (_25251_, _25250_, _25248_);
  or (_25252_, _25251_, _25203_);
  and (_25253_, _25252_, _03521_);
  nor (_25254_, _13184_, _09753_);
  nor (_25255_, _25254_, _25199_);
  nor (_25256_, _25255_, _03521_);
  or (_25258_, _25256_, _08905_);
  or (_25259_, _25258_, _25253_);
  and (_25260_, _13198_, _05303_);
  or (_25261_, _25199_, _04527_);
  or (_25262_, _25261_, _25260_);
  and (_25263_, _06295_, _05303_);
  nor (_25264_, _25263_, _25199_);
  and (_25265_, _25264_, _03624_);
  nor (_25266_, _25265_, _03744_);
  and (_25267_, _25266_, _25262_);
  and (_25269_, _25267_, _25259_);
  and (_25270_, _13204_, _05303_);
  nor (_25271_, _25270_, _25199_);
  nor (_25272_, _25271_, _03745_);
  nor (_25273_, _25272_, _25269_);
  nor (_25274_, _25273_, _03611_);
  nor (_25275_, _25199_, _05576_);
  not (_25276_, _25275_);
  nor (_25277_, _25264_, _04523_);
  and (_25278_, _25277_, _25276_);
  nor (_25280_, _25278_, _25274_);
  nor (_25281_, _25280_, _03733_);
  nor (_25282_, _25205_, _03734_);
  and (_25283_, _25282_, _25276_);
  nor (_25284_, _25283_, _03618_);
  not (_25285_, _25284_);
  nor (_25286_, _25285_, _25281_);
  nor (_25287_, _13197_, _09753_);
  or (_25288_, _25199_, _06453_);
  nor (_25289_, _25288_, _25287_);
  or (_25291_, _25289_, _03741_);
  nor (_25292_, _25291_, _25286_);
  nor (_25293_, _13203_, _09753_);
  nor (_25294_, _25293_, _25199_);
  nor (_25295_, _25294_, _06458_);
  or (_25296_, _25295_, _25292_);
  and (_25297_, _25296_, _03948_);
  nor (_25298_, _25211_, _03948_);
  or (_25299_, _25298_, _25297_);
  and (_25300_, _25299_, _03446_);
  nor (_25302_, _25232_, _03446_);
  or (_25303_, _25302_, _25300_);
  and (_25304_, _25303_, _03474_);
  and (_25305_, _13253_, _05303_);
  nor (_25306_, _25305_, _25199_);
  nor (_25307_, _25306_, _03474_);
  or (_25308_, _25307_, _25304_);
  or (_25309_, _25308_, _43193_);
  or (_25310_, _43189_, \oc8051_golden_model_1.PSW [5]);
  and (_25311_, _25310_, _42003_);
  and (_43828_, _25311_, _25309_);
  and (_25313_, _07920_, _07910_);
  not (_25314_, _08694_);
  nor (_25315_, _25314_, _08639_);
  nor (_25316_, _25315_, _03732_);
  nor (_25317_, _08564_, _08209_);
  and (_25318_, _25317_, _08582_);
  nor (_25319_, _05303_, _15890_);
  nor (_25320_, _05417_, _09753_);
  nor (_25321_, _25320_, _25319_);
  and (_25323_, _25321_, _07454_);
  nor (_25324_, _08088_, _08038_);
  nor (_25325_, _25324_, _08024_);
  nor (_25326_, _05932_, _15890_);
  and (_25327_, _13304_, _05932_);
  nor (_25328_, _25327_, _25326_);
  nor (_25329_, _25328_, _03466_);
  and (_25330_, _05303_, \oc8051_golden_model_1.ACC [6]);
  nor (_25331_, _25330_, _25319_);
  nor (_25332_, _25331_, _04437_);
  nor (_25334_, _04436_, _15890_);
  or (_25335_, _25334_, _25332_);
  and (_25336_, _25335_, _04432_);
  nor (_25337_, _13293_, _09753_);
  nor (_25338_, _25337_, _25319_);
  nor (_25339_, _25338_, _04432_);
  or (_25340_, _25339_, _25336_);
  and (_25341_, _25340_, _03470_);
  and (_25342_, _13280_, _05932_);
  nor (_25343_, _25342_, _25326_);
  nor (_25345_, _25343_, _03470_);
  or (_25346_, _25345_, _03527_);
  or (_25347_, _25346_, _25341_);
  nand (_25348_, _25321_, _03527_);
  and (_25349_, _25348_, _25347_);
  and (_25350_, _25349_, _03531_);
  nor (_25351_, _25331_, _03531_);
  or (_25352_, _25351_, _25350_);
  and (_25353_, _25352_, _03466_);
  nor (_25354_, _25353_, _25329_);
  nor (_25356_, _25354_, _03458_);
  nor (_25357_, _25326_, _13311_);
  or (_25358_, _25357_, _03459_);
  or (_25359_, _25358_, _25343_);
  and (_25360_, _25359_, _08191_);
  not (_25361_, _25360_);
  nor (_25362_, _25361_, _25356_);
  nor (_25363_, _08209_, _08191_);
  and (_25364_, _25363_, _08250_);
  or (_25365_, _25364_, _04066_);
  nor (_25366_, _25365_, _25362_);
  or (_25367_, _25366_, _25325_);
  and (_25368_, _25367_, _03599_);
  or (_25369_, _08639_, _07940_);
  or (_25370_, _25369_, _10314_);
  and (_25371_, _25370_, _08267_);
  nor (_25372_, _25371_, _25368_);
  or (_25373_, _07943_, _07941_);
  nor (_25374_, _25373_, _08012_);
  or (_25375_, _25374_, _03452_);
  nor (_25378_, _25375_, _25372_);
  nor (_25379_, _13329_, _24659_);
  nor (_25380_, _25379_, _25326_);
  nor (_25381_, _25380_, _03453_);
  nor (_25382_, _25381_, _07454_);
  not (_25383_, _25382_);
  nor (_25384_, _25383_, _25378_);
  nor (_25385_, _25384_, _25323_);
  nor (_25386_, _25385_, _04082_);
  and (_25387_, _06526_, _05303_);
  nor (_25389_, _25319_, _04500_);
  not (_25390_, _25389_);
  nor (_25391_, _25390_, _25387_);
  nor (_25392_, _25391_, _03224_);
  not (_25393_, _25392_);
  nor (_25394_, _25393_, _25386_);
  nor (_25395_, _13387_, _09753_);
  nor (_25396_, _25395_, _25319_);
  nor (_25397_, _25396_, _03521_);
  or (_25398_, _25397_, _08905_);
  or (_25400_, _25398_, _25394_);
  and (_25401_, _13402_, _05303_);
  or (_25402_, _25319_, _04527_);
  or (_25403_, _25402_, _25401_);
  and (_25404_, _14949_, _05303_);
  nor (_25405_, _25404_, _25319_);
  and (_25406_, _25405_, _03624_);
  nor (_25407_, _25406_, _03744_);
  and (_25408_, _25407_, _25403_);
  and (_25409_, _25408_, _25400_);
  and (_25411_, _13407_, _05303_);
  nor (_25412_, _25411_, _25319_);
  nor (_25413_, _25412_, _03745_);
  nor (_25414_, _25413_, _25409_);
  nor (_25415_, _25414_, _03611_);
  nor (_25416_, _25319_, _05469_);
  not (_25417_, _25416_);
  nor (_25418_, _25405_, _04523_);
  and (_25419_, _25418_, _25417_);
  nor (_25420_, _25419_, _25415_);
  nor (_25422_, _25420_, _03733_);
  nor (_25423_, _25331_, _03734_);
  and (_25424_, _25423_, _25417_);
  or (_25425_, _25424_, _25422_);
  and (_25426_, _25425_, _06453_);
  nor (_25427_, _13400_, _09753_);
  nor (_25428_, _25427_, _25319_);
  nor (_25429_, _25428_, _06453_);
  or (_25430_, _25429_, _25426_);
  and (_25431_, _25430_, _06458_);
  nor (_25433_, _13406_, _09753_);
  nor (_25434_, _25433_, _25319_);
  nor (_25435_, _25434_, _06458_);
  nor (_25436_, _25435_, _15728_);
  not (_25437_, _25436_);
  nor (_25438_, _25437_, _25431_);
  nor (_25439_, _25438_, _25318_);
  nor (_25440_, _25439_, _08595_);
  nor (_25441_, _08038_, _08599_);
  nand (_25442_, _25441_, _08614_);
  and (_25444_, _25442_, _03732_);
  not (_25445_, _25444_);
  nor (_25446_, _25445_, _25440_);
  nor (_25447_, _25446_, _25316_);
  nor (_25448_, _25447_, _08627_);
  not (_25449_, _07943_);
  and (_25450_, _08724_, _25449_);
  nor (_25451_, _25450_, _08709_);
  nor (_25452_, _25451_, _07920_);
  not (_25453_, _25452_);
  nor (_25455_, _25453_, _25448_);
  nor (_25456_, _25455_, _25313_);
  nor (_25457_, _25456_, _04184_);
  nor (_25458_, _08770_, _08742_);
  nor (_25459_, _25458_, _03478_);
  not (_25460_, _25459_);
  nor (_25461_, _25460_, _25457_);
  or (_25462_, _08802_, _08783_);
  and (_25463_, _25462_, _08785_);
  nor (_25464_, _25463_, _25461_);
  nor (_25466_, _08837_, _08786_);
  nor (_25467_, _25466_, _25464_);
  and (_25468_, _25467_, _03948_);
  nor (_25469_, _25338_, _03948_);
  or (_25470_, _25469_, _25468_);
  and (_25471_, _25470_, _03446_);
  nor (_25472_, _25328_, _03446_);
  or (_25473_, _25472_, _25471_);
  and (_25474_, _25473_, _03474_);
  and (_25475_, _13456_, _05303_);
  nor (_25477_, _25319_, _25475_);
  nor (_25478_, _25477_, _03474_);
  or (_25479_, _25478_, _25474_);
  or (_25480_, _25479_, _43193_);
  or (_25481_, _43189_, \oc8051_golden_model_1.PSW [6]);
  and (_25482_, _25481_, _42003_);
  and (_43829_, _25482_, _25480_);
  not (_25483_, \oc8051_golden_model_1.PCON [0]);
  nor (_25484_, _05261_, _25483_);
  nor (_25485_, _05722_, _10456_);
  nor (_25487_, _25485_, _25484_);
  and (_25488_, _25487_, _17198_);
  and (_25489_, _05261_, \oc8051_golden_model_1.ACC [0]);
  nor (_25490_, _25489_, _25484_);
  nor (_25491_, _25490_, _03531_);
  nor (_25492_, _25490_, _04437_);
  nor (_25493_, _04436_, _25483_);
  or (_25494_, _25493_, _25492_);
  and (_25495_, _25494_, _04432_);
  nor (_25496_, _25487_, _04432_);
  or (_25498_, _25496_, _25495_);
  and (_25499_, _25498_, _04457_);
  and (_25500_, _05261_, _04429_);
  nor (_25501_, _25500_, _25484_);
  nor (_25502_, _25501_, _04457_);
  nor (_25503_, _25502_, _25499_);
  nor (_25504_, _25503_, _03530_);
  or (_25505_, _25504_, _07454_);
  nor (_25506_, _25505_, _25491_);
  and (_25507_, _25501_, _07454_);
  nor (_25509_, _25507_, _25506_);
  nor (_25510_, _25509_, _04082_);
  and (_25511_, _06617_, _05261_);
  nor (_25512_, _25484_, _04500_);
  not (_25513_, _25512_);
  nor (_25514_, _25513_, _25511_);
  nor (_25515_, _25514_, _25510_);
  nor (_25516_, _25515_, _03224_);
  nor (_25517_, _12164_, _10456_);
  or (_25518_, _25484_, _03521_);
  nor (_25520_, _25518_, _25517_);
  or (_25521_, _25520_, _03624_);
  nor (_25522_, _25521_, _25516_);
  and (_25523_, _05261_, _06350_);
  nor (_25524_, _25523_, _25484_);
  nand (_25525_, _25524_, _04527_);
  and (_25526_, _25525_, _08905_);
  nor (_25527_, _25526_, _25522_);
  and (_25528_, _12177_, _05261_);
  nor (_25529_, _25528_, _25484_);
  and (_25531_, _25529_, _03623_);
  nor (_25532_, _25531_, _25527_);
  nor (_25533_, _25532_, _03744_);
  and (_25534_, _12183_, _05261_);
  or (_25535_, _25484_, _03745_);
  nor (_25536_, _25535_, _25534_);
  or (_25537_, _25536_, _03611_);
  nor (_25538_, _25537_, _25533_);
  or (_25539_, _25524_, _04523_);
  nor (_25540_, _25539_, _25485_);
  nor (_25541_, _25540_, _25538_);
  nor (_25542_, _25541_, _03733_);
  and (_25543_, _12182_, _05261_);
  or (_25544_, _25543_, _25484_);
  and (_25545_, _25544_, _03733_);
  or (_25546_, _25545_, _25542_);
  and (_25547_, _25546_, _06453_);
  nor (_25548_, _12057_, _10456_);
  nor (_25549_, _25548_, _25484_);
  nor (_25550_, _25549_, _06453_);
  or (_25553_, _25550_, _25547_);
  and (_25554_, _25553_, _06458_);
  nor (_25555_, _12181_, _10456_);
  nor (_25556_, _25555_, _25484_);
  nor (_25557_, _25556_, _06458_);
  nor (_25558_, _25557_, _17198_);
  not (_25559_, _25558_);
  nor (_25560_, _25559_, _25554_);
  nor (_25561_, _25560_, _25488_);
  or (_25562_, _25561_, _43193_);
  or (_25564_, _43189_, \oc8051_golden_model_1.PCON [0]);
  and (_25565_, _25564_, _42003_);
  and (_43830_, _25565_, _25562_);
  and (_25566_, _06572_, _05261_);
  not (_25567_, \oc8051_golden_model_1.PCON [1]);
  nor (_25568_, _05261_, _25567_);
  nor (_25569_, _25568_, _04500_);
  not (_25570_, _25569_);
  nor (_25571_, _25570_, _25566_);
  not (_25572_, _25571_);
  nor (_25574_, _10456_, _04635_);
  nor (_25575_, _25574_, _25568_);
  and (_25576_, _25575_, _07454_);
  nor (_25577_, _05261_, \oc8051_golden_model_1.PCON [1]);
  and (_25578_, _05261_, _03269_);
  nor (_25579_, _25578_, _25577_);
  and (_25580_, _25579_, _04436_);
  nor (_25581_, _04436_, _25567_);
  or (_25582_, _25581_, _25580_);
  and (_25583_, _25582_, _04432_);
  and (_25585_, _12265_, _05261_);
  nor (_25586_, _25585_, _25577_);
  and (_25587_, _25586_, _03534_);
  or (_25588_, _25587_, _25583_);
  and (_25589_, _25588_, _04457_);
  nor (_25590_, _25575_, _04457_);
  nor (_25591_, _25590_, _25589_);
  nor (_25592_, _25591_, _03530_);
  and (_25593_, _25579_, _03530_);
  nor (_25594_, _25593_, _07454_);
  not (_25596_, _25594_);
  nor (_25597_, _25596_, _25592_);
  nor (_25598_, _25597_, _25576_);
  nor (_25599_, _25598_, _04082_);
  nor (_25600_, _25599_, _03224_);
  and (_25601_, _25600_, _25572_);
  not (_25602_, _25577_);
  and (_25603_, _12360_, _05261_);
  nor (_25604_, _25603_, _03521_);
  and (_25605_, _25604_, _25602_);
  nor (_25607_, _25605_, _25601_);
  nor (_25608_, _25607_, _08905_);
  nor (_25609_, _12375_, _10456_);
  nor (_25610_, _25609_, _04527_);
  and (_25611_, _05261_, _04325_);
  nor (_25612_, _25611_, _04509_);
  or (_25613_, _25612_, _25610_);
  and (_25614_, _25613_, _25602_);
  nor (_25615_, _25614_, _25608_);
  nor (_25616_, _25615_, _03744_);
  nor (_25618_, _12381_, _10456_);
  nor (_25619_, _25618_, _03745_);
  and (_25620_, _25619_, _25602_);
  nor (_25621_, _25620_, _25616_);
  nor (_25622_, _25621_, _03611_);
  nor (_25623_, _12374_, _10456_);
  nor (_25624_, _25623_, _04523_);
  and (_25625_, _25624_, _25602_);
  nor (_25626_, _25625_, _25622_);
  nor (_25627_, _25626_, _03733_);
  nor (_25629_, _25568_, _05674_);
  nor (_25630_, _25629_, _03734_);
  and (_25631_, _25630_, _25579_);
  nor (_25632_, _25631_, _25627_);
  or (_25633_, _25632_, _18526_);
  and (_25634_, _25611_, _05673_);
  or (_25635_, _25577_, _06453_);
  or (_25636_, _25635_, _25634_);
  and (_25637_, _25578_, _05673_);
  or (_25638_, _25577_, _06458_);
  or (_25640_, _25638_, _25637_);
  and (_25641_, _25640_, _03948_);
  and (_25642_, _25641_, _25636_);
  and (_25643_, _25642_, _25633_);
  nor (_25644_, _25586_, _03948_);
  nor (_25645_, _25644_, _25643_);
  and (_25646_, _25645_, _03474_);
  nor (_25647_, _25585_, _25568_);
  nor (_25648_, _25647_, _03474_);
  or (_25649_, _25648_, _25646_);
  or (_25651_, _25649_, _43193_);
  or (_25652_, _43189_, \oc8051_golden_model_1.PCON [1]);
  and (_25653_, _25652_, _42003_);
  and (_43831_, _25653_, _25651_);
  not (_25654_, \oc8051_golden_model_1.PCON [2]);
  nor (_25655_, _05261_, _25654_);
  nor (_25656_, _12587_, _10456_);
  nor (_25657_, _25656_, _25655_);
  nor (_25658_, _25657_, _06458_);
  nor (_25659_, _10456_, _05073_);
  nor (_25661_, _25659_, _25655_);
  and (_25662_, _25661_, _07454_);
  nor (_25663_, _12467_, _10456_);
  nor (_25664_, _25663_, _25655_);
  nor (_25665_, _25664_, _04432_);
  nor (_25666_, _04436_, _25654_);
  and (_25667_, _05261_, \oc8051_golden_model_1.ACC [2]);
  nor (_25668_, _25667_, _25655_);
  nor (_25669_, _25668_, _04437_);
  nor (_25670_, _25669_, _25666_);
  nor (_25672_, _25670_, _03534_);
  or (_25673_, _25672_, _25665_);
  and (_25674_, _25673_, _04457_);
  nor (_25675_, _25661_, _04457_);
  or (_25676_, _25675_, _25674_);
  and (_25677_, _25676_, _03531_);
  nor (_25678_, _25668_, _03531_);
  nor (_25679_, _25678_, _07454_);
  not (_25680_, _25679_);
  nor (_25681_, _25680_, _25677_);
  nor (_25683_, _25681_, _25662_);
  nor (_25684_, _25683_, _04082_);
  and (_25685_, _06710_, _05261_);
  nor (_25686_, _25655_, _04500_);
  not (_25687_, _25686_);
  nor (_25688_, _25687_, _25685_);
  nor (_25689_, _25688_, _25684_);
  nor (_25690_, _25689_, _03224_);
  nor (_25691_, _12568_, _10456_);
  or (_25692_, _25655_, _03521_);
  nor (_25694_, _25692_, _25691_);
  or (_25695_, _25694_, _03624_);
  nor (_25696_, _25695_, _25690_);
  and (_25697_, _05261_, _06399_);
  nor (_25698_, _25697_, _25655_);
  nand (_25699_, _25698_, _04527_);
  and (_25700_, _25699_, _08905_);
  nor (_25701_, _25700_, _25696_);
  and (_25702_, _12582_, _05261_);
  nor (_25703_, _25702_, _25655_);
  and (_25705_, _25703_, _03623_);
  nor (_25706_, _25705_, _25701_);
  nor (_25707_, _25706_, _03744_);
  and (_25708_, _12588_, _05261_);
  or (_25709_, _25655_, _03745_);
  nor (_25710_, _25709_, _25708_);
  or (_25711_, _25710_, _03611_);
  nor (_25712_, _25711_, _25707_);
  nor (_25713_, _25655_, _05772_);
  not (_25714_, _25713_);
  nor (_25716_, _25698_, _04523_);
  and (_25717_, _25716_, _25714_);
  nor (_25718_, _25717_, _25712_);
  nor (_25719_, _25718_, _03733_);
  nor (_25720_, _25668_, _03734_);
  and (_25721_, _25720_, _25714_);
  nor (_25722_, _25721_, _03618_);
  not (_25723_, _25722_);
  nor (_25724_, _25723_, _25719_);
  nor (_25725_, _12581_, _10456_);
  or (_25727_, _25655_, _06453_);
  nor (_25728_, _25727_, _25725_);
  or (_25729_, _25728_, _03741_);
  nor (_25730_, _25729_, _25724_);
  nor (_25731_, _25730_, _25658_);
  nor (_25732_, _25731_, _03767_);
  nor (_25733_, _25664_, _03948_);
  or (_25734_, _25733_, _03473_);
  nor (_25735_, _25734_, _25732_);
  and (_25736_, _12638_, _05261_);
  or (_25737_, _25655_, _03474_);
  nor (_25738_, _25737_, _25736_);
  nor (_25739_, _25738_, _25735_);
  or (_25740_, _25739_, _43193_);
  or (_25741_, _43189_, \oc8051_golden_model_1.PCON [2]);
  and (_25742_, _25741_, _42003_);
  and (_43832_, _25742_, _25740_);
  not (_25743_, \oc8051_golden_model_1.PCON [3]);
  nor (_25744_, _05261_, _25743_);
  nor (_25745_, _12792_, _10456_);
  nor (_25748_, _25745_, _25744_);
  nor (_25749_, _25748_, _06458_);
  and (_25750_, _12793_, _05261_);
  nor (_25751_, _25750_, _25744_);
  nor (_25752_, _25751_, _03745_);
  and (_25753_, _06664_, _05261_);
  or (_25754_, _25753_, _25744_);
  and (_25755_, _25754_, _04082_);
  and (_25756_, _05261_, \oc8051_golden_model_1.ACC [3]);
  nor (_25757_, _25756_, _25744_);
  nor (_25759_, _25757_, _03531_);
  nor (_25760_, _25757_, _04437_);
  nor (_25761_, _04436_, _25743_);
  or (_25762_, _25761_, _25760_);
  and (_25763_, _25762_, _04432_);
  nor (_25764_, _12652_, _10456_);
  nor (_25765_, _25764_, _25744_);
  nor (_25766_, _25765_, _04432_);
  or (_25767_, _25766_, _25763_);
  and (_25768_, _25767_, _04457_);
  nor (_25770_, _10456_, _04885_);
  nor (_25771_, _25770_, _25744_);
  nor (_25772_, _25771_, _04457_);
  nor (_25773_, _25772_, _25768_);
  nor (_25774_, _25773_, _03530_);
  or (_25775_, _25774_, _07454_);
  nor (_25776_, _25775_, _25759_);
  and (_25777_, _25771_, _07454_);
  or (_25778_, _25777_, _04082_);
  nor (_25779_, _25778_, _25776_);
  or (_25781_, _25779_, _25755_);
  and (_25782_, _25781_, _03521_);
  nor (_25783_, _12773_, _10456_);
  nor (_25784_, _25783_, _25744_);
  nor (_25785_, _25784_, _03521_);
  or (_25786_, _25785_, _08905_);
  or (_25787_, _25786_, _25782_);
  and (_25788_, _12787_, _05261_);
  or (_25789_, _25744_, _04527_);
  or (_25790_, _25789_, _25788_);
  and (_25792_, _05261_, _06356_);
  nor (_25793_, _25792_, _25744_);
  and (_25794_, _25793_, _03624_);
  nor (_25795_, _25794_, _03744_);
  and (_25796_, _25795_, _25790_);
  and (_25797_, _25796_, _25787_);
  nor (_25798_, _25797_, _25752_);
  nor (_25799_, _25798_, _03611_);
  nor (_25800_, _25744_, _05625_);
  not (_25801_, _25800_);
  nor (_25803_, _25793_, _04523_);
  and (_25804_, _25803_, _25801_);
  nor (_25805_, _25804_, _25799_);
  nor (_25806_, _25805_, _03733_);
  nor (_25807_, _25757_, _03734_);
  and (_25808_, _25807_, _25801_);
  or (_25809_, _25808_, _25806_);
  and (_25810_, _25809_, _06453_);
  nor (_25811_, _12786_, _10456_);
  nor (_25812_, _25811_, _25744_);
  nor (_25814_, _25812_, _06453_);
  or (_25815_, _25814_, _25810_);
  and (_25816_, _25815_, _06458_);
  nor (_25817_, _25816_, _25749_);
  nor (_25818_, _25817_, _03767_);
  nor (_25819_, _25765_, _03948_);
  or (_25820_, _25819_, _03473_);
  nor (_25821_, _25820_, _25818_);
  and (_25822_, _12843_, _05261_);
  nor (_25823_, _25822_, _25744_);
  and (_25825_, _25823_, _03473_);
  nor (_25826_, _25825_, _25821_);
  or (_25827_, _25826_, _43193_);
  or (_25828_, _43189_, \oc8051_golden_model_1.PCON [3]);
  and (_25829_, _25828_, _42003_);
  and (_43833_, _25829_, _25827_);
  not (_25830_, \oc8051_golden_model_1.PCON [4]);
  nor (_25831_, _05261_, _25830_);
  nor (_25832_, _12991_, _10456_);
  nor (_25833_, _25832_, _25831_);
  nor (_25835_, _25833_, _06458_);
  and (_25836_, _12992_, _05261_);
  nor (_25837_, _25836_, _25831_);
  nor (_25838_, _25837_, _03745_);
  and (_25839_, _06337_, _05261_);
  nor (_25840_, _25839_, _25831_);
  and (_25841_, _25840_, _03624_);
  nor (_25842_, _05831_, _10456_);
  nor (_25843_, _25842_, _25831_);
  and (_25844_, _25843_, _07454_);
  and (_25846_, _05261_, \oc8051_golden_model_1.ACC [4]);
  nor (_25847_, _25846_, _25831_);
  nor (_25848_, _25847_, _04437_);
  nor (_25849_, _04436_, _25830_);
  or (_25850_, _25849_, _25848_);
  and (_25851_, _25850_, _04432_);
  nor (_25852_, _12856_, _10456_);
  nor (_25853_, _25852_, _25831_);
  nor (_25854_, _25853_, _04432_);
  or (_25855_, _25854_, _25851_);
  and (_25857_, _25855_, _04457_);
  nor (_25858_, _25843_, _04457_);
  nor (_25859_, _25858_, _25857_);
  nor (_25860_, _25859_, _03530_);
  nor (_25861_, _25847_, _03531_);
  nor (_25862_, _25861_, _07454_);
  not (_25863_, _25862_);
  nor (_25864_, _25863_, _25860_);
  nor (_25865_, _25864_, _25844_);
  nor (_25866_, _25865_, _04082_);
  and (_25868_, _06802_, _05261_);
  nor (_25869_, _25831_, _04500_);
  not (_25870_, _25869_);
  nor (_25871_, _25870_, _25868_);
  or (_25872_, _25871_, _03224_);
  nor (_25873_, _25872_, _25866_);
  nor (_25874_, _12972_, _10456_);
  nor (_25875_, _25874_, _25831_);
  nor (_25876_, _25875_, _03521_);
  or (_25877_, _25876_, _03624_);
  nor (_25879_, _25877_, _25873_);
  nor (_25880_, _25879_, _25841_);
  or (_25881_, _25880_, _03623_);
  and (_25882_, _12986_, _05261_);
  or (_25883_, _25882_, _25831_);
  or (_25884_, _25883_, _04527_);
  and (_25885_, _25884_, _03745_);
  and (_25886_, _25885_, _25881_);
  nor (_25887_, _25886_, _25838_);
  nor (_25888_, _25887_, _03611_);
  nor (_25890_, _25831_, _05880_);
  not (_25891_, _25890_);
  nor (_25892_, _25840_, _04523_);
  and (_25893_, _25892_, _25891_);
  nor (_25894_, _25893_, _25888_);
  nor (_25895_, _25894_, _03733_);
  nor (_25896_, _25847_, _03734_);
  and (_25897_, _25896_, _25891_);
  or (_25898_, _25897_, _25895_);
  and (_25899_, _25898_, _06453_);
  nor (_25901_, _12985_, _10456_);
  nor (_25902_, _25901_, _25831_);
  nor (_25903_, _25902_, _06453_);
  or (_25904_, _25903_, _25899_);
  and (_25905_, _25904_, _06458_);
  nor (_25906_, _25905_, _25835_);
  nor (_25907_, _25906_, _03767_);
  nor (_25908_, _25853_, _03948_);
  or (_25909_, _25908_, _03473_);
  nor (_25910_, _25909_, _25907_);
  and (_25912_, _13051_, _05261_);
  or (_25913_, _25831_, _03474_);
  nor (_25914_, _25913_, _25912_);
  nor (_25915_, _25914_, _25910_);
  or (_25916_, _25915_, _43193_);
  or (_25917_, _43189_, \oc8051_golden_model_1.PCON [4]);
  and (_25918_, _25917_, _42003_);
  and (_43834_, _25918_, _25916_);
  not (_25919_, \oc8051_golden_model_1.PCON [5]);
  nor (_25920_, _05261_, _25919_);
  nor (_25922_, _13203_, _10456_);
  nor (_25923_, _25922_, _25920_);
  nor (_25924_, _25923_, _06458_);
  and (_25925_, _13204_, _05261_);
  nor (_25926_, _25925_, _25920_);
  nor (_25927_, _25926_, _03745_);
  and (_25928_, _06757_, _05261_);
  or (_25929_, _25928_, _25920_);
  and (_25930_, _25929_, _04082_);
  and (_25931_, _05261_, \oc8051_golden_model_1.ACC [5]);
  nor (_25933_, _25931_, _25920_);
  nor (_25934_, _25933_, _04437_);
  nor (_25935_, _04436_, _25919_);
  or (_25936_, _25935_, _25934_);
  and (_25937_, _25936_, _04432_);
  nor (_25938_, _13070_, _10456_);
  nor (_25939_, _25938_, _25920_);
  nor (_25940_, _25939_, _04432_);
  or (_25941_, _25940_, _25937_);
  and (_25942_, _25941_, _04457_);
  nor (_25944_, _05526_, _10456_);
  nor (_25945_, _25944_, _25920_);
  nor (_25946_, _25945_, _04457_);
  nor (_25947_, _25946_, _25942_);
  nor (_25948_, _25947_, _03530_);
  nor (_25949_, _25933_, _03531_);
  nor (_25950_, _25949_, _07454_);
  not (_25951_, _25950_);
  nor (_25952_, _25951_, _25948_);
  and (_25953_, _25945_, _07454_);
  or (_25955_, _25953_, _04082_);
  nor (_25956_, _25955_, _25952_);
  or (_25957_, _25956_, _25930_);
  and (_25958_, _25957_, _03521_);
  nor (_25959_, _13184_, _10456_);
  nor (_25960_, _25959_, _25920_);
  nor (_25961_, _25960_, _03521_);
  or (_25962_, _25961_, _08905_);
  or (_25963_, _25962_, _25958_);
  and (_25964_, _13198_, _05261_);
  or (_25966_, _25920_, _04527_);
  or (_25967_, _25966_, _25964_);
  and (_25968_, _06295_, _05261_);
  nor (_25969_, _25968_, _25920_);
  and (_25970_, _25969_, _03624_);
  nor (_25971_, _25970_, _03744_);
  and (_25972_, _25971_, _25967_);
  and (_25973_, _25972_, _25963_);
  nor (_25974_, _25973_, _25927_);
  nor (_25975_, _25974_, _03611_);
  nor (_25977_, _25920_, _05576_);
  not (_25978_, _25977_);
  nor (_25979_, _25969_, _04523_);
  and (_25980_, _25979_, _25978_);
  nor (_25981_, _25980_, _25975_);
  nor (_25982_, _25981_, _03733_);
  nor (_25983_, _25933_, _03734_);
  and (_25984_, _25983_, _25978_);
  nor (_25985_, _25984_, _03618_);
  not (_25986_, _25985_);
  nor (_25988_, _25986_, _25982_);
  nor (_25989_, _13197_, _10456_);
  or (_25990_, _25920_, _06453_);
  nor (_25991_, _25990_, _25989_);
  or (_25992_, _25991_, _03741_);
  nor (_25993_, _25992_, _25988_);
  nor (_25994_, _25993_, _25924_);
  nor (_25995_, _25994_, _03767_);
  nor (_25996_, _25939_, _03948_);
  or (_25997_, _25996_, _03473_);
  nor (_25999_, _25997_, _25995_);
  and (_26000_, _13253_, _05261_);
  or (_26001_, _25920_, _03474_);
  nor (_26002_, _26001_, _26000_);
  nor (_26003_, _26002_, _25999_);
  or (_26004_, _26003_, _43193_);
  or (_26005_, _43189_, \oc8051_golden_model_1.PCON [5]);
  and (_26006_, _26005_, _42003_);
  and (_43835_, _26006_, _26004_);
  not (_26007_, \oc8051_golden_model_1.PCON [6]);
  nor (_26009_, _05261_, _26007_);
  nor (_26010_, _13406_, _10456_);
  nor (_26011_, _26010_, _26009_);
  nor (_26012_, _26011_, _06458_);
  and (_26013_, _13407_, _05261_);
  nor (_26014_, _26013_, _26009_);
  nor (_26015_, _26014_, _03745_);
  and (_26016_, _06526_, _05261_);
  or (_26017_, _26016_, _26009_);
  and (_26018_, _26017_, _04082_);
  and (_26020_, _05261_, \oc8051_golden_model_1.ACC [6]);
  nor (_26021_, _26020_, _26009_);
  nor (_26022_, _26021_, _04437_);
  nor (_26023_, _04436_, _26007_);
  or (_26024_, _26023_, _26022_);
  and (_26025_, _26024_, _04432_);
  nor (_26026_, _13293_, _10456_);
  nor (_26027_, _26026_, _26009_);
  nor (_26028_, _26027_, _04432_);
  or (_26029_, _26028_, _26025_);
  and (_26031_, _26029_, _04457_);
  nor (_26032_, _05417_, _10456_);
  nor (_26033_, _26032_, _26009_);
  nor (_26034_, _26033_, _04457_);
  nor (_26035_, _26034_, _26031_);
  nor (_26036_, _26035_, _03530_);
  nor (_26037_, _26021_, _03531_);
  nor (_26038_, _26037_, _07454_);
  not (_26039_, _26038_);
  nor (_26040_, _26039_, _26036_);
  and (_26042_, _26033_, _07454_);
  or (_26043_, _26042_, _04082_);
  nor (_26044_, _26043_, _26040_);
  or (_26045_, _26044_, _26018_);
  and (_26046_, _26045_, _03521_);
  nor (_26047_, _13387_, _10456_);
  nor (_26048_, _26047_, _26009_);
  nor (_26049_, _26048_, _03521_);
  or (_26050_, _26049_, _08905_);
  or (_26051_, _26050_, _26046_);
  and (_26053_, _13402_, _05261_);
  or (_26054_, _26009_, _04527_);
  or (_26055_, _26054_, _26053_);
  and (_26056_, _14949_, _05261_);
  nor (_26057_, _26056_, _26009_);
  and (_26058_, _26057_, _03624_);
  nor (_26059_, _26058_, _03744_);
  and (_26060_, _26059_, _26055_);
  and (_26061_, _26060_, _26051_);
  nor (_26062_, _26061_, _26015_);
  nor (_26064_, _26062_, _03611_);
  nor (_26065_, _26009_, _05469_);
  not (_26066_, _26065_);
  nor (_26067_, _26057_, _04523_);
  and (_26068_, _26067_, _26066_);
  nor (_26069_, _26068_, _26064_);
  nor (_26070_, _26069_, _03733_);
  nor (_26071_, _26021_, _03734_);
  and (_26072_, _26071_, _26066_);
  or (_26073_, _26072_, _26070_);
  and (_26075_, _26073_, _06453_);
  nor (_26076_, _13400_, _10456_);
  nor (_26077_, _26076_, _26009_);
  nor (_26078_, _26077_, _06453_);
  or (_26079_, _26078_, _26075_);
  and (_26080_, _26079_, _06458_);
  nor (_26081_, _26080_, _26012_);
  nor (_26082_, _26081_, _03767_);
  nor (_26083_, _26027_, _03948_);
  or (_26084_, _26083_, _03473_);
  nor (_26085_, _26084_, _26082_);
  and (_26086_, _13456_, _05261_);
  or (_26087_, _26009_, _03474_);
  nor (_26088_, _26087_, _26086_);
  nor (_26089_, _26088_, _26085_);
  or (_26090_, _26089_, _43193_);
  or (_26091_, _43189_, \oc8051_golden_model_1.PCON [6]);
  and (_26092_, _26091_, _42003_);
  and (_43836_, _26092_, _26090_);
  not (_26093_, \oc8051_golden_model_1.SBUF [0]);
  nor (_26096_, _05270_, _26093_);
  nor (_26097_, _05722_, _10537_);
  nor (_26098_, _26097_, _26096_);
  and (_26099_, _26098_, _17198_);
  and (_26100_, _05270_, \oc8051_golden_model_1.ACC [0]);
  nor (_26101_, _26100_, _26096_);
  nor (_26102_, _26101_, _03531_);
  nor (_26103_, _26102_, _07454_);
  nor (_26104_, _26098_, _04432_);
  nor (_26105_, _04436_, _26093_);
  nor (_26107_, _26101_, _04437_);
  nor (_26108_, _26107_, _26105_);
  nor (_26109_, _26108_, _03534_);
  or (_26110_, _26109_, _03527_);
  nor (_26111_, _26110_, _26104_);
  or (_26112_, _26111_, _03530_);
  and (_26113_, _26112_, _26103_);
  and (_26114_, _05270_, _04429_);
  and (_26115_, _06903_, _04457_);
  or (_26116_, _26115_, _26096_);
  nor (_26118_, _26116_, _26114_);
  nor (_26119_, _26118_, _26113_);
  nor (_26120_, _26119_, _04082_);
  and (_26121_, _06617_, _05270_);
  nor (_26122_, _26096_, _04500_);
  not (_26123_, _26122_);
  nor (_26124_, _26123_, _26121_);
  nor (_26125_, _26124_, _26120_);
  nor (_26126_, _26125_, _03224_);
  nor (_26127_, _12164_, _10537_);
  or (_26129_, _26096_, _03521_);
  nor (_26130_, _26129_, _26127_);
  or (_26131_, _26130_, _03624_);
  nor (_26132_, _26131_, _26126_);
  and (_26133_, _05270_, _06350_);
  nor (_26134_, _26133_, _26096_);
  nand (_26135_, _26134_, _04527_);
  and (_26136_, _26135_, _08905_);
  nor (_26137_, _26136_, _26132_);
  and (_26138_, _12177_, _05270_);
  nor (_26140_, _26138_, _26096_);
  and (_26141_, _26140_, _03623_);
  nor (_26142_, _26141_, _26137_);
  nor (_26143_, _26142_, _03744_);
  and (_26144_, _12183_, _05270_);
  or (_26145_, _26096_, _03745_);
  nor (_26146_, _26145_, _26144_);
  or (_26147_, _26146_, _03611_);
  nor (_26148_, _26147_, _26143_);
  or (_26149_, _26134_, _04523_);
  nor (_26151_, _26149_, _26097_);
  nor (_26152_, _26151_, _26148_);
  nor (_26153_, _26152_, _03733_);
  nor (_26154_, _26096_, _05722_);
  or (_26155_, _26154_, _03734_);
  nor (_26156_, _26155_, _26101_);
  or (_26157_, _26156_, _26153_);
  and (_26158_, _26157_, _06453_);
  nor (_26159_, _12057_, _10537_);
  nor (_26160_, _26159_, _26096_);
  nor (_26162_, _26160_, _06453_);
  or (_26163_, _26162_, _26158_);
  and (_26164_, _26163_, _06458_);
  nor (_26165_, _12181_, _10537_);
  nor (_26166_, _26165_, _26096_);
  nor (_26167_, _26166_, _06458_);
  nor (_26168_, _26167_, _17198_);
  not (_26169_, _26168_);
  nor (_26170_, _26169_, _26164_);
  nor (_26171_, _26170_, _26099_);
  or (_26173_, _26171_, _43193_);
  or (_26174_, _43189_, \oc8051_golden_model_1.SBUF [0]);
  and (_26175_, _26174_, _42003_);
  and (_43839_, _26175_, _26173_);
  and (_26176_, _06572_, _05270_);
  not (_26177_, \oc8051_golden_model_1.SBUF [1]);
  nor (_26178_, _05270_, _26177_);
  nor (_26179_, _26178_, _04500_);
  not (_26180_, _26179_);
  nor (_26181_, _26180_, _26176_);
  not (_26183_, _26181_);
  nor (_26184_, _10537_, _04635_);
  nor (_26185_, _26184_, _26178_);
  and (_26186_, _26185_, _07454_);
  nor (_26187_, _05270_, \oc8051_golden_model_1.SBUF [1]);
  and (_26188_, _05270_, _03269_);
  nor (_26189_, _26188_, _26187_);
  and (_26190_, _26189_, _04436_);
  nor (_26191_, _04436_, _26177_);
  or (_26192_, _26191_, _26190_);
  and (_26193_, _26192_, _04432_);
  and (_26194_, _12265_, _05270_);
  nor (_26195_, _26194_, _26187_);
  and (_26196_, _26195_, _03534_);
  or (_26197_, _26196_, _26193_);
  and (_26198_, _26197_, _04457_);
  nor (_26199_, _26185_, _04457_);
  nor (_26200_, _26199_, _26198_);
  nor (_26201_, _26200_, _03530_);
  and (_26202_, _26189_, _03530_);
  nor (_26205_, _26202_, _07454_);
  not (_26206_, _26205_);
  nor (_26207_, _26206_, _26201_);
  nor (_26208_, _26207_, _26186_);
  nor (_26209_, _26208_, _04082_);
  nor (_26210_, _26209_, _03224_);
  and (_26211_, _26210_, _26183_);
  not (_26212_, _26187_);
  and (_26213_, _12360_, _05270_);
  nor (_26214_, _26213_, _03521_);
  and (_26216_, _26214_, _26212_);
  nor (_26217_, _26216_, _26211_);
  nor (_26218_, _26217_, _08905_);
  nor (_26219_, _12375_, _10537_);
  nor (_26220_, _26219_, _04527_);
  and (_26221_, _05270_, _04325_);
  nor (_26222_, _26221_, _04509_);
  nor (_26223_, _26222_, _26220_);
  nor (_26224_, _26223_, _26187_);
  nor (_26225_, _26224_, _26218_);
  nor (_26227_, _26225_, _03744_);
  nor (_26228_, _12381_, _10537_);
  nor (_26229_, _26228_, _03745_);
  and (_26230_, _26229_, _26212_);
  nor (_26231_, _26230_, _26227_);
  nor (_26232_, _26231_, _03611_);
  nor (_26233_, _12374_, _10537_);
  nor (_26234_, _26233_, _04523_);
  and (_26235_, _26234_, _26212_);
  nor (_26236_, _26235_, _26232_);
  nor (_26238_, _26236_, _03733_);
  nor (_26239_, _26178_, _05674_);
  nor (_26240_, _26239_, _03734_);
  and (_26241_, _26240_, _26189_);
  nor (_26242_, _26241_, _26238_);
  or (_26243_, _26242_, _18526_);
  and (_26244_, _26221_, _05673_);
  nor (_26245_, _26244_, _06453_);
  and (_26246_, _26245_, _26212_);
  nand (_26247_, _26188_, _05673_);
  nor (_26249_, _26187_, _06458_);
  and (_26250_, _26249_, _26247_);
  or (_26251_, _26250_, _03767_);
  nor (_26252_, _26251_, _26246_);
  and (_26253_, _26252_, _26243_);
  nor (_26254_, _26195_, _03948_);
  nor (_26255_, _26254_, _26253_);
  and (_26256_, _26255_, _03474_);
  nor (_26257_, _26194_, _26178_);
  nor (_26258_, _26257_, _03474_);
  or (_26260_, _26258_, _26256_);
  or (_26261_, _26260_, _43193_);
  or (_26262_, _43189_, \oc8051_golden_model_1.SBUF [1]);
  and (_26263_, _26262_, _42003_);
  and (_43840_, _26263_, _26261_);
  not (_26264_, \oc8051_golden_model_1.SBUF [2]);
  nor (_26265_, _05270_, _26264_);
  nor (_26266_, _12587_, _10537_);
  nor (_26267_, _26266_, _26265_);
  nor (_26268_, _26267_, _06458_);
  nor (_26270_, _10537_, _05073_);
  nor (_26271_, _26270_, _26265_);
  and (_26272_, _26271_, _07454_);
  nor (_26273_, _12467_, _10537_);
  nor (_26274_, _26273_, _26265_);
  nor (_26275_, _26274_, _04432_);
  nor (_26276_, _04436_, _26264_);
  and (_26277_, _05270_, \oc8051_golden_model_1.ACC [2]);
  nor (_26278_, _26277_, _26265_);
  nor (_26279_, _26278_, _04437_);
  nor (_26281_, _26279_, _26276_);
  nor (_26282_, _26281_, _03534_);
  or (_26283_, _26282_, _26275_);
  and (_26284_, _26283_, _04457_);
  nor (_26285_, _26271_, _04457_);
  or (_26286_, _26285_, _26284_);
  and (_26287_, _26286_, _03531_);
  nor (_26288_, _26278_, _03531_);
  nor (_26289_, _26288_, _07454_);
  not (_26290_, _26289_);
  nor (_26292_, _26290_, _26287_);
  nor (_26293_, _26292_, _26272_);
  nor (_26294_, _26293_, _04082_);
  and (_26295_, _06710_, _05270_);
  nor (_26296_, _26265_, _04500_);
  not (_26297_, _26296_);
  nor (_26298_, _26297_, _26295_);
  nor (_26299_, _26298_, _26294_);
  nor (_26300_, _26299_, _03224_);
  nor (_26301_, _12568_, _10537_);
  or (_26303_, _26265_, _03521_);
  nor (_26304_, _26303_, _26301_);
  or (_26305_, _26304_, _03624_);
  nor (_26306_, _26305_, _26300_);
  and (_26307_, _05270_, _06399_);
  nor (_26308_, _26307_, _26265_);
  nand (_26309_, _26308_, _04527_);
  and (_26310_, _26309_, _08905_);
  nor (_26311_, _26310_, _26306_);
  and (_26312_, _12582_, _05270_);
  nor (_26314_, _26312_, _26265_);
  and (_26315_, _26314_, _03623_);
  nor (_26316_, _26315_, _26311_);
  nor (_26317_, _26316_, _03744_);
  and (_26318_, _12588_, _05270_);
  or (_26319_, _26265_, _03745_);
  nor (_26320_, _26319_, _26318_);
  or (_26321_, _26320_, _03611_);
  nor (_26322_, _26321_, _26317_);
  nor (_26323_, _26265_, _05772_);
  not (_26325_, _26323_);
  nor (_26326_, _26308_, _04523_);
  and (_26327_, _26326_, _26325_);
  nor (_26328_, _26327_, _26322_);
  nor (_26329_, _26328_, _03733_);
  nor (_26330_, _26278_, _03734_);
  and (_26331_, _26330_, _26325_);
  nor (_26332_, _26331_, _03618_);
  not (_26333_, _26332_);
  nor (_26334_, _26333_, _26329_);
  nor (_26336_, _12581_, _10537_);
  or (_26337_, _26265_, _06453_);
  nor (_26338_, _26337_, _26336_);
  or (_26339_, _26338_, _03741_);
  nor (_26340_, _26339_, _26334_);
  nor (_26341_, _26340_, _26268_);
  nor (_26342_, _26341_, _03767_);
  nor (_26343_, _26274_, _03948_);
  or (_26344_, _26343_, _03473_);
  nor (_26345_, _26344_, _26342_);
  and (_26347_, _12638_, _05270_);
  or (_26348_, _26265_, _03474_);
  nor (_26349_, _26348_, _26347_);
  nor (_26350_, _26349_, _26345_);
  or (_26351_, _26350_, _43193_);
  or (_26352_, _43189_, \oc8051_golden_model_1.SBUF [2]);
  and (_26353_, _26352_, _42003_);
  and (_43841_, _26353_, _26351_);
  not (_26354_, \oc8051_golden_model_1.SBUF [3]);
  nor (_26355_, _05270_, _26354_);
  nor (_26357_, _12792_, _10537_);
  nor (_26358_, _26357_, _26355_);
  nor (_26359_, _26358_, _06458_);
  and (_26360_, _12793_, _05270_);
  nor (_26361_, _26360_, _26355_);
  nor (_26362_, _26361_, _03745_);
  and (_26363_, _06664_, _05270_);
  or (_26364_, _26363_, _26355_);
  and (_26365_, _26364_, _04082_);
  and (_26366_, _05270_, \oc8051_golden_model_1.ACC [3]);
  nor (_26368_, _26366_, _26355_);
  nor (_26369_, _26368_, _04437_);
  nor (_26370_, _04436_, _26354_);
  or (_26371_, _26370_, _26369_);
  and (_26372_, _26371_, _04432_);
  nor (_26373_, _12652_, _10537_);
  nor (_26374_, _26373_, _26355_);
  nor (_26375_, _26374_, _04432_);
  or (_26376_, _26375_, _26372_);
  and (_26377_, _26376_, _04457_);
  nor (_26379_, _10537_, _04885_);
  nor (_26380_, _26379_, _26355_);
  nor (_26381_, _26380_, _04457_);
  nor (_26382_, _26381_, _26377_);
  nor (_26383_, _26382_, _03530_);
  nor (_26384_, _26368_, _03531_);
  nor (_26385_, _26384_, _07454_);
  not (_26386_, _26385_);
  nor (_26387_, _26386_, _26383_);
  and (_26388_, _26380_, _07454_);
  or (_26390_, _26388_, _04082_);
  nor (_26391_, _26390_, _26387_);
  or (_26392_, _26391_, _26365_);
  and (_26393_, _26392_, _03521_);
  nor (_26394_, _12773_, _10537_);
  nor (_26395_, _26394_, _26355_);
  nor (_26396_, _26395_, _03521_);
  or (_26397_, _26396_, _08905_);
  or (_26398_, _26397_, _26393_);
  and (_26399_, _12787_, _05270_);
  or (_26401_, _26355_, _04527_);
  or (_26402_, _26401_, _26399_);
  and (_26403_, _05270_, _06356_);
  nor (_26404_, _26403_, _26355_);
  and (_26405_, _26404_, _03624_);
  nor (_26406_, _26405_, _03744_);
  and (_26407_, _26406_, _26402_);
  and (_26408_, _26407_, _26398_);
  nor (_26409_, _26408_, _26362_);
  nor (_26410_, _26409_, _03611_);
  nor (_26412_, _26355_, _05625_);
  not (_26413_, _26412_);
  nor (_26414_, _26404_, _04523_);
  and (_26415_, _26414_, _26413_);
  nor (_26416_, _26415_, _26410_);
  nor (_26417_, _26416_, _03733_);
  nor (_26418_, _26368_, _03734_);
  and (_26419_, _26418_, _26413_);
  nor (_26420_, _26419_, _03618_);
  not (_26421_, _26420_);
  nor (_26423_, _26421_, _26417_);
  nor (_26424_, _12786_, _10537_);
  or (_26425_, _26355_, _06453_);
  nor (_26426_, _26425_, _26424_);
  or (_26427_, _26426_, _03741_);
  nor (_26428_, _26427_, _26423_);
  nor (_26429_, _26428_, _26359_);
  nor (_26430_, _26429_, _03767_);
  nor (_26431_, _26374_, _03948_);
  or (_26432_, _26431_, _03473_);
  nor (_26434_, _26432_, _26430_);
  and (_26435_, _12843_, _05270_);
  or (_26436_, _26355_, _03474_);
  nor (_26437_, _26436_, _26435_);
  nor (_26438_, _26437_, _26434_);
  or (_26439_, _26438_, _43193_);
  or (_26440_, _43189_, \oc8051_golden_model_1.SBUF [3]);
  and (_26441_, _26440_, _42003_);
  and (_43842_, _26441_, _26439_);
  not (_26442_, \oc8051_golden_model_1.SBUF [4]);
  nor (_26444_, _05270_, _26442_);
  nor (_26445_, _12991_, _10537_);
  nor (_26446_, _26445_, _26444_);
  nor (_26447_, _26446_, _06458_);
  and (_26448_, _12992_, _05270_);
  nor (_26449_, _26448_, _26444_);
  nor (_26450_, _26449_, _03745_);
  and (_26451_, _06337_, _05270_);
  nor (_26452_, _26451_, _26444_);
  and (_26453_, _26452_, _03624_);
  nor (_26455_, _05831_, _10537_);
  nor (_26456_, _26455_, _26444_);
  and (_26457_, _26456_, _07454_);
  and (_26458_, _05270_, \oc8051_golden_model_1.ACC [4]);
  nor (_26459_, _26458_, _26444_);
  nor (_26460_, _26459_, _04437_);
  nor (_26461_, _04436_, _26442_);
  or (_26462_, _26461_, _26460_);
  and (_26463_, _26462_, _04432_);
  nor (_26464_, _12856_, _10537_);
  nor (_26466_, _26464_, _26444_);
  nor (_26467_, _26466_, _04432_);
  or (_26468_, _26467_, _26463_);
  and (_26469_, _26468_, _04457_);
  nor (_26470_, _26456_, _04457_);
  nor (_26471_, _26470_, _26469_);
  nor (_26472_, _26471_, _03530_);
  nor (_26473_, _26459_, _03531_);
  nor (_26474_, _26473_, _07454_);
  not (_26475_, _26474_);
  nor (_26477_, _26475_, _26472_);
  nor (_26478_, _26477_, _26457_);
  nor (_26479_, _26478_, _04082_);
  and (_26480_, _06802_, _05270_);
  nor (_26481_, _26444_, _04500_);
  not (_26482_, _26481_);
  nor (_26483_, _26482_, _26480_);
  or (_26484_, _26483_, _03224_);
  nor (_26485_, _26484_, _26479_);
  nor (_26486_, _12972_, _10537_);
  nor (_26488_, _26486_, _26444_);
  nor (_26489_, _26488_, _03521_);
  or (_26490_, _26489_, _03624_);
  nor (_26491_, _26490_, _26485_);
  nor (_26492_, _26491_, _26453_);
  or (_26493_, _26492_, _03623_);
  and (_26494_, _12986_, _05270_);
  or (_26495_, _26494_, _26444_);
  or (_26496_, _26495_, _04527_);
  and (_26497_, _26496_, _03745_);
  and (_26499_, _26497_, _26493_);
  nor (_26500_, _26499_, _26450_);
  nor (_26501_, _26500_, _03611_);
  nor (_26502_, _26444_, _05880_);
  not (_26503_, _26502_);
  nor (_26504_, _26452_, _04523_);
  and (_26505_, _26504_, _26503_);
  nor (_26506_, _26505_, _26501_);
  nor (_26507_, _26506_, _03733_);
  nor (_26508_, _26459_, _03734_);
  and (_26510_, _26508_, _26503_);
  nor (_26511_, _26510_, _03618_);
  not (_26512_, _26511_);
  nor (_26513_, _26512_, _26507_);
  nor (_26514_, _12985_, _10537_);
  or (_26515_, _26444_, _06453_);
  nor (_26516_, _26515_, _26514_);
  or (_26517_, _26516_, _03741_);
  nor (_26518_, _26517_, _26513_);
  nor (_26519_, _26518_, _26447_);
  nor (_26521_, _26519_, _03767_);
  nor (_26522_, _26466_, _03948_);
  or (_26523_, _26522_, _03473_);
  nor (_26524_, _26523_, _26521_);
  and (_26525_, _13051_, _05270_);
  or (_26526_, _26444_, _03474_);
  nor (_26527_, _26526_, _26525_);
  nor (_26528_, _26527_, _26524_);
  or (_26529_, _26528_, _43193_);
  or (_26530_, _43189_, \oc8051_golden_model_1.SBUF [4]);
  and (_26532_, _26530_, _42003_);
  and (_43845_, _26532_, _26529_);
  not (_26533_, \oc8051_golden_model_1.SBUF [5]);
  nor (_26534_, _05270_, _26533_);
  nor (_26535_, _13203_, _10537_);
  nor (_26536_, _26535_, _26534_);
  nor (_26537_, _26536_, _06458_);
  and (_26538_, _13204_, _05270_);
  nor (_26539_, _26538_, _26534_);
  nor (_26540_, _26539_, _03745_);
  and (_26542_, _06757_, _05270_);
  or (_26543_, _26542_, _26534_);
  and (_26544_, _26543_, _04082_);
  and (_26545_, _05270_, \oc8051_golden_model_1.ACC [5]);
  nor (_26546_, _26545_, _26534_);
  nor (_26547_, _26546_, _03531_);
  nor (_26548_, _26546_, _04437_);
  nor (_26549_, _04436_, _26533_);
  or (_26550_, _26549_, _26548_);
  and (_26551_, _26550_, _04432_);
  nor (_26553_, _13070_, _10537_);
  nor (_26554_, _26553_, _26534_);
  nor (_26555_, _26554_, _04432_);
  or (_26556_, _26555_, _26551_);
  and (_26557_, _26556_, _04457_);
  nor (_26558_, _05526_, _10537_);
  nor (_26559_, _26558_, _26534_);
  nor (_26560_, _26559_, _04457_);
  nor (_26561_, _26560_, _26557_);
  nor (_26562_, _26561_, _03530_);
  or (_26564_, _26562_, _07454_);
  nor (_26565_, _26564_, _26547_);
  and (_26566_, _26559_, _07454_);
  or (_26567_, _26566_, _04082_);
  nor (_26568_, _26567_, _26565_);
  or (_26569_, _26568_, _26544_);
  and (_26570_, _26569_, _03521_);
  nor (_26571_, _13184_, _10537_);
  nor (_26572_, _26571_, _26534_);
  nor (_26573_, _26572_, _03521_);
  or (_26575_, _26573_, _08905_);
  or (_26576_, _26575_, _26570_);
  and (_26577_, _13198_, _05270_);
  or (_26578_, _26534_, _04527_);
  or (_26579_, _26578_, _26577_);
  and (_26580_, _06295_, _05270_);
  nor (_26581_, _26580_, _26534_);
  and (_26582_, _26581_, _03624_);
  nor (_26583_, _26582_, _03744_);
  and (_26584_, _26583_, _26579_);
  and (_26586_, _26584_, _26576_);
  nor (_26587_, _26586_, _26540_);
  nor (_26588_, _26587_, _03611_);
  nor (_26589_, _26534_, _05576_);
  not (_26590_, _26589_);
  nor (_26591_, _26581_, _04523_);
  and (_26592_, _26591_, _26590_);
  nor (_26593_, _26592_, _26588_);
  nor (_26594_, _26593_, _03733_);
  nor (_26595_, _26546_, _03734_);
  and (_26597_, _26595_, _26590_);
  nor (_26598_, _26597_, _03618_);
  not (_26599_, _26598_);
  nor (_26600_, _26599_, _26594_);
  nor (_26601_, _13197_, _10537_);
  or (_26602_, _26534_, _06453_);
  nor (_26603_, _26602_, _26601_);
  or (_26604_, _26603_, _03741_);
  nor (_26605_, _26604_, _26600_);
  nor (_26606_, _26605_, _26537_);
  nor (_26608_, _26606_, _03767_);
  nor (_26609_, _26554_, _03948_);
  or (_26610_, _26609_, _03473_);
  nor (_26611_, _26610_, _26608_);
  and (_26612_, _13253_, _05270_);
  or (_26613_, _26534_, _03474_);
  nor (_26614_, _26613_, _26612_);
  nor (_26615_, _26614_, _26611_);
  or (_26616_, _26615_, _43193_);
  or (_26617_, _43189_, \oc8051_golden_model_1.SBUF [5]);
  and (_26619_, _26617_, _42003_);
  and (_43846_, _26619_, _26616_);
  not (_26620_, \oc8051_golden_model_1.SBUF [6]);
  nor (_26621_, _05270_, _26620_);
  nor (_26622_, _13406_, _10537_);
  nor (_26623_, _26622_, _26621_);
  nor (_26624_, _26623_, _06458_);
  and (_26625_, _13407_, _05270_);
  nor (_26626_, _26625_, _26621_);
  nor (_26627_, _26626_, _03745_);
  and (_26629_, _06526_, _05270_);
  or (_26630_, _26629_, _26621_);
  and (_26631_, _26630_, _04082_);
  and (_26632_, _05270_, \oc8051_golden_model_1.ACC [6]);
  nor (_26633_, _26632_, _26621_);
  nor (_26634_, _26633_, _04437_);
  nor (_26635_, _04436_, _26620_);
  or (_26636_, _26635_, _26634_);
  and (_26637_, _26636_, _04432_);
  nor (_26638_, _13293_, _10537_);
  nor (_26639_, _26638_, _26621_);
  nor (_26640_, _26639_, _04432_);
  or (_26641_, _26640_, _26637_);
  and (_26642_, _26641_, _04457_);
  nor (_26643_, _05417_, _10537_);
  nor (_26644_, _26643_, _26621_);
  nor (_26645_, _26644_, _04457_);
  nor (_26646_, _26645_, _26642_);
  nor (_26647_, _26646_, _03530_);
  nor (_26648_, _26633_, _03531_);
  nor (_26651_, _26648_, _07454_);
  not (_26652_, _26651_);
  nor (_26653_, _26652_, _26647_);
  and (_26654_, _26644_, _07454_);
  or (_26655_, _26654_, _04082_);
  nor (_26656_, _26655_, _26653_);
  or (_26657_, _26656_, _26631_);
  and (_26658_, _26657_, _03521_);
  nor (_26659_, _13387_, _10537_);
  nor (_26660_, _26659_, _26621_);
  nor (_26662_, _26660_, _03521_);
  or (_26663_, _26662_, _08905_);
  or (_26664_, _26663_, _26658_);
  and (_26665_, _13402_, _05270_);
  or (_26666_, _26621_, _04527_);
  or (_26667_, _26666_, _26665_);
  and (_26668_, _14949_, _05270_);
  nor (_26669_, _26668_, _26621_);
  and (_26670_, _26669_, _03624_);
  nor (_26671_, _26670_, _03744_);
  and (_26673_, _26671_, _26667_);
  and (_26674_, _26673_, _26664_);
  nor (_26675_, _26674_, _26627_);
  nor (_26676_, _26675_, _03611_);
  nor (_26677_, _26621_, _05469_);
  not (_26678_, _26677_);
  nor (_26679_, _26669_, _04523_);
  and (_26680_, _26679_, _26678_);
  nor (_26681_, _26680_, _26676_);
  nor (_26682_, _26681_, _03733_);
  nor (_26684_, _26633_, _03734_);
  and (_26685_, _26684_, _26678_);
  nor (_26686_, _26685_, _03618_);
  not (_26687_, _26686_);
  nor (_26688_, _26687_, _26682_);
  nor (_26689_, _13400_, _10537_);
  or (_26690_, _26621_, _06453_);
  nor (_26691_, _26690_, _26689_);
  or (_26692_, _26691_, _03741_);
  nor (_26693_, _26692_, _26688_);
  nor (_26695_, _26693_, _26624_);
  nor (_26696_, _26695_, _03767_);
  nor (_26697_, _26639_, _03948_);
  or (_26698_, _26697_, _03473_);
  nor (_26699_, _26698_, _26696_);
  and (_26700_, _13456_, _05270_);
  or (_26701_, _26621_, _03474_);
  nor (_26702_, _26701_, _26700_);
  nor (_26703_, _26702_, _26699_);
  or (_26704_, _26703_, _43193_);
  or (_26706_, _43189_, \oc8051_golden_model_1.SBUF [6]);
  and (_26707_, _26706_, _42003_);
  and (_43847_, _26707_, _26704_);
  not (_26708_, \oc8051_golden_model_1.SCON [0]);
  nor (_26709_, _05333_, _26708_);
  and (_26710_, _12183_, _05333_);
  nor (_26711_, _26710_, _26709_);
  nor (_26712_, _26711_, _03745_);
  and (_26713_, _05333_, _06350_);
  nor (_26714_, _26713_, _26709_);
  and (_26716_, _26714_, _03624_);
  and (_26717_, _05333_, _04429_);
  nor (_26718_, _26717_, _26709_);
  and (_26719_, _26718_, _07454_);
  and (_26720_, _05333_, \oc8051_golden_model_1.ACC [0]);
  nor (_26721_, _26720_, _26709_);
  nor (_26722_, _26721_, _04437_);
  nor (_26723_, _04436_, _26708_);
  or (_26724_, _26723_, _26722_);
  and (_26725_, _26724_, _04432_);
  nor (_26727_, _05722_, _10618_);
  nor (_26728_, _26727_, _26709_);
  nor (_26729_, _26728_, _04432_);
  or (_26730_, _26729_, _26725_);
  and (_26731_, _26730_, _03470_);
  nor (_26732_, _05942_, _26708_);
  and (_26733_, _12075_, _05942_);
  nor (_26734_, _26733_, _26732_);
  nor (_26735_, _26734_, _03470_);
  nor (_26736_, _26735_, _26731_);
  nor (_26738_, _26736_, _03527_);
  nor (_26739_, _26718_, _04457_);
  or (_26740_, _26739_, _26738_);
  and (_26741_, _26740_, _03531_);
  nor (_26742_, _26721_, _03531_);
  or (_26743_, _26742_, _26741_);
  and (_26744_, _26743_, _03466_);
  and (_26745_, _26709_, _03465_);
  or (_26746_, _26745_, _26744_);
  and (_26747_, _26746_, _03459_);
  nor (_26749_, _26728_, _03459_);
  or (_26750_, _26749_, _26747_);
  and (_26751_, _26750_, _03453_);
  nor (_26752_, _12106_, _10655_);
  nor (_26753_, _26752_, _26732_);
  nor (_26754_, _26753_, _03453_);
  or (_26755_, _26754_, _07454_);
  nor (_26756_, _26755_, _26751_);
  nor (_26757_, _26756_, _26719_);
  nor (_26758_, _26757_, _04082_);
  and (_26760_, _06617_, _05333_);
  nor (_26761_, _26709_, _04500_);
  not (_26762_, _26761_);
  nor (_26763_, _26762_, _26760_);
  or (_26764_, _26763_, _03224_);
  nor (_26765_, _26764_, _26758_);
  nor (_26766_, _12164_, _10618_);
  nor (_26767_, _26766_, _26709_);
  nor (_26768_, _26767_, _03521_);
  or (_26769_, _26768_, _03624_);
  nor (_26771_, _26769_, _26765_);
  nor (_26772_, _26771_, _26716_);
  or (_26773_, _26772_, _03623_);
  and (_26774_, _12177_, _05333_);
  or (_26775_, _26774_, _26709_);
  or (_26776_, _26775_, _04527_);
  and (_26777_, _26776_, _03745_);
  and (_26778_, _26777_, _26773_);
  nor (_26779_, _26778_, _26712_);
  nor (_26780_, _26779_, _03611_);
  or (_26782_, _26714_, _04523_);
  nor (_26783_, _26782_, _26727_);
  nor (_26784_, _26783_, _26780_);
  nor (_26785_, _26784_, _03733_);
  and (_26786_, _12182_, _05333_);
  or (_26787_, _26786_, _26709_);
  and (_26788_, _26787_, _03733_);
  or (_26789_, _26788_, _26785_);
  and (_26790_, _26789_, _06453_);
  nor (_26791_, _12057_, _10618_);
  nor (_26793_, _26791_, _26709_);
  nor (_26794_, _26793_, _06453_);
  or (_26795_, _26794_, _26790_);
  and (_26796_, _26795_, _06458_);
  nor (_26797_, _12181_, _10618_);
  nor (_26798_, _26797_, _26709_);
  nor (_26799_, _26798_, _06458_);
  or (_26800_, _26799_, _26796_);
  and (_26801_, _26800_, _03948_);
  nor (_26802_, _26728_, _03948_);
  or (_26804_, _26802_, _26801_);
  and (_26805_, _26804_, _03446_);
  and (_26806_, _26709_, _03445_);
  or (_26807_, _26806_, _26805_);
  and (_26808_, _26807_, _03474_);
  nor (_26809_, _26728_, _03474_);
  or (_26810_, _26809_, _26808_);
  or (_26811_, _26810_, _43193_);
  or (_26812_, _43189_, \oc8051_golden_model_1.SCON [0]);
  and (_26813_, _26812_, _42003_);
  and (_43848_, _26813_, _26811_);
  not (_26815_, \oc8051_golden_model_1.SCON [1]);
  nor (_26816_, _05333_, _26815_);
  and (_26817_, _06572_, _05333_);
  or (_26818_, _26817_, _26816_);
  and (_26819_, _26818_, _04082_);
  nor (_26820_, _05333_, \oc8051_golden_model_1.SCON [1]);
  and (_26821_, _05333_, _03269_);
  nor (_26822_, _26821_, _26820_);
  and (_26823_, _26822_, _04436_);
  nor (_26825_, _04436_, _26815_);
  or (_26826_, _26825_, _26823_);
  and (_26827_, _26826_, _04432_);
  and (_26828_, _12265_, _05333_);
  nor (_26829_, _26828_, _26820_);
  and (_26830_, _26829_, _03534_);
  or (_26831_, _26830_, _26827_);
  and (_26832_, _26831_, _03470_);
  and (_26833_, _12269_, _05942_);
  nor (_26834_, _05942_, _26815_);
  or (_26836_, _26834_, _03527_);
  or (_26837_, _26836_, _26833_);
  and (_26838_, _26837_, _03533_);
  nor (_26839_, _26838_, _26832_);
  nor (_26840_, _10618_, _04635_);
  nor (_26841_, _26840_, _26816_);
  and (_26842_, _26841_, _03527_);
  nor (_26843_, _26842_, _26839_);
  and (_26844_, _26843_, _03531_);
  and (_26845_, _26822_, _03530_);
  or (_26847_, _26845_, _26844_);
  and (_26848_, _26847_, _03466_);
  and (_26849_, _12256_, _05942_);
  nor (_26850_, _26849_, _26834_);
  nor (_26851_, _26850_, _03466_);
  or (_26852_, _26851_, _26848_);
  and (_26853_, _26852_, _03459_);
  and (_26854_, _26833_, _12284_);
  or (_26855_, _26854_, _26834_);
  and (_26856_, _26855_, _03458_);
  or (_26858_, _26856_, _26853_);
  and (_26859_, _26858_, _03453_);
  nor (_26860_, _12301_, _10655_);
  nor (_26861_, _26834_, _26860_);
  nor (_26862_, _26861_, _03453_);
  or (_26863_, _26862_, _07454_);
  nor (_26864_, _26863_, _26859_);
  and (_26865_, _26841_, _07454_);
  or (_26866_, _26865_, _04082_);
  nor (_26867_, _26866_, _26864_);
  or (_26869_, _26867_, _26819_);
  and (_26870_, _26869_, _03521_);
  nor (_26871_, _12360_, _10618_);
  nor (_26872_, _26871_, _26816_);
  nor (_26873_, _26872_, _03521_);
  nor (_26874_, _26873_, _26870_);
  nor (_26875_, _26874_, _08905_);
  not (_26876_, _26820_);
  nor (_26877_, _12375_, _10618_);
  nor (_26878_, _26877_, _04527_);
  and (_26880_, _05333_, _04325_);
  nor (_26881_, _26880_, _04509_);
  or (_26882_, _26881_, _26878_);
  and (_26883_, _26882_, _26876_);
  nor (_26884_, _26883_, _26875_);
  nor (_26885_, _26884_, _03744_);
  nor (_26886_, _12381_, _10618_);
  nor (_26887_, _26886_, _03745_);
  and (_26888_, _26887_, _26876_);
  nor (_26889_, _26888_, _26885_);
  nor (_26891_, _26889_, _03611_);
  nor (_26892_, _12374_, _10618_);
  nor (_26893_, _26892_, _04523_);
  and (_26894_, _26893_, _26876_);
  nor (_26895_, _26894_, _26891_);
  nor (_26896_, _26895_, _03733_);
  nor (_26897_, _26816_, _05674_);
  nor (_26898_, _26897_, _03734_);
  and (_26899_, _26898_, _26822_);
  nor (_26900_, _26899_, _26896_);
  or (_26902_, _26900_, _18526_);
  and (_26903_, _26821_, _05673_);
  nor (_26904_, _26903_, _06458_);
  and (_26905_, _26904_, _26876_);
  nor (_26906_, _26905_, _03767_);
  and (_26907_, _26880_, _05673_);
  or (_26908_, _26820_, _06453_);
  or (_26909_, _26908_, _26907_);
  and (_26910_, _26909_, _26906_);
  and (_26911_, _26910_, _26902_);
  nor (_26913_, _26829_, _03948_);
  or (_26914_, _26913_, _03445_);
  nor (_26915_, _26914_, _26911_);
  nor (_26916_, _26850_, _03446_);
  or (_26917_, _26916_, _03473_);
  nor (_26918_, _26917_, _26915_);
  nor (_26919_, _26828_, _26816_);
  and (_26920_, _26919_, _03473_);
  nor (_26921_, _26920_, _26918_);
  or (_26922_, _26921_, _43193_);
  or (_26924_, _43189_, \oc8051_golden_model_1.SCON [1]);
  and (_26925_, _26924_, _42003_);
  and (_43849_, _26925_, _26922_);
  not (_26926_, \oc8051_golden_model_1.SCON [2]);
  nor (_26927_, _05333_, _26926_);
  and (_26928_, _05333_, _06399_);
  nor (_26929_, _26928_, _26927_);
  and (_26930_, _26929_, _03624_);
  nor (_26931_, _10618_, _05073_);
  nor (_26932_, _26931_, _26927_);
  and (_26933_, _26932_, _07454_);
  and (_26934_, _05333_, \oc8051_golden_model_1.ACC [2]);
  nor (_26935_, _26934_, _26927_);
  nor (_26936_, _26935_, _04437_);
  nor (_26937_, _04436_, _26926_);
  or (_26938_, _26937_, _26936_);
  and (_26939_, _26938_, _04432_);
  nor (_26940_, _12467_, _10618_);
  nor (_26941_, _26940_, _26927_);
  nor (_26942_, _26941_, _04432_);
  or (_26945_, _26942_, _26939_);
  and (_26946_, _26945_, _03470_);
  nor (_26947_, _05942_, _26926_);
  and (_26948_, _12462_, _05942_);
  nor (_26949_, _26948_, _26947_);
  nor (_26950_, _26949_, _03470_);
  or (_26951_, _26950_, _26946_);
  and (_26952_, _26951_, _04457_);
  nor (_26953_, _26932_, _04457_);
  or (_26954_, _26953_, _26952_);
  and (_26956_, _26954_, _03531_);
  nor (_26957_, _26935_, _03531_);
  or (_26958_, _26957_, _26956_);
  and (_26959_, _26958_, _03466_);
  and (_26960_, _12460_, _05942_);
  nor (_26961_, _26960_, _26947_);
  nor (_26962_, _26961_, _03466_);
  or (_26963_, _26962_, _26959_);
  and (_26964_, _26963_, _03459_);
  and (_26965_, _26948_, _12491_);
  or (_26967_, _26965_, _26947_);
  and (_26968_, _26967_, _03458_);
  or (_26969_, _26968_, _26964_);
  and (_26970_, _26969_, _03453_);
  nor (_26971_, _12509_, _10655_);
  nor (_26972_, _26971_, _26947_);
  nor (_26973_, _26972_, _03453_);
  nor (_26974_, _26973_, _07454_);
  not (_26975_, _26974_);
  nor (_26976_, _26975_, _26970_);
  nor (_26978_, _26976_, _26933_);
  nor (_26979_, _26978_, _04082_);
  and (_26980_, _06710_, _05333_);
  nor (_26981_, _26927_, _04500_);
  not (_26982_, _26981_);
  nor (_26983_, _26982_, _26980_);
  or (_26984_, _26983_, _03224_);
  nor (_26985_, _26984_, _26979_);
  nor (_26986_, _12568_, _10618_);
  nor (_26987_, _26927_, _26986_);
  nor (_26989_, _26987_, _03521_);
  or (_26990_, _26989_, _03624_);
  nor (_26991_, _26990_, _26985_);
  nor (_26992_, _26991_, _26930_);
  or (_26993_, _26992_, _03623_);
  and (_26994_, _12582_, _05333_);
  or (_26995_, _26994_, _26927_);
  or (_26996_, _26995_, _04527_);
  and (_26997_, _26996_, _03745_);
  and (_26998_, _26997_, _26993_);
  and (_27000_, _12588_, _05333_);
  nor (_27001_, _27000_, _26927_);
  nor (_27002_, _27001_, _03745_);
  nor (_27003_, _27002_, _26998_);
  nor (_27004_, _27003_, _03611_);
  nor (_27005_, _26927_, _05772_);
  not (_27006_, _27005_);
  nor (_27007_, _26929_, _04523_);
  and (_27008_, _27007_, _27006_);
  nor (_27009_, _27008_, _27004_);
  nor (_27011_, _27009_, _03733_);
  nor (_27012_, _26935_, _03734_);
  and (_27013_, _27012_, _27006_);
  or (_27014_, _27013_, _27011_);
  and (_27015_, _27014_, _06453_);
  nor (_27016_, _12581_, _10618_);
  nor (_27017_, _27016_, _26927_);
  nor (_27018_, _27017_, _06453_);
  or (_27019_, _27018_, _27015_);
  and (_27020_, _27019_, _06458_);
  nor (_27022_, _12587_, _10618_);
  nor (_27023_, _27022_, _26927_);
  nor (_27024_, _27023_, _06458_);
  or (_27025_, _27024_, _27020_);
  and (_27026_, _27025_, _03948_);
  nor (_27027_, _26941_, _03948_);
  or (_27028_, _27027_, _27026_);
  and (_27029_, _27028_, _03446_);
  nor (_27030_, _26961_, _03446_);
  or (_27031_, _27030_, _27029_);
  and (_27033_, _27031_, _03474_);
  and (_27034_, _12638_, _05333_);
  nor (_27035_, _27034_, _26927_);
  nor (_27036_, _27035_, _03474_);
  or (_27037_, _27036_, _27033_);
  or (_27038_, _27037_, _43193_);
  or (_27039_, _43189_, \oc8051_golden_model_1.SCON [2]);
  and (_27040_, _27039_, _42003_);
  and (_43850_, _27040_, _27038_);
  not (_27041_, \oc8051_golden_model_1.SCON [3]);
  nor (_27042_, _05333_, _27041_);
  and (_27043_, _05333_, _06356_);
  nor (_27044_, _27043_, _27042_);
  and (_27045_, _27044_, _03624_);
  nor (_27046_, _10618_, _04885_);
  nor (_27047_, _27046_, _27042_);
  and (_27048_, _27047_, _07454_);
  and (_27049_, _05333_, \oc8051_golden_model_1.ACC [3]);
  nor (_27050_, _27049_, _27042_);
  nor (_27051_, _27050_, _04437_);
  nor (_27054_, _04436_, _27041_);
  or (_27055_, _27054_, _27051_);
  and (_27056_, _27055_, _04432_);
  nor (_27057_, _12652_, _10618_);
  nor (_27058_, _27057_, _27042_);
  nor (_27059_, _27058_, _04432_);
  or (_27060_, _27059_, _27056_);
  and (_27061_, _27060_, _03470_);
  nor (_27062_, _05942_, _27041_);
  and (_27063_, _12664_, _05942_);
  nor (_27065_, _27063_, _27062_);
  nor (_27066_, _27065_, _03470_);
  or (_27067_, _27066_, _03527_);
  or (_27068_, _27067_, _27061_);
  nand (_27069_, _27047_, _03527_);
  and (_27070_, _27069_, _27068_);
  and (_27071_, _27070_, _03531_);
  nor (_27072_, _27050_, _03531_);
  or (_27073_, _27072_, _27071_);
  and (_27074_, _27073_, _03466_);
  and (_27076_, _12662_, _05942_);
  nor (_27077_, _27076_, _27062_);
  nor (_27078_, _27077_, _03466_);
  or (_27079_, _27078_, _03458_);
  or (_27080_, _27079_, _27074_);
  nor (_27081_, _27062_, _12691_);
  nor (_27082_, _27081_, _27065_);
  or (_27083_, _27082_, _03459_);
  and (_27084_, _27083_, _03453_);
  and (_27085_, _27084_, _27080_);
  nor (_27087_, _12709_, _10655_);
  nor (_27088_, _27087_, _27062_);
  nor (_27089_, _27088_, _03453_);
  nor (_27090_, _27089_, _07454_);
  not (_27091_, _27090_);
  nor (_27092_, _27091_, _27085_);
  nor (_27093_, _27092_, _27048_);
  nor (_27094_, _27093_, _04082_);
  and (_27095_, _06664_, _05333_);
  nor (_27096_, _27042_, _04500_);
  not (_27098_, _27096_);
  nor (_27099_, _27098_, _27095_);
  or (_27100_, _27099_, _03224_);
  nor (_27101_, _27100_, _27094_);
  nor (_27102_, _12773_, _10618_);
  nor (_27103_, _27042_, _27102_);
  nor (_27104_, _27103_, _03521_);
  or (_27105_, _27104_, _03624_);
  nor (_27106_, _27105_, _27101_);
  nor (_27107_, _27106_, _27045_);
  or (_27109_, _27107_, _03623_);
  and (_27110_, _12787_, _05333_);
  or (_27111_, _27110_, _27042_);
  or (_27112_, _27111_, _04527_);
  and (_27113_, _27112_, _03745_);
  and (_27114_, _27113_, _27109_);
  and (_27115_, _12793_, _05333_);
  nor (_27116_, _27115_, _27042_);
  nor (_27117_, _27116_, _03745_);
  nor (_27118_, _27117_, _27114_);
  nor (_27120_, _27118_, _03611_);
  nor (_27121_, _27042_, _05625_);
  not (_27122_, _27121_);
  nor (_27123_, _27044_, _04523_);
  and (_27124_, _27123_, _27122_);
  nor (_27125_, _27124_, _27120_);
  nor (_27126_, _27125_, _03733_);
  nor (_27127_, _27050_, _03734_);
  and (_27128_, _27127_, _27122_);
  nor (_27129_, _27128_, _03618_);
  not (_27131_, _27129_);
  nor (_27132_, _27131_, _27126_);
  nor (_27133_, _12786_, _10618_);
  or (_27134_, _27042_, _06453_);
  nor (_27135_, _27134_, _27133_);
  or (_27136_, _27135_, _03741_);
  nor (_27137_, _27136_, _27132_);
  nor (_27138_, _12792_, _10618_);
  nor (_27139_, _27138_, _27042_);
  nor (_27140_, _27139_, _06458_);
  or (_27142_, _27140_, _27137_);
  and (_27143_, _27142_, _03948_);
  nor (_27144_, _27058_, _03948_);
  or (_27145_, _27144_, _27143_);
  and (_27146_, _27145_, _03446_);
  nor (_27147_, _27077_, _03446_);
  or (_27148_, _27147_, _27146_);
  and (_27149_, _27148_, _03474_);
  and (_27150_, _12843_, _05333_);
  nor (_27151_, _27150_, _27042_);
  nor (_27153_, _27151_, _03474_);
  or (_27154_, _27153_, _27149_);
  or (_27155_, _27154_, _43193_);
  or (_27156_, _43189_, \oc8051_golden_model_1.SCON [3]);
  and (_27157_, _27156_, _42003_);
  and (_43851_, _27157_, _27155_);
  not (_27158_, \oc8051_golden_model_1.SCON [4]);
  nor (_27159_, _05333_, _27158_);
  nor (_27160_, _05831_, _10618_);
  nor (_27161_, _27160_, _27159_);
  and (_27163_, _27161_, _07454_);
  nor (_27164_, _05942_, _27158_);
  and (_27165_, _12864_, _05942_);
  nor (_27166_, _27165_, _27164_);
  nor (_27167_, _27166_, _03466_);
  and (_27168_, _05333_, \oc8051_golden_model_1.ACC [4]);
  nor (_27169_, _27168_, _27159_);
  nor (_27170_, _27169_, _04437_);
  nor (_27171_, _04436_, _27158_);
  or (_27172_, _27171_, _27170_);
  and (_27174_, _27172_, _04432_);
  nor (_27175_, _12856_, _10618_);
  nor (_27176_, _27175_, _27159_);
  nor (_27177_, _27176_, _04432_);
  or (_27178_, _27177_, _27174_);
  and (_27179_, _27178_, _03470_);
  and (_27180_, _12866_, _05942_);
  nor (_27181_, _27180_, _27164_);
  nor (_27182_, _27181_, _03470_);
  or (_27183_, _27182_, _03527_);
  or (_27185_, _27183_, _27179_);
  nand (_27186_, _27161_, _03527_);
  and (_27187_, _27186_, _27185_);
  and (_27188_, _27187_, _03531_);
  nor (_27189_, _27169_, _03531_);
  or (_27190_, _27189_, _27188_);
  and (_27191_, _27190_, _03466_);
  nor (_27192_, _27191_, _27167_);
  nor (_27193_, _27192_, _03458_);
  nor (_27194_, _27164_, _12894_);
  or (_27196_, _27181_, _03459_);
  nor (_27197_, _27196_, _27194_);
  nor (_27198_, _27197_, _27193_);
  nor (_27199_, _27198_, _03452_);
  nor (_27200_, _12912_, _10655_);
  nor (_27201_, _27200_, _27164_);
  nor (_27202_, _27201_, _03453_);
  nor (_27203_, _27202_, _07454_);
  not (_27204_, _27203_);
  nor (_27205_, _27204_, _27199_);
  nor (_27207_, _27205_, _27163_);
  nor (_27208_, _27207_, _04082_);
  and (_27209_, _06802_, _05333_);
  nor (_27210_, _27159_, _04500_);
  not (_27211_, _27210_);
  nor (_27212_, _27211_, _27209_);
  nor (_27213_, _27212_, _03224_);
  not (_27214_, _27213_);
  nor (_27215_, _27214_, _27208_);
  nor (_27216_, _12972_, _10618_);
  nor (_27218_, _27216_, _27159_);
  nor (_27219_, _27218_, _03521_);
  or (_27220_, _27219_, _08905_);
  or (_27221_, _27220_, _27215_);
  and (_27222_, _12986_, _05333_);
  or (_27223_, _27159_, _04527_);
  or (_27224_, _27223_, _27222_);
  and (_27225_, _06337_, _05333_);
  nor (_27226_, _27225_, _27159_);
  and (_27227_, _27226_, _03624_);
  nor (_27229_, _27227_, _03744_);
  and (_27230_, _27229_, _27224_);
  and (_27231_, _27230_, _27221_);
  and (_27232_, _12992_, _05333_);
  nor (_27233_, _27232_, _27159_);
  nor (_27234_, _27233_, _03745_);
  nor (_27235_, _27234_, _27231_);
  nor (_27236_, _27235_, _03611_);
  nor (_27237_, _27159_, _05880_);
  not (_27238_, _27237_);
  nor (_27240_, _27226_, _04523_);
  and (_27241_, _27240_, _27238_);
  nor (_27242_, _27241_, _27236_);
  nor (_27243_, _27242_, _03733_);
  nor (_27244_, _27169_, _03734_);
  and (_27245_, _27244_, _27238_);
  nor (_27246_, _27245_, _03618_);
  not (_27247_, _27246_);
  nor (_27248_, _27247_, _27243_);
  nor (_27249_, _12985_, _10618_);
  or (_27251_, _27159_, _06453_);
  nor (_27252_, _27251_, _27249_);
  or (_27253_, _27252_, _03741_);
  nor (_27254_, _27253_, _27248_);
  nor (_27255_, _12991_, _10618_);
  nor (_27256_, _27255_, _27159_);
  nor (_27257_, _27256_, _06458_);
  or (_27258_, _27257_, _27254_);
  and (_27259_, _27258_, _03948_);
  nor (_27260_, _27176_, _03948_);
  or (_27261_, _27260_, _27259_);
  and (_27262_, _27261_, _03446_);
  nor (_27263_, _27166_, _03446_);
  or (_27264_, _27263_, _27262_);
  and (_27265_, _27264_, _03474_);
  and (_27266_, _13051_, _05333_);
  nor (_27267_, _27266_, _27159_);
  nor (_27268_, _27267_, _03474_);
  or (_27269_, _27268_, _27265_);
  or (_27270_, _27269_, _43193_);
  or (_27273_, _43189_, \oc8051_golden_model_1.SCON [4]);
  and (_27274_, _27273_, _42003_);
  and (_43852_, _27274_, _27270_);
  not (_27275_, \oc8051_golden_model_1.SCON [5]);
  nor (_27276_, _05333_, _27275_);
  and (_27277_, _06757_, _05333_);
  or (_27278_, _27277_, _27276_);
  and (_27279_, _27278_, _04082_);
  and (_27280_, _05333_, \oc8051_golden_model_1.ACC [5]);
  nor (_27281_, _27280_, _27276_);
  nor (_27283_, _27281_, _04437_);
  nor (_27284_, _04436_, _27275_);
  or (_27285_, _27284_, _27283_);
  and (_27286_, _27285_, _04432_);
  nor (_27287_, _13070_, _10618_);
  nor (_27288_, _27287_, _27276_);
  nor (_27289_, _27288_, _04432_);
  or (_27290_, _27289_, _27286_);
  and (_27291_, _27290_, _03470_);
  nor (_27292_, _05942_, _27275_);
  and (_27294_, _13095_, _05942_);
  nor (_27295_, _27294_, _27292_);
  nor (_27296_, _27295_, _03470_);
  or (_27297_, _27296_, _03527_);
  or (_27298_, _27297_, _27291_);
  nor (_27299_, _05526_, _10618_);
  nor (_27300_, _27299_, _27276_);
  nand (_27301_, _27300_, _03527_);
  and (_27302_, _27301_, _27298_);
  and (_27303_, _27302_, _03531_);
  nor (_27305_, _27281_, _03531_);
  or (_27306_, _27305_, _27303_);
  and (_27307_, _27306_, _03466_);
  and (_27308_, _13078_, _05942_);
  nor (_27309_, _27308_, _27292_);
  nor (_27310_, _27309_, _03466_);
  or (_27311_, _27310_, _27307_);
  and (_27312_, _27311_, _03459_);
  nor (_27313_, _27292_, _13110_);
  nor (_27314_, _27313_, _27295_);
  and (_27316_, _27314_, _03458_);
  or (_27317_, _27316_, _27312_);
  and (_27318_, _27317_, _03453_);
  nor (_27319_, _13076_, _10655_);
  nor (_27320_, _27319_, _27292_);
  nor (_27321_, _27320_, _03453_);
  nor (_27322_, _27321_, _07454_);
  not (_27323_, _27322_);
  nor (_27324_, _27323_, _27318_);
  and (_27325_, _27300_, _07454_);
  or (_27327_, _27325_, _04082_);
  nor (_27328_, _27327_, _27324_);
  or (_27329_, _27328_, _27279_);
  and (_27330_, _27329_, _03521_);
  nor (_27331_, _13184_, _10618_);
  nor (_27332_, _27331_, _27276_);
  nor (_27333_, _27332_, _03521_);
  or (_27334_, _27333_, _08905_);
  or (_27335_, _27334_, _27330_);
  and (_27336_, _13198_, _05333_);
  or (_27338_, _27276_, _04527_);
  or (_27339_, _27338_, _27336_);
  and (_27340_, _06295_, _05333_);
  nor (_27341_, _27340_, _27276_);
  and (_27342_, _27341_, _03624_);
  nor (_27343_, _27342_, _03744_);
  and (_27344_, _27343_, _27339_);
  and (_27345_, _27344_, _27335_);
  and (_27346_, _13204_, _05333_);
  nor (_27347_, _27346_, _27276_);
  nor (_27349_, _27347_, _03745_);
  nor (_27350_, _27349_, _27345_);
  nor (_27351_, _27350_, _03611_);
  nor (_27352_, _27276_, _05576_);
  not (_27353_, _27352_);
  nor (_27354_, _27341_, _04523_);
  and (_27355_, _27354_, _27353_);
  nor (_27356_, _27355_, _27351_);
  nor (_27357_, _27356_, _03733_);
  nor (_27358_, _27281_, _03734_);
  and (_27360_, _27358_, _27353_);
  nor (_27361_, _27360_, _03618_);
  not (_27362_, _27361_);
  nor (_27363_, _27362_, _27357_);
  nor (_27364_, _13197_, _10618_);
  or (_27365_, _27276_, _06453_);
  nor (_27366_, _27365_, _27364_);
  or (_27367_, _27366_, _03741_);
  nor (_27368_, _27367_, _27363_);
  nor (_27369_, _13203_, _10618_);
  nor (_27371_, _27369_, _27276_);
  nor (_27372_, _27371_, _06458_);
  or (_27373_, _27372_, _27368_);
  and (_27374_, _27373_, _03948_);
  nor (_27375_, _27288_, _03948_);
  or (_27376_, _27375_, _27374_);
  and (_27377_, _27376_, _03446_);
  nor (_27378_, _27309_, _03446_);
  or (_27379_, _27378_, _27377_);
  and (_27380_, _27379_, _03474_);
  and (_27382_, _13253_, _05333_);
  nor (_27383_, _27382_, _27276_);
  nor (_27384_, _27383_, _03474_);
  or (_27385_, _27384_, _27380_);
  or (_27386_, _27385_, _43193_);
  or (_27387_, _43189_, \oc8051_golden_model_1.SCON [5]);
  and (_27388_, _27387_, _42003_);
  and (_43853_, _27388_, _27386_);
  not (_27389_, \oc8051_golden_model_1.SCON [6]);
  nor (_27390_, _05333_, _27389_);
  and (_27392_, _06526_, _05333_);
  or (_27393_, _27392_, _27390_);
  and (_27394_, _27393_, _04082_);
  and (_27395_, _05333_, \oc8051_golden_model_1.ACC [6]);
  nor (_27396_, _27395_, _27390_);
  nor (_27397_, _27396_, _04437_);
  nor (_27398_, _04436_, _27389_);
  or (_27399_, _27398_, _27397_);
  and (_27400_, _27399_, _04432_);
  nor (_27401_, _13293_, _10618_);
  nor (_27403_, _27401_, _27390_);
  nor (_27404_, _27403_, _04432_);
  or (_27405_, _27404_, _27400_);
  and (_27406_, _27405_, _03470_);
  nor (_27407_, _05942_, _27389_);
  and (_27408_, _13280_, _05942_);
  nor (_27409_, _27408_, _27407_);
  nor (_27410_, _27409_, _03470_);
  or (_27411_, _27410_, _03527_);
  or (_27412_, _27411_, _27406_);
  nor (_27414_, _05417_, _10618_);
  nor (_27415_, _27414_, _27390_);
  nand (_27416_, _27415_, _03527_);
  and (_27417_, _27416_, _27412_);
  and (_27418_, _27417_, _03531_);
  nor (_27419_, _27396_, _03531_);
  or (_27420_, _27419_, _27418_);
  and (_27421_, _27420_, _03466_);
  and (_27422_, _13304_, _05942_);
  nor (_27423_, _27422_, _27407_);
  nor (_27425_, _27423_, _03466_);
  or (_27426_, _27425_, _03458_);
  or (_27427_, _27426_, _27421_);
  nor (_27428_, _27407_, _13311_);
  nor (_27429_, _27428_, _27409_);
  or (_27430_, _27429_, _03459_);
  and (_27431_, _27430_, _03453_);
  and (_27432_, _27431_, _27427_);
  nor (_27433_, _13329_, _10655_);
  nor (_27434_, _27433_, _27407_);
  nor (_27436_, _27434_, _03453_);
  nor (_27437_, _27436_, _07454_);
  not (_27438_, _27437_);
  nor (_27439_, _27438_, _27432_);
  and (_27440_, _27415_, _07454_);
  or (_27441_, _27440_, _04082_);
  nor (_27442_, _27441_, _27439_);
  or (_27443_, _27442_, _27394_);
  and (_27444_, _27443_, _03521_);
  nor (_27445_, _13387_, _10618_);
  nor (_27447_, _27445_, _27390_);
  nor (_27448_, _27447_, _03521_);
  or (_27449_, _27448_, _08905_);
  or (_27450_, _27449_, _27444_);
  and (_27451_, _13402_, _05333_);
  or (_27452_, _27390_, _04527_);
  or (_27453_, _27452_, _27451_);
  and (_27454_, _14949_, _05333_);
  nor (_27455_, _27454_, _27390_);
  and (_27456_, _27455_, _03624_);
  nor (_27458_, _27456_, _03744_);
  and (_27459_, _27458_, _27453_);
  and (_27460_, _27459_, _27450_);
  and (_27461_, _13407_, _05333_);
  nor (_27462_, _27461_, _27390_);
  nor (_27463_, _27462_, _03745_);
  nor (_27464_, _27463_, _27460_);
  nor (_27465_, _27464_, _03611_);
  nor (_27466_, _27390_, _05469_);
  not (_27467_, _27466_);
  nor (_27469_, _27455_, _04523_);
  and (_27470_, _27469_, _27467_);
  nor (_27471_, _27470_, _27465_);
  nor (_27472_, _27471_, _03733_);
  nor (_27473_, _27396_, _03734_);
  and (_27474_, _27473_, _27467_);
  nor (_27475_, _27474_, _03618_);
  not (_27476_, _27475_);
  nor (_27477_, _27476_, _27472_);
  nor (_27478_, _13400_, _10618_);
  or (_27480_, _27390_, _06453_);
  nor (_27481_, _27480_, _27478_);
  or (_27482_, _27481_, _03741_);
  nor (_27483_, _27482_, _27477_);
  nor (_27484_, _13406_, _10618_);
  nor (_27485_, _27484_, _27390_);
  nor (_27486_, _27485_, _06458_);
  or (_27487_, _27486_, _27483_);
  and (_27488_, _27487_, _03948_);
  nor (_27489_, _27403_, _03948_);
  or (_27491_, _27489_, _27488_);
  and (_27492_, _27491_, _03446_);
  nor (_27493_, _27423_, _03446_);
  or (_27494_, _27493_, _27492_);
  and (_27495_, _27494_, _03474_);
  and (_27496_, _13456_, _05333_);
  nor (_27497_, _27496_, _27390_);
  nor (_27498_, _27497_, _03474_);
  or (_27499_, _27498_, _27495_);
  or (_27500_, _27499_, _43193_);
  or (_27502_, _43189_, \oc8051_golden_model_1.SCON [6]);
  and (_27503_, _27502_, _42003_);
  and (_43854_, _27503_, _27500_);
  nor (_27504_, _05323_, _03455_);
  nor (_27505_, _05722_, _10741_);
  nor (_27506_, _27505_, _27504_);
  and (_27507_, _27506_, _17198_);
  and (_27508_, _05323_, \oc8051_golden_model_1.ACC [0]);
  nor (_27509_, _27508_, _27504_);
  nor (_27510_, _27509_, _04437_);
  nor (_27512_, _04436_, _03455_);
  or (_27513_, _27512_, _27510_);
  and (_27514_, _27513_, _04432_);
  nor (_27515_, _27506_, _04432_);
  or (_27516_, _27515_, _27514_);
  and (_27517_, _27516_, _04457_);
  or (_27518_, _27517_, _04027_);
  and (_27519_, _27518_, _03531_);
  nor (_27520_, _27509_, _03531_);
  or (_27521_, _27520_, _27519_);
  and (_27522_, _27521_, _04577_);
  nor (_27523_, _07454_, _04473_);
  not (_27524_, _27523_);
  nor (_27525_, _27524_, _27522_);
  not (_27526_, _27504_);
  and (_27527_, _05323_, _04429_);
  nor (_27528_, _27527_, _06903_);
  and (_27529_, _27528_, _27526_);
  nor (_27530_, _27529_, _27525_);
  nor (_27531_, _27530_, _04082_);
  and (_27534_, _06617_, _05323_);
  nor (_27535_, _27504_, _04500_);
  not (_27536_, _27535_);
  nor (_27537_, _27536_, _27534_);
  nor (_27538_, _27537_, _27531_);
  nor (_27539_, _27538_, _03224_);
  nor (_27540_, _12164_, _10741_);
  or (_27541_, _27504_, _03521_);
  nor (_27542_, _27541_, _27540_);
  or (_27543_, _27542_, _03624_);
  nor (_27545_, _27543_, _27539_);
  and (_27546_, _05323_, _06350_);
  nor (_27547_, _27546_, _27504_);
  nand (_27548_, _27547_, _04527_);
  and (_27549_, _27548_, _08905_);
  nor (_27550_, _27549_, _27545_);
  and (_27551_, _12177_, _05323_);
  nor (_27552_, _27551_, _27504_);
  and (_27553_, _27552_, _03623_);
  nor (_27554_, _27553_, _27550_);
  nor (_27556_, _27554_, _03744_);
  and (_27557_, _12183_, _05323_);
  or (_27558_, _27504_, _03745_);
  nor (_27559_, _27558_, _27557_);
  or (_27560_, _27559_, _03611_);
  nor (_27561_, _27560_, _27556_);
  or (_27562_, _27547_, _04523_);
  nor (_27563_, _27562_, _27505_);
  nor (_27564_, _27563_, _27561_);
  nor (_27565_, _27564_, _03733_);
  and (_27567_, _12182_, _05323_);
  or (_27568_, _27567_, _27504_);
  and (_27569_, _27568_, _03733_);
  or (_27570_, _27569_, _27565_);
  and (_27571_, _27570_, _06453_);
  nor (_27572_, _12057_, _10741_);
  nor (_27573_, _27572_, _27504_);
  nor (_27574_, _27573_, _06453_);
  or (_27575_, _27574_, _27571_);
  and (_27576_, _27575_, _06458_);
  nor (_27578_, _12181_, _10741_);
  nor (_27579_, _27578_, _27504_);
  nor (_27580_, _27579_, _06458_);
  nor (_27581_, _27580_, _17198_);
  not (_27582_, _27581_);
  nor (_27583_, _27582_, _27576_);
  nor (_27584_, _27583_, _27507_);
  and (_27585_, _27584_, _43189_);
  nor (_27586_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27587_, _27586_, _00001_);
  or (_43857_, _27587_, _27585_);
  nor (_27589_, _05323_, _04342_);
  and (_27590_, _12265_, _05323_);
  nor (_27591_, _27590_, _27589_);
  nor (_27592_, _27591_, _03474_);
  nor (_27593_, _10848_, _04342_);
  and (_27594_, _03168_, _04342_);
  not (_27595_, _03168_);
  nor (_27596_, _05323_, \oc8051_golden_model_1.SP [1]);
  and (_27597_, _05323_, _03269_);
  nor (_27599_, _27597_, _27596_);
  nor (_27600_, _27599_, _04437_);
  nor (_27601_, _10754_, \oc8051_golden_model_1.SP [1]);
  and (_27602_, _03204_, \oc8051_golden_model_1.SP [1]);
  nor (_27603_, _27602_, _27601_);
  nor (_27604_, _27603_, _27600_);
  and (_27605_, _27604_, _04432_);
  nor (_27606_, _27596_, _27590_);
  and (_27607_, _27606_, _03534_);
  or (_27608_, _27607_, _27605_);
  and (_27610_, _27608_, _03202_);
  nor (_27611_, _03202_, \oc8051_golden_model_1.SP [1]);
  or (_27612_, _27611_, _03527_);
  or (_27613_, _27612_, _27610_);
  nand (_27614_, _04572_, _03527_);
  and (_27615_, _27614_, _27613_);
  and (_27616_, _27615_, _03531_);
  and (_27617_, _27599_, _03530_);
  or (_27618_, _27617_, _27616_);
  and (_27619_, _27618_, _04577_);
  or (_27621_, _27619_, _04756_);
  nor (_27622_, _27621_, _04576_);
  and (_27623_, _04756_, \oc8051_golden_model_1.SP [1]);
  or (_27624_, _27623_, _07454_);
  nor (_27625_, _27624_, _27622_);
  nand (_27626_, _05323_, _04635_);
  nor (_27627_, _27596_, _06903_);
  and (_27628_, _27627_, _27626_);
  nor (_27629_, _27628_, _04082_);
  not (_27630_, _27629_);
  nor (_27632_, _27630_, _27625_);
  and (_27633_, _06572_, _05323_);
  nor (_27634_, _27589_, _04500_);
  not (_27635_, _27634_);
  nor (_27636_, _27635_, _27633_);
  nor (_27637_, _27636_, _03224_);
  not (_27638_, _27637_);
  nor (_27639_, _27638_, _27632_);
  nor (_27640_, _12360_, _10741_);
  or (_27641_, _27640_, _27589_);
  and (_27643_, _27641_, _03224_);
  nor (_27644_, _27643_, _27639_);
  nor (_27645_, _27644_, _03624_);
  and (_27646_, _05323_, _06354_);
  or (_27647_, _27646_, _27589_);
  and (_27648_, _27647_, _03624_);
  or (_27649_, _27648_, _27645_);
  and (_27650_, _27649_, _27595_);
  or (_27651_, _27650_, _27594_);
  and (_27652_, _27651_, _04527_);
  nor (_27654_, _12375_, _10741_);
  or (_27655_, _27654_, _04527_);
  nor (_27656_, _27655_, _27596_);
  nor (_27657_, _27656_, _27652_);
  nor (_27658_, _27657_, _03744_);
  nor (_27659_, _12381_, _10741_);
  or (_27660_, _27659_, _03745_);
  nor (_27661_, _27660_, _27596_);
  nor (_27662_, _27661_, _27658_);
  nor (_27663_, _27662_, _03611_);
  nor (_27665_, _12374_, _10741_);
  or (_27666_, _27665_, _04523_);
  nor (_27667_, _27666_, _27596_);
  nor (_27668_, _27667_, _27663_);
  nor (_27669_, _27668_, _10829_);
  and (_27670_, _03182_, _04342_);
  nor (_27671_, _27589_, _05674_);
  nor (_27672_, _27671_, _03734_);
  and (_27673_, _27672_, _27599_);
  nor (_27674_, _27673_, _27670_);
  not (_27676_, _27674_);
  nor (_27677_, _27676_, _27669_);
  or (_27678_, _27677_, _18526_);
  nor (_27679_, _12380_, _10741_);
  or (_27680_, _27679_, _27589_);
  and (_27681_, _27680_, _03741_);
  not (_27682_, _10848_);
  nor (_27683_, _12373_, _10741_);
  or (_27684_, _27683_, _27589_);
  and (_27685_, _27684_, _03618_);
  or (_27687_, _27685_, _27682_);
  nor (_27688_, _27687_, _27681_);
  and (_27689_, _27688_, _27678_);
  nor (_27690_, _27689_, _27593_);
  and (_27691_, _27690_, _03476_);
  and (_27692_, _03475_, _04342_);
  or (_27693_, _27692_, _27691_);
  and (_27694_, _27693_, _03948_);
  and (_27695_, _27606_, _03767_);
  nor (_27696_, _27695_, _04986_);
  not (_27698_, _27696_);
  nor (_27699_, _27698_, _27694_);
  nor (_27700_, _04553_, _04342_);
  nor (_27701_, _27700_, _03473_);
  not (_27702_, _27701_);
  nor (_27703_, _27702_, _27699_);
  nor (_27704_, _27703_, _27592_);
  nor (_27705_, _27704_, _43193_);
  nor (_27706_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27707_, _27706_, _00001_);
  or (_43858_, _27707_, _27705_);
  and (_27709_, _05169_, _03191_);
  nor (_27710_, _05323_, _03857_);
  and (_27711_, _12588_, _05323_);
  nor (_27712_, _27711_, _27710_);
  nor (_27713_, _27712_, _03745_);
  and (_27714_, _13839_, _03168_);
  not (_27715_, _27710_);
  nor (_27716_, _10741_, _05073_);
  nor (_27717_, _27716_, _06903_);
  and (_27719_, _27717_, _27715_);
  nor (_27720_, _12467_, _10741_);
  nor (_27721_, _27720_, _27710_);
  and (_27722_, _27721_, _03534_);
  and (_27723_, _05323_, \oc8051_golden_model_1.ACC [2]);
  nor (_27724_, _27723_, _27710_);
  or (_27725_, _27724_, _04437_);
  nand (_27726_, _10754_, \oc8051_golden_model_1.SP [2]);
  nor (_27727_, _13839_, _03204_);
  nor (_27728_, _27727_, _03534_);
  and (_27730_, _27728_, _27726_);
  and (_27731_, _27730_, _27725_);
  nor (_27732_, _27731_, _05977_);
  not (_27733_, _27732_);
  nor (_27734_, _27733_, _27722_);
  nor (_27735_, _13839_, _03202_);
  or (_27736_, _27735_, _03527_);
  nor (_27737_, _27736_, _27734_);
  and (_27738_, _06035_, _03527_);
  nor (_27739_, _27738_, _27737_);
  and (_27741_, _27739_, _03531_);
  nor (_27742_, _27724_, _03531_);
  or (_27743_, _27742_, _27741_);
  and (_27744_, _27743_, _04577_);
  nor (_27745_, _27744_, _05014_);
  nor (_27746_, _27745_, _04756_);
  and (_27747_, _05169_, _04756_);
  nor (_27748_, _27747_, _07454_);
  not (_27749_, _27748_);
  nor (_27750_, _27749_, _27746_);
  nor (_27752_, _27750_, _27719_);
  nor (_27753_, _27752_, _04082_);
  and (_27754_, _06710_, _05323_);
  nor (_27755_, _27710_, _04500_);
  not (_27756_, _27755_);
  nor (_27757_, _27756_, _27754_);
  or (_27758_, _27757_, _03224_);
  nor (_27759_, _27758_, _27753_);
  nor (_27760_, _12568_, _10741_);
  nor (_27761_, _27760_, _27710_);
  nor (_27763_, _27761_, _03521_);
  or (_27764_, _27763_, _03624_);
  or (_27765_, _27764_, _27759_);
  and (_27766_, _05323_, _06399_);
  nor (_27767_, _27766_, _27710_);
  nand (_27768_, _27767_, _03624_);
  and (_27769_, _27768_, _27765_);
  nor (_27770_, _27769_, _03168_);
  nor (_27771_, _27770_, _27714_);
  nor (_27772_, _27771_, _03623_);
  and (_27774_, _12582_, _05323_);
  or (_27775_, _27710_, _04527_);
  nor (_27776_, _27775_, _27774_);
  or (_27777_, _27776_, _03744_);
  nor (_27778_, _27777_, _27772_);
  nor (_27779_, _27778_, _27713_);
  nor (_27780_, _27779_, _03611_);
  and (_27781_, _27715_, _05771_);
  not (_27782_, _27781_);
  nor (_27783_, _27767_, _04523_);
  and (_27785_, _27783_, _27782_);
  nor (_27786_, _27785_, _27780_);
  nor (_27787_, _27786_, _10829_);
  nor (_27788_, _27724_, _03734_);
  and (_27789_, _27788_, _27782_);
  and (_27790_, _05169_, _03182_);
  nor (_27791_, _27790_, _27789_);
  and (_27792_, _27791_, _06453_);
  not (_27793_, _27792_);
  nor (_27794_, _27793_, _27787_);
  nor (_27796_, _12581_, _10741_);
  nor (_27797_, _27796_, _27710_);
  and (_27798_, _27797_, _03618_);
  nor (_27799_, _27798_, _27794_);
  nor (_27800_, _27799_, _03741_);
  nor (_27801_, _12587_, _10741_);
  or (_27802_, _27710_, _06458_);
  nor (_27803_, _27802_, _27801_);
  or (_27804_, _27803_, _03752_);
  nor (_27805_, _27804_, _27800_);
  and (_27806_, _13839_, _03752_);
  or (_27807_, _27806_, _27805_);
  and (_27808_, _27807_, _04803_);
  or (_27809_, _27808_, _27709_);
  and (_27810_, _27809_, _03476_);
  and (_27811_, _13839_, _03475_);
  or (_27812_, _27811_, _03767_);
  nor (_27813_, _27812_, _27810_);
  and (_27814_, _27721_, _03767_);
  nor (_27815_, _27814_, _04986_);
  not (_27818_, _27815_);
  nor (_27819_, _27818_, _27813_);
  nor (_27820_, _13839_, _04553_);
  nor (_27821_, _27820_, _03473_);
  not (_27822_, _27821_);
  nor (_27823_, _27822_, _27819_);
  and (_27824_, _12638_, _05323_);
  nor (_27825_, _27824_, _27710_);
  and (_27826_, _27825_, _03473_);
  nor (_27827_, _27826_, _27823_);
  and (_27829_, _27827_, _43189_);
  nor (_27830_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27831_, _27830_, _00001_);
  or (_43859_, _27831_, _27829_);
  nor (_27832_, _05172_, _04553_);
  and (_27833_, _05172_, _03191_);
  nor (_27834_, _05323_, _03526_);
  and (_27835_, _12793_, _05323_);
  nor (_27836_, _27835_, _27834_);
  nor (_27837_, _27836_, _03745_);
  and (_27839_, _13636_, _03168_);
  nor (_27840_, _10741_, _04885_);
  nor (_27841_, _27840_, _27834_);
  nor (_27842_, _27841_, _06903_);
  or (_27843_, _27842_, _04082_);
  nor (_27844_, _12652_, _10741_);
  nor (_27845_, _27844_, _27834_);
  and (_27846_, _27845_, _03534_);
  and (_27847_, _05323_, \oc8051_golden_model_1.ACC [3]);
  nor (_27848_, _27847_, _27834_);
  or (_27850_, _27848_, _04437_);
  nand (_27851_, _10754_, \oc8051_golden_model_1.SP [3]);
  nor (_27852_, _13636_, _03204_);
  nor (_27853_, _27852_, _03534_);
  and (_27854_, _27853_, _27851_);
  and (_27855_, _27854_, _27850_);
  nor (_27856_, _27855_, _05977_);
  not (_27857_, _27856_);
  nor (_27858_, _27857_, _27846_);
  nor (_27859_, _13636_, _03202_);
  or (_27861_, _27859_, _03527_);
  nor (_27862_, _27861_, _27858_);
  and (_27863_, _06018_, _03527_);
  nor (_27864_, _27863_, _27862_);
  and (_27865_, _27864_, _03531_);
  nor (_27866_, _27848_, _03531_);
  or (_27867_, _27866_, _27865_);
  and (_27868_, _27867_, _04577_);
  or (_27869_, _27868_, _04756_);
  nor (_27870_, _27869_, _04934_);
  and (_27872_, _13636_, _04756_);
  or (_27873_, _27872_, _07454_);
  nor (_27874_, _27873_, _27870_);
  nor (_27875_, _27874_, _27843_);
  and (_27876_, _06664_, _05323_);
  nor (_27877_, _27834_, _04500_);
  not (_27878_, _27877_);
  nor (_27879_, _27878_, _27876_);
  or (_27880_, _27879_, _03224_);
  nor (_27881_, _27880_, _27875_);
  nor (_27883_, _12773_, _10741_);
  nor (_27884_, _27883_, _27834_);
  nor (_27885_, _27884_, _03521_);
  or (_27886_, _27885_, _03624_);
  or (_27887_, _27886_, _27881_);
  and (_27888_, _05323_, _06356_);
  nor (_27889_, _27888_, _27834_);
  nand (_27890_, _27889_, _03624_);
  and (_27891_, _27890_, _27887_);
  nor (_27892_, _27891_, _03168_);
  nor (_27894_, _27892_, _27839_);
  nor (_27895_, _27894_, _03623_);
  and (_27896_, _12787_, _05323_);
  or (_27897_, _27834_, _04527_);
  nor (_27898_, _27897_, _27896_);
  or (_27899_, _27898_, _03744_);
  nor (_27900_, _27899_, _27895_);
  nor (_27901_, _27900_, _27837_);
  nor (_27902_, _27901_, _03611_);
  nor (_27903_, _27834_, _05625_);
  not (_27905_, _27903_);
  nor (_27906_, _27889_, _04523_);
  and (_27907_, _27906_, _27905_);
  nor (_27908_, _27907_, _27902_);
  nor (_27909_, _27908_, _10829_);
  nor (_27910_, _27848_, _03734_);
  and (_27911_, _27910_, _27905_);
  and (_27912_, _05172_, _03182_);
  nor (_27913_, _27912_, _27911_);
  and (_27914_, _27913_, _06453_);
  not (_27916_, _27914_);
  nor (_27917_, _27916_, _27909_);
  nor (_27918_, _12786_, _10741_);
  nor (_27919_, _27918_, _27834_);
  and (_27920_, _27919_, _03618_);
  nor (_27921_, _27920_, _27917_);
  nor (_27922_, _27921_, _03741_);
  nor (_27923_, _12792_, _10741_);
  or (_27924_, _27834_, _06458_);
  nor (_27925_, _27924_, _27923_);
  or (_27927_, _27925_, _03752_);
  nor (_27928_, _27927_, _27922_);
  nor (_27929_, _06014_, _03526_);
  nor (_27930_, _27929_, _06015_);
  nor (_27931_, _27930_, _10735_);
  or (_27932_, _27931_, _27928_);
  and (_27933_, _27932_, _04803_);
  or (_27934_, _27933_, _27833_);
  and (_27935_, _27934_, _03476_);
  nor (_27936_, _27930_, _03476_);
  or (_27938_, _27936_, _27935_);
  and (_27939_, _27938_, _03948_);
  nor (_27940_, _27845_, _03948_);
  nor (_27941_, _27940_, _04986_);
  not (_27942_, _27941_);
  nor (_27943_, _27942_, _27939_);
  nor (_27944_, _27943_, _27832_);
  and (_27945_, _27944_, _03474_);
  and (_27946_, _12843_, _05323_);
  nor (_27947_, _27946_, _27834_);
  nor (_27949_, _27947_, _03474_);
  or (_27950_, _27949_, _27945_);
  or (_27951_, _27950_, _43193_);
  or (_27952_, _43189_, \oc8051_golden_model_1.SP [3]);
  and (_27953_, _27952_, _42003_);
  and (_43860_, _27953_, _27951_);
  nor (_27954_, _04891_, \oc8051_golden_model_1.SP [4]);
  nor (_27955_, _27954_, _10727_);
  nor (_27956_, _27955_, _04553_);
  nor (_27957_, _05323_, _10770_);
  and (_27959_, _12992_, _05323_);
  nor (_27960_, _27959_, _27957_);
  nor (_27961_, _27960_, _03745_);
  nor (_27962_, _05831_, _10741_);
  nor (_27963_, _27962_, _27957_);
  nor (_27964_, _27963_, _06903_);
  or (_27965_, _27964_, _04082_);
  nor (_27966_, _12856_, _10741_);
  nor (_27967_, _27966_, _27957_);
  and (_27968_, _27967_, _03534_);
  and (_27970_, _05323_, \oc8051_golden_model_1.ACC [4]);
  nor (_27971_, _27970_, _27957_);
  or (_27972_, _27971_, _04437_);
  nand (_27973_, _10754_, \oc8051_golden_model_1.SP [4]);
  not (_27974_, _27955_);
  nor (_27975_, _27974_, _03204_);
  nor (_27976_, _27975_, _03534_);
  and (_27977_, _27976_, _27973_);
  and (_27978_, _27977_, _27972_);
  nor (_27979_, _27978_, _05977_);
  not (_27981_, _27979_);
  nor (_27982_, _27981_, _27968_);
  nor (_27983_, _27974_, _03202_);
  or (_27984_, _27983_, _03527_);
  nor (_27985_, _27984_, _27982_);
  and (_27986_, _10771_, _03455_);
  nor (_27987_, _06017_, _10770_);
  nor (_27988_, _27987_, _27986_);
  and (_27989_, _27988_, _03527_);
  nor (_27990_, _27989_, _27985_);
  and (_27992_, _27990_, _03531_);
  nor (_27993_, _27971_, _03531_);
  or (_27994_, _27993_, _27992_);
  and (_27995_, _27994_, _04577_);
  nor (_27996_, _04892_, _10770_);
  and (_27997_, _04892_, _10770_);
  nor (_27998_, _27997_, _27996_);
  and (_27999_, _27998_, _03464_);
  nor (_28000_, _27999_, _04756_);
  not (_28001_, _28000_);
  nor (_28003_, _28001_, _27995_);
  and (_28004_, _27974_, _04756_);
  or (_28005_, _28004_, _07454_);
  nor (_28006_, _28005_, _28003_);
  nor (_28007_, _28006_, _27965_);
  and (_28008_, _06802_, _05323_);
  nor (_28009_, _27957_, _04500_);
  not (_28010_, _28009_);
  nor (_28011_, _28010_, _28008_);
  or (_28012_, _28011_, _03224_);
  nor (_28014_, _28012_, _28007_);
  nor (_28015_, _12972_, _10741_);
  nor (_28016_, _28015_, _27957_);
  nor (_28017_, _28016_, _03521_);
  or (_28018_, _28017_, _03624_);
  or (_28019_, _28018_, _28014_);
  and (_28020_, _06337_, _05323_);
  nor (_28021_, _28020_, _27957_);
  nand (_28022_, _28021_, _03624_);
  and (_28023_, _28022_, _28019_);
  nor (_28025_, _28023_, _03168_);
  and (_28026_, _27974_, _03168_);
  nor (_28027_, _28026_, _28025_);
  nor (_28028_, _28027_, _03623_);
  and (_28029_, _12986_, _05323_);
  or (_28030_, _27957_, _04527_);
  nor (_28031_, _28030_, _28029_);
  or (_28032_, _28031_, _03744_);
  nor (_28033_, _28032_, _28028_);
  nor (_28034_, _28033_, _27961_);
  nor (_28036_, _28034_, _03611_);
  nor (_28037_, _27957_, _05880_);
  not (_28038_, _28037_);
  nor (_28039_, _28021_, _04523_);
  and (_28040_, _28039_, _28038_);
  nor (_28041_, _28040_, _28036_);
  nor (_28042_, _28041_, _10829_);
  nor (_28043_, _27971_, _03734_);
  and (_28044_, _28043_, _28038_);
  and (_28045_, _27955_, _03182_);
  nor (_28047_, _28045_, _28044_);
  and (_28048_, _28047_, _06453_);
  not (_28049_, _28048_);
  nor (_28050_, _28049_, _28042_);
  nor (_28051_, _12985_, _10741_);
  nor (_28052_, _28051_, _27957_);
  and (_28053_, _28052_, _03618_);
  nor (_28054_, _28053_, _28050_);
  nor (_28055_, _28054_, _03741_);
  nor (_28056_, _12991_, _10741_);
  or (_28058_, _27957_, _06458_);
  nor (_28059_, _28058_, _28056_);
  or (_28060_, _28059_, _03752_);
  nor (_28061_, _28060_, _28055_);
  nor (_28062_, _06015_, _10770_);
  nor (_28063_, _28062_, _10771_);
  nor (_28064_, _28063_, _10735_);
  or (_28065_, _28064_, _28061_);
  and (_28066_, _28065_, _04803_);
  and (_28067_, _27955_, _03191_);
  or (_28069_, _28067_, _28066_);
  and (_28070_, _28069_, _03476_);
  nor (_28071_, _28063_, _03476_);
  or (_28072_, _28071_, _28070_);
  and (_28073_, _28072_, _03948_);
  nor (_28074_, _27967_, _03948_);
  nor (_28075_, _28074_, _04986_);
  not (_28076_, _28075_);
  nor (_28077_, _28076_, _28073_);
  nor (_28078_, _28077_, _27956_);
  and (_28080_, _28078_, _03474_);
  and (_28081_, _13051_, _05323_);
  nor (_28082_, _28081_, _27957_);
  nor (_28083_, _28082_, _03474_);
  or (_28084_, _28083_, _28080_);
  or (_28085_, _28084_, _43193_);
  or (_28086_, _43189_, \oc8051_golden_model_1.SP [4]);
  and (_28087_, _28086_, _42003_);
  and (_43861_, _28087_, _28085_);
  nor (_28088_, _10727_, \oc8051_golden_model_1.SP [5]);
  nor (_28090_, _28088_, _10728_);
  nor (_28091_, _28090_, _04553_);
  nor (_28092_, _05323_, _10769_);
  and (_28093_, _13204_, _05323_);
  nor (_28094_, _28093_, _28092_);
  nor (_28095_, _28094_, _03745_);
  nor (_28096_, _05526_, _10741_);
  nor (_28097_, _28096_, _28092_);
  nor (_28098_, _28097_, _06903_);
  or (_28099_, _28098_, _04082_);
  nor (_28101_, _13070_, _10741_);
  nor (_28102_, _28101_, _28092_);
  and (_28103_, _28102_, _03534_);
  and (_28104_, _05323_, \oc8051_golden_model_1.ACC [5]);
  nor (_28105_, _28104_, _28092_);
  or (_28106_, _28105_, _04437_);
  nand (_28107_, _10754_, \oc8051_golden_model_1.SP [5]);
  not (_28108_, _28090_);
  nor (_28109_, _28108_, _03204_);
  nor (_28110_, _28109_, _03534_);
  and (_28112_, _28110_, _28107_);
  and (_28113_, _28112_, _28106_);
  nor (_28114_, _28113_, _05977_);
  not (_28115_, _28114_);
  nor (_28116_, _28115_, _28103_);
  nor (_28117_, _28108_, _03202_);
  or (_28118_, _28117_, _03527_);
  nor (_28119_, _28118_, _28116_);
  and (_28120_, _10772_, _03455_);
  nor (_28121_, _27986_, _10769_);
  nor (_28123_, _28121_, _28120_);
  and (_28124_, _28123_, _03527_);
  nor (_28125_, _28124_, _28119_);
  and (_28126_, _28125_, _03531_);
  nor (_28127_, _28105_, _03531_);
  or (_28128_, _28127_, _28126_);
  and (_28129_, _28128_, _04577_);
  and (_28130_, _10728_, \oc8051_golden_model_1.SP [0]);
  nor (_28131_, _27996_, \oc8051_golden_model_1.SP [5]);
  nor (_28132_, _28131_, _28130_);
  and (_28134_, _28132_, _03464_);
  nor (_28135_, _28134_, _04756_);
  not (_28136_, _28135_);
  nor (_28137_, _28136_, _28129_);
  and (_28138_, _28108_, _04756_);
  or (_28139_, _28138_, _07454_);
  nor (_28140_, _28139_, _28137_);
  nor (_28141_, _28140_, _28099_);
  and (_28142_, _06757_, _05323_);
  nor (_28143_, _28092_, _04500_);
  not (_28145_, _28143_);
  nor (_28146_, _28145_, _28142_);
  or (_28147_, _28146_, _03224_);
  nor (_28148_, _28147_, _28141_);
  nor (_28149_, _13184_, _10741_);
  nor (_28150_, _28149_, _28092_);
  nor (_28151_, _28150_, _03521_);
  or (_28152_, _28151_, _03624_);
  or (_28153_, _28152_, _28148_);
  and (_28154_, _06295_, _05323_);
  nor (_28156_, _28154_, _28092_);
  nand (_28157_, _28156_, _03624_);
  and (_28158_, _28157_, _28153_);
  nor (_28159_, _28158_, _03168_);
  and (_28160_, _28108_, _03168_);
  nor (_28161_, _28160_, _28159_);
  nor (_28162_, _28161_, _03623_);
  and (_28163_, _13198_, _05323_);
  or (_28164_, _28092_, _04527_);
  nor (_28165_, _28164_, _28163_);
  or (_28167_, _28165_, _03744_);
  nor (_28168_, _28167_, _28162_);
  nor (_28169_, _28168_, _28095_);
  nor (_28170_, _28169_, _03611_);
  nor (_28171_, _28092_, _05576_);
  not (_28172_, _28171_);
  nor (_28173_, _28156_, _04523_);
  and (_28174_, _28173_, _28172_);
  nor (_28175_, _28174_, _28170_);
  nor (_28176_, _28175_, _10829_);
  nor (_28178_, _28105_, _03734_);
  and (_28179_, _28178_, _28172_);
  and (_28180_, _28090_, _03182_);
  nor (_28181_, _28180_, _28179_);
  and (_28182_, _28181_, _06453_);
  not (_28183_, _28182_);
  nor (_28184_, _28183_, _28176_);
  nor (_28185_, _13197_, _10741_);
  nor (_28186_, _28185_, _28092_);
  and (_28187_, _28186_, _03618_);
  nor (_28189_, _28187_, _28184_);
  nor (_28190_, _28189_, _03741_);
  nor (_28191_, _13203_, _10741_);
  or (_28192_, _28092_, _06458_);
  nor (_28193_, _28192_, _28191_);
  or (_28194_, _28193_, _03752_);
  nor (_28195_, _28194_, _28190_);
  nor (_28196_, _10771_, _10769_);
  nor (_28197_, _28196_, _10772_);
  nor (_28198_, _28197_, _10735_);
  or (_28200_, _28198_, _28195_);
  and (_28201_, _28200_, _04803_);
  and (_28202_, _28090_, _03191_);
  or (_28203_, _28202_, _28201_);
  and (_28204_, _28203_, _03476_);
  nor (_28205_, _28197_, _03476_);
  or (_28206_, _28205_, _28204_);
  and (_28207_, _28206_, _03948_);
  nor (_28208_, _28102_, _03948_);
  nor (_28209_, _28208_, _04986_);
  not (_28211_, _28209_);
  nor (_28212_, _28211_, _28207_);
  nor (_28213_, _28212_, _28091_);
  nor (_28214_, _28213_, _03473_);
  and (_28215_, _13253_, _05323_);
  nor (_28216_, _28215_, _28092_);
  and (_28217_, _28216_, _03473_);
  nor (_28218_, _28217_, _28214_);
  or (_28219_, _28218_, _43193_);
  or (_28220_, _43189_, \oc8051_golden_model_1.SP [5]);
  and (_28222_, _28220_, _42003_);
  and (_43862_, _28222_, _28219_);
  nor (_28223_, _05323_, _10768_);
  and (_28224_, _13407_, _05323_);
  or (_28225_, _28224_, _28223_);
  and (_28226_, _28225_, _03744_);
  nor (_28227_, _13293_, _10741_);
  or (_28228_, _28227_, _28223_);
  or (_28229_, _28228_, _04432_);
  and (_28230_, _05323_, \oc8051_golden_model_1.ACC [6]);
  or (_28232_, _28230_, _28223_);
  and (_28233_, _28232_, _04436_);
  and (_28234_, _10754_, \oc8051_golden_model_1.SP [6]);
  nor (_28235_, _10728_, \oc8051_golden_model_1.SP [6]);
  nor (_28236_, _28235_, _10729_);
  and (_28237_, _28236_, _04435_);
  or (_28238_, _28237_, _03534_);
  or (_28239_, _28238_, _28234_);
  or (_28240_, _28239_, _28233_);
  and (_28241_, _28240_, _03202_);
  and (_28242_, _28241_, _28229_);
  and (_28243_, _28236_, _05977_);
  or (_28244_, _28243_, _03527_);
  or (_28245_, _28244_, _28242_);
  nor (_28246_, _28120_, _10768_);
  nor (_28247_, _28246_, _10774_);
  nand (_28248_, _28247_, _03527_);
  and (_28249_, _28248_, _28245_);
  or (_28250_, _28249_, _03530_);
  or (_28251_, _28232_, _03531_);
  and (_28254_, _28251_, _04577_);
  and (_28255_, _28254_, _28250_);
  nor (_28256_, _28130_, \oc8051_golden_model_1.SP [6]);
  nor (_28257_, _28256_, _10784_);
  and (_28258_, _28257_, _03464_);
  or (_28259_, _28258_, _28255_);
  and (_28260_, _28259_, _04757_);
  nand (_28261_, _28236_, _04756_);
  nand (_28262_, _28261_, _06903_);
  or (_28263_, _28262_, _28260_);
  nor (_28265_, _05417_, _10741_);
  or (_28266_, _28223_, _06903_);
  or (_28267_, _28266_, _28265_);
  and (_28268_, _28267_, _28263_);
  or (_28269_, _28268_, _04082_);
  and (_28270_, _06526_, _05323_);
  or (_28271_, _28223_, _04500_);
  or (_28272_, _28271_, _28270_);
  and (_28273_, _28272_, _03521_);
  and (_28274_, _28273_, _28269_);
  nor (_28276_, _13387_, _10741_);
  or (_28277_, _28276_, _28223_);
  and (_28278_, _28277_, _03224_);
  or (_28279_, _28278_, _03624_);
  or (_28280_, _28279_, _28274_);
  and (_28281_, _14949_, _05323_);
  or (_28282_, _28281_, _28223_);
  or (_28283_, _28282_, _04509_);
  and (_28284_, _28283_, _28280_);
  or (_28285_, _28284_, _03168_);
  or (_28287_, _28236_, _27595_);
  and (_28288_, _28287_, _28285_);
  or (_28289_, _28288_, _03623_);
  and (_28290_, _13402_, _05323_);
  or (_28291_, _28290_, _28223_);
  or (_28292_, _28291_, _04527_);
  and (_28293_, _28292_, _03745_);
  and (_28294_, _28293_, _28289_);
  or (_28295_, _28294_, _28226_);
  and (_28296_, _28295_, _04523_);
  or (_28298_, _28223_, _05469_);
  and (_28299_, _28282_, _03611_);
  and (_28300_, _28299_, _28298_);
  or (_28301_, _28300_, _28296_);
  and (_28302_, _28301_, _10828_);
  and (_28303_, _28232_, _03733_);
  and (_28304_, _28303_, _28298_);
  and (_28305_, _28236_, _03182_);
  or (_28306_, _28305_, _03618_);
  or (_28307_, _28306_, _28304_);
  or (_28309_, _28307_, _28302_);
  nor (_28310_, _13400_, _10741_);
  or (_28311_, _28310_, _28223_);
  or (_28312_, _28311_, _06453_);
  and (_28313_, _28312_, _28309_);
  or (_28314_, _28313_, _03741_);
  nor (_28315_, _13406_, _10741_);
  or (_28316_, _28223_, _06458_);
  or (_28317_, _28316_, _28315_);
  and (_28318_, _28317_, _10735_);
  and (_28320_, _28318_, _28314_);
  nor (_28321_, _10772_, _10768_);
  or (_28322_, _28321_, _10773_);
  and (_28323_, _28322_, _03752_);
  or (_28324_, _28323_, _03191_);
  or (_28325_, _28324_, _28320_);
  or (_28326_, _28236_, _04803_);
  and (_28327_, _28326_, _03476_);
  and (_28328_, _28327_, _28325_);
  and (_28329_, _28322_, _03475_);
  or (_28331_, _28329_, _03767_);
  or (_28332_, _28331_, _28328_);
  or (_28333_, _28228_, _03948_);
  and (_28334_, _28333_, _04553_);
  and (_28335_, _28334_, _28332_);
  and (_28336_, _28236_, _04986_);
  or (_28337_, _28336_, _03473_);
  or (_28338_, _28337_, _28335_);
  and (_28339_, _13456_, _05323_);
  or (_28340_, _28223_, _03474_);
  or (_28342_, _28340_, _28339_);
  and (_28343_, _28342_, _28338_);
  or (_28344_, _28343_, _43193_);
  or (_28345_, _43189_, \oc8051_golden_model_1.SP [6]);
  and (_28346_, _28345_, _42003_);
  and (_43865_, _28346_, _28344_);
  not (_28347_, \oc8051_golden_model_1.TCON [0]);
  nor (_28348_, _05286_, _28347_);
  and (_28349_, _12183_, _05286_);
  nor (_28350_, _28349_, _28348_);
  nor (_28352_, _28350_, _03745_);
  and (_28353_, _05286_, _06350_);
  nor (_28354_, _28353_, _28348_);
  and (_28355_, _28354_, _03624_);
  and (_28356_, _05286_, _04429_);
  nor (_28357_, _28356_, _28348_);
  and (_28358_, _28357_, _07454_);
  and (_28359_, _05286_, \oc8051_golden_model_1.ACC [0]);
  nor (_28360_, _28359_, _28348_);
  nor (_28361_, _28360_, _04437_);
  nor (_28363_, _04436_, _28347_);
  or (_28364_, _28363_, _28361_);
  and (_28365_, _28364_, _04432_);
  nor (_28366_, _05722_, _10876_);
  nor (_28367_, _28366_, _28348_);
  nor (_28368_, _28367_, _04432_);
  or (_28369_, _28368_, _28365_);
  and (_28370_, _28369_, _03470_);
  nor (_28371_, _05924_, _28347_);
  and (_28372_, _12075_, _05924_);
  nor (_28374_, _28372_, _28371_);
  nor (_28375_, _28374_, _03470_);
  nor (_28376_, _28375_, _28370_);
  nor (_28377_, _28376_, _03527_);
  nor (_28378_, _28357_, _04457_);
  or (_28379_, _28378_, _28377_);
  and (_28380_, _28379_, _03531_);
  nor (_28381_, _28360_, _03531_);
  or (_28382_, _28381_, _28380_);
  and (_28383_, _28382_, _03466_);
  and (_28385_, _28348_, _03465_);
  or (_28386_, _28385_, _28383_);
  and (_28387_, _28386_, _03459_);
  nor (_28388_, _28367_, _03459_);
  or (_28389_, _28388_, _28387_);
  and (_28390_, _28389_, _03453_);
  nor (_28391_, _12106_, _10913_);
  nor (_28392_, _28391_, _28371_);
  nor (_28393_, _28392_, _03453_);
  or (_28394_, _28393_, _07454_);
  nor (_28396_, _28394_, _28390_);
  nor (_28397_, _28396_, _28358_);
  nor (_28398_, _28397_, _04082_);
  and (_28399_, _06617_, _05286_);
  nor (_28400_, _28348_, _04500_);
  not (_28401_, _28400_);
  nor (_28402_, _28401_, _28399_);
  or (_28403_, _28402_, _03224_);
  nor (_28404_, _28403_, _28398_);
  nor (_28405_, _12164_, _10876_);
  nor (_28407_, _28405_, _28348_);
  nor (_28408_, _28407_, _03521_);
  or (_28409_, _28408_, _03624_);
  nor (_28410_, _28409_, _28404_);
  nor (_28411_, _28410_, _28355_);
  or (_28412_, _28411_, _03623_);
  and (_28413_, _12177_, _05286_);
  or (_28414_, _28413_, _28348_);
  or (_28415_, _28414_, _04527_);
  and (_28416_, _28415_, _03745_);
  and (_28418_, _28416_, _28412_);
  nor (_28419_, _28418_, _28352_);
  nor (_28420_, _28419_, _03611_);
  or (_28421_, _28354_, _04523_);
  nor (_28422_, _28421_, _28366_);
  nor (_28423_, _28422_, _28420_);
  nor (_28424_, _28423_, _03733_);
  and (_28425_, _12182_, _05286_);
  or (_28426_, _28425_, _28348_);
  and (_28427_, _28426_, _03733_);
  or (_28428_, _28427_, _28424_);
  and (_28429_, _28428_, _06453_);
  nor (_28430_, _12057_, _10876_);
  nor (_28431_, _28430_, _28348_);
  nor (_28432_, _28431_, _06453_);
  or (_28433_, _28432_, _28429_);
  and (_28434_, _28433_, _06458_);
  nor (_28435_, _12181_, _10876_);
  nor (_28436_, _28435_, _28348_);
  nor (_28437_, _28436_, _06458_);
  or (_28440_, _28437_, _28434_);
  and (_28441_, _28440_, _03948_);
  nor (_28442_, _28367_, _03948_);
  or (_28443_, _28442_, _28441_);
  and (_28444_, _28443_, _03446_);
  and (_28445_, _28348_, _03445_);
  nor (_28446_, _28445_, _03473_);
  not (_28447_, _28446_);
  nor (_28448_, _28447_, _28444_);
  and (_28449_, _28367_, _03473_);
  or (_28451_, _28449_, _28448_);
  nand (_28452_, _28451_, _43189_);
  or (_28453_, _43189_, \oc8051_golden_model_1.TCON [0]);
  and (_28454_, _28453_, _42003_);
  and (_43866_, _28454_, _28452_);
  or (_28455_, _05286_, \oc8051_golden_model_1.TCON [1]);
  and (_28456_, _12265_, _05286_);
  not (_28457_, _28456_);
  and (_28458_, _28457_, _28455_);
  or (_28459_, _28458_, _04432_);
  nand (_28461_, _05286_, _03269_);
  and (_28462_, _28461_, _28455_);
  and (_28463_, _28462_, _04436_);
  and (_28464_, _04437_, \oc8051_golden_model_1.TCON [1]);
  or (_28465_, _28464_, _03534_);
  or (_28466_, _28465_, _28463_);
  and (_28467_, _28466_, _03470_);
  and (_28468_, _28467_, _28459_);
  and (_28469_, _12269_, _05924_);
  and (_28470_, _10913_, \oc8051_golden_model_1.TCON [1]);
  or (_28472_, _28470_, _03527_);
  or (_28473_, _28472_, _28469_);
  and (_28474_, _28473_, _03533_);
  or (_28475_, _28474_, _28468_);
  and (_28476_, _10876_, \oc8051_golden_model_1.TCON [1]);
  nor (_28477_, _10876_, _04635_);
  or (_28478_, _28477_, _28476_);
  or (_28479_, _28478_, _04457_);
  and (_28480_, _28479_, _28475_);
  or (_28481_, _28480_, _03530_);
  or (_28483_, _28462_, _03531_);
  and (_28484_, _28483_, _03466_);
  and (_28485_, _28484_, _28481_);
  and (_28486_, _12256_, _05924_);
  or (_28487_, _28486_, _28470_);
  and (_28488_, _28487_, _03465_);
  or (_28489_, _28488_, _03458_);
  or (_28490_, _28489_, _28485_);
  and (_28491_, _28469_, _12284_);
  or (_28492_, _28470_, _03459_);
  or (_28494_, _28492_, _28491_);
  and (_28495_, _28494_, _28490_);
  and (_28496_, _28495_, _03453_);
  nor (_28497_, _12301_, _10913_);
  or (_28498_, _28470_, _28497_);
  and (_28499_, _28498_, _03452_);
  or (_28500_, _28499_, _07454_);
  or (_28501_, _28500_, _28496_);
  or (_28502_, _28478_, _06903_);
  and (_28503_, _28502_, _28501_);
  or (_28505_, _28503_, _04082_);
  and (_28506_, _06572_, _05286_);
  or (_28507_, _28476_, _04500_);
  or (_28508_, _28507_, _28506_);
  and (_28509_, _28508_, _03521_);
  and (_28510_, _28509_, _28505_);
  nor (_28511_, _12360_, _10876_);
  or (_28512_, _28511_, _28476_);
  and (_28513_, _28512_, _03224_);
  or (_28514_, _28513_, _28510_);
  and (_28516_, _28514_, _03625_);
  or (_28517_, _12375_, _10876_);
  and (_28518_, _28517_, _03623_);
  nand (_28519_, _05286_, _04325_);
  and (_28520_, _28519_, _03624_);
  or (_28521_, _28520_, _28518_);
  and (_28522_, _28521_, _28455_);
  or (_28523_, _28522_, _28516_);
  and (_28524_, _28523_, _03745_);
  or (_28525_, _12381_, _10876_);
  and (_28527_, _28455_, _03744_);
  and (_28528_, _28527_, _28525_);
  or (_28529_, _28528_, _28524_);
  and (_28530_, _28529_, _04523_);
  or (_28531_, _12374_, _10876_);
  and (_28532_, _28455_, _03611_);
  and (_28533_, _28532_, _28531_);
  or (_28534_, _28533_, _28530_);
  and (_28535_, _28534_, _03734_);
  or (_28536_, _28476_, _05674_);
  and (_28538_, _28462_, _03733_);
  and (_28539_, _28538_, _28536_);
  or (_28540_, _28539_, _28535_);
  and (_28541_, _28540_, _03742_);
  or (_28542_, _28519_, _05674_);
  and (_28543_, _28455_, _03618_);
  and (_28544_, _28543_, _28542_);
  or (_28545_, _28461_, _05674_);
  and (_28546_, _28455_, _03741_);
  and (_28547_, _28546_, _28545_);
  or (_28549_, _28547_, _03767_);
  or (_28550_, _28549_, _28544_);
  or (_28551_, _28550_, _28541_);
  or (_28552_, _28458_, _03948_);
  and (_28553_, _28552_, _03446_);
  and (_28554_, _28553_, _28551_);
  and (_28555_, _28487_, _03445_);
  or (_28556_, _28555_, _03473_);
  or (_28557_, _28556_, _28554_);
  or (_28558_, _28476_, _03474_);
  or (_28560_, _28558_, _28456_);
  and (_28561_, _28560_, _28557_);
  and (_28562_, _28561_, _43189_);
  nor (_28563_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_28564_, _28563_, _00001_);
  or (_43867_, _28564_, _28562_);
  not (_28565_, \oc8051_golden_model_1.TCON [2]);
  nor (_28566_, _05286_, _28565_);
  and (_28567_, _05286_, _06399_);
  nor (_28568_, _28567_, _28566_);
  and (_28570_, _28568_, _03624_);
  nor (_28571_, _10876_, _05073_);
  nor (_28572_, _28571_, _28566_);
  and (_28573_, _28572_, _07454_);
  and (_28574_, _05286_, \oc8051_golden_model_1.ACC [2]);
  nor (_28575_, _28574_, _28566_);
  nor (_28576_, _28575_, _04437_);
  nor (_28577_, _04436_, _28565_);
  or (_28578_, _28577_, _28576_);
  and (_28579_, _28578_, _04432_);
  nor (_28581_, _12467_, _10876_);
  nor (_28582_, _28581_, _28566_);
  nor (_28583_, _28582_, _04432_);
  or (_28584_, _28583_, _28579_);
  and (_28585_, _28584_, _03470_);
  nor (_28586_, _05924_, _28565_);
  and (_28587_, _12462_, _05924_);
  nor (_28588_, _28587_, _28586_);
  nor (_28589_, _28588_, _03470_);
  or (_28590_, _28589_, _28585_);
  and (_28592_, _28590_, _04457_);
  nor (_28593_, _28572_, _04457_);
  or (_28594_, _28593_, _28592_);
  and (_28595_, _28594_, _03531_);
  nor (_28596_, _28575_, _03531_);
  or (_28597_, _28596_, _28595_);
  and (_28598_, _28597_, _03466_);
  and (_28599_, _12460_, _05924_);
  nor (_28600_, _28599_, _28586_);
  nor (_28601_, _28600_, _03466_);
  or (_28603_, _28601_, _03458_);
  or (_28604_, _28603_, _28598_);
  and (_28605_, _28587_, _12491_);
  or (_28606_, _28586_, _03459_);
  or (_28607_, _28606_, _28605_);
  and (_28608_, _28607_, _03453_);
  and (_28609_, _28608_, _28604_);
  nor (_28610_, _12509_, _10913_);
  nor (_28611_, _28610_, _28586_);
  nor (_28612_, _28611_, _03453_);
  nor (_28614_, _28612_, _07454_);
  not (_28615_, _28614_);
  nor (_28616_, _28615_, _28609_);
  nor (_28617_, _28616_, _28573_);
  nor (_28618_, _28617_, _04082_);
  and (_28619_, _06710_, _05286_);
  nor (_28620_, _28566_, _04500_);
  not (_28621_, _28620_);
  nor (_28622_, _28621_, _28619_);
  or (_28623_, _28622_, _03224_);
  nor (_28625_, _28623_, _28618_);
  nor (_28626_, _12568_, _10876_);
  nor (_28627_, _28566_, _28626_);
  nor (_28628_, _28627_, _03521_);
  or (_28629_, _28628_, _03624_);
  nor (_28630_, _28629_, _28625_);
  nor (_28631_, _28630_, _28570_);
  or (_28632_, _28631_, _03623_);
  and (_28633_, _12582_, _05286_);
  or (_28634_, _28633_, _28566_);
  or (_28636_, _28634_, _04527_);
  and (_28637_, _28636_, _03745_);
  and (_28638_, _28637_, _28632_);
  and (_28639_, _12588_, _05286_);
  nor (_28640_, _28639_, _28566_);
  nor (_28641_, _28640_, _03745_);
  nor (_28642_, _28641_, _28638_);
  nor (_28643_, _28642_, _03611_);
  nor (_28644_, _28566_, _05772_);
  not (_28645_, _28644_);
  nor (_28647_, _28568_, _04523_);
  and (_28648_, _28647_, _28645_);
  nor (_28649_, _28648_, _28643_);
  nor (_28650_, _28649_, _03733_);
  nor (_28651_, _28575_, _03734_);
  and (_28652_, _28651_, _28645_);
  or (_28653_, _28652_, _28650_);
  and (_28654_, _28653_, _06453_);
  nor (_28655_, _12581_, _10876_);
  nor (_28656_, _28655_, _28566_);
  nor (_28658_, _28656_, _06453_);
  or (_28659_, _28658_, _28654_);
  and (_28660_, _28659_, _06458_);
  nor (_28661_, _12587_, _10876_);
  nor (_28662_, _28661_, _28566_);
  nor (_28663_, _28662_, _06458_);
  or (_28664_, _28663_, _28660_);
  and (_28665_, _28664_, _03948_);
  nor (_28666_, _28582_, _03948_);
  or (_28667_, _28666_, _28665_);
  and (_28669_, _28667_, _03446_);
  nor (_28670_, _28600_, _03446_);
  nor (_28671_, _28670_, _03473_);
  not (_28672_, _28671_);
  nor (_28673_, _28672_, _28669_);
  and (_28674_, _12638_, _05286_);
  or (_28675_, _28566_, _03474_);
  nor (_28676_, _28675_, _28674_);
  nor (_28677_, _28676_, _28673_);
  or (_28678_, _28677_, _43193_);
  or (_28680_, _43189_, \oc8051_golden_model_1.TCON [2]);
  and (_28681_, _28680_, _42003_);
  and (_43868_, _28681_, _28678_);
  not (_28682_, \oc8051_golden_model_1.TCON [3]);
  nor (_28683_, _05286_, _28682_);
  and (_28684_, _05286_, _06356_);
  nor (_28685_, _28684_, _28683_);
  and (_28686_, _28685_, _03624_);
  nor (_28687_, _10876_, _04885_);
  nor (_28688_, _28687_, _28683_);
  and (_28690_, _28688_, _07454_);
  and (_28691_, _05286_, \oc8051_golden_model_1.ACC [3]);
  nor (_28692_, _28691_, _28683_);
  nor (_28693_, _28692_, _04437_);
  nor (_28694_, _04436_, _28682_);
  or (_28695_, _28694_, _28693_);
  and (_28696_, _28695_, _04432_);
  nor (_28697_, _12652_, _10876_);
  nor (_28698_, _28697_, _28683_);
  nor (_28699_, _28698_, _04432_);
  or (_28701_, _28699_, _28696_);
  and (_28702_, _28701_, _03470_);
  nor (_28703_, _05924_, _28682_);
  and (_28704_, _12664_, _05924_);
  nor (_28705_, _28704_, _28703_);
  nor (_28706_, _28705_, _03470_);
  or (_28707_, _28706_, _03527_);
  or (_28708_, _28707_, _28702_);
  nand (_28709_, _28688_, _03527_);
  and (_28710_, _28709_, _28708_);
  and (_28712_, _28710_, _03531_);
  nor (_28713_, _28692_, _03531_);
  or (_28714_, _28713_, _28712_);
  and (_28715_, _28714_, _03466_);
  and (_28716_, _12662_, _05924_);
  nor (_28717_, _28716_, _28703_);
  nor (_28718_, _28717_, _03466_);
  or (_28719_, _28718_, _28715_);
  and (_28720_, _28719_, _03459_);
  nor (_28721_, _28703_, _12691_);
  nor (_28723_, _28721_, _28705_);
  and (_28724_, _28723_, _03458_);
  or (_28725_, _28724_, _28720_);
  and (_28726_, _28725_, _03453_);
  nor (_28727_, _12709_, _10913_);
  nor (_28728_, _28727_, _28703_);
  nor (_28729_, _28728_, _03453_);
  nor (_28730_, _28729_, _07454_);
  not (_28731_, _28730_);
  nor (_28732_, _28731_, _28726_);
  nor (_28734_, _28732_, _28690_);
  nor (_28735_, _28734_, _04082_);
  and (_28736_, _06664_, _05286_);
  nor (_28737_, _28683_, _04500_);
  not (_28738_, _28737_);
  nor (_28739_, _28738_, _28736_);
  or (_28740_, _28739_, _03224_);
  nor (_28741_, _28740_, _28735_);
  nor (_28742_, _12773_, _10876_);
  nor (_28743_, _28683_, _28742_);
  nor (_28745_, _28743_, _03521_);
  or (_28746_, _28745_, _03624_);
  nor (_28747_, _28746_, _28741_);
  nor (_28748_, _28747_, _28686_);
  or (_28749_, _28748_, _03623_);
  and (_28750_, _12787_, _05286_);
  or (_28751_, _28750_, _28683_);
  or (_28752_, _28751_, _04527_);
  and (_28753_, _28752_, _03745_);
  and (_28754_, _28753_, _28749_);
  and (_28756_, _12793_, _05286_);
  nor (_28757_, _28756_, _28683_);
  nor (_28758_, _28757_, _03745_);
  nor (_28759_, _28758_, _28754_);
  nor (_28760_, _28759_, _03611_);
  nor (_28761_, _28683_, _05625_);
  not (_28762_, _28761_);
  nor (_28763_, _28685_, _04523_);
  and (_28764_, _28763_, _28762_);
  nor (_28765_, _28764_, _28760_);
  nor (_28767_, _28765_, _03733_);
  nor (_28768_, _28692_, _03734_);
  and (_28769_, _28768_, _28762_);
  or (_28770_, _28769_, _28767_);
  and (_28771_, _28770_, _06453_);
  nor (_28772_, _12786_, _10876_);
  nor (_28773_, _28772_, _28683_);
  nor (_28774_, _28773_, _06453_);
  or (_28775_, _28774_, _28771_);
  and (_28776_, _28775_, _06458_);
  nor (_28778_, _12792_, _10876_);
  nor (_28779_, _28778_, _28683_);
  nor (_28780_, _28779_, _06458_);
  or (_28781_, _28780_, _28776_);
  and (_28782_, _28781_, _03948_);
  nor (_28783_, _28698_, _03948_);
  or (_28784_, _28783_, _28782_);
  and (_28785_, _28784_, _03446_);
  nor (_28786_, _28717_, _03446_);
  nor (_28787_, _28786_, _03473_);
  not (_28789_, _28787_);
  nor (_28790_, _28789_, _28785_);
  and (_28791_, _12843_, _05286_);
  or (_28792_, _28683_, _03474_);
  nor (_28793_, _28792_, _28791_);
  nor (_28794_, _28793_, _28790_);
  or (_28795_, _28794_, _43193_);
  or (_28796_, _43189_, \oc8051_golden_model_1.TCON [3]);
  and (_28797_, _28796_, _42003_);
  and (_43869_, _28797_, _28795_);
  not (_28799_, \oc8051_golden_model_1.TCON [4]);
  nor (_28800_, _05286_, _28799_);
  nor (_28801_, _05831_, _10876_);
  nor (_28802_, _28801_, _28800_);
  and (_28803_, _28802_, _07454_);
  nor (_28804_, _05924_, _28799_);
  and (_28805_, _12864_, _05924_);
  nor (_28806_, _28805_, _28804_);
  nor (_28807_, _28806_, _03466_);
  and (_28808_, _05286_, \oc8051_golden_model_1.ACC [4]);
  nor (_28810_, _28808_, _28800_);
  nor (_28811_, _28810_, _04437_);
  nor (_28812_, _04436_, _28799_);
  or (_28813_, _28812_, _28811_);
  and (_28814_, _28813_, _04432_);
  nor (_28815_, _12856_, _10876_);
  nor (_28816_, _28815_, _28800_);
  nor (_28817_, _28816_, _04432_);
  or (_28818_, _28817_, _28814_);
  and (_28819_, _28818_, _03470_);
  and (_28821_, _12866_, _05924_);
  nor (_28822_, _28821_, _28804_);
  nor (_28823_, _28822_, _03470_);
  or (_28824_, _28823_, _03527_);
  or (_28825_, _28824_, _28819_);
  nand (_28826_, _28802_, _03527_);
  and (_28827_, _28826_, _28825_);
  and (_28828_, _28827_, _03531_);
  nor (_28829_, _28810_, _03531_);
  or (_28830_, _28829_, _28828_);
  and (_28832_, _28830_, _03466_);
  nor (_28833_, _28832_, _28807_);
  nor (_28834_, _28833_, _03458_);
  nor (_28835_, _28804_, _12894_);
  or (_28836_, _28822_, _03459_);
  nor (_28837_, _28836_, _28835_);
  nor (_28838_, _28837_, _28834_);
  nor (_28839_, _28838_, _03452_);
  nor (_28840_, _12912_, _10913_);
  nor (_28841_, _28840_, _28804_);
  nor (_28843_, _28841_, _03453_);
  nor (_28844_, _28843_, _07454_);
  not (_28845_, _28844_);
  nor (_28846_, _28845_, _28839_);
  nor (_28847_, _28846_, _28803_);
  nor (_28848_, _28847_, _04082_);
  and (_28849_, _06802_, _05286_);
  nor (_28850_, _28800_, _04500_);
  not (_28851_, _28850_);
  nor (_28852_, _28851_, _28849_);
  nor (_28854_, _28852_, _03224_);
  not (_28855_, _28854_);
  nor (_28856_, _28855_, _28848_);
  nor (_28857_, _12972_, _10876_);
  nor (_28858_, _28857_, _28800_);
  nor (_28859_, _28858_, _03521_);
  or (_28860_, _28859_, _08905_);
  or (_28861_, _28860_, _28856_);
  and (_28862_, _12986_, _05286_);
  or (_28863_, _28800_, _04527_);
  or (_28865_, _28863_, _28862_);
  and (_28866_, _06337_, _05286_);
  nor (_28867_, _28866_, _28800_);
  and (_28868_, _28867_, _03624_);
  nor (_28869_, _28868_, _03744_);
  and (_28870_, _28869_, _28865_);
  and (_28871_, _28870_, _28861_);
  and (_28872_, _12992_, _05286_);
  nor (_28873_, _28872_, _28800_);
  nor (_28874_, _28873_, _03745_);
  nor (_28876_, _28874_, _28871_);
  nor (_28877_, _28876_, _03611_);
  nor (_28878_, _28800_, _05880_);
  not (_28879_, _28878_);
  nor (_28880_, _28867_, _04523_);
  and (_28881_, _28880_, _28879_);
  nor (_28882_, _28881_, _28877_);
  nor (_28883_, _28882_, _03733_);
  nor (_28884_, _28810_, _03734_);
  and (_28885_, _28884_, _28879_);
  or (_28887_, _28885_, _28883_);
  and (_28888_, _28887_, _06453_);
  nor (_28889_, _12985_, _10876_);
  nor (_28890_, _28889_, _28800_);
  nor (_28891_, _28890_, _06453_);
  or (_28892_, _28891_, _28888_);
  and (_28893_, _28892_, _06458_);
  nor (_28894_, _12991_, _10876_);
  nor (_28895_, _28894_, _28800_);
  nor (_28896_, _28895_, _06458_);
  or (_28897_, _28896_, _28893_);
  and (_28898_, _28897_, _03948_);
  nor (_28899_, _28816_, _03948_);
  or (_28900_, _28899_, _28898_);
  and (_28901_, _28900_, _03446_);
  nor (_28902_, _28806_, _03446_);
  nor (_28903_, _28902_, _03473_);
  not (_28904_, _28903_);
  nor (_28905_, _28904_, _28901_);
  and (_28906_, _13051_, _05286_);
  or (_28908_, _28800_, _03474_);
  nor (_28909_, _28908_, _28906_);
  nor (_28910_, _28909_, _28905_);
  or (_28911_, _28910_, _43193_);
  or (_28912_, _43189_, \oc8051_golden_model_1.TCON [4]);
  and (_28913_, _28912_, _42003_);
  and (_43870_, _28913_, _28911_);
  not (_28914_, \oc8051_golden_model_1.TCON [5]);
  nor (_28915_, _05286_, _28914_);
  and (_28916_, _06757_, _05286_);
  or (_28918_, _28916_, _28915_);
  and (_28919_, _28918_, _04082_);
  and (_28920_, _05286_, \oc8051_golden_model_1.ACC [5]);
  nor (_28921_, _28920_, _28915_);
  nor (_28922_, _28921_, _04437_);
  nor (_28923_, _04436_, _28914_);
  or (_28924_, _28923_, _28922_);
  and (_28925_, _28924_, _04432_);
  nor (_28926_, _13070_, _10876_);
  nor (_28927_, _28926_, _28915_);
  nor (_28929_, _28927_, _04432_);
  or (_28930_, _28929_, _28925_);
  and (_28931_, _28930_, _03470_);
  nor (_28932_, _05924_, _28914_);
  and (_28933_, _13095_, _05924_);
  nor (_28934_, _28933_, _28932_);
  nor (_28935_, _28934_, _03470_);
  or (_28936_, _28935_, _03527_);
  or (_28937_, _28936_, _28931_);
  nor (_28938_, _05526_, _10876_);
  nor (_28940_, _28938_, _28915_);
  nand (_28941_, _28940_, _03527_);
  and (_28942_, _28941_, _28937_);
  and (_28943_, _28942_, _03531_);
  nor (_28944_, _28921_, _03531_);
  or (_28945_, _28944_, _28943_);
  and (_28946_, _28945_, _03466_);
  and (_28947_, _13078_, _05924_);
  nor (_28948_, _28947_, _28932_);
  nor (_28949_, _28948_, _03466_);
  or (_28951_, _28949_, _03458_);
  or (_28952_, _28951_, _28946_);
  nor (_28953_, _28932_, _13110_);
  nor (_28954_, _28953_, _28934_);
  or (_28955_, _28954_, _03459_);
  and (_28956_, _28955_, _03453_);
  and (_28957_, _28956_, _28952_);
  nor (_28958_, _13076_, _10913_);
  nor (_28959_, _28958_, _28932_);
  nor (_28960_, _28959_, _03453_);
  nor (_28961_, _28960_, _07454_);
  not (_28962_, _28961_);
  nor (_28963_, _28962_, _28957_);
  and (_28964_, _28940_, _07454_);
  or (_28965_, _28964_, _04082_);
  nor (_28966_, _28965_, _28963_);
  or (_28967_, _28966_, _28919_);
  and (_28968_, _28967_, _03521_);
  nor (_28969_, _13184_, _10876_);
  nor (_28970_, _28969_, _28915_);
  nor (_28973_, _28970_, _03521_);
  or (_28974_, _28973_, _08905_);
  or (_28975_, _28974_, _28968_);
  and (_28976_, _13198_, _05286_);
  or (_28977_, _28915_, _04527_);
  or (_28978_, _28977_, _28976_);
  and (_28979_, _06295_, _05286_);
  nor (_28980_, _28979_, _28915_);
  and (_28981_, _28980_, _03624_);
  nor (_28982_, _28981_, _03744_);
  and (_28984_, _28982_, _28978_);
  and (_28985_, _28984_, _28975_);
  and (_28986_, _13204_, _05286_);
  nor (_28987_, _28986_, _28915_);
  nor (_28988_, _28987_, _03745_);
  nor (_28989_, _28988_, _28985_);
  nor (_28990_, _28989_, _03611_);
  nor (_28991_, _28915_, _05576_);
  not (_28992_, _28991_);
  nor (_28993_, _28980_, _04523_);
  and (_28995_, _28993_, _28992_);
  nor (_28996_, _28995_, _28990_);
  nor (_28997_, _28996_, _03733_);
  nor (_28998_, _28921_, _03734_);
  and (_28999_, _28998_, _28992_);
  nor (_29000_, _28999_, _03618_);
  not (_29001_, _29000_);
  nor (_29002_, _29001_, _28997_);
  nor (_29003_, _13197_, _10876_);
  or (_29004_, _28915_, _06453_);
  nor (_29006_, _29004_, _29003_);
  or (_29007_, _29006_, _03741_);
  nor (_29008_, _29007_, _29002_);
  nor (_29009_, _13203_, _10876_);
  nor (_29010_, _29009_, _28915_);
  nor (_29011_, _29010_, _06458_);
  or (_29012_, _29011_, _29008_);
  and (_29013_, _29012_, _03948_);
  nor (_29014_, _28927_, _03948_);
  or (_29015_, _29014_, _29013_);
  and (_29017_, _29015_, _03446_);
  nor (_29018_, _28948_, _03446_);
  or (_29019_, _29018_, _29017_);
  and (_29020_, _29019_, _03474_);
  and (_29021_, _13253_, _05286_);
  nor (_29022_, _29021_, _28915_);
  nor (_29023_, _29022_, _03474_);
  or (_29024_, _29023_, _29020_);
  or (_29025_, _29024_, _43193_);
  or (_29026_, _43189_, \oc8051_golden_model_1.TCON [5]);
  and (_29028_, _29026_, _42003_);
  and (_43871_, _29028_, _29025_);
  not (_29029_, \oc8051_golden_model_1.TCON [6]);
  nor (_29030_, _05286_, _29029_);
  and (_29031_, _06526_, _05286_);
  or (_29032_, _29031_, _29030_);
  and (_29033_, _29032_, _04082_);
  and (_29034_, _05286_, \oc8051_golden_model_1.ACC [6]);
  nor (_29035_, _29034_, _29030_);
  nor (_29036_, _29035_, _04437_);
  nor (_29038_, _04436_, _29029_);
  or (_29039_, _29038_, _29036_);
  and (_29040_, _29039_, _04432_);
  nor (_29041_, _13293_, _10876_);
  nor (_29042_, _29041_, _29030_);
  nor (_29043_, _29042_, _04432_);
  or (_29044_, _29043_, _29040_);
  and (_29045_, _29044_, _03470_);
  nor (_29046_, _05924_, _29029_);
  and (_29047_, _13280_, _05924_);
  nor (_29049_, _29047_, _29046_);
  nor (_29050_, _29049_, _03470_);
  or (_29051_, _29050_, _03527_);
  or (_29052_, _29051_, _29045_);
  nor (_29053_, _05417_, _10876_);
  nor (_29054_, _29053_, _29030_);
  nand (_29055_, _29054_, _03527_);
  and (_29056_, _29055_, _29052_);
  and (_29057_, _29056_, _03531_);
  nor (_29058_, _29035_, _03531_);
  or (_29060_, _29058_, _29057_);
  and (_29061_, _29060_, _03466_);
  and (_29062_, _13304_, _05924_);
  nor (_29063_, _29062_, _29046_);
  nor (_29064_, _29063_, _03466_);
  or (_29065_, _29064_, _29061_);
  and (_29066_, _29065_, _03459_);
  nor (_29067_, _29046_, _13311_);
  nor (_29068_, _29067_, _29049_);
  and (_29069_, _29068_, _03458_);
  or (_29071_, _29069_, _29066_);
  and (_29072_, _29071_, _03453_);
  nor (_29073_, _13329_, _10913_);
  nor (_29074_, _29073_, _29046_);
  nor (_29075_, _29074_, _03453_);
  nor (_29076_, _29075_, _07454_);
  not (_29077_, _29076_);
  nor (_29078_, _29077_, _29072_);
  and (_29079_, _29054_, _07454_);
  or (_29080_, _29079_, _04082_);
  nor (_29082_, _29080_, _29078_);
  or (_29083_, _29082_, _29033_);
  and (_29084_, _29083_, _03521_);
  nor (_29085_, _13387_, _10876_);
  nor (_29086_, _29085_, _29030_);
  nor (_29087_, _29086_, _03521_);
  or (_29088_, _29087_, _08905_);
  or (_29089_, _29088_, _29084_);
  and (_29090_, _13402_, _05286_);
  or (_29091_, _29030_, _04527_);
  or (_29093_, _29091_, _29090_);
  and (_29094_, _14949_, _05286_);
  nor (_29095_, _29094_, _29030_);
  and (_29096_, _29095_, _03624_);
  nor (_29097_, _29096_, _03744_);
  and (_29098_, _29097_, _29093_);
  and (_29099_, _29098_, _29089_);
  and (_29100_, _13407_, _05286_);
  nor (_29101_, _29100_, _29030_);
  nor (_29102_, _29101_, _03745_);
  nor (_29104_, _29102_, _29099_);
  nor (_29105_, _29104_, _03611_);
  nor (_29106_, _29030_, _05469_);
  not (_29107_, _29106_);
  nor (_29108_, _29095_, _04523_);
  and (_29109_, _29108_, _29107_);
  nor (_29110_, _29109_, _29105_);
  nor (_29111_, _29110_, _03733_);
  nor (_29112_, _29035_, _03734_);
  and (_29113_, _29112_, _29107_);
  nor (_29115_, _29113_, _03618_);
  not (_29116_, _29115_);
  nor (_29117_, _29116_, _29111_);
  nor (_29118_, _13400_, _10876_);
  or (_29119_, _29030_, _06453_);
  nor (_29120_, _29119_, _29118_);
  or (_29121_, _29120_, _03741_);
  nor (_29122_, _29121_, _29117_);
  nor (_29123_, _13406_, _10876_);
  nor (_29124_, _29123_, _29030_);
  nor (_29126_, _29124_, _06458_);
  or (_29127_, _29126_, _29122_);
  and (_29128_, _29127_, _03948_);
  nor (_29129_, _29042_, _03948_);
  or (_29130_, _29129_, _29128_);
  and (_29131_, _29130_, _03446_);
  nor (_29132_, _29063_, _03446_);
  or (_29133_, _29132_, _29131_);
  and (_29134_, _29133_, _03474_);
  and (_29135_, _13456_, _05286_);
  nor (_29137_, _29135_, _29030_);
  nor (_29138_, _29137_, _03474_);
  or (_29139_, _29138_, _29134_);
  or (_29140_, _29139_, _43193_);
  or (_29141_, _43189_, \oc8051_golden_model_1.TCON [6]);
  and (_29142_, _29141_, _42003_);
  and (_43872_, _29142_, _29140_);
  not (_29143_, \oc8051_golden_model_1.TH0 [0]);
  nor (_29144_, _05339_, _29143_);
  nor (_29145_, _05722_, _10983_);
  nor (_29147_, _29145_, _29144_);
  and (_29148_, _29147_, _17198_);
  and (_29149_, _05339_, \oc8051_golden_model_1.ACC [0]);
  nor (_29150_, _29149_, _29144_);
  nor (_29151_, _29150_, _03531_);
  nor (_29152_, _29151_, _07454_);
  nor (_29153_, _29147_, _04432_);
  nor (_29154_, _04436_, _29143_);
  nor (_29155_, _29150_, _04437_);
  nor (_29156_, _29155_, _29154_);
  nor (_29158_, _29156_, _03534_);
  or (_29159_, _29158_, _03527_);
  nor (_29160_, _29159_, _29153_);
  or (_29161_, _29160_, _03530_);
  and (_29162_, _29161_, _29152_);
  and (_29163_, _05339_, _04429_);
  or (_29164_, _29144_, _26115_);
  nor (_29165_, _29164_, _29163_);
  nor (_29166_, _29165_, _29162_);
  nor (_29167_, _29166_, _04082_);
  and (_29169_, _06617_, _05339_);
  nor (_29170_, _29144_, _04500_);
  not (_29171_, _29170_);
  nor (_29172_, _29171_, _29169_);
  nor (_29173_, _29172_, _29167_);
  nor (_29174_, _29173_, _03224_);
  nor (_29175_, _12164_, _10983_);
  or (_29176_, _29144_, _03521_);
  nor (_29177_, _29176_, _29175_);
  or (_29178_, _29177_, _03624_);
  nor (_29180_, _29178_, _29174_);
  and (_29181_, _05339_, _06350_);
  nor (_29182_, _29181_, _29144_);
  nand (_29183_, _29182_, _04527_);
  and (_29184_, _29183_, _08905_);
  nor (_29185_, _29184_, _29180_);
  and (_29186_, _12177_, _05339_);
  nor (_29187_, _29186_, _29144_);
  and (_29188_, _29187_, _03623_);
  nor (_29189_, _29188_, _29185_);
  nor (_29191_, _29189_, _03744_);
  and (_29192_, _12183_, _05339_);
  or (_29193_, _29144_, _03745_);
  nor (_29194_, _29193_, _29192_);
  or (_29195_, _29194_, _03611_);
  nor (_29196_, _29195_, _29191_);
  or (_29197_, _29182_, _04523_);
  nor (_29198_, _29197_, _29145_);
  nor (_29199_, _29198_, _29196_);
  nor (_29200_, _29199_, _03733_);
  and (_29202_, _12182_, _05339_);
  or (_29203_, _29202_, _29144_);
  and (_29204_, _29203_, _03733_);
  or (_29205_, _29204_, _29200_);
  and (_29206_, _29205_, _06453_);
  nor (_29207_, _12057_, _10983_);
  nor (_29208_, _29207_, _29144_);
  nor (_29209_, _29208_, _06453_);
  or (_29210_, _29209_, _29206_);
  and (_29211_, _29210_, _06458_);
  nor (_29213_, _12181_, _10983_);
  nor (_29214_, _29213_, _29144_);
  nor (_29215_, _29214_, _06458_);
  nor (_29216_, _29215_, _17198_);
  not (_29217_, _29216_);
  nor (_29218_, _29217_, _29211_);
  nor (_29219_, _29218_, _29148_);
  or (_29220_, _29219_, _43193_);
  or (_29221_, _43189_, \oc8051_golden_model_1.TH0 [0]);
  and (_29222_, _29221_, _42003_);
  and (_43875_, _29222_, _29220_);
  and (_29224_, _06572_, _05339_);
  not (_29225_, \oc8051_golden_model_1.TH0 [1]);
  nor (_29226_, _05339_, _29225_);
  nor (_29227_, _29226_, _04500_);
  not (_29228_, _29227_);
  nor (_29229_, _29228_, _29224_);
  not (_29230_, _29229_);
  nor (_29231_, _05339_, \oc8051_golden_model_1.TH0 [1]);
  and (_29232_, _05339_, _03269_);
  nor (_29234_, _29232_, _29231_);
  and (_29235_, _29234_, _03530_);
  and (_29236_, _29234_, _04436_);
  nor (_29237_, _04436_, _29225_);
  or (_29238_, _29237_, _29236_);
  and (_29239_, _29238_, _04432_);
  and (_29240_, _12265_, _05339_);
  nor (_29241_, _29240_, _29231_);
  and (_29242_, _29241_, _03534_);
  or (_29243_, _29242_, _29239_);
  and (_29245_, _29243_, _04457_);
  nor (_29246_, _10983_, _04635_);
  nor (_29247_, _29246_, _29226_);
  nor (_29248_, _29247_, _04457_);
  nor (_29249_, _29248_, _29245_);
  nor (_29250_, _29249_, _03530_);
  or (_29251_, _29250_, _07454_);
  nor (_29252_, _29251_, _29235_);
  and (_29253_, _29247_, _07454_);
  nor (_29254_, _29253_, _29252_);
  nor (_29256_, _29254_, _04082_);
  nor (_29257_, _29256_, _03224_);
  and (_29258_, _29257_, _29230_);
  not (_29259_, _29231_);
  and (_29260_, _12360_, _05339_);
  nor (_29261_, _29260_, _03521_);
  and (_29262_, _29261_, _29259_);
  nor (_29263_, _29262_, _29258_);
  nor (_29264_, _29263_, _08905_);
  nor (_29265_, _12375_, _10983_);
  nor (_29267_, _29265_, _04527_);
  and (_29268_, _05339_, _04325_);
  nor (_29269_, _29268_, _04509_);
  nor (_29270_, _29269_, _29267_);
  nor (_29271_, _29270_, _29231_);
  nor (_29272_, _29271_, _29264_);
  nor (_29273_, _29272_, _03744_);
  nor (_29274_, _12381_, _10983_);
  nor (_29275_, _29274_, _03745_);
  and (_29276_, _29275_, _29259_);
  nor (_29278_, _29276_, _29273_);
  nor (_29279_, _29278_, _03611_);
  nor (_29280_, _12374_, _10983_);
  nor (_29281_, _29280_, _04523_);
  and (_29282_, _29281_, _29259_);
  nor (_29283_, _29282_, _29279_);
  nor (_29284_, _29283_, _03733_);
  nor (_29285_, _29226_, _05674_);
  nor (_29286_, _29285_, _03734_);
  and (_29287_, _29286_, _29234_);
  nor (_29289_, _29287_, _29284_);
  or (_29290_, _29289_, _18526_);
  and (_29291_, _29268_, _05673_);
  nor (_29292_, _29291_, _06453_);
  and (_29293_, _29292_, _29259_);
  nand (_29294_, _29232_, _05673_);
  nor (_29295_, _29231_, _06458_);
  and (_29296_, _29295_, _29294_);
  or (_29297_, _29296_, _03767_);
  nor (_29298_, _29297_, _29293_);
  and (_29300_, _29298_, _29290_);
  nor (_29301_, _29241_, _03948_);
  nor (_29302_, _29301_, _29300_);
  and (_29303_, _29302_, _03474_);
  nor (_29304_, _29240_, _29226_);
  nor (_29305_, _29304_, _03474_);
  or (_29306_, _29305_, _29303_);
  or (_29307_, _29306_, _43193_);
  or (_29308_, _43189_, \oc8051_golden_model_1.TH0 [1]);
  and (_29309_, _29308_, _42003_);
  and (_43876_, _29309_, _29307_);
  not (_29311_, \oc8051_golden_model_1.TH0 [2]);
  nor (_29312_, _05339_, _29311_);
  nor (_29313_, _12587_, _10983_);
  nor (_29314_, _29313_, _29312_);
  nor (_29315_, _29314_, _06458_);
  and (_29316_, _06710_, _05339_);
  nor (_29317_, _29316_, _29312_);
  or (_29318_, _29317_, _04500_);
  and (_29319_, _05339_, \oc8051_golden_model_1.ACC [2]);
  nor (_29321_, _29319_, _29312_);
  nor (_29322_, _29321_, _04437_);
  nor (_29323_, _04436_, _29311_);
  or (_29324_, _29323_, _29322_);
  and (_29325_, _29324_, _04432_);
  nor (_29326_, _12467_, _10983_);
  nor (_29327_, _29326_, _29312_);
  nor (_29328_, _29327_, _04432_);
  or (_29329_, _29328_, _29325_);
  and (_29330_, _29329_, _04457_);
  nor (_29332_, _10983_, _05073_);
  nor (_29333_, _29332_, _29312_);
  nor (_29334_, _29333_, _04457_);
  nor (_29335_, _29334_, _29330_);
  nor (_29336_, _29335_, _03530_);
  nor (_29337_, _29321_, _03531_);
  nor (_29338_, _29337_, _07454_);
  not (_29339_, _29338_);
  nor (_29340_, _29339_, _29336_);
  and (_29341_, _29333_, _07454_);
  or (_29343_, _29341_, _04082_);
  or (_29344_, _29343_, _29340_);
  and (_29345_, _29344_, _03521_);
  and (_29346_, _29345_, _29318_);
  nor (_29347_, _12568_, _10983_);
  or (_29348_, _29312_, _03521_);
  nor (_29349_, _29348_, _29347_);
  or (_29350_, _29349_, _03624_);
  nor (_29351_, _29350_, _29346_);
  and (_29352_, _05339_, _06399_);
  nor (_29354_, _29352_, _29312_);
  nand (_29355_, _29354_, _04527_);
  and (_29356_, _29355_, _08905_);
  nor (_29357_, _29356_, _29351_);
  and (_29358_, _12582_, _05339_);
  nor (_29359_, _29358_, _29312_);
  and (_29360_, _29359_, _03623_);
  nor (_29361_, _29360_, _29357_);
  nor (_29362_, _29361_, _03744_);
  and (_29363_, _12588_, _05339_);
  or (_29365_, _29312_, _03745_);
  nor (_29366_, _29365_, _29363_);
  or (_29367_, _29366_, _03611_);
  nor (_29368_, _29367_, _29362_);
  nor (_29369_, _29312_, _05772_);
  not (_29370_, _29369_);
  nor (_29371_, _29354_, _04523_);
  and (_29372_, _29371_, _29370_);
  nor (_29373_, _29372_, _29368_);
  nor (_29374_, _29373_, _03733_);
  nor (_29376_, _29321_, _03734_);
  and (_29377_, _29376_, _29370_);
  or (_29378_, _29377_, _29374_);
  and (_29379_, _29378_, _06453_);
  nor (_29380_, _12581_, _10983_);
  nor (_29381_, _29380_, _29312_);
  nor (_29382_, _29381_, _06453_);
  or (_29383_, _29382_, _29379_);
  and (_29384_, _29383_, _06458_);
  nor (_29385_, _29384_, _29315_);
  nor (_29387_, _29385_, _03767_);
  nor (_29388_, _29327_, _03948_);
  or (_29389_, _29388_, _03473_);
  nor (_29390_, _29389_, _29387_);
  and (_29391_, _12638_, _05339_);
  or (_29392_, _29312_, _03474_);
  nor (_29393_, _29392_, _29391_);
  nor (_29394_, _29393_, _29390_);
  or (_29395_, _29394_, _43193_);
  or (_29396_, _43189_, \oc8051_golden_model_1.TH0 [2]);
  and (_29398_, _29396_, _42003_);
  and (_43877_, _29398_, _29395_);
  not (_29399_, \oc8051_golden_model_1.TH0 [3]);
  nor (_29400_, _05339_, _29399_);
  nor (_29401_, _12792_, _10983_);
  nor (_29402_, _29401_, _29400_);
  nor (_29403_, _29402_, _06458_);
  and (_29404_, _12793_, _05339_);
  nor (_29405_, _29404_, _29400_);
  nor (_29406_, _29405_, _03745_);
  and (_29408_, _06664_, _05339_);
  or (_29409_, _29408_, _29400_);
  and (_29410_, _29409_, _04082_);
  and (_29411_, _05339_, \oc8051_golden_model_1.ACC [3]);
  nor (_29412_, _29411_, _29400_);
  nor (_29413_, _29412_, _03531_);
  nor (_29414_, _29412_, _04437_);
  nor (_29415_, _04436_, _29399_);
  or (_29416_, _29415_, _29414_);
  and (_29417_, _29416_, _04432_);
  nor (_29419_, _12652_, _10983_);
  nor (_29420_, _29419_, _29400_);
  nor (_29421_, _29420_, _04432_);
  or (_29422_, _29421_, _29417_);
  and (_29423_, _29422_, _04457_);
  nor (_29424_, _10983_, _04885_);
  nor (_29425_, _29424_, _29400_);
  nor (_29426_, _29425_, _04457_);
  nor (_29427_, _29426_, _29423_);
  nor (_29428_, _29427_, _03530_);
  or (_29430_, _29428_, _07454_);
  nor (_29431_, _29430_, _29413_);
  and (_29432_, _29425_, _07454_);
  or (_29433_, _29432_, _04082_);
  nor (_29434_, _29433_, _29431_);
  or (_29435_, _29434_, _29410_);
  and (_29436_, _29435_, _03521_);
  nor (_29437_, _12773_, _10983_);
  nor (_29438_, _29437_, _29400_);
  nor (_29439_, _29438_, _03521_);
  or (_29440_, _29439_, _08905_);
  or (_29441_, _29440_, _29436_);
  and (_29442_, _12787_, _05339_);
  or (_29443_, _29400_, _04527_);
  or (_29444_, _29443_, _29442_);
  and (_29445_, _05339_, _06356_);
  nor (_29446_, _29445_, _29400_);
  and (_29447_, _29446_, _03624_);
  nor (_29448_, _29447_, _03744_);
  and (_29449_, _29448_, _29444_);
  and (_29451_, _29449_, _29441_);
  nor (_29452_, _29451_, _29406_);
  nor (_29453_, _29452_, _03611_);
  nor (_29454_, _29400_, _05625_);
  not (_29455_, _29454_);
  nor (_29456_, _29446_, _04523_);
  and (_29457_, _29456_, _29455_);
  nor (_29458_, _29457_, _29453_);
  nor (_29459_, _29458_, _03733_);
  nor (_29460_, _29412_, _03734_);
  and (_29462_, _29460_, _29455_);
  nor (_29463_, _29462_, _03618_);
  not (_29464_, _29463_);
  nor (_29465_, _29464_, _29459_);
  nor (_29466_, _12786_, _10983_);
  or (_29467_, _29400_, _06453_);
  nor (_29468_, _29467_, _29466_);
  or (_29469_, _29468_, _03741_);
  nor (_29470_, _29469_, _29465_);
  nor (_29471_, _29470_, _29403_);
  nor (_29473_, _29471_, _03767_);
  nor (_29474_, _29420_, _03948_);
  or (_29475_, _29474_, _03473_);
  nor (_29476_, _29475_, _29473_);
  and (_29477_, _12843_, _05339_);
  or (_29478_, _29400_, _03474_);
  nor (_29479_, _29478_, _29477_);
  nor (_29480_, _29479_, _29476_);
  or (_29481_, _29480_, _43193_);
  or (_29482_, _43189_, \oc8051_golden_model_1.TH0 [3]);
  and (_29484_, _29482_, _42003_);
  and (_43878_, _29484_, _29481_);
  not (_29485_, \oc8051_golden_model_1.TH0 [4]);
  nor (_29486_, _05339_, _29485_);
  nor (_29487_, _12991_, _10983_);
  nor (_29488_, _29487_, _29486_);
  nor (_29489_, _29488_, _06458_);
  and (_29490_, _12992_, _05339_);
  nor (_29491_, _29490_, _29486_);
  nor (_29492_, _29491_, _03745_);
  and (_29494_, _06337_, _05339_);
  nor (_29495_, _29494_, _29486_);
  and (_29496_, _29495_, _03624_);
  and (_29497_, _05339_, \oc8051_golden_model_1.ACC [4]);
  nor (_29498_, _29497_, _29486_);
  nor (_29499_, _29498_, _03531_);
  nor (_29500_, _29498_, _04437_);
  nor (_29501_, _04436_, _29485_);
  or (_29502_, _29501_, _29500_);
  and (_29503_, _29502_, _04432_);
  nor (_29504_, _12856_, _10983_);
  nor (_29505_, _29504_, _29486_);
  nor (_29506_, _29505_, _04432_);
  or (_29507_, _29506_, _29503_);
  and (_29508_, _29507_, _04457_);
  nor (_29509_, _05831_, _10983_);
  nor (_29510_, _29509_, _29486_);
  nor (_29511_, _29510_, _04457_);
  nor (_29512_, _29511_, _29508_);
  nor (_29513_, _29512_, _03530_);
  or (_29516_, _29513_, _07454_);
  nor (_29517_, _29516_, _29499_);
  and (_29518_, _29510_, _07454_);
  nor (_29519_, _29518_, _29517_);
  nor (_29520_, _29519_, _04082_);
  and (_29521_, _06802_, _05339_);
  nor (_29522_, _29486_, _04500_);
  not (_29523_, _29522_);
  nor (_29524_, _29523_, _29521_);
  or (_29525_, _29524_, _03224_);
  nor (_29527_, _29525_, _29520_);
  nor (_29528_, _12972_, _10983_);
  nor (_29529_, _29528_, _29486_);
  nor (_29530_, _29529_, _03521_);
  or (_29531_, _29530_, _03624_);
  nor (_29532_, _29531_, _29527_);
  nor (_29533_, _29532_, _29496_);
  or (_29534_, _29533_, _03623_);
  and (_29535_, _12986_, _05339_);
  or (_29536_, _29535_, _29486_);
  or (_29538_, _29536_, _04527_);
  and (_29539_, _29538_, _03745_);
  and (_29540_, _29539_, _29534_);
  nor (_29541_, _29540_, _29492_);
  nor (_29542_, _29541_, _03611_);
  nor (_29543_, _29486_, _05880_);
  not (_29544_, _29543_);
  nor (_29545_, _29495_, _04523_);
  and (_29546_, _29545_, _29544_);
  nor (_29547_, _29546_, _29542_);
  nor (_29549_, _29547_, _03733_);
  nor (_29550_, _29498_, _03734_);
  and (_29551_, _29550_, _29544_);
  nor (_29552_, _29551_, _03618_);
  not (_29553_, _29552_);
  nor (_29554_, _29553_, _29549_);
  nor (_29555_, _12985_, _10983_);
  or (_29556_, _29486_, _06453_);
  nor (_29557_, _29556_, _29555_);
  or (_29558_, _29557_, _03741_);
  nor (_29560_, _29558_, _29554_);
  nor (_29561_, _29560_, _29489_);
  nor (_29562_, _29561_, _03767_);
  nor (_29563_, _29505_, _03948_);
  or (_29564_, _29563_, _03473_);
  nor (_29565_, _29564_, _29562_);
  and (_29566_, _13051_, _05339_);
  or (_29567_, _29486_, _03474_);
  nor (_29568_, _29567_, _29566_);
  nor (_29569_, _29568_, _29565_);
  or (_29571_, _29569_, _43193_);
  or (_29572_, _43189_, \oc8051_golden_model_1.TH0 [4]);
  and (_29573_, _29572_, _42003_);
  and (_43879_, _29573_, _29571_);
  not (_29574_, \oc8051_golden_model_1.TH0 [5]);
  nor (_29575_, _05339_, _29574_);
  nor (_29576_, _13203_, _10983_);
  nor (_29577_, _29576_, _29575_);
  nor (_29578_, _29577_, _06458_);
  and (_29579_, _13204_, _05339_);
  nor (_29581_, _29579_, _29575_);
  nor (_29582_, _29581_, _03745_);
  and (_29583_, _06757_, _05339_);
  or (_29584_, _29583_, _29575_);
  and (_29585_, _29584_, _04082_);
  and (_29586_, _05339_, \oc8051_golden_model_1.ACC [5]);
  nor (_29587_, _29586_, _29575_);
  nor (_29588_, _29587_, _03531_);
  nor (_29589_, _29587_, _04437_);
  nor (_29590_, _04436_, _29574_);
  or (_29592_, _29590_, _29589_);
  and (_29593_, _29592_, _04432_);
  nor (_29594_, _13070_, _10983_);
  nor (_29595_, _29594_, _29575_);
  nor (_29596_, _29595_, _04432_);
  or (_29597_, _29596_, _29593_);
  and (_29598_, _29597_, _04457_);
  nor (_29599_, _05526_, _10983_);
  nor (_29600_, _29599_, _29575_);
  nor (_29601_, _29600_, _04457_);
  nor (_29603_, _29601_, _29598_);
  nor (_29604_, _29603_, _03530_);
  or (_29605_, _29604_, _07454_);
  nor (_29606_, _29605_, _29588_);
  and (_29607_, _29600_, _07454_);
  or (_29608_, _29607_, _04082_);
  nor (_29609_, _29608_, _29606_);
  or (_29610_, _29609_, _29585_);
  and (_29611_, _29610_, _03521_);
  nor (_29612_, _13184_, _10983_);
  nor (_29614_, _29612_, _29575_);
  nor (_29615_, _29614_, _03521_);
  or (_29616_, _29615_, _08905_);
  or (_29617_, _29616_, _29611_);
  and (_29618_, _13198_, _05339_);
  or (_29619_, _29575_, _04527_);
  or (_29620_, _29619_, _29618_);
  and (_29621_, _06295_, _05339_);
  nor (_29622_, _29621_, _29575_);
  and (_29623_, _29622_, _03624_);
  nor (_29625_, _29623_, _03744_);
  and (_29626_, _29625_, _29620_);
  and (_29627_, _29626_, _29617_);
  nor (_29628_, _29627_, _29582_);
  nor (_29629_, _29628_, _03611_);
  nor (_29630_, _29575_, _05576_);
  not (_29631_, _29630_);
  nor (_29632_, _29622_, _04523_);
  and (_29633_, _29632_, _29631_);
  nor (_29634_, _29633_, _29629_);
  nor (_29636_, _29634_, _03733_);
  nor (_29637_, _29587_, _03734_);
  and (_29638_, _29637_, _29631_);
  or (_29639_, _29638_, _29636_);
  and (_29640_, _29639_, _06453_);
  nor (_29641_, _13197_, _10983_);
  nor (_29642_, _29641_, _29575_);
  nor (_29643_, _29642_, _06453_);
  or (_29644_, _29643_, _29640_);
  and (_29645_, _29644_, _06458_);
  nor (_29647_, _29645_, _29578_);
  nor (_29648_, _29647_, _03767_);
  nor (_29649_, _29595_, _03948_);
  or (_29650_, _29649_, _03473_);
  nor (_29651_, _29650_, _29648_);
  and (_29652_, _13253_, _05339_);
  or (_29653_, _29575_, _03474_);
  nor (_29654_, _29653_, _29652_);
  nor (_29655_, _29654_, _29651_);
  or (_29656_, _29655_, _43193_);
  or (_29658_, _43189_, \oc8051_golden_model_1.TH0 [5]);
  and (_29659_, _29658_, _42003_);
  and (_43880_, _29659_, _29656_);
  not (_29660_, \oc8051_golden_model_1.TH0 [6]);
  nor (_29661_, _05339_, _29660_);
  nor (_29662_, _13406_, _10983_);
  nor (_29663_, _29662_, _29661_);
  nor (_29664_, _29663_, _06458_);
  and (_29665_, _13407_, _05339_);
  nor (_29666_, _29665_, _29661_);
  nor (_29668_, _29666_, _03745_);
  and (_29669_, _06526_, _05339_);
  or (_29670_, _29669_, _29661_);
  and (_29671_, _29670_, _04082_);
  and (_29672_, _05339_, \oc8051_golden_model_1.ACC [6]);
  nor (_29673_, _29672_, _29661_);
  nor (_29674_, _29673_, _04437_);
  nor (_29675_, _04436_, _29660_);
  or (_29676_, _29675_, _29674_);
  and (_29677_, _29676_, _04432_);
  nor (_29679_, _13293_, _10983_);
  nor (_29680_, _29679_, _29661_);
  nor (_29681_, _29680_, _04432_);
  or (_29682_, _29681_, _29677_);
  and (_29683_, _29682_, _04457_);
  nor (_29684_, _05417_, _10983_);
  nor (_29685_, _29684_, _29661_);
  nor (_29686_, _29685_, _04457_);
  nor (_29687_, _29686_, _29683_);
  nor (_29688_, _29687_, _03530_);
  nor (_29690_, _29673_, _03531_);
  nor (_29691_, _29690_, _07454_);
  not (_29692_, _29691_);
  nor (_29693_, _29692_, _29688_);
  and (_29694_, _29685_, _07454_);
  or (_29695_, _29694_, _04082_);
  nor (_29696_, _29695_, _29693_);
  or (_29697_, _29696_, _29671_);
  and (_29698_, _29697_, _03521_);
  nor (_29699_, _13387_, _10983_);
  nor (_29701_, _29699_, _29661_);
  nor (_29702_, _29701_, _03521_);
  or (_29703_, _29702_, _08905_);
  or (_29704_, _29703_, _29698_);
  and (_29705_, _13402_, _05339_);
  or (_29706_, _29661_, _04527_);
  or (_29707_, _29706_, _29705_);
  and (_29708_, _14949_, _05339_);
  nor (_29709_, _29708_, _29661_);
  and (_29710_, _29709_, _03624_);
  nor (_29712_, _29710_, _03744_);
  and (_29713_, _29712_, _29707_);
  and (_29714_, _29713_, _29704_);
  nor (_29715_, _29714_, _29668_);
  nor (_29716_, _29715_, _03611_);
  nor (_29717_, _29661_, _05469_);
  not (_29718_, _29717_);
  nor (_29719_, _29709_, _04523_);
  and (_29720_, _29719_, _29718_);
  nor (_29721_, _29720_, _29716_);
  nor (_29723_, _29721_, _03733_);
  nor (_29724_, _29673_, _03734_);
  and (_29725_, _29724_, _29718_);
  nor (_29726_, _29725_, _03618_);
  not (_29727_, _29726_);
  nor (_29728_, _29727_, _29723_);
  nor (_29729_, _13400_, _10983_);
  or (_29730_, _29661_, _06453_);
  nor (_29731_, _29730_, _29729_);
  or (_29732_, _29731_, _03741_);
  nor (_29734_, _29732_, _29728_);
  nor (_29735_, _29734_, _29664_);
  nor (_29736_, _29735_, _03767_);
  nor (_29737_, _29680_, _03948_);
  or (_29738_, _29737_, _03473_);
  nor (_29739_, _29738_, _29736_);
  and (_29740_, _13456_, _05339_);
  or (_29741_, _29661_, _03474_);
  nor (_29742_, _29741_, _29740_);
  nor (_29743_, _29742_, _29739_);
  or (_29745_, _29743_, _43193_);
  or (_29746_, _43189_, \oc8051_golden_model_1.TH0 [6]);
  and (_29747_, _29746_, _42003_);
  and (_43881_, _29747_, _29745_);
  not (_29748_, \oc8051_golden_model_1.TH1 [0]);
  nor (_29749_, _05342_, _29748_);
  nor (_29750_, _05722_, _11066_);
  nor (_29751_, _29750_, _29749_);
  and (_29752_, _29751_, _17198_);
  and (_29753_, _05342_, \oc8051_golden_model_1.ACC [0]);
  nor (_29755_, _29753_, _29749_);
  nor (_29756_, _29755_, _03531_);
  nor (_29757_, _29755_, _04437_);
  nor (_29758_, _04436_, _29748_);
  or (_29759_, _29758_, _29757_);
  and (_29760_, _29759_, _04432_);
  nor (_29761_, _29751_, _04432_);
  or (_29762_, _29761_, _29760_);
  and (_29763_, _29762_, _04457_);
  and (_29764_, _05342_, _04429_);
  nor (_29765_, _29764_, _29749_);
  nor (_29766_, _29765_, _04457_);
  nor (_29767_, _29766_, _29763_);
  nor (_29768_, _29767_, _03530_);
  or (_29769_, _29768_, _07454_);
  nor (_29770_, _29769_, _29756_);
  and (_29771_, _29765_, _07454_);
  nor (_29772_, _29771_, _29770_);
  nor (_29773_, _29772_, _04082_);
  and (_29774_, _06617_, _05342_);
  nor (_29777_, _29749_, _04500_);
  not (_29778_, _29777_);
  nor (_29779_, _29778_, _29774_);
  nor (_29780_, _29779_, _29773_);
  nor (_29781_, _29780_, _03224_);
  nor (_29782_, _12164_, _11066_);
  or (_29783_, _29749_, _03521_);
  nor (_29784_, _29783_, _29782_);
  or (_29785_, _29784_, _03624_);
  nor (_29786_, _29785_, _29781_);
  and (_29788_, _05342_, _06350_);
  nor (_29789_, _29788_, _29749_);
  nand (_29790_, _29789_, _04527_);
  and (_29791_, _29790_, _08905_);
  nor (_29792_, _29791_, _29786_);
  and (_29793_, _12177_, _05342_);
  nor (_29794_, _29793_, _29749_);
  and (_29795_, _29794_, _03623_);
  nor (_29796_, _29795_, _29792_);
  nor (_29797_, _29796_, _03744_);
  and (_29799_, _12183_, _05342_);
  or (_29800_, _29749_, _03745_);
  nor (_29801_, _29800_, _29799_);
  or (_29802_, _29801_, _03611_);
  nor (_29803_, _29802_, _29797_);
  or (_29804_, _29789_, _04523_);
  nor (_29805_, _29804_, _29750_);
  nor (_29806_, _29805_, _29803_);
  nor (_29807_, _29806_, _03733_);
  nor (_29808_, _29749_, _05722_);
  or (_29810_, _29808_, _03734_);
  nor (_29811_, _29810_, _29755_);
  or (_29812_, _29811_, _29807_);
  and (_29813_, _29812_, _06453_);
  nor (_29814_, _12057_, _11066_);
  nor (_29815_, _29814_, _29749_);
  nor (_29816_, _29815_, _06453_);
  or (_29817_, _29816_, _29813_);
  and (_29818_, _29817_, _06458_);
  nor (_29819_, _12181_, _11066_);
  nor (_29821_, _29819_, _29749_);
  nor (_29822_, _29821_, _06458_);
  nor (_29823_, _29822_, _17198_);
  not (_29824_, _29823_);
  nor (_29825_, _29824_, _29818_);
  nor (_29826_, _29825_, _29752_);
  or (_29827_, _29826_, _43193_);
  or (_29828_, _43189_, \oc8051_golden_model_1.TH1 [0]);
  and (_29829_, _29828_, _42003_);
  and (_43884_, _29829_, _29827_);
  and (_29831_, _06572_, _05342_);
  not (_29832_, \oc8051_golden_model_1.TH1 [1]);
  nor (_29833_, _05342_, _29832_);
  nor (_29834_, _29833_, _04500_);
  not (_29835_, _29834_);
  nor (_29836_, _29835_, _29831_);
  not (_29837_, _29836_);
  nor (_29838_, _11066_, _04635_);
  nor (_29839_, _29838_, _29833_);
  and (_29840_, _29839_, _07454_);
  nor (_29842_, _05342_, \oc8051_golden_model_1.TH1 [1]);
  and (_29843_, _05342_, _03269_);
  nor (_29844_, _29843_, _29842_);
  and (_29845_, _29844_, _04436_);
  nor (_29846_, _04436_, _29832_);
  or (_29847_, _29846_, _29845_);
  and (_29848_, _29847_, _04432_);
  and (_29849_, _12265_, _05342_);
  nor (_29850_, _29849_, _29842_);
  and (_29851_, _29850_, _03534_);
  or (_29853_, _29851_, _29848_);
  and (_29854_, _29853_, _04457_);
  nor (_29855_, _29839_, _04457_);
  nor (_29856_, _29855_, _29854_);
  nor (_29857_, _29856_, _03530_);
  and (_29858_, _29844_, _03530_);
  nor (_29859_, _29858_, _07454_);
  not (_29860_, _29859_);
  nor (_29861_, _29860_, _29857_);
  nor (_29862_, _29861_, _29840_);
  nor (_29864_, _29862_, _04082_);
  nor (_29865_, _29864_, _03224_);
  and (_29866_, _29865_, _29837_);
  not (_29867_, _29842_);
  and (_29868_, _12360_, _05342_);
  nor (_29869_, _29868_, _03521_);
  and (_29870_, _29869_, _29867_);
  nor (_29871_, _29870_, _29866_);
  nor (_29872_, _29871_, _08905_);
  nor (_29873_, _12375_, _11066_);
  nor (_29875_, _29873_, _04527_);
  and (_29876_, _05342_, _04325_);
  nor (_29877_, _29876_, _04509_);
  or (_29878_, _29877_, _29875_);
  and (_29879_, _29878_, _29867_);
  nor (_29880_, _29879_, _29872_);
  nor (_29881_, _29880_, _03744_);
  nor (_29882_, _12381_, _11066_);
  nor (_29883_, _29882_, _03745_);
  and (_29884_, _29883_, _29867_);
  nor (_29886_, _29884_, _29881_);
  nor (_29887_, _29886_, _03611_);
  nor (_29888_, _12374_, _11066_);
  nor (_29889_, _29888_, _04523_);
  and (_29890_, _29889_, _29867_);
  nor (_29891_, _29890_, _29887_);
  nor (_29892_, _29891_, _03733_);
  nor (_29893_, _29833_, _05674_);
  nor (_29894_, _29893_, _03734_);
  and (_29895_, _29894_, _29844_);
  nor (_29897_, _29895_, _29892_);
  or (_29898_, _29897_, _18526_);
  nand (_29899_, _12380_, _05342_);
  and (_29900_, _29899_, _03741_);
  and (_29901_, _29900_, _29867_);
  nor (_29902_, _29901_, _03767_);
  and (_29903_, _29876_, _05673_);
  or (_29904_, _29842_, _06453_);
  or (_29905_, _29904_, _29903_);
  and (_29906_, _29905_, _29902_);
  and (_29908_, _29906_, _29898_);
  nor (_29909_, _29850_, _03948_);
  nor (_29910_, _29909_, _29908_);
  and (_29911_, _29910_, _03474_);
  nor (_29912_, _29849_, _29833_);
  nor (_29913_, _29912_, _03474_);
  or (_29914_, _29913_, _29911_);
  or (_29915_, _29914_, _43193_);
  or (_29916_, _43189_, \oc8051_golden_model_1.TH1 [1]);
  and (_29917_, _29916_, _42003_);
  and (_43885_, _29917_, _29915_);
  not (_29919_, \oc8051_golden_model_1.TH1 [2]);
  nor (_29920_, _05342_, _29919_);
  nor (_29921_, _12587_, _11066_);
  nor (_29922_, _29921_, _29920_);
  nor (_29923_, _29922_, _06458_);
  and (_29924_, _12588_, _05342_);
  nor (_29925_, _29924_, _29920_);
  nor (_29926_, _29925_, _03745_);
  nor (_29927_, _11066_, _05073_);
  nor (_29929_, _29927_, _29920_);
  and (_29930_, _29929_, _07454_);
  and (_29931_, _05342_, \oc8051_golden_model_1.ACC [2]);
  nor (_29932_, _29931_, _29920_);
  nor (_29933_, _29932_, _03531_);
  nor (_29934_, _29932_, _04437_);
  nor (_29935_, _04436_, _29919_);
  or (_29936_, _29935_, _29934_);
  and (_29937_, _29936_, _04432_);
  nor (_29938_, _12467_, _11066_);
  nor (_29940_, _29938_, _29920_);
  nor (_29941_, _29940_, _04432_);
  or (_29942_, _29941_, _29937_);
  and (_29943_, _29942_, _04457_);
  nor (_29944_, _29929_, _04457_);
  nor (_29945_, _29944_, _29943_);
  nor (_29946_, _29945_, _03530_);
  or (_29947_, _29946_, _07454_);
  nor (_29948_, _29947_, _29933_);
  nor (_29949_, _29948_, _29930_);
  nor (_29951_, _29949_, _04082_);
  and (_29952_, _06710_, _05342_);
  nor (_29953_, _29920_, _04500_);
  not (_29954_, _29953_);
  nor (_29955_, _29954_, _29952_);
  nor (_29956_, _29955_, _03224_);
  not (_29957_, _29956_);
  nor (_29958_, _29957_, _29951_);
  nor (_29959_, _12568_, _11066_);
  nor (_29960_, _29959_, _29920_);
  nor (_29962_, _29960_, _03521_);
  or (_29963_, _29962_, _08905_);
  or (_29964_, _29963_, _29958_);
  and (_29965_, _12582_, _05342_);
  or (_29966_, _29920_, _04527_);
  or (_29967_, _29966_, _29965_);
  and (_29968_, _05342_, _06399_);
  nor (_29969_, _29968_, _29920_);
  and (_29970_, _29969_, _03624_);
  nor (_29971_, _29970_, _03744_);
  and (_29973_, _29971_, _29967_);
  and (_29974_, _29973_, _29964_);
  nor (_29975_, _29974_, _29926_);
  nor (_29976_, _29975_, _03611_);
  nor (_29977_, _29920_, _05772_);
  not (_29978_, _29977_);
  nor (_29979_, _29969_, _04523_);
  and (_29980_, _29979_, _29978_);
  nor (_29981_, _29980_, _29976_);
  nor (_29982_, _29981_, _03733_);
  nor (_29984_, _29932_, _03734_);
  and (_29985_, _29984_, _29978_);
  or (_29986_, _29985_, _29982_);
  and (_29987_, _29986_, _06453_);
  nor (_29988_, _12581_, _11066_);
  nor (_29989_, _29988_, _29920_);
  nor (_29990_, _29989_, _06453_);
  or (_29991_, _29990_, _29987_);
  and (_29992_, _29991_, _06458_);
  nor (_29993_, _29992_, _29923_);
  nor (_29995_, _29993_, _03767_);
  nor (_29996_, _29940_, _03948_);
  or (_29997_, _29996_, _03473_);
  nor (_29998_, _29997_, _29995_);
  and (_29999_, _12638_, _05342_);
  or (_30000_, _29920_, _03474_);
  nor (_30001_, _30000_, _29999_);
  nor (_30002_, _30001_, _29998_);
  or (_30003_, _30002_, _43193_);
  or (_30004_, _43189_, \oc8051_golden_model_1.TH1 [2]);
  and (_30006_, _30004_, _42003_);
  and (_43886_, _30006_, _30003_);
  not (_30007_, \oc8051_golden_model_1.TH1 [3]);
  nor (_30008_, _05342_, _30007_);
  nor (_30009_, _12792_, _11066_);
  nor (_30010_, _30009_, _30008_);
  nor (_30011_, _30010_, _06458_);
  and (_30012_, _12793_, _05342_);
  nor (_30013_, _30012_, _30008_);
  nor (_30014_, _30013_, _03745_);
  and (_30016_, _06664_, _05342_);
  or (_30017_, _30016_, _30008_);
  and (_30018_, _30017_, _04082_);
  and (_30019_, _05342_, \oc8051_golden_model_1.ACC [3]);
  nor (_30020_, _30019_, _30008_);
  nor (_30021_, _30020_, _04437_);
  nor (_30022_, _04436_, _30007_);
  or (_30023_, _30022_, _30021_);
  and (_30024_, _30023_, _04432_);
  nor (_30025_, _12652_, _11066_);
  nor (_30027_, _30025_, _30008_);
  nor (_30028_, _30027_, _04432_);
  or (_30029_, _30028_, _30024_);
  and (_30030_, _30029_, _04457_);
  nor (_30031_, _11066_, _04885_);
  nor (_30032_, _30031_, _30008_);
  nor (_30033_, _30032_, _04457_);
  nor (_30034_, _30033_, _30030_);
  nor (_30035_, _30034_, _03530_);
  nor (_30036_, _30020_, _03531_);
  nor (_30038_, _30036_, _07454_);
  not (_30039_, _30038_);
  nor (_30040_, _30039_, _30035_);
  and (_30041_, _30032_, _07454_);
  or (_30042_, _30041_, _04082_);
  nor (_30043_, _30042_, _30040_);
  or (_30044_, _30043_, _30018_);
  and (_30045_, _30044_, _03521_);
  nor (_30046_, _12773_, _11066_);
  nor (_30047_, _30046_, _30008_);
  nor (_30049_, _30047_, _03521_);
  or (_30050_, _30049_, _08905_);
  or (_30051_, _30050_, _30045_);
  and (_30052_, _12787_, _05342_);
  or (_30053_, _30008_, _04527_);
  or (_30054_, _30053_, _30052_);
  and (_30055_, _05342_, _06356_);
  nor (_30056_, _30055_, _30008_);
  and (_30057_, _30056_, _03624_);
  nor (_30058_, _30057_, _03744_);
  and (_30060_, _30058_, _30054_);
  and (_30061_, _30060_, _30051_);
  nor (_30062_, _30061_, _30014_);
  nor (_30063_, _30062_, _03611_);
  nor (_30064_, _30008_, _05625_);
  not (_30065_, _30064_);
  nor (_30066_, _30056_, _04523_);
  and (_30067_, _30066_, _30065_);
  nor (_30068_, _30067_, _30063_);
  nor (_30069_, _30068_, _03733_);
  nor (_30070_, _30020_, _03734_);
  and (_30071_, _30070_, _30065_);
  or (_30072_, _30071_, _30069_);
  and (_30073_, _30072_, _06453_);
  nor (_30074_, _12786_, _11066_);
  nor (_30075_, _30074_, _30008_);
  nor (_30076_, _30075_, _06453_);
  or (_30077_, _30076_, _30073_);
  and (_30078_, _30077_, _06458_);
  nor (_30079_, _30078_, _30011_);
  nor (_30082_, _30079_, _03767_);
  nor (_30083_, _30027_, _03948_);
  or (_30084_, _30083_, _03473_);
  nor (_30085_, _30084_, _30082_);
  and (_30086_, _12843_, _05342_);
  or (_30087_, _30008_, _03474_);
  nor (_30088_, _30087_, _30086_);
  nor (_30089_, _30088_, _30085_);
  or (_30090_, _30089_, _43193_);
  or (_30091_, _43189_, \oc8051_golden_model_1.TH1 [3]);
  and (_30093_, _30091_, _42003_);
  and (_43887_, _30093_, _30090_);
  not (_30094_, \oc8051_golden_model_1.TH1 [4]);
  nor (_30095_, _05342_, _30094_);
  nor (_30096_, _12991_, _11066_);
  nor (_30097_, _30096_, _30095_);
  nor (_30098_, _30097_, _06458_);
  and (_30099_, _12992_, _05342_);
  nor (_30100_, _30099_, _30095_);
  nor (_30101_, _30100_, _03745_);
  and (_30103_, _06337_, _05342_);
  nor (_30104_, _30103_, _30095_);
  and (_30105_, _30104_, _03624_);
  nor (_30106_, _05831_, _11066_);
  nor (_30107_, _30106_, _30095_);
  and (_30108_, _30107_, _07454_);
  and (_30109_, _05342_, \oc8051_golden_model_1.ACC [4]);
  nor (_30110_, _30109_, _30095_);
  nor (_30111_, _30110_, _03531_);
  nor (_30112_, _30110_, _04437_);
  nor (_30114_, _04436_, _30094_);
  or (_30115_, _30114_, _30112_);
  and (_30116_, _30115_, _04432_);
  nor (_30117_, _12856_, _11066_);
  nor (_30118_, _30117_, _30095_);
  nor (_30119_, _30118_, _04432_);
  or (_30120_, _30119_, _30116_);
  and (_30121_, _30120_, _04457_);
  nor (_30122_, _30107_, _04457_);
  nor (_30123_, _30122_, _30121_);
  nor (_30125_, _30123_, _03530_);
  or (_30126_, _30125_, _07454_);
  nor (_30127_, _30126_, _30111_);
  nor (_30128_, _30127_, _30108_);
  nor (_30129_, _30128_, _04082_);
  and (_30130_, _06802_, _05342_);
  nor (_30131_, _30095_, _04500_);
  not (_30132_, _30131_);
  nor (_30133_, _30132_, _30130_);
  or (_30134_, _30133_, _03224_);
  nor (_30136_, _30134_, _30129_);
  nor (_30137_, _12972_, _11066_);
  nor (_30138_, _30137_, _30095_);
  nor (_30139_, _30138_, _03521_);
  or (_30140_, _30139_, _03624_);
  nor (_30141_, _30140_, _30136_);
  nor (_30142_, _30141_, _30105_);
  or (_30143_, _30142_, _03623_);
  and (_30144_, _12986_, _05342_);
  or (_30145_, _30144_, _30095_);
  or (_30147_, _30145_, _04527_);
  and (_30148_, _30147_, _03745_);
  and (_30149_, _30148_, _30143_);
  nor (_30150_, _30149_, _30101_);
  nor (_30151_, _30150_, _03611_);
  nor (_30152_, _30095_, _05880_);
  not (_30153_, _30152_);
  nor (_30154_, _30104_, _04523_);
  and (_30155_, _30154_, _30153_);
  nor (_30156_, _30155_, _30151_);
  nor (_30157_, _30156_, _03733_);
  nor (_30158_, _30110_, _03734_);
  and (_30159_, _30158_, _30153_);
  nor (_30160_, _30159_, _03618_);
  not (_30161_, _30160_);
  nor (_30162_, _30161_, _30157_);
  nor (_30163_, _12985_, _11066_);
  or (_30164_, _30095_, _06453_);
  nor (_30165_, _30164_, _30163_);
  or (_30166_, _30165_, _03741_);
  nor (_30168_, _30166_, _30162_);
  nor (_30169_, _30168_, _30098_);
  nor (_30170_, _30169_, _03767_);
  nor (_30171_, _30118_, _03948_);
  or (_30172_, _30171_, _03473_);
  nor (_30173_, _30172_, _30170_);
  and (_30174_, _13051_, _05342_);
  or (_30175_, _30095_, _03474_);
  nor (_30176_, _30175_, _30174_);
  nor (_30177_, _30176_, _30173_);
  or (_30179_, _30177_, _43193_);
  or (_30180_, _43189_, \oc8051_golden_model_1.TH1 [4]);
  and (_30181_, _30180_, _42003_);
  and (_43888_, _30181_, _30179_);
  not (_30182_, \oc8051_golden_model_1.TH1 [5]);
  nor (_30183_, _05342_, _30182_);
  nor (_30184_, _13203_, _11066_);
  nor (_30185_, _30184_, _30183_);
  nor (_30186_, _30185_, _06458_);
  and (_30187_, _13204_, _05342_);
  nor (_30189_, _30187_, _30183_);
  nor (_30190_, _30189_, _03745_);
  and (_30191_, _06757_, _05342_);
  or (_30192_, _30191_, _30183_);
  and (_30193_, _30192_, _04082_);
  and (_30194_, _05342_, \oc8051_golden_model_1.ACC [5]);
  nor (_30195_, _30194_, _30183_);
  nor (_30196_, _30195_, _03531_);
  nor (_30197_, _30195_, _04437_);
  nor (_30198_, _04436_, _30182_);
  or (_30200_, _30198_, _30197_);
  and (_30201_, _30200_, _04432_);
  nor (_30202_, _13070_, _11066_);
  nor (_30203_, _30202_, _30183_);
  nor (_30204_, _30203_, _04432_);
  or (_30205_, _30204_, _30201_);
  and (_30206_, _30205_, _04457_);
  nor (_30207_, _05526_, _11066_);
  nor (_30208_, _30207_, _30183_);
  nor (_30209_, _30208_, _04457_);
  nor (_30211_, _30209_, _30206_);
  nor (_30212_, _30211_, _03530_);
  or (_30213_, _30212_, _07454_);
  nor (_30214_, _30213_, _30196_);
  and (_30215_, _30208_, _07454_);
  or (_30216_, _30215_, _04082_);
  nor (_30217_, _30216_, _30214_);
  or (_30218_, _30217_, _30193_);
  and (_30219_, _30218_, _03521_);
  nor (_30220_, _13184_, _11066_);
  nor (_30222_, _30220_, _30183_);
  nor (_30223_, _30222_, _03521_);
  or (_30224_, _30223_, _08905_);
  or (_30225_, _30224_, _30219_);
  and (_30226_, _13198_, _05342_);
  or (_30227_, _30183_, _04527_);
  or (_30228_, _30227_, _30226_);
  and (_30229_, _06295_, _05342_);
  nor (_30230_, _30229_, _30183_);
  and (_30231_, _30230_, _03624_);
  nor (_30233_, _30231_, _03744_);
  and (_30234_, _30233_, _30228_);
  and (_30235_, _30234_, _30225_);
  nor (_30236_, _30235_, _30190_);
  nor (_30237_, _30236_, _03611_);
  nor (_30238_, _30183_, _05576_);
  not (_30239_, _30238_);
  nor (_30240_, _30230_, _04523_);
  and (_30241_, _30240_, _30239_);
  nor (_30242_, _30241_, _30237_);
  nor (_30244_, _30242_, _03733_);
  nor (_30245_, _30195_, _03734_);
  and (_30246_, _30245_, _30239_);
  nor (_30247_, _30246_, _03618_);
  not (_30248_, _30247_);
  nor (_30249_, _30248_, _30244_);
  nor (_30250_, _13197_, _11066_);
  or (_30251_, _30183_, _06453_);
  nor (_30252_, _30251_, _30250_);
  or (_30253_, _30252_, _03741_);
  nor (_30255_, _30253_, _30249_);
  nor (_30256_, _30255_, _30186_);
  nor (_30257_, _30256_, _03767_);
  nor (_30258_, _30203_, _03948_);
  or (_30259_, _30258_, _03473_);
  nor (_30260_, _30259_, _30257_);
  and (_30261_, _13253_, _05342_);
  or (_30262_, _30183_, _03474_);
  nor (_30263_, _30262_, _30261_);
  nor (_30264_, _30263_, _30260_);
  or (_30266_, _30264_, _43193_);
  or (_30267_, _43189_, \oc8051_golden_model_1.TH1 [5]);
  and (_30268_, _30267_, _42003_);
  and (_43889_, _30268_, _30266_);
  not (_30269_, \oc8051_golden_model_1.TH1 [6]);
  nor (_30270_, _05342_, _30269_);
  nor (_30271_, _13406_, _11066_);
  nor (_30272_, _30271_, _30270_);
  nor (_30273_, _30272_, _06458_);
  and (_30274_, _13407_, _05342_);
  nor (_30276_, _30274_, _30270_);
  nor (_30277_, _30276_, _03745_);
  and (_30278_, _06526_, _05342_);
  or (_30279_, _30278_, _30270_);
  and (_30280_, _30279_, _04082_);
  and (_30281_, _05342_, \oc8051_golden_model_1.ACC [6]);
  nor (_30282_, _30281_, _30270_);
  nor (_30283_, _30282_, _03531_);
  nor (_30284_, _30282_, _04437_);
  nor (_30285_, _04436_, _30269_);
  or (_30287_, _30285_, _30284_);
  and (_30288_, _30287_, _04432_);
  nor (_30289_, _13293_, _11066_);
  nor (_30290_, _30289_, _30270_);
  nor (_30291_, _30290_, _04432_);
  or (_30292_, _30291_, _30288_);
  and (_30293_, _30292_, _04457_);
  nor (_30294_, _05417_, _11066_);
  nor (_30295_, _30294_, _30270_);
  nor (_30296_, _30295_, _04457_);
  nor (_30298_, _30296_, _30293_);
  nor (_30299_, _30298_, _03530_);
  or (_30300_, _30299_, _07454_);
  nor (_30301_, _30300_, _30283_);
  and (_30302_, _30295_, _07454_);
  or (_30303_, _30302_, _04082_);
  nor (_30304_, _30303_, _30301_);
  or (_30305_, _30304_, _30280_);
  and (_30306_, _30305_, _03521_);
  nor (_30307_, _13387_, _11066_);
  nor (_30309_, _30307_, _30270_);
  nor (_30310_, _30309_, _03521_);
  or (_30311_, _30310_, _08905_);
  or (_30312_, _30311_, _30306_);
  and (_30313_, _13402_, _05342_);
  or (_30314_, _30270_, _04527_);
  or (_30315_, _30314_, _30313_);
  and (_30316_, _14949_, _05342_);
  nor (_30317_, _30316_, _30270_);
  and (_30318_, _30317_, _03624_);
  nor (_30320_, _30318_, _03744_);
  and (_30321_, _30320_, _30315_);
  and (_30322_, _30321_, _30312_);
  nor (_30323_, _30322_, _30277_);
  nor (_30324_, _30323_, _03611_);
  nor (_30325_, _30270_, _05469_);
  not (_30326_, _30325_);
  nor (_30327_, _30317_, _04523_);
  and (_30328_, _30327_, _30326_);
  nor (_30329_, _30328_, _30324_);
  nor (_30331_, _30329_, _03733_);
  nor (_30332_, _30282_, _03734_);
  and (_30333_, _30332_, _30326_);
  or (_30334_, _30333_, _30331_);
  and (_30335_, _30334_, _06453_);
  nor (_30336_, _13400_, _11066_);
  nor (_30337_, _30336_, _30270_);
  nor (_30338_, _30337_, _06453_);
  or (_30339_, _30338_, _30335_);
  and (_30340_, _30339_, _06458_);
  nor (_30342_, _30340_, _30273_);
  nor (_30343_, _30342_, _03767_);
  nor (_30344_, _30290_, _03948_);
  or (_30345_, _30344_, _03473_);
  nor (_30346_, _30345_, _30343_);
  and (_30347_, _13456_, _05342_);
  or (_30348_, _30270_, _03474_);
  nor (_30349_, _30348_, _30347_);
  nor (_30350_, _30349_, _30346_);
  or (_30351_, _30350_, _43193_);
  or (_30353_, _43189_, \oc8051_golden_model_1.TH1 [6]);
  and (_30354_, _30353_, _42003_);
  and (_43890_, _30354_, _30351_);
  not (_30355_, \oc8051_golden_model_1.TL0 [0]);
  nor (_30356_, _05348_, _30355_);
  nor (_30357_, _05722_, _11147_);
  nor (_30358_, _30357_, _30356_);
  and (_30359_, _30358_, _17198_);
  and (_30360_, _05348_, \oc8051_golden_model_1.ACC [0]);
  nor (_30361_, _30360_, _30356_);
  nor (_30363_, _30361_, _03531_);
  nor (_30364_, _30361_, _04437_);
  nor (_30365_, _04436_, _30355_);
  or (_30366_, _30365_, _30364_);
  and (_30367_, _30366_, _04432_);
  nor (_30368_, _30358_, _04432_);
  or (_30369_, _30368_, _30367_);
  and (_30370_, _30369_, _04457_);
  and (_30371_, _05348_, _04429_);
  nor (_30372_, _30371_, _30356_);
  nor (_30374_, _30372_, _04457_);
  nor (_30375_, _30374_, _30370_);
  nor (_30376_, _30375_, _03530_);
  or (_30377_, _30376_, _07454_);
  nor (_30378_, _30377_, _30363_);
  and (_30379_, _30372_, _07454_);
  nor (_30380_, _30379_, _30378_);
  nor (_30381_, _30380_, _04082_);
  and (_30382_, _06617_, _05348_);
  nor (_30383_, _30356_, _04500_);
  not (_30385_, _30383_);
  nor (_30386_, _30385_, _30382_);
  nor (_30387_, _30386_, _30381_);
  nor (_30388_, _30387_, _03224_);
  nor (_30389_, _12164_, _11147_);
  or (_30390_, _30356_, _03521_);
  nor (_30391_, _30390_, _30389_);
  or (_30392_, _30391_, _03624_);
  nor (_30393_, _30392_, _30388_);
  and (_30394_, _05348_, _06350_);
  nor (_30395_, _30394_, _30356_);
  nor (_30396_, _30395_, _04509_);
  or (_30397_, _30396_, _30393_);
  and (_30398_, _30397_, _04527_);
  and (_30399_, _12177_, _05348_);
  nor (_30400_, _30399_, _30356_);
  nor (_30401_, _30400_, _04527_);
  or (_30402_, _30401_, _30398_);
  nor (_30403_, _30402_, _03744_);
  and (_30404_, _12183_, _05348_);
  or (_30407_, _30356_, _03745_);
  nor (_30408_, _30407_, _30404_);
  or (_30409_, _30408_, _03611_);
  nor (_30410_, _30409_, _30403_);
  or (_30411_, _30395_, _04523_);
  nor (_30412_, _30411_, _30357_);
  nor (_30413_, _30412_, _30410_);
  nor (_30414_, _30413_, _03733_);
  nor (_30415_, _30356_, _05722_);
  or (_30416_, _30415_, _03734_);
  nor (_30418_, _30416_, _30361_);
  or (_30419_, _30418_, _30414_);
  and (_30420_, _30419_, _06453_);
  nor (_30421_, _12057_, _11147_);
  nor (_30422_, _30421_, _30356_);
  nor (_30423_, _30422_, _06453_);
  or (_30424_, _30423_, _30420_);
  and (_30425_, _30424_, _06458_);
  nor (_30426_, _12181_, _11147_);
  nor (_30427_, _30426_, _30356_);
  nor (_30429_, _30427_, _06458_);
  nor (_30430_, _30429_, _17198_);
  not (_30431_, _30430_);
  nor (_30432_, _30431_, _30425_);
  nor (_30433_, _30432_, _30359_);
  or (_30434_, _30433_, _43193_);
  or (_30435_, _43189_, \oc8051_golden_model_1.TL0 [0]);
  and (_30436_, _30435_, _42003_);
  and (_43893_, _30436_, _30434_);
  and (_30437_, _06572_, _05348_);
  not (_30439_, \oc8051_golden_model_1.TL0 [1]);
  nor (_30440_, _05348_, _30439_);
  nor (_30441_, _30440_, _04500_);
  not (_30442_, _30441_);
  nor (_30443_, _30442_, _30437_);
  not (_30444_, _30443_);
  nor (_30445_, _11147_, _04635_);
  nor (_30446_, _30445_, _30440_);
  and (_30447_, _30446_, _07454_);
  nor (_30448_, _05348_, \oc8051_golden_model_1.TL0 [1]);
  and (_30450_, _05348_, _03269_);
  nor (_30451_, _30450_, _30448_);
  and (_30452_, _30451_, _04436_);
  nor (_30453_, _04436_, _30439_);
  or (_30454_, _30453_, _30452_);
  and (_30455_, _30454_, _04432_);
  and (_30456_, _12265_, _05348_);
  nor (_30457_, _30456_, _30448_);
  and (_30458_, _30457_, _03534_);
  or (_30459_, _30458_, _30455_);
  and (_30461_, _30459_, _04457_);
  nor (_30462_, _30446_, _04457_);
  nor (_30463_, _30462_, _30461_);
  nor (_30464_, _30463_, _03530_);
  and (_30465_, _30451_, _03530_);
  nor (_30466_, _30465_, _07454_);
  not (_30467_, _30466_);
  nor (_30468_, _30467_, _30464_);
  nor (_30469_, _30468_, _30447_);
  nor (_30471_, _30469_, _04082_);
  nor (_30474_, _30471_, _03224_);
  and (_30476_, _30474_, _30444_);
  not (_30478_, _30448_);
  and (_30480_, _12360_, _05348_);
  nor (_30482_, _30480_, _03521_);
  and (_30484_, _30482_, _30478_);
  nor (_30486_, _30484_, _30476_);
  nor (_30488_, _30486_, _08905_);
  nor (_30490_, _12375_, _11147_);
  nor (_30492_, _30490_, _04527_);
  and (_30494_, _05348_, _04325_);
  nor (_30495_, _30494_, _04509_);
  or (_30496_, _30495_, _30492_);
  and (_30497_, _30496_, _30478_);
  nor (_30498_, _30497_, _30488_);
  nor (_30499_, _30498_, _03744_);
  nor (_30500_, _12381_, _11147_);
  nor (_30501_, _30500_, _03745_);
  and (_30502_, _30501_, _30478_);
  nor (_30503_, _30502_, _30499_);
  nor (_30505_, _30503_, _03611_);
  nor (_30506_, _12374_, _11147_);
  nor (_30507_, _30506_, _04523_);
  and (_30508_, _30507_, _30478_);
  nor (_30509_, _30508_, _30505_);
  nor (_30510_, _30509_, _03733_);
  nor (_30511_, _30440_, _05674_);
  nor (_30512_, _30511_, _03734_);
  and (_30513_, _30512_, _30451_);
  nor (_30514_, _30513_, _30510_);
  or (_30516_, _30514_, _18526_);
  and (_30517_, _30450_, _05673_);
  nor (_30518_, _30517_, _06458_);
  and (_30519_, _30518_, _30478_);
  nor (_30520_, _30519_, _03767_);
  and (_30521_, _30494_, _05673_);
  or (_30522_, _30448_, _06453_);
  or (_30523_, _30522_, _30521_);
  and (_30524_, _30523_, _30520_);
  and (_30525_, _30524_, _30516_);
  nor (_30527_, _30457_, _03948_);
  nor (_30528_, _30527_, _30525_);
  and (_30529_, _30528_, _03474_);
  nor (_30530_, _30456_, _30440_);
  nor (_30531_, _30530_, _03474_);
  or (_30532_, _30531_, _30529_);
  or (_30533_, _30532_, _43193_);
  or (_30534_, _43189_, \oc8051_golden_model_1.TL0 [1]);
  and (_30535_, _30534_, _42003_);
  and (_43894_, _30535_, _30533_);
  not (_30537_, \oc8051_golden_model_1.TL0 [2]);
  nor (_30538_, _05348_, _30537_);
  nor (_30539_, _12587_, _11147_);
  nor (_30540_, _30539_, _30538_);
  nor (_30541_, _30540_, _06458_);
  and (_30542_, _12588_, _05348_);
  nor (_30543_, _30542_, _30538_);
  nor (_30544_, _30543_, _03745_);
  nor (_30545_, _11147_, _05073_);
  nor (_30546_, _30545_, _30538_);
  and (_30548_, _30546_, _07454_);
  and (_30549_, _05348_, \oc8051_golden_model_1.ACC [2]);
  nor (_30550_, _30549_, _30538_);
  nor (_30551_, _30550_, _03531_);
  nor (_30552_, _30550_, _04437_);
  nor (_30553_, _04436_, _30537_);
  or (_30554_, _30553_, _30552_);
  and (_30555_, _30554_, _04432_);
  nor (_30556_, _12467_, _11147_);
  nor (_30557_, _30556_, _30538_);
  nor (_30559_, _30557_, _04432_);
  or (_30560_, _30559_, _30555_);
  and (_30561_, _30560_, _04457_);
  nor (_30562_, _30546_, _04457_);
  nor (_30563_, _30562_, _30561_);
  nor (_30564_, _30563_, _03530_);
  or (_30565_, _30564_, _07454_);
  nor (_30566_, _30565_, _30551_);
  nor (_30567_, _30566_, _30548_);
  nor (_30568_, _30567_, _04082_);
  and (_30570_, _06710_, _05348_);
  nor (_30571_, _30538_, _04500_);
  not (_30572_, _30571_);
  nor (_30573_, _30572_, _30570_);
  nor (_30574_, _30573_, _03224_);
  not (_30575_, _30574_);
  nor (_30576_, _30575_, _30568_);
  nor (_30577_, _12568_, _11147_);
  nor (_30578_, _30577_, _30538_);
  nor (_30579_, _30578_, _03521_);
  or (_30581_, _30579_, _08905_);
  or (_30582_, _30581_, _30576_);
  and (_30583_, _12582_, _05348_);
  or (_30584_, _30538_, _04527_);
  or (_30585_, _30584_, _30583_);
  and (_30586_, _05348_, _06399_);
  nor (_30587_, _30586_, _30538_);
  and (_30588_, _30587_, _03624_);
  nor (_30589_, _30588_, _03744_);
  and (_30590_, _30589_, _30585_);
  and (_30592_, _30590_, _30582_);
  nor (_30593_, _30592_, _30544_);
  nor (_30594_, _30593_, _03611_);
  nor (_30595_, _30538_, _05772_);
  not (_30596_, _30595_);
  nor (_30597_, _30587_, _04523_);
  and (_30598_, _30597_, _30596_);
  nor (_30599_, _30598_, _30594_);
  nor (_30600_, _30599_, _03733_);
  nor (_30601_, _30550_, _03734_);
  and (_30603_, _30601_, _30596_);
  nor (_30604_, _30603_, _03618_);
  not (_30605_, _30604_);
  nor (_30606_, _30605_, _30600_);
  nor (_30607_, _12581_, _11147_);
  or (_30608_, _30538_, _06453_);
  nor (_30609_, _30608_, _30607_);
  or (_30610_, _30609_, _03741_);
  nor (_30611_, _30610_, _30606_);
  nor (_30612_, _30611_, _30541_);
  nor (_30614_, _30612_, _03767_);
  nor (_30615_, _30557_, _03948_);
  or (_30616_, _30615_, _03473_);
  nor (_30617_, _30616_, _30614_);
  and (_30618_, _12638_, _05348_);
  or (_30619_, _30538_, _03474_);
  nor (_30620_, _30619_, _30618_);
  nor (_30621_, _30620_, _30617_);
  or (_30622_, _30621_, _43193_);
  or (_30623_, _43189_, \oc8051_golden_model_1.TL0 [2]);
  and (_30625_, _30623_, _42003_);
  and (_43895_, _30625_, _30622_);
  not (_30626_, \oc8051_golden_model_1.TL0 [3]);
  nor (_30627_, _05348_, _30626_);
  nor (_30628_, _12792_, _11147_);
  nor (_30629_, _30628_, _30627_);
  nor (_30630_, _30629_, _06458_);
  and (_30631_, _12793_, _05348_);
  nor (_30632_, _30631_, _30627_);
  nor (_30633_, _30632_, _03745_);
  and (_30635_, _06664_, _05348_);
  or (_30636_, _30635_, _30627_);
  and (_30637_, _30636_, _04082_);
  and (_30638_, _05348_, \oc8051_golden_model_1.ACC [3]);
  nor (_30639_, _30638_, _30627_);
  nor (_30640_, _30639_, _03531_);
  nor (_30641_, _30639_, _04437_);
  nor (_30642_, _04436_, _30626_);
  or (_30643_, _30642_, _30641_);
  and (_30644_, _30643_, _04432_);
  nor (_30646_, _12652_, _11147_);
  nor (_30647_, _30646_, _30627_);
  nor (_30648_, _30647_, _04432_);
  or (_30649_, _30648_, _30644_);
  and (_30650_, _30649_, _04457_);
  nor (_30651_, _11147_, _04885_);
  nor (_30652_, _30651_, _30627_);
  nor (_30653_, _30652_, _04457_);
  nor (_30654_, _30653_, _30650_);
  nor (_30655_, _30654_, _03530_);
  or (_30657_, _30655_, _07454_);
  nor (_30658_, _30657_, _30640_);
  and (_30659_, _30652_, _07454_);
  or (_30660_, _30659_, _04082_);
  nor (_30661_, _30660_, _30658_);
  or (_30662_, _30661_, _30637_);
  and (_30663_, _30662_, _03521_);
  nor (_30664_, _12773_, _11147_);
  nor (_30665_, _30664_, _30627_);
  nor (_30666_, _30665_, _03521_);
  or (_30668_, _30666_, _08905_);
  or (_30669_, _30668_, _30663_);
  and (_30670_, _12787_, _05348_);
  or (_30671_, _30627_, _04527_);
  or (_30672_, _30671_, _30670_);
  and (_30673_, _05348_, _06356_);
  nor (_30674_, _30673_, _30627_);
  and (_30675_, _30674_, _03624_);
  nor (_30676_, _30675_, _03744_);
  and (_30677_, _30676_, _30672_);
  and (_30679_, _30677_, _30669_);
  nor (_30680_, _30679_, _30633_);
  nor (_30681_, _30680_, _03611_);
  nor (_30682_, _30627_, _05625_);
  not (_30683_, _30682_);
  nor (_30684_, _30674_, _04523_);
  and (_30685_, _30684_, _30683_);
  nor (_30686_, _30685_, _30681_);
  nor (_30687_, _30686_, _03733_);
  nor (_30688_, _30639_, _03734_);
  and (_30690_, _30688_, _30683_);
  or (_30691_, _30690_, _30687_);
  and (_30692_, _30691_, _06453_);
  nor (_30693_, _12786_, _11147_);
  nor (_30694_, _30693_, _30627_);
  nor (_30695_, _30694_, _06453_);
  or (_30696_, _30695_, _30692_);
  and (_30697_, _30696_, _06458_);
  nor (_30698_, _30697_, _30630_);
  nor (_30699_, _30698_, _03767_);
  nor (_30701_, _30647_, _03948_);
  or (_30702_, _30701_, _03473_);
  nor (_30703_, _30702_, _30699_);
  and (_30704_, _12843_, _05348_);
  or (_30705_, _30627_, _03474_);
  nor (_30706_, _30705_, _30704_);
  nor (_30707_, _30706_, _30703_);
  or (_30708_, _30707_, _43193_);
  or (_30709_, _43189_, \oc8051_golden_model_1.TL0 [3]);
  and (_30710_, _30709_, _42003_);
  and (_43896_, _30710_, _30708_);
  not (_30712_, \oc8051_golden_model_1.TL0 [4]);
  nor (_30713_, _05348_, _30712_);
  nor (_30714_, _12991_, _11147_);
  nor (_30715_, _30714_, _30713_);
  nor (_30716_, _30715_, _06458_);
  and (_30717_, _12992_, _05348_);
  nor (_30718_, _30717_, _30713_);
  nor (_30719_, _30718_, _03745_);
  and (_30720_, _06337_, _05348_);
  nor (_30722_, _30720_, _30713_);
  and (_30723_, _30722_, _03624_);
  and (_30724_, _05348_, \oc8051_golden_model_1.ACC [4]);
  nor (_30725_, _30724_, _30713_);
  nor (_30726_, _30725_, _03531_);
  nor (_30727_, _30725_, _04437_);
  nor (_30728_, _04436_, _30712_);
  or (_30729_, _30728_, _30727_);
  and (_30730_, _30729_, _04432_);
  nor (_30731_, _12856_, _11147_);
  nor (_30733_, _30731_, _30713_);
  nor (_30734_, _30733_, _04432_);
  or (_30735_, _30734_, _30730_);
  and (_30736_, _30735_, _04457_);
  nor (_30737_, _05831_, _11147_);
  nor (_30738_, _30737_, _30713_);
  nor (_30739_, _30738_, _04457_);
  nor (_30740_, _30739_, _30736_);
  nor (_30741_, _30740_, _03530_);
  or (_30742_, _30741_, _07454_);
  nor (_30744_, _30742_, _30726_);
  and (_30745_, _30738_, _07454_);
  nor (_30746_, _30745_, _30744_);
  nor (_30747_, _30746_, _04082_);
  and (_30748_, _06802_, _05348_);
  nor (_30749_, _30713_, _04500_);
  not (_30750_, _30749_);
  nor (_30751_, _30750_, _30748_);
  or (_30752_, _30751_, _03224_);
  nor (_30753_, _30752_, _30747_);
  nor (_30755_, _12972_, _11147_);
  nor (_30756_, _30755_, _30713_);
  nor (_30757_, _30756_, _03521_);
  or (_30758_, _30757_, _03624_);
  nor (_30759_, _30758_, _30753_);
  nor (_30760_, _30759_, _30723_);
  or (_30761_, _30760_, _03623_);
  and (_30762_, _12986_, _05348_);
  or (_30763_, _30762_, _30713_);
  or (_30764_, _30763_, _04527_);
  and (_30766_, _30764_, _03745_);
  and (_30767_, _30766_, _30761_);
  nor (_30768_, _30767_, _30719_);
  nor (_30769_, _30768_, _03611_);
  nor (_30770_, _30713_, _05880_);
  not (_30771_, _30770_);
  nor (_30772_, _30722_, _04523_);
  and (_30773_, _30772_, _30771_);
  nor (_30774_, _30773_, _30769_);
  nor (_30775_, _30774_, _03733_);
  nor (_30777_, _30725_, _03734_);
  and (_30778_, _30777_, _30771_);
  or (_30779_, _30778_, _30775_);
  and (_30780_, _30779_, _06453_);
  nor (_30781_, _12985_, _11147_);
  nor (_30782_, _30781_, _30713_);
  nor (_30783_, _30782_, _06453_);
  or (_30784_, _30783_, _30780_);
  and (_30785_, _30784_, _06458_);
  nor (_30786_, _30785_, _30716_);
  nor (_30788_, _30786_, _03767_);
  nor (_30789_, _30733_, _03948_);
  or (_30790_, _30789_, _03473_);
  nor (_30791_, _30790_, _30788_);
  and (_30792_, _13051_, _05348_);
  or (_30793_, _30713_, _03474_);
  nor (_30794_, _30793_, _30792_);
  nor (_30795_, _30794_, _30791_);
  or (_30796_, _30795_, _43193_);
  or (_30797_, _43189_, \oc8051_golden_model_1.TL0 [4]);
  and (_30799_, _30797_, _42003_);
  and (_43897_, _30799_, _30796_);
  not (_30800_, \oc8051_golden_model_1.TL0 [5]);
  nor (_30801_, _05348_, _30800_);
  nor (_30802_, _13203_, _11147_);
  nor (_30803_, _30802_, _30801_);
  nor (_30804_, _30803_, _06458_);
  and (_30805_, _13204_, _05348_);
  nor (_30806_, _30805_, _30801_);
  nor (_30807_, _30806_, _03745_);
  and (_30809_, _06757_, _05348_);
  or (_30810_, _30809_, _30801_);
  and (_30811_, _30810_, _04082_);
  and (_30812_, _05348_, \oc8051_golden_model_1.ACC [5]);
  nor (_30813_, _30812_, _30801_);
  nor (_30814_, _30813_, _03531_);
  nor (_30815_, _30813_, _04437_);
  nor (_30816_, _04436_, _30800_);
  or (_30817_, _30816_, _30815_);
  and (_30818_, _30817_, _04432_);
  nor (_30820_, _13070_, _11147_);
  nor (_30821_, _30820_, _30801_);
  nor (_30822_, _30821_, _04432_);
  or (_30823_, _30822_, _30818_);
  and (_30824_, _30823_, _04457_);
  nor (_30825_, _05526_, _11147_);
  nor (_30826_, _30825_, _30801_);
  nor (_30827_, _30826_, _04457_);
  nor (_30828_, _30827_, _30824_);
  nor (_30829_, _30828_, _03530_);
  or (_30831_, _30829_, _07454_);
  nor (_30832_, _30831_, _30814_);
  and (_30833_, _30826_, _07454_);
  or (_30834_, _30833_, _04082_);
  nor (_30835_, _30834_, _30832_);
  or (_30836_, _30835_, _30811_);
  and (_30837_, _30836_, _03521_);
  nor (_30838_, _13184_, _11147_);
  nor (_30839_, _30838_, _30801_);
  nor (_30840_, _30839_, _03521_);
  or (_30842_, _30840_, _08905_);
  or (_30843_, _30842_, _30837_);
  and (_30844_, _13198_, _05348_);
  or (_30845_, _30801_, _04527_);
  or (_30846_, _30845_, _30844_);
  and (_30847_, _06295_, _05348_);
  nor (_30848_, _30847_, _30801_);
  and (_30849_, _30848_, _03624_);
  nor (_30850_, _30849_, _03744_);
  and (_30851_, _30850_, _30846_);
  and (_30853_, _30851_, _30843_);
  nor (_30854_, _30853_, _30807_);
  nor (_30855_, _30854_, _03611_);
  nor (_30856_, _30801_, _05576_);
  not (_30857_, _30856_);
  nor (_30858_, _30848_, _04523_);
  and (_30859_, _30858_, _30857_);
  nor (_30860_, _30859_, _30855_);
  nor (_30861_, _30860_, _03733_);
  nor (_30862_, _30813_, _03734_);
  and (_30864_, _30862_, _30857_);
  nor (_30865_, _30864_, _03618_);
  not (_30866_, _30865_);
  nor (_30867_, _30866_, _30861_);
  nor (_30868_, _13197_, _11147_);
  or (_30869_, _30801_, _06453_);
  nor (_30870_, _30869_, _30868_);
  or (_30871_, _30870_, _03741_);
  nor (_30872_, _30871_, _30867_);
  nor (_30873_, _30872_, _30804_);
  nor (_30875_, _30873_, _03767_);
  nor (_30876_, _30821_, _03948_);
  or (_30877_, _30876_, _03473_);
  nor (_30878_, _30877_, _30875_);
  and (_30879_, _13253_, _05348_);
  or (_30880_, _30801_, _03474_);
  nor (_30881_, _30880_, _30879_);
  nor (_30882_, _30881_, _30878_);
  or (_30883_, _30882_, _43193_);
  or (_30884_, _43189_, \oc8051_golden_model_1.TL0 [5]);
  and (_30885_, _30884_, _42003_);
  and (_43898_, _30885_, _30883_);
  not (_30886_, \oc8051_golden_model_1.TL0 [6]);
  nor (_30887_, _05348_, _30886_);
  nor (_30888_, _13406_, _11147_);
  nor (_30889_, _30888_, _30887_);
  nor (_30890_, _30889_, _06458_);
  and (_30891_, _13407_, _05348_);
  nor (_30892_, _30891_, _30887_);
  nor (_30893_, _30892_, _03745_);
  and (_30896_, _06526_, _05348_);
  or (_30897_, _30896_, _30887_);
  and (_30898_, _30897_, _04082_);
  and (_30899_, _05348_, \oc8051_golden_model_1.ACC [6]);
  nor (_30900_, _30899_, _30887_);
  nor (_30901_, _30900_, _04437_);
  nor (_30902_, _04436_, _30886_);
  or (_30903_, _30902_, _30901_);
  and (_30904_, _30903_, _04432_);
  nor (_30905_, _13293_, _11147_);
  nor (_30906_, _30905_, _30887_);
  nor (_30907_, _30906_, _04432_);
  or (_30908_, _30907_, _30904_);
  and (_30909_, _30908_, _04457_);
  nor (_30910_, _05417_, _11147_);
  nor (_30911_, _30910_, _30887_);
  nor (_30912_, _30911_, _04457_);
  nor (_30913_, _30912_, _30909_);
  nor (_30914_, _30913_, _03530_);
  nor (_30915_, _30900_, _03531_);
  nor (_30917_, _30915_, _07454_);
  not (_30918_, _30917_);
  nor (_30919_, _30918_, _30914_);
  and (_30920_, _30911_, _07454_);
  or (_30921_, _30920_, _04082_);
  nor (_30922_, _30921_, _30919_);
  or (_30923_, _30922_, _30898_);
  and (_30924_, _30923_, _03521_);
  nor (_30925_, _13387_, _11147_);
  nor (_30926_, _30925_, _30887_);
  nor (_30928_, _30926_, _03521_);
  or (_30929_, _30928_, _08905_);
  or (_30930_, _30929_, _30924_);
  and (_30931_, _13402_, _05348_);
  or (_30932_, _30887_, _04527_);
  or (_30933_, _30932_, _30931_);
  and (_30934_, _14949_, _05348_);
  nor (_30935_, _30934_, _30887_);
  and (_30936_, _30935_, _03624_);
  nor (_30937_, _30936_, _03744_);
  and (_30939_, _30937_, _30933_);
  and (_30940_, _30939_, _30930_);
  nor (_30941_, _30940_, _30893_);
  nor (_30942_, _30941_, _03611_);
  nor (_30943_, _30887_, _05469_);
  not (_30944_, _30943_);
  nor (_30945_, _30935_, _04523_);
  and (_30946_, _30945_, _30944_);
  nor (_30947_, _30946_, _30942_);
  nor (_30948_, _30947_, _03733_);
  nor (_30950_, _30900_, _03734_);
  and (_30951_, _30950_, _30944_);
  nor (_30952_, _30951_, _03618_);
  not (_30953_, _30952_);
  nor (_30954_, _30953_, _30948_);
  nor (_30955_, _13400_, _11147_);
  or (_30956_, _30887_, _06453_);
  nor (_30957_, _30956_, _30955_);
  or (_30958_, _30957_, _03741_);
  nor (_30959_, _30958_, _30954_);
  nor (_30961_, _30959_, _30890_);
  nor (_30962_, _30961_, _03767_);
  nor (_30963_, _30906_, _03948_);
  or (_30964_, _30963_, _03473_);
  nor (_30965_, _30964_, _30962_);
  and (_30966_, _13456_, _05348_);
  or (_30967_, _30887_, _03474_);
  nor (_30968_, _30967_, _30966_);
  nor (_30969_, _30968_, _30965_);
  or (_30970_, _30969_, _43193_);
  or (_30972_, _43189_, \oc8051_golden_model_1.TL0 [6]);
  and (_30973_, _30972_, _42003_);
  and (_43899_, _30973_, _30970_);
  not (_30974_, \oc8051_golden_model_1.TL1 [0]);
  nor (_30975_, _05444_, _30974_);
  nor (_30976_, _05722_, _11229_);
  nor (_30977_, _30976_, _30975_);
  and (_30978_, _30977_, _17198_);
  and (_30979_, _05444_, \oc8051_golden_model_1.ACC [0]);
  nor (_30980_, _30979_, _30975_);
  nor (_30982_, _30980_, _03531_);
  nor (_30983_, _30980_, _04437_);
  nor (_30984_, _04436_, _30974_);
  or (_30985_, _30984_, _30983_);
  and (_30986_, _30985_, _04432_);
  nor (_30987_, _30977_, _04432_);
  or (_30988_, _30987_, _30986_);
  and (_30989_, _30988_, _04457_);
  and (_30990_, _05350_, _04429_);
  nor (_30991_, _30990_, _30975_);
  nor (_30993_, _30991_, _04457_);
  nor (_30994_, _30993_, _30989_);
  nor (_30995_, _30994_, _03530_);
  or (_30996_, _30995_, _07454_);
  nor (_30997_, _30996_, _30982_);
  and (_30998_, _30991_, _07454_);
  nor (_30999_, _30998_, _30997_);
  nor (_31000_, _30999_, _04082_);
  nor (_31001_, _30975_, _04500_);
  nand (_31002_, _06617_, _05350_);
  and (_31004_, _31002_, _31001_);
  nor (_31005_, _31004_, _31000_);
  nor (_31006_, _31005_, _03224_);
  or (_31007_, _12164_, _11229_);
  nor (_31008_, _30975_, _03521_);
  and (_31009_, _31008_, _31007_);
  or (_31010_, _31009_, _03624_);
  nor (_31011_, _31010_, _31006_);
  and (_31012_, _05444_, _06350_);
  nor (_31013_, _31012_, _30975_);
  nor (_31015_, _31013_, _04509_);
  or (_31016_, _31015_, _31011_);
  and (_31017_, _31016_, _04527_);
  and (_31018_, _12177_, _05444_);
  nor (_31019_, _31018_, _30975_);
  nor (_31020_, _31019_, _04527_);
  or (_31021_, _31020_, _31017_);
  nor (_31022_, _31021_, _03744_);
  nand (_31023_, _12183_, _05350_);
  nor (_31024_, _30975_, _03745_);
  and (_31026_, _31024_, _31023_);
  or (_31027_, _31026_, _03611_);
  nor (_31028_, _31027_, _31022_);
  nor (_31029_, _31013_, _04523_);
  not (_31030_, _31029_);
  nor (_31031_, _31030_, _30976_);
  nor (_31032_, _31031_, _31028_);
  nor (_31033_, _31032_, _03733_);
  nor (_31034_, _30975_, _05722_);
  or (_31035_, _31034_, _03734_);
  nor (_31037_, _31035_, _30980_);
  or (_31038_, _31037_, _31033_);
  and (_31039_, _31038_, _06453_);
  nor (_31040_, _12057_, _11263_);
  nor (_31041_, _31040_, _30975_);
  nor (_31042_, _31041_, _06453_);
  or (_31043_, _31042_, _31039_);
  and (_31044_, _31043_, _06458_);
  nor (_31045_, _12181_, _11229_);
  nor (_31046_, _31045_, _30975_);
  nor (_31048_, _31046_, _06458_);
  nor (_31049_, _31048_, _17198_);
  not (_31050_, _31049_);
  nor (_31051_, _31050_, _31044_);
  nor (_31052_, _31051_, _30978_);
  or (_31053_, _31052_, _43193_);
  or (_31054_, _43189_, \oc8051_golden_model_1.TL1 [0]);
  and (_31055_, _31054_, _42003_);
  and (_43902_, _31055_, _31053_);
  not (_31056_, \oc8051_golden_model_1.TL1 [1]);
  nor (_31058_, _05444_, _31056_);
  nor (_31059_, _11229_, _04635_);
  nor (_31060_, _31059_, _31058_);
  and (_31061_, _31060_, _07454_);
  nor (_31062_, _05444_, \oc8051_golden_model_1.TL1 [1]);
  and (_31063_, _05350_, _03269_);
  nor (_31064_, _31063_, _31062_);
  and (_31065_, _31064_, _03530_);
  and (_31066_, _31064_, _04436_);
  nor (_31067_, _04436_, _31056_);
  or (_31069_, _31067_, _31066_);
  and (_31070_, _31069_, _04432_);
  and (_31071_, _12265_, _05444_);
  nor (_31072_, _31071_, _31062_);
  and (_31073_, _31072_, _03534_);
  or (_31074_, _31073_, _31070_);
  and (_31075_, _31074_, _04457_);
  nor (_31076_, _31060_, _04457_);
  nor (_31077_, _31076_, _31075_);
  nor (_31078_, _31077_, _03530_);
  or (_31080_, _31078_, _07454_);
  nor (_31081_, _31080_, _31065_);
  nor (_31082_, _31081_, _31061_);
  nor (_31083_, _31082_, _04082_);
  nor (_31084_, _31083_, _03224_);
  nor (_31085_, _31058_, _04500_);
  nand (_31086_, _06572_, _05350_);
  nand (_31087_, _31086_, _31085_);
  and (_31088_, _31087_, _31084_);
  and (_31089_, _12360_, _05444_);
  or (_31091_, _31089_, _03521_);
  nor (_31092_, _31091_, _31062_);
  nor (_31093_, _31092_, _31088_);
  nor (_31094_, _31093_, _08905_);
  nor (_31095_, _12375_, _11229_);
  nor (_31096_, _31095_, _04527_);
  and (_31097_, _05350_, _04325_);
  nor (_31098_, _31097_, _04509_);
  nor (_31099_, _31098_, _31096_);
  nor (_31100_, _31099_, _31062_);
  nor (_31102_, _31100_, _31094_);
  nor (_31103_, _31102_, _03744_);
  nor (_31104_, _12381_, _11263_);
  or (_31105_, _31104_, _03745_);
  nor (_31106_, _31105_, _31062_);
  nor (_31107_, _31106_, _31103_);
  nor (_31108_, _31107_, _03611_);
  nor (_31109_, _12374_, _11263_);
  or (_31110_, _31109_, _04523_);
  nor (_31111_, _31110_, _31062_);
  nor (_31112_, _31111_, _31108_);
  nor (_31113_, _31112_, _03733_);
  nor (_31114_, _31058_, _05674_);
  nor (_31115_, _31114_, _03734_);
  and (_31116_, _31115_, _31064_);
  nor (_31117_, _31116_, _31113_);
  or (_31118_, _31117_, _18526_);
  nand (_31119_, _31097_, _05673_);
  nor (_31120_, _31062_, _06453_);
  and (_31121_, _31120_, _31119_);
  not (_31124_, _31121_);
  and (_31125_, _12380_, _05444_);
  or (_31126_, _31125_, _06458_);
  nor (_31127_, _31126_, _31062_);
  nor (_31128_, _31127_, _03767_);
  and (_31129_, _31128_, _31124_);
  and (_31130_, _31129_, _31118_);
  nor (_31131_, _31072_, _03948_);
  nor (_31132_, _31131_, _31130_);
  and (_31133_, _31132_, _03474_);
  nor (_31135_, _31071_, _31058_);
  nor (_31136_, _31135_, _03474_);
  or (_31137_, _31136_, _31133_);
  or (_31138_, _31137_, _43193_);
  or (_31139_, _43189_, \oc8051_golden_model_1.TL1 [1]);
  and (_31140_, _31139_, _42003_);
  and (_43903_, _31140_, _31138_);
  not (_31141_, \oc8051_golden_model_1.TL1 [2]);
  nor (_31142_, _05444_, _31141_);
  nor (_31143_, _12587_, _11229_);
  nor (_31145_, _31143_, _31142_);
  nor (_31146_, _31145_, _06458_);
  and (_31147_, _12588_, _05350_);
  nor (_31148_, _31147_, _31142_);
  nor (_31149_, _31148_, _03745_);
  and (_31150_, _05444_, \oc8051_golden_model_1.ACC [2]);
  nor (_31151_, _31150_, _31142_);
  nor (_31152_, _31151_, _03531_);
  nor (_31153_, _31151_, _04437_);
  nor (_31154_, _04436_, _31141_);
  or (_31156_, _31154_, _31153_);
  and (_31157_, _31156_, _04432_);
  nor (_31158_, _12467_, _11229_);
  nor (_31159_, _31158_, _31142_);
  nor (_31160_, _31159_, _04432_);
  or (_31161_, _31160_, _31157_);
  and (_31162_, _31161_, _04457_);
  nor (_31163_, _11229_, _05073_);
  nor (_31164_, _31163_, _31142_);
  nor (_31165_, _31164_, _04457_);
  nor (_31167_, _31165_, _31162_);
  nor (_31168_, _31167_, _03530_);
  or (_31169_, _31168_, _07454_);
  nor (_31170_, _31169_, _31152_);
  and (_31171_, _31164_, _07454_);
  nor (_31172_, _31171_, _31170_);
  nor (_31173_, _31172_, _04082_);
  nor (_31174_, _31142_, _04500_);
  nand (_31175_, _06710_, _05350_);
  and (_31176_, _31175_, _31174_);
  or (_31178_, _31176_, _03224_);
  nor (_31179_, _31178_, _31173_);
  nor (_31180_, _12568_, _11229_);
  nor (_31181_, _31180_, _31142_);
  nor (_31182_, _31181_, _03521_);
  or (_31183_, _31182_, _08905_);
  or (_31184_, _31183_, _31179_);
  and (_31185_, _12582_, _05350_);
  or (_31186_, _31142_, _04527_);
  or (_31187_, _31186_, _31185_);
  and (_31189_, _05444_, _06399_);
  nor (_31190_, _31189_, _31142_);
  and (_31191_, _31190_, _03624_);
  nor (_31192_, _31191_, _03744_);
  and (_31193_, _31192_, _31187_);
  and (_31194_, _31193_, _31184_);
  nor (_31195_, _31194_, _31149_);
  nor (_31196_, _31195_, _03611_);
  nor (_31197_, _31142_, _05772_);
  not (_31198_, _31197_);
  nor (_31200_, _31190_, _04523_);
  and (_31201_, _31200_, _31198_);
  nor (_31202_, _31201_, _31196_);
  nor (_31203_, _31202_, _03733_);
  nor (_31204_, _31151_, _03734_);
  and (_31205_, _31204_, _31198_);
  nor (_31206_, _31205_, _03618_);
  not (_31207_, _31206_);
  nor (_31208_, _31207_, _31203_);
  or (_31209_, _12581_, _11229_);
  nor (_31211_, _31142_, _06453_);
  and (_31212_, _31211_, _31209_);
  or (_31213_, _31212_, _03741_);
  nor (_31214_, _31213_, _31208_);
  nor (_31215_, _31214_, _31146_);
  nor (_31216_, _31215_, _03767_);
  nor (_31217_, _31159_, _03948_);
  or (_31218_, _31217_, _03473_);
  nor (_31219_, _31218_, _31216_);
  nand (_31220_, _12638_, _05350_);
  nor (_31222_, _31142_, _03474_);
  and (_31223_, _31222_, _31220_);
  nor (_31224_, _31223_, _31219_);
  or (_31225_, _31224_, _43193_);
  or (_31226_, _43189_, \oc8051_golden_model_1.TL1 [2]);
  and (_31227_, _31226_, _42003_);
  and (_43904_, _31227_, _31225_);
  not (_31228_, \oc8051_golden_model_1.TL1 [3]);
  nor (_31229_, _05444_, _31228_);
  nor (_31230_, _12792_, _11229_);
  nor (_31232_, _31230_, _31229_);
  nor (_31233_, _31232_, _06458_);
  and (_31234_, _12793_, _05350_);
  nor (_31235_, _31234_, _31229_);
  nor (_31236_, _31235_, _03745_);
  and (_31237_, _06664_, _05444_);
  or (_31238_, _31237_, _31229_);
  and (_31239_, _31238_, _04082_);
  and (_31240_, _05444_, \oc8051_golden_model_1.ACC [3]);
  nor (_31241_, _31240_, _31229_);
  nor (_31243_, _31241_, _03531_);
  nor (_31244_, _31241_, _04437_);
  nor (_31245_, _04436_, _31228_);
  or (_31246_, _31245_, _31244_);
  and (_31247_, _31246_, _04432_);
  nor (_31248_, _12652_, _11229_);
  nor (_31249_, _31248_, _31229_);
  nor (_31250_, _31249_, _04432_);
  or (_31251_, _31250_, _31247_);
  and (_31252_, _31251_, _04457_);
  nor (_31254_, _11229_, _04885_);
  nor (_31255_, _31254_, _31229_);
  nor (_31256_, _31255_, _04457_);
  nor (_31257_, _31256_, _31252_);
  nor (_31258_, _31257_, _03530_);
  or (_31259_, _31258_, _07454_);
  nor (_31260_, _31259_, _31243_);
  and (_31261_, _31255_, _07454_);
  or (_31262_, _31261_, _04082_);
  nor (_31263_, _31262_, _31260_);
  or (_31265_, _31263_, _31239_);
  and (_31266_, _31265_, _03521_);
  nor (_31267_, _12773_, _11229_);
  nor (_31268_, _31267_, _31229_);
  nor (_31269_, _31268_, _03521_);
  or (_31270_, _31269_, _08905_);
  or (_31271_, _31270_, _31266_);
  and (_31272_, _12787_, _05350_);
  or (_31273_, _31229_, _04527_);
  or (_31274_, _31273_, _31272_);
  and (_31276_, _05444_, _06356_);
  nor (_31277_, _31276_, _31229_);
  and (_31278_, _31277_, _03624_);
  nor (_31279_, _31278_, _03744_);
  and (_31280_, _31279_, _31274_);
  and (_31281_, _31280_, _31271_);
  nor (_31282_, _31281_, _31236_);
  nor (_31283_, _31282_, _03611_);
  nor (_31284_, _31229_, _05625_);
  not (_31285_, _31284_);
  nor (_31287_, _31277_, _04523_);
  and (_31288_, _31287_, _31285_);
  nor (_31289_, _31288_, _31283_);
  nor (_31290_, _31289_, _03733_);
  nor (_31291_, _31241_, _03734_);
  and (_31292_, _31291_, _31285_);
  nor (_31293_, _31292_, _03618_);
  not (_31294_, _31293_);
  nor (_31295_, _31294_, _31290_);
  or (_31296_, _12786_, _11229_);
  nor (_31298_, _31229_, _06453_);
  and (_31299_, _31298_, _31296_);
  or (_31300_, _31299_, _03741_);
  nor (_31301_, _31300_, _31295_);
  nor (_31302_, _31301_, _31233_);
  nor (_31303_, _31302_, _03767_);
  nor (_31304_, _31249_, _03948_);
  or (_31305_, _31304_, _03473_);
  nor (_31306_, _31305_, _31303_);
  nand (_31307_, _12843_, _05350_);
  nor (_31309_, _31229_, _03474_);
  and (_31310_, _31309_, _31307_);
  nor (_31311_, _31310_, _31306_);
  or (_31312_, _31311_, _43193_);
  or (_31313_, _43189_, \oc8051_golden_model_1.TL1 [3]);
  and (_31314_, _31313_, _42003_);
  and (_43905_, _31314_, _31312_);
  not (_31315_, \oc8051_golden_model_1.TL1 [4]);
  nor (_31316_, _05444_, _31315_);
  nor (_31317_, _12991_, _11229_);
  nor (_31319_, _31317_, _31316_);
  nor (_31320_, _31319_, _06458_);
  and (_31321_, _12992_, _05350_);
  nor (_31322_, _31321_, _31316_);
  nor (_31323_, _31322_, _03745_);
  and (_31324_, _06337_, _05444_);
  nor (_31325_, _31324_, _31316_);
  and (_31326_, _31325_, _03624_);
  nor (_31327_, _05831_, _11229_);
  nor (_31328_, _31327_, _31316_);
  and (_31330_, _31328_, _07454_);
  and (_31331_, _05444_, \oc8051_golden_model_1.ACC [4]);
  nor (_31332_, _31331_, _31316_);
  nor (_31333_, _31332_, _03531_);
  nor (_31334_, _31332_, _04437_);
  nor (_31335_, _04436_, _31315_);
  or (_31336_, _31335_, _31334_);
  and (_31337_, _31336_, _04432_);
  nor (_31338_, _12856_, _11229_);
  nor (_31339_, _31338_, _31316_);
  nor (_31341_, _31339_, _04432_);
  or (_31342_, _31341_, _31337_);
  and (_31343_, _31342_, _04457_);
  nor (_31344_, _31328_, _04457_);
  nor (_31345_, _31344_, _31343_);
  nor (_31346_, _31345_, _03530_);
  or (_31347_, _31346_, _07454_);
  nor (_31348_, _31347_, _31333_);
  nor (_31349_, _31348_, _31330_);
  nor (_31350_, _31349_, _04082_);
  nor (_31352_, _31316_, _04500_);
  nand (_31353_, _06802_, _05350_);
  and (_31354_, _31353_, _31352_);
  or (_31355_, _31354_, _03224_);
  nor (_31356_, _31355_, _31350_);
  nor (_31357_, _12972_, _11263_);
  nor (_31358_, _31357_, _31316_);
  nor (_31359_, _31358_, _03521_);
  or (_31360_, _31359_, _03624_);
  nor (_31361_, _31360_, _31356_);
  nor (_31363_, _31361_, _31326_);
  or (_31364_, _31363_, _03623_);
  and (_31365_, _12986_, _05444_);
  or (_31366_, _31365_, _31316_);
  or (_31367_, _31366_, _04527_);
  and (_31368_, _31367_, _03745_);
  and (_31369_, _31368_, _31364_);
  nor (_31370_, _31369_, _31323_);
  nor (_31371_, _31370_, _03611_);
  nor (_31372_, _31316_, _05880_);
  not (_31374_, _31372_);
  nor (_31375_, _31325_, _04523_);
  and (_31376_, _31375_, _31374_);
  nor (_31377_, _31376_, _31371_);
  nor (_31378_, _31377_, _03733_);
  nor (_31379_, _31332_, _03734_);
  and (_31380_, _31379_, _31374_);
  nor (_31381_, _31380_, _03618_);
  not (_31382_, _31381_);
  nor (_31383_, _31382_, _31378_);
  or (_31385_, _12985_, _11229_);
  nor (_31386_, _31316_, _06453_);
  and (_31387_, _31386_, _31385_);
  or (_31388_, _31387_, _03741_);
  nor (_31389_, _31388_, _31383_);
  nor (_31390_, _31389_, _31320_);
  nor (_31391_, _31390_, _03767_);
  nor (_31392_, _31339_, _03948_);
  or (_31393_, _31392_, _03473_);
  nor (_31394_, _31393_, _31391_);
  nand (_31396_, _13051_, _05350_);
  nor (_31397_, _31316_, _03474_);
  and (_31398_, _31397_, _31396_);
  nor (_31399_, _31398_, _31394_);
  or (_31400_, _31399_, _43193_);
  or (_31401_, _43189_, \oc8051_golden_model_1.TL1 [4]);
  and (_31402_, _31401_, _42003_);
  and (_43906_, _31402_, _31400_);
  not (_31403_, \oc8051_golden_model_1.TL1 [5]);
  nor (_31404_, _05444_, _31403_);
  nor (_31406_, _13203_, _11229_);
  nor (_31407_, _31406_, _31404_);
  nor (_31408_, _31407_, _06458_);
  and (_31409_, _13204_, _05350_);
  nor (_31410_, _31409_, _31404_);
  nor (_31411_, _31410_, _03745_);
  and (_31412_, _06757_, _05444_);
  or (_31413_, _31412_, _31404_);
  and (_31414_, _31413_, _04082_);
  and (_31415_, _05444_, \oc8051_golden_model_1.ACC [5]);
  nor (_31417_, _31415_, _31404_);
  nor (_31418_, _31417_, _03531_);
  nor (_31419_, _31417_, _04437_);
  nor (_31420_, _04436_, _31403_);
  or (_31421_, _31420_, _31419_);
  and (_31422_, _31421_, _04432_);
  nor (_31423_, _13070_, _11229_);
  nor (_31424_, _31423_, _31404_);
  nor (_31425_, _31424_, _04432_);
  or (_31426_, _31425_, _31422_);
  and (_31428_, _31426_, _04457_);
  nor (_31429_, _05526_, _11229_);
  nor (_31430_, _31429_, _31404_);
  nor (_31431_, _31430_, _04457_);
  nor (_31432_, _31431_, _31428_);
  nor (_31433_, _31432_, _03530_);
  or (_31434_, _31433_, _07454_);
  nor (_31435_, _31434_, _31418_);
  and (_31436_, _31430_, _07454_);
  or (_31437_, _31436_, _04082_);
  nor (_31439_, _31437_, _31435_);
  or (_31440_, _31439_, _31414_);
  and (_31441_, _31440_, _03521_);
  nor (_31442_, _13184_, _11229_);
  nor (_31443_, _31442_, _31404_);
  nor (_31444_, _31443_, _03521_);
  or (_31445_, _31444_, _08905_);
  or (_31446_, _31445_, _31441_);
  and (_31447_, _13198_, _05350_);
  or (_31448_, _31404_, _04527_);
  or (_31450_, _31448_, _31447_);
  and (_31451_, _06295_, _05444_);
  nor (_31452_, _31451_, _31404_);
  and (_31453_, _31452_, _03624_);
  nor (_31454_, _31453_, _03744_);
  and (_31455_, _31454_, _31450_);
  and (_31456_, _31455_, _31446_);
  nor (_31457_, _31456_, _31411_);
  nor (_31458_, _31457_, _03611_);
  nor (_31459_, _31404_, _05576_);
  not (_31461_, _31459_);
  nor (_31462_, _31452_, _04523_);
  and (_31463_, _31462_, _31461_);
  nor (_31464_, _31463_, _31458_);
  nor (_31465_, _31464_, _03733_);
  nor (_31466_, _31417_, _03734_);
  and (_31467_, _31466_, _31461_);
  nor (_31468_, _31467_, _03618_);
  not (_31469_, _31468_);
  nor (_31470_, _31469_, _31465_);
  or (_31472_, _13197_, _11229_);
  nor (_31473_, _31404_, _06453_);
  and (_31474_, _31473_, _31472_);
  or (_31475_, _31474_, _03741_);
  nor (_31476_, _31475_, _31470_);
  nor (_31477_, _31476_, _31408_);
  nor (_31478_, _31477_, _03767_);
  nor (_31479_, _31424_, _03948_);
  or (_31480_, _31479_, _03473_);
  nor (_31481_, _31480_, _31478_);
  nand (_31483_, _13253_, _05350_);
  nor (_31484_, _31404_, _03474_);
  and (_31485_, _31484_, _31483_);
  nor (_31486_, _31485_, _31481_);
  or (_31487_, _31486_, _43193_);
  or (_31488_, _43189_, \oc8051_golden_model_1.TL1 [5]);
  and (_31489_, _31488_, _42003_);
  and (_43907_, _31489_, _31487_);
  not (_31490_, \oc8051_golden_model_1.TL1 [6]);
  nor (_31491_, _05444_, _31490_);
  nor (_31493_, _13406_, _11229_);
  nor (_31494_, _31493_, _31491_);
  nor (_31495_, _31494_, _06458_);
  and (_31496_, _13407_, _05350_);
  nor (_31497_, _31496_, _31491_);
  nor (_31498_, _31497_, _03745_);
  and (_31499_, _06526_, _05444_);
  or (_31500_, _31499_, _31491_);
  and (_31501_, _31500_, _04082_);
  and (_31502_, _05444_, \oc8051_golden_model_1.ACC [6]);
  nor (_31504_, _31502_, _31491_);
  nor (_31505_, _31504_, _03531_);
  nor (_31506_, _31504_, _04437_);
  nor (_31507_, _04436_, _31490_);
  or (_31508_, _31507_, _31506_);
  and (_31509_, _31508_, _04432_);
  nor (_31510_, _13293_, _11229_);
  nor (_31511_, _31510_, _31491_);
  nor (_31512_, _31511_, _04432_);
  or (_31513_, _31512_, _31509_);
  and (_31515_, _31513_, _04457_);
  nor (_31516_, _05417_, _11229_);
  nor (_31517_, _31516_, _31491_);
  nor (_31518_, _31517_, _04457_);
  nor (_31519_, _31518_, _31515_);
  nor (_31520_, _31519_, _03530_);
  or (_31521_, _31520_, _07454_);
  nor (_31522_, _31521_, _31505_);
  and (_31523_, _31517_, _07454_);
  or (_31524_, _31523_, _04082_);
  nor (_31526_, _31524_, _31522_);
  or (_31527_, _31526_, _31501_);
  and (_31528_, _31527_, _03521_);
  nor (_31529_, _13387_, _11229_);
  nor (_31530_, _31529_, _31491_);
  nor (_31531_, _31530_, _03521_);
  or (_31532_, _31531_, _08905_);
  or (_31533_, _31532_, _31528_);
  and (_31534_, _13402_, _05350_);
  or (_31535_, _31491_, _04527_);
  or (_31537_, _31535_, _31534_);
  and (_31538_, _14949_, _05444_);
  nor (_31539_, _31538_, _31491_);
  and (_31540_, _31539_, _03624_);
  nor (_31541_, _31540_, _03744_);
  and (_31542_, _31541_, _31537_);
  and (_31543_, _31542_, _31533_);
  nor (_31544_, _31543_, _31498_);
  nor (_31545_, _31544_, _03611_);
  nor (_31546_, _31491_, _05469_);
  not (_31548_, _31546_);
  nor (_31549_, _31539_, _04523_);
  and (_31550_, _31549_, _31548_);
  nor (_31551_, _31550_, _31545_);
  nor (_31552_, _31551_, _03733_);
  nor (_31553_, _31504_, _03734_);
  and (_31554_, _31553_, _31548_);
  or (_31555_, _31554_, _31552_);
  and (_31556_, _31555_, _06453_);
  nor (_31557_, _13400_, _11263_);
  nor (_31559_, _31557_, _31491_);
  nor (_31560_, _31559_, _06453_);
  or (_31561_, _31560_, _31556_);
  and (_31562_, _31561_, _06458_);
  nor (_31563_, _31562_, _31495_);
  nor (_31564_, _31563_, _03767_);
  nor (_31565_, _31511_, _03948_);
  or (_31566_, _31565_, _03473_);
  nor (_31567_, _31566_, _31564_);
  nand (_31568_, _13456_, _05350_);
  nor (_31570_, _31491_, _03474_);
  and (_31571_, _31570_, _31568_);
  nor (_31572_, _31571_, _31567_);
  or (_31573_, _31572_, _43193_);
  or (_31574_, _43189_, \oc8051_golden_model_1.TL1 [6]);
  and (_31575_, _31574_, _42003_);
  and (_43909_, _31575_, _31573_);
  not (_31576_, \oc8051_golden_model_1.TMOD [0]);
  nor (_31577_, _05331_, _31576_);
  nor (_31578_, _05722_, _11311_);
  nor (_31580_, _31578_, _31577_);
  and (_31581_, _31580_, _17198_);
  and (_31582_, _05331_, \oc8051_golden_model_1.ACC [0]);
  nor (_31583_, _31582_, _31577_);
  nor (_31584_, _31583_, _03531_);
  nor (_31585_, _31583_, _04437_);
  nor (_31586_, _04436_, _31576_);
  or (_31587_, _31586_, _31585_);
  and (_31588_, _31587_, _04432_);
  nor (_31589_, _31580_, _04432_);
  or (_31591_, _31589_, _31588_);
  and (_31592_, _31591_, _04457_);
  and (_31593_, _05331_, _04429_);
  nor (_31594_, _31593_, _31577_);
  nor (_31595_, _31594_, _04457_);
  nor (_31596_, _31595_, _31592_);
  nor (_31597_, _31596_, _03530_);
  or (_31598_, _31597_, _07454_);
  nor (_31599_, _31598_, _31584_);
  and (_31600_, _31594_, _07454_);
  nor (_31602_, _31600_, _31599_);
  nor (_31603_, _31602_, _04082_);
  and (_31604_, _06617_, _05331_);
  nor (_31605_, _31577_, _04500_);
  not (_31606_, _31605_);
  nor (_31607_, _31606_, _31604_);
  nor (_31608_, _31607_, _31603_);
  nor (_31609_, _31608_, _03224_);
  nor (_31610_, _12164_, _11311_);
  or (_31611_, _31577_, _03521_);
  nor (_31613_, _31611_, _31610_);
  or (_31614_, _31613_, _03624_);
  nor (_31615_, _31614_, _31609_);
  and (_31616_, _05331_, _06350_);
  nor (_31617_, _31616_, _31577_);
  nor (_31618_, _31617_, _04509_);
  or (_31619_, _31618_, _31615_);
  and (_31620_, _31619_, _04527_);
  and (_31621_, _12177_, _05331_);
  nor (_31622_, _31621_, _31577_);
  nor (_31624_, _31622_, _04527_);
  or (_31625_, _31624_, _31620_);
  nor (_31626_, _31625_, _03744_);
  and (_31627_, _12183_, _05331_);
  or (_31628_, _31577_, _03745_);
  nor (_31629_, _31628_, _31627_);
  or (_31630_, _31629_, _03611_);
  nor (_31631_, _31630_, _31626_);
  or (_31632_, _31617_, _04523_);
  nor (_31633_, _31632_, _31578_);
  nor (_31634_, _31633_, _31631_);
  nor (_31635_, _31634_, _03733_);
  and (_31636_, _12182_, _05331_);
  or (_31637_, _31636_, _31577_);
  and (_31638_, _31637_, _03733_);
  or (_31639_, _31638_, _31635_);
  and (_31640_, _31639_, _06453_);
  nor (_31641_, _12057_, _11311_);
  nor (_31642_, _31641_, _31577_);
  nor (_31643_, _31642_, _06453_);
  or (_31645_, _31643_, _31640_);
  and (_31646_, _31645_, _06458_);
  nor (_31647_, _12181_, _11311_);
  nor (_31648_, _31647_, _31577_);
  nor (_31649_, _31648_, _06458_);
  nor (_31650_, _31649_, _17198_);
  not (_31651_, _31650_);
  nor (_31652_, _31651_, _31646_);
  nor (_31653_, _31652_, _31581_);
  or (_31654_, _31653_, _43193_);
  or (_31656_, _43189_, \oc8051_golden_model_1.TMOD [0]);
  and (_31657_, _31656_, _42003_);
  and (_43910_, _31657_, _31654_);
  and (_31658_, _06572_, _05331_);
  not (_31659_, \oc8051_golden_model_1.TMOD [1]);
  nor (_31660_, _05331_, _31659_);
  nor (_31661_, _31660_, _04500_);
  not (_31662_, _31661_);
  nor (_31663_, _31662_, _31658_);
  not (_31664_, _31663_);
  nor (_31666_, _11311_, _04635_);
  nor (_31667_, _31666_, _31660_);
  and (_31668_, _31667_, _07454_);
  nor (_31669_, _05331_, \oc8051_golden_model_1.TMOD [1]);
  and (_31670_, _05331_, _03269_);
  nor (_31671_, _31670_, _31669_);
  and (_31672_, _31671_, _03530_);
  and (_31673_, _31671_, _04436_);
  nor (_31674_, _04436_, _31659_);
  or (_31675_, _31674_, _31673_);
  and (_31677_, _31675_, _04432_);
  and (_31678_, _12265_, _05331_);
  nor (_31679_, _31678_, _31669_);
  and (_31680_, _31679_, _03534_);
  or (_31681_, _31680_, _31677_);
  and (_31682_, _31681_, _04457_);
  nor (_31683_, _31667_, _04457_);
  nor (_31684_, _31683_, _31682_);
  nor (_31685_, _31684_, _03530_);
  or (_31686_, _31685_, _07454_);
  nor (_31687_, _31686_, _31672_);
  nor (_31688_, _31687_, _31668_);
  nor (_31689_, _31688_, _04082_);
  nor (_31690_, _31689_, _03224_);
  and (_31691_, _31690_, _31664_);
  not (_31692_, _31669_);
  and (_31693_, _12360_, _05331_);
  nor (_31694_, _31693_, _03521_);
  and (_31695_, _31694_, _31692_);
  nor (_31696_, _31695_, _31691_);
  nor (_31699_, _31696_, _08905_);
  nor (_31700_, _12375_, _11311_);
  nor (_31701_, _31700_, _04527_);
  and (_31702_, _05331_, _04325_);
  nor (_31703_, _31702_, _04509_);
  nor (_31704_, _31703_, _31701_);
  nor (_31705_, _31704_, _31669_);
  nor (_31706_, _31705_, _31699_);
  nor (_31707_, _31706_, _03744_);
  nor (_31708_, _12381_, _11311_);
  nor (_31710_, _31708_, _03745_);
  and (_31711_, _31710_, _31692_);
  nor (_31712_, _31711_, _31707_);
  nor (_31713_, _31712_, _03611_);
  nor (_31714_, _12374_, _11311_);
  nor (_31715_, _31714_, _04523_);
  and (_31716_, _31715_, _31692_);
  nor (_31717_, _31716_, _31713_);
  nor (_31718_, _31717_, _03733_);
  nor (_31719_, _31660_, _05674_);
  nor (_31721_, _31719_, _03734_);
  and (_31722_, _31721_, _31671_);
  nor (_31723_, _31722_, _31718_);
  or (_31724_, _31723_, _18526_);
  and (_31725_, _31702_, _05673_);
  nor (_31726_, _31725_, _06453_);
  and (_31727_, _31726_, _31692_);
  nand (_31728_, _31670_, _05673_);
  nor (_31729_, _31669_, _06458_);
  and (_31730_, _31729_, _31728_);
  or (_31732_, _31730_, _03767_);
  nor (_31733_, _31732_, _31727_);
  and (_31734_, _31733_, _31724_);
  nor (_31735_, _31679_, _03948_);
  nor (_31736_, _31735_, _31734_);
  and (_31737_, _31736_, _03474_);
  nor (_31738_, _31678_, _31660_);
  nor (_31739_, _31738_, _03474_);
  or (_31740_, _31739_, _31737_);
  or (_31741_, _31740_, _43193_);
  or (_31743_, _43189_, \oc8051_golden_model_1.TMOD [1]);
  and (_31744_, _31743_, _42003_);
  and (_43911_, _31744_, _31741_);
  not (_31745_, \oc8051_golden_model_1.TMOD [2]);
  nor (_31746_, _05331_, _31745_);
  nor (_31747_, _12587_, _11311_);
  nor (_31748_, _31747_, _31746_);
  nor (_31749_, _31748_, _06458_);
  and (_31750_, _12588_, _05331_);
  nor (_31751_, _31750_, _31746_);
  nor (_31753_, _31751_, _03745_);
  nor (_31754_, _11311_, _05073_);
  nor (_31755_, _31754_, _31746_);
  and (_31756_, _31755_, _07454_);
  and (_31757_, _05331_, \oc8051_golden_model_1.ACC [2]);
  nor (_31758_, _31757_, _31746_);
  nor (_31759_, _31758_, _03531_);
  nor (_31760_, _31758_, _04437_);
  nor (_31761_, _04436_, _31745_);
  or (_31762_, _31761_, _31760_);
  and (_31764_, _31762_, _04432_);
  nor (_31765_, _12467_, _11311_);
  nor (_31766_, _31765_, _31746_);
  nor (_31767_, _31766_, _04432_);
  or (_31768_, _31767_, _31764_);
  and (_31769_, _31768_, _04457_);
  nor (_31770_, _31755_, _04457_);
  nor (_31771_, _31770_, _31769_);
  nor (_31772_, _31771_, _03530_);
  or (_31773_, _31772_, _07454_);
  nor (_31775_, _31773_, _31759_);
  nor (_31776_, _31775_, _31756_);
  nor (_31777_, _31776_, _04082_);
  and (_31778_, _06710_, _05331_);
  nor (_31779_, _31746_, _04500_);
  not (_31780_, _31779_);
  nor (_31781_, _31780_, _31778_);
  nor (_31782_, _31781_, _03224_);
  not (_31783_, _31782_);
  nor (_31784_, _31783_, _31777_);
  nor (_31786_, _12568_, _11311_);
  nor (_31787_, _31786_, _31746_);
  nor (_31788_, _31787_, _03521_);
  or (_31789_, _31788_, _08905_);
  or (_31790_, _31789_, _31784_);
  and (_31791_, _12582_, _05331_);
  or (_31792_, _31746_, _04527_);
  or (_31793_, _31792_, _31791_);
  and (_31794_, _05331_, _06399_);
  nor (_31795_, _31794_, _31746_);
  and (_31797_, _31795_, _03624_);
  nor (_31798_, _31797_, _03744_);
  and (_31799_, _31798_, _31793_);
  and (_31800_, _31799_, _31790_);
  nor (_31801_, _31800_, _31753_);
  nor (_31802_, _31801_, _03611_);
  nor (_31803_, _31746_, _05772_);
  not (_31804_, _31803_);
  nor (_31805_, _31795_, _04523_);
  and (_31806_, _31805_, _31804_);
  nor (_31808_, _31806_, _31802_);
  nor (_31809_, _31808_, _03733_);
  nor (_31810_, _31758_, _03734_);
  and (_31811_, _31810_, _31804_);
  nor (_31812_, _31811_, _03618_);
  not (_31813_, _31812_);
  nor (_31814_, _31813_, _31809_);
  nor (_31815_, _12581_, _11311_);
  or (_31816_, _31746_, _06453_);
  nor (_31817_, _31816_, _31815_);
  or (_31819_, _31817_, _03741_);
  nor (_31820_, _31819_, _31814_);
  nor (_31821_, _31820_, _31749_);
  nor (_31822_, _31821_, _03767_);
  nor (_31823_, _31766_, _03948_);
  or (_31824_, _31823_, _03473_);
  nor (_31825_, _31824_, _31822_);
  and (_31826_, _12638_, _05331_);
  or (_31827_, _31746_, _03474_);
  nor (_31828_, _31827_, _31826_);
  nor (_31830_, _31828_, _31825_);
  or (_31831_, _31830_, _43193_);
  or (_31832_, _43189_, \oc8051_golden_model_1.TMOD [2]);
  and (_31833_, _31832_, _42003_);
  and (_43914_, _31833_, _31831_);
  not (_31834_, \oc8051_golden_model_1.TMOD [3]);
  nor (_31835_, _05331_, _31834_);
  nor (_31836_, _12792_, _11311_);
  nor (_31837_, _31836_, _31835_);
  nor (_31838_, _31837_, _06458_);
  and (_31840_, _12793_, _05331_);
  nor (_31841_, _31840_, _31835_);
  nor (_31842_, _31841_, _03745_);
  and (_31843_, _06664_, _05331_);
  or (_31844_, _31843_, _31835_);
  and (_31845_, _31844_, _04082_);
  and (_31846_, _05331_, \oc8051_golden_model_1.ACC [3]);
  nor (_31847_, _31846_, _31835_);
  nor (_31848_, _31847_, _03531_);
  nor (_31849_, _31847_, _04437_);
  nor (_31851_, _04436_, _31834_);
  or (_31852_, _31851_, _31849_);
  and (_31853_, _31852_, _04432_);
  nor (_31854_, _12652_, _11311_);
  nor (_31855_, _31854_, _31835_);
  nor (_31856_, _31855_, _04432_);
  or (_31857_, _31856_, _31853_);
  and (_31858_, _31857_, _04457_);
  nor (_31859_, _11311_, _04885_);
  nor (_31860_, _31859_, _31835_);
  nor (_31862_, _31860_, _04457_);
  nor (_31863_, _31862_, _31858_);
  nor (_31864_, _31863_, _03530_);
  or (_31865_, _31864_, _07454_);
  nor (_31866_, _31865_, _31848_);
  and (_31867_, _31860_, _07454_);
  or (_31868_, _31867_, _04082_);
  nor (_31869_, _31868_, _31866_);
  or (_31870_, _31869_, _31845_);
  and (_31871_, _31870_, _03521_);
  nor (_31873_, _12773_, _11311_);
  nor (_31874_, _31873_, _31835_);
  nor (_31875_, _31874_, _03521_);
  or (_31876_, _31875_, _08905_);
  or (_31877_, _31876_, _31871_);
  and (_31878_, _12787_, _05331_);
  or (_31879_, _31835_, _04527_);
  or (_31880_, _31879_, _31878_);
  and (_31881_, _05331_, _06356_);
  nor (_31882_, _31881_, _31835_);
  and (_31884_, _31882_, _03624_);
  nor (_31885_, _31884_, _03744_);
  and (_31886_, _31885_, _31880_);
  and (_31887_, _31886_, _31877_);
  nor (_31888_, _31887_, _31842_);
  nor (_31889_, _31888_, _03611_);
  nor (_31890_, _31835_, _05625_);
  not (_31891_, _31890_);
  nor (_31892_, _31882_, _04523_);
  and (_31893_, _31892_, _31891_);
  nor (_31895_, _31893_, _31889_);
  nor (_31896_, _31895_, _03733_);
  nor (_31897_, _31847_, _03734_);
  and (_31898_, _31897_, _31891_);
  or (_31899_, _31898_, _31896_);
  and (_31900_, _31899_, _06453_);
  nor (_31901_, _12786_, _11311_);
  nor (_31902_, _31901_, _31835_);
  nor (_31903_, _31902_, _06453_);
  or (_31904_, _31903_, _31900_);
  and (_31906_, _31904_, _06458_);
  nor (_31907_, _31906_, _31838_);
  nor (_31908_, _31907_, _03767_);
  nor (_31909_, _31855_, _03948_);
  or (_31910_, _31909_, _03473_);
  nor (_31911_, _31910_, _31908_);
  and (_31912_, _12843_, _05331_);
  or (_31913_, _31835_, _03474_);
  nor (_31914_, _31913_, _31912_);
  nor (_31915_, _31914_, _31911_);
  or (_31917_, _31915_, _43193_);
  or (_31918_, _43189_, \oc8051_golden_model_1.TMOD [3]);
  and (_31919_, _31918_, _42003_);
  and (_43915_, _31919_, _31917_);
  not (_31920_, \oc8051_golden_model_1.TMOD [4]);
  nor (_31921_, _05331_, _31920_);
  nor (_31922_, _12991_, _11311_);
  nor (_31923_, _31922_, _31921_);
  nor (_31924_, _31923_, _06458_);
  and (_31925_, _12992_, _05331_);
  nor (_31927_, _31925_, _31921_);
  nor (_31928_, _31927_, _03745_);
  and (_31929_, _06337_, _05331_);
  nor (_31930_, _31929_, _31921_);
  and (_31931_, _31930_, _03624_);
  and (_31932_, _05331_, \oc8051_golden_model_1.ACC [4]);
  nor (_31933_, _31932_, _31921_);
  nor (_31934_, _31933_, _03531_);
  nor (_31935_, _31933_, _04437_);
  nor (_31936_, _04436_, _31920_);
  or (_31938_, _31936_, _31935_);
  and (_31939_, _31938_, _04432_);
  nor (_31940_, _12856_, _11311_);
  nor (_31941_, _31940_, _31921_);
  nor (_31942_, _31941_, _04432_);
  or (_31943_, _31942_, _31939_);
  and (_31944_, _31943_, _04457_);
  nor (_31945_, _05831_, _11311_);
  nor (_31946_, _31945_, _31921_);
  nor (_31947_, _31946_, _04457_);
  nor (_31949_, _31947_, _31944_);
  nor (_31950_, _31949_, _03530_);
  or (_31951_, _31950_, _07454_);
  nor (_31952_, _31951_, _31934_);
  and (_31953_, _31946_, _07454_);
  nor (_31954_, _31953_, _31952_);
  nor (_31955_, _31954_, _04082_);
  and (_31956_, _06802_, _05331_);
  nor (_31957_, _31921_, _04500_);
  not (_31958_, _31957_);
  nor (_31960_, _31958_, _31956_);
  or (_31961_, _31960_, _03224_);
  nor (_31962_, _31961_, _31955_);
  nor (_31963_, _12972_, _11311_);
  nor (_31964_, _31963_, _31921_);
  nor (_31965_, _31964_, _03521_);
  or (_31966_, _31965_, _03624_);
  nor (_31967_, _31966_, _31962_);
  nor (_31968_, _31967_, _31931_);
  or (_31969_, _31968_, _03623_);
  and (_31971_, _12986_, _05331_);
  or (_31972_, _31971_, _31921_);
  or (_31973_, _31972_, _04527_);
  and (_31974_, _31973_, _03745_);
  and (_31975_, _31974_, _31969_);
  nor (_31976_, _31975_, _31928_);
  nor (_31977_, _31976_, _03611_);
  nor (_31978_, _31921_, _05880_);
  not (_31979_, _31978_);
  nor (_31980_, _31930_, _04523_);
  and (_31982_, _31980_, _31979_);
  nor (_31983_, _31982_, _31977_);
  nor (_31984_, _31983_, _03733_);
  nor (_31985_, _31933_, _03734_);
  and (_31986_, _31985_, _31979_);
  nor (_31987_, _31986_, _03618_);
  not (_31988_, _31987_);
  nor (_31989_, _31988_, _31984_);
  nor (_31990_, _12985_, _11311_);
  or (_31991_, _31921_, _06453_);
  nor (_31993_, _31991_, _31990_);
  or (_31994_, _31993_, _03741_);
  nor (_31995_, _31994_, _31989_);
  nor (_31996_, _31995_, _31924_);
  nor (_31997_, _31996_, _03767_);
  nor (_31998_, _31941_, _03948_);
  or (_31999_, _31998_, _03473_);
  nor (_32000_, _31999_, _31997_);
  and (_32001_, _13051_, _05331_);
  or (_32002_, _31921_, _03474_);
  nor (_32004_, _32002_, _32001_);
  nor (_32005_, _32004_, _32000_);
  or (_32006_, _32005_, _43193_);
  or (_32007_, _43189_, \oc8051_golden_model_1.TMOD [4]);
  and (_32008_, _32007_, _42003_);
  and (_43916_, _32008_, _32006_);
  not (_32009_, \oc8051_golden_model_1.TMOD [5]);
  nor (_32010_, _05331_, _32009_);
  nor (_32011_, _13203_, _11311_);
  nor (_32012_, _32011_, _32010_);
  nor (_32014_, _32012_, _06458_);
  and (_32015_, _13204_, _05331_);
  nor (_32016_, _32015_, _32010_);
  nor (_32017_, _32016_, _03745_);
  and (_32018_, _06757_, _05331_);
  or (_32019_, _32018_, _32010_);
  and (_32020_, _32019_, _04082_);
  and (_32021_, _05331_, \oc8051_golden_model_1.ACC [5]);
  nor (_32022_, _32021_, _32010_);
  nor (_32023_, _32022_, _03531_);
  nor (_32025_, _32022_, _04437_);
  nor (_32026_, _04436_, _32009_);
  or (_32027_, _32026_, _32025_);
  and (_32028_, _32027_, _04432_);
  nor (_32029_, _13070_, _11311_);
  nor (_32030_, _32029_, _32010_);
  nor (_32031_, _32030_, _04432_);
  or (_32032_, _32031_, _32028_);
  and (_32033_, _32032_, _04457_);
  nor (_32034_, _05526_, _11311_);
  nor (_32036_, _32034_, _32010_);
  nor (_32037_, _32036_, _04457_);
  nor (_32038_, _32037_, _32033_);
  nor (_32039_, _32038_, _03530_);
  or (_32040_, _32039_, _07454_);
  nor (_32041_, _32040_, _32023_);
  and (_32042_, _32036_, _07454_);
  or (_32043_, _32042_, _04082_);
  nor (_32044_, _32043_, _32041_);
  or (_32045_, _32044_, _32020_);
  and (_32047_, _32045_, _03521_);
  nor (_32048_, _13184_, _11311_);
  nor (_32049_, _32048_, _32010_);
  nor (_32050_, _32049_, _03521_);
  or (_32051_, _32050_, _08905_);
  or (_32052_, _32051_, _32047_);
  and (_32053_, _13198_, _05331_);
  or (_32054_, _32010_, _04527_);
  or (_32055_, _32054_, _32053_);
  and (_32056_, _06295_, _05331_);
  nor (_32058_, _32056_, _32010_);
  and (_32059_, _32058_, _03624_);
  nor (_32060_, _32059_, _03744_);
  and (_32061_, _32060_, _32055_);
  and (_32062_, _32061_, _32052_);
  nor (_32063_, _32062_, _32017_);
  nor (_32064_, _32063_, _03611_);
  nor (_32065_, _32010_, _05576_);
  not (_32066_, _32065_);
  nor (_32067_, _32058_, _04523_);
  and (_32069_, _32067_, _32066_);
  nor (_32070_, _32069_, _32064_);
  nor (_32071_, _32070_, _03733_);
  nor (_32072_, _32022_, _03734_);
  and (_32073_, _32072_, _32066_);
  or (_32074_, _32073_, _32071_);
  and (_32075_, _32074_, _06453_);
  nor (_32076_, _13197_, _11311_);
  nor (_32077_, _32076_, _32010_);
  nor (_32078_, _32077_, _06453_);
  or (_32080_, _32078_, _32075_);
  and (_32081_, _32080_, _06458_);
  nor (_32082_, _32081_, _32014_);
  nor (_32083_, _32082_, _03767_);
  nor (_32084_, _32030_, _03948_);
  or (_32085_, _32084_, _03473_);
  nor (_32086_, _32085_, _32083_);
  and (_32087_, _13253_, _05331_);
  or (_32088_, _32010_, _03474_);
  nor (_32089_, _32088_, _32087_);
  nor (_32091_, _32089_, _32086_);
  or (_32092_, _32091_, _43193_);
  or (_32093_, _43189_, \oc8051_golden_model_1.TMOD [5]);
  and (_32094_, _32093_, _42003_);
  and (_43917_, _32094_, _32092_);
  not (_32095_, \oc8051_golden_model_1.TMOD [6]);
  nor (_32096_, _05331_, _32095_);
  nor (_32097_, _13406_, _11311_);
  nor (_32098_, _32097_, _32096_);
  nor (_32099_, _32098_, _06458_);
  and (_32101_, _13407_, _05331_);
  nor (_32102_, _32101_, _32096_);
  nor (_32103_, _32102_, _03745_);
  and (_32104_, _06526_, _05331_);
  or (_32105_, _32104_, _32096_);
  and (_32106_, _32105_, _04082_);
  and (_32107_, _05331_, \oc8051_golden_model_1.ACC [6]);
  nor (_32108_, _32107_, _32096_);
  nor (_32109_, _32108_, _03531_);
  nor (_32110_, _32108_, _04437_);
  nor (_32112_, _04436_, _32095_);
  or (_32113_, _32112_, _32110_);
  and (_32114_, _32113_, _04432_);
  nor (_32115_, _13293_, _11311_);
  nor (_32116_, _32115_, _32096_);
  nor (_32117_, _32116_, _04432_);
  or (_32118_, _32117_, _32114_);
  and (_32119_, _32118_, _04457_);
  nor (_32120_, _05417_, _11311_);
  nor (_32121_, _32120_, _32096_);
  nor (_32123_, _32121_, _04457_);
  nor (_32124_, _32123_, _32119_);
  nor (_32125_, _32124_, _03530_);
  or (_32126_, _32125_, _07454_);
  nor (_32127_, _32126_, _32109_);
  and (_32128_, _32121_, _07454_);
  or (_32129_, _32128_, _04082_);
  nor (_32130_, _32129_, _32127_);
  or (_32131_, _32130_, _32106_);
  and (_32132_, _32131_, _03521_);
  nor (_32134_, _13387_, _11311_);
  nor (_32135_, _32134_, _32096_);
  nor (_32136_, _32135_, _03521_);
  or (_32137_, _32136_, _08905_);
  or (_32138_, _32137_, _32132_);
  and (_32139_, _13402_, _05331_);
  or (_32140_, _32096_, _04527_);
  or (_32141_, _32140_, _32139_);
  and (_32142_, _14949_, _05331_);
  nor (_32143_, _32142_, _32096_);
  and (_32145_, _32143_, _03624_);
  nor (_32146_, _32145_, _03744_);
  and (_32147_, _32146_, _32141_);
  and (_32148_, _32147_, _32138_);
  nor (_32149_, _32148_, _32103_);
  nor (_32150_, _32149_, _03611_);
  nor (_32151_, _32096_, _05469_);
  not (_32152_, _32151_);
  nor (_32153_, _32143_, _04523_);
  and (_32154_, _32153_, _32152_);
  nor (_32156_, _32154_, _32150_);
  nor (_32157_, _32156_, _03733_);
  nor (_32158_, _32108_, _03734_);
  and (_32159_, _32158_, _32152_);
  or (_32160_, _32159_, _32157_);
  and (_32161_, _32160_, _06453_);
  nor (_32162_, _13400_, _11311_);
  nor (_32163_, _32162_, _32096_);
  nor (_32164_, _32163_, _06453_);
  or (_32165_, _32164_, _32161_);
  and (_32167_, _32165_, _06458_);
  nor (_32168_, _32167_, _32099_);
  nor (_32169_, _32168_, _03767_);
  nor (_32170_, _32116_, _03948_);
  or (_32171_, _32170_, _03473_);
  nor (_32172_, _32171_, _32169_);
  and (_32173_, _13456_, _05331_);
  or (_32174_, _32096_, _03474_);
  nor (_32175_, _32174_, _32173_);
  nor (_32176_, _32175_, _32172_);
  or (_32178_, _32176_, _43193_);
  or (_32179_, _43189_, \oc8051_golden_model_1.TMOD [6]);
  and (_32180_, _32179_, _42003_);
  and (_43918_, _32180_, _32178_);
  not (_32181_, _24605_);
  and (_32182_, _32181_, _04118_);
  and (_32183_, _11991_, _11998_);
  nor (_32184_, _32183_, _02897_);
  and (_32185_, _11406_, _08816_);
  nor (_32186_, _32185_, _02897_);
  nor (_32188_, _07983_, _02897_);
  and (_32189_, _07983_, _02897_);
  nor (_32190_, _32189_, _32188_);
  nor (_32191_, _32190_, _11942_);
  not (_32192_, _03178_);
  and (_32193_, _11413_, _06453_);
  nor (_32194_, _32193_, _02897_);
  not (_32195_, _03182_);
  nor (_32196_, _11901_, _03611_);
  nor (_32197_, _32196_, _02897_);
  not (_32199_, _03172_);
  and (_32200_, _11416_, _04527_);
  nor (_32201_, _32200_, _02897_);
  and (_32202_, _03624_, _02897_);
  nor (_32203_, _04118_, _03214_);
  nor (_32204_, _11424_, _02897_);
  nor (_32205_, _04118_, _03207_);
  and (_32206_, _10163_, \oc8051_golden_model_1.PC [0]);
  and (_32207_, _10122_, _02897_);
  and (_32208_, _04118_, \oc8051_golden_model_1.PC [0]);
  nor (_32210_, _32208_, _11507_);
  nor (_32211_, _32210_, _10163_);
  nor (_32212_, _32211_, _10158_);
  nor (_32213_, _32212_, _32207_);
  nor (_32214_, _32213_, _32206_);
  nor (_32215_, _04118_, _03212_);
  and (_32216_, _03209_, _03204_);
  nor (_32217_, _32216_, _04118_);
  nor (_32218_, _11687_, _02897_);
  nor (_32219_, _32218_, _11677_);
  nor (_32221_, _11683_, _02897_);
  and (_32222_, _11683_, _02897_);
  nor (_32223_, _32222_, _32221_);
  and (_32224_, _32223_, _03204_);
  not (_32225_, _32224_);
  nand (_32226_, _32225_, _11687_);
  and (_32227_, _32226_, _32219_);
  or (_32228_, _32227_, _05998_);
  nor (_32229_, _32228_, _32217_);
  and (_32230_, _11566_, \oc8051_golden_model_1.PC [0]);
  nand (_32232_, _11565_, _11563_);
  and (_32233_, _03989_, _02897_);
  nor (_32234_, _32233_, _11621_);
  and (_32235_, _32234_, _32232_);
  or (_32236_, _32235_, _32230_);
  nor (_32237_, _32236_, _05997_);
  nor (_32238_, _32237_, _32229_);
  nor (_32239_, _32238_, _04012_);
  and (_32240_, _04012_, \oc8051_golden_model_1.PC [0]);
  nor (_32241_, _32240_, _03534_);
  not (_32243_, _32241_);
  nor (_32244_, _32243_, _32239_);
  not (_32245_, _32244_);
  not (_32246_, _32210_);
  and (_32247_, _32246_, _11439_);
  and (_32248_, _05722_, _05624_);
  and (_32249_, _32248_, _11436_);
  nand (_32250_, _32249_, _12464_);
  nor (_32251_, _32250_, _02897_);
  or (_32252_, _32251_, _04432_);
  or (_32254_, _32252_, _32247_);
  and (_32255_, _32254_, _11430_);
  and (_32256_, _32255_, _32245_);
  nor (_32257_, _11430_, _02897_);
  nor (_32258_, _32257_, _05977_);
  not (_32259_, _32258_);
  nor (_32260_, _32259_, _32256_);
  nor (_32261_, _04118_, _03202_);
  and (_32262_, _11723_, _11715_);
  not (_32263_, _32262_);
  nor (_32265_, _32263_, _32261_);
  not (_32266_, _32265_);
  nor (_32267_, _32266_, _32260_);
  nor (_32268_, _32262_, _02897_);
  nor (_32269_, _32268_, _11727_);
  not (_32270_, _32269_);
  nor (_32271_, _32270_, _32267_);
  nor (_32272_, _32271_, _32215_);
  nor (_32273_, _32272_, _10021_);
  and (_32274_, _10055_, \oc8051_golden_model_1.PC [0]);
  nor (_32276_, _32210_, _10055_);
  or (_32277_, _32276_, _10017_);
  nor (_32278_, _32277_, _32274_);
  or (_32279_, _32278_, _10020_);
  nor (_32280_, _32279_, _32273_);
  and (_32281_, _10116_, _02897_);
  and (_32282_, _32210_, _11743_);
  nor (_32283_, _32282_, _32281_);
  and (_32284_, _32283_, _10020_);
  nor (_32285_, _32284_, _32280_);
  and (_32287_, _32285_, _03994_);
  nor (_32288_, _32246_, _09975_);
  and (_32289_, _09975_, _02897_);
  nor (_32290_, _32289_, _32288_);
  nor (_32291_, _32290_, _03994_);
  nor (_32292_, _32291_, _32287_);
  nor (_32293_, _32292_, _10124_);
  nor (_32294_, _32293_, _32214_);
  nor (_32295_, _32294_, _04755_);
  or (_32296_, _32295_, _11425_);
  nor (_32298_, _32296_, _32205_);
  or (_32299_, _32298_, _11776_);
  nor (_32300_, _32299_, _32204_);
  and (_32301_, _11419_, _03233_);
  not (_32302_, _32301_);
  or (_32303_, _32302_, _32300_);
  nor (_32304_, _32303_, _32203_);
  nor (_32305_, _32301_, _02897_);
  nor (_32306_, _32305_, _03219_);
  not (_32307_, _32306_);
  nor (_32309_, _32307_, _32304_);
  nor (_32310_, _04118_, _05919_);
  nor (_32311_, _03621_, _03224_);
  and (_32312_, _32311_, _11806_);
  not (_32313_, _32312_);
  nor (_32314_, _32313_, _32310_);
  not (_32315_, _32314_);
  nor (_32316_, _32315_, _32309_);
  nor (_32317_, _32312_, _02897_);
  nor (_32318_, _32317_, _03159_);
  not (_32319_, _32318_);
  nor (_32320_, _32319_, _32316_);
  nor (_32321_, _04118_, _03160_);
  or (_32322_, _32321_, _11813_);
  nor (_32323_, _32322_, _32320_);
  nor (_32324_, _32234_, _11814_);
  nor (_32325_, _32324_, _32323_);
  and (_32326_, _32325_, _04509_);
  or (_32327_, _32326_, _32202_);
  and (_32328_, _32327_, _23814_);
  and (_32331_, _11828_, _03336_);
  or (_32332_, _32331_, _32328_);
  and (_32333_, _32332_, _27595_);
  nor (_32334_, _04118_, _27595_);
  or (_32335_, _32334_, _32333_);
  and (_32336_, _32335_, _23819_);
  not (_32337_, _32200_);
  and (_32338_, _08864_, \oc8051_golden_model_1.PC [0]);
  and (_32339_, _32234_, _11894_);
  or (_32340_, _32339_, _32338_);
  and (_32342_, _32340_, _11868_);
  nor (_32343_, _32342_, _32337_);
  not (_32344_, _32343_);
  nor (_32345_, _32344_, _32336_);
  nor (_32346_, _32345_, _32201_);
  and (_32347_, _32346_, _32199_);
  nor (_32348_, _04118_, _32199_);
  or (_32349_, _32348_, _32347_);
  and (_32350_, _32349_, _11893_);
  not (_32351_, _32196_);
  nor (_32353_, _32234_, _11894_);
  nor (_32354_, _08864_, \oc8051_golden_model_1.PC [0]);
  nor (_32355_, _32354_, _11893_);
  not (_32356_, _32355_);
  nor (_32357_, _32356_, _32353_);
  nor (_32358_, _32357_, _32351_);
  not (_32359_, _32358_);
  nor (_32360_, _32359_, _32350_);
  nor (_32361_, _32360_, _32197_);
  and (_32362_, _32361_, _32195_);
  nor (_32364_, _04118_, _32195_);
  or (_32365_, _32364_, _32362_);
  and (_32366_, _32365_, _24078_);
  not (_32367_, _32193_);
  and (_32368_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and (_32369_, _32234_, _07982_);
  or (_32370_, _32369_, _32368_);
  and (_32371_, _32370_, _11915_);
  nor (_32372_, _32371_, _32367_);
  not (_32373_, _32372_);
  nor (_32374_, _32373_, _32366_);
  nor (_32375_, _32374_, _32194_);
  and (_32376_, _32375_, _32192_);
  nor (_32377_, _04118_, _32192_);
  or (_32378_, _32377_, _32376_);
  and (_32379_, _32378_, _11942_);
  and (_32380_, _11408_, _08708_);
  not (_32381_, _32380_);
  or (_32382_, _32381_, _32379_);
  nor (_32383_, _32382_, _32191_);
  nor (_32385_, _32380_, _02897_);
  nor (_32386_, _32385_, _03752_);
  not (_32387_, _32386_);
  nor (_32388_, _32387_, _32383_);
  and (_32389_, _06617_, _03752_);
  or (_32390_, _32389_, _32388_);
  and (_32391_, _32390_, _04803_);
  nor (_32392_, _04118_, _04803_);
  or (_32393_, _32392_, _32391_);
  and (_32394_, _32393_, _03814_);
  and (_32396_, _32246_, _09953_);
  nor (_32397_, _09953_, _02897_);
  or (_32398_, _32397_, _03814_);
  or (_32399_, _32398_, _32396_);
  and (_32400_, _32399_, _32185_);
  not (_32401_, _32400_);
  nor (_32402_, _32401_, _32394_);
  nor (_32403_, _32402_, _32186_);
  and (_32404_, _32403_, _03476_);
  and (_32405_, _06617_, _03475_);
  or (_32407_, _32405_, _32404_);
  and (_32408_, _32407_, _11405_);
  nor (_32409_, _04118_, _11405_);
  nor (_32410_, _32409_, _32408_);
  nor (_32411_, _32410_, _03644_);
  not (_32412_, _32183_);
  and (_32413_, _09953_, \oc8051_golden_model_1.PC [0]);
  nor (_32414_, _32210_, _09953_);
  nor (_32415_, _32414_, _32413_);
  and (_32416_, _32415_, _03644_);
  nor (_32418_, _32416_, _32412_);
  not (_32419_, _32418_);
  nor (_32420_, _32419_, _32411_);
  nor (_32421_, _32420_, _32184_);
  nor (_32422_, _32421_, _04986_);
  and (_32423_, _04986_, _04118_);
  nor (_32424_, _32423_, _03445_);
  not (_32425_, _32424_);
  nor (_32426_, _32425_, _32422_);
  and (_32427_, _32415_, _03445_);
  and (_32429_, _12015_, _11392_);
  not (_32430_, _32429_);
  nor (_32431_, _32430_, _32427_);
  not (_32432_, _32431_);
  nor (_32433_, _32432_, _32426_);
  nor (_32434_, _32429_, _02897_);
  nor (_32435_, _32434_, _32433_);
  nor (_32436_, _32435_, _32181_);
  or (_32437_, _32436_, _12031_);
  nor (_32438_, _32437_, _32182_);
  and (_32440_, _12031_, _02897_);
  nor (_32441_, _32440_, _32438_);
  nand (_32442_, _32441_, _43189_);
  or (_32443_, _43189_, \oc8051_golden_model_1.PC [0]);
  and (_32444_, _32443_, _42003_);
  and (_43920_, _32444_, _32442_);
  and (_32445_, _03473_, _02860_);
  and (_32446_, _04736_, _06838_);
  nor (_32447_, _11998_, _03313_);
  and (_32448_, _07927_, _03270_);
  and (_32450_, _11901_, _03270_);
  nor (_32451_, _08493_, _02860_);
  nor (_32452_, _15828_, _03313_);
  nor (_32453_, _11723_, _03313_);
  or (_32454_, _32250_, _03313_);
  nor (_32455_, _11509_, _11507_);
  nor (_32456_, _32455_, _11510_);
  not (_32457_, _32456_);
  or (_32458_, _32457_, _11437_);
  and (_32459_, _32458_, _03534_);
  nand (_32461_, _32459_, _32454_);
  nor (_32462_, _11623_, _11621_);
  nor (_32463_, _32462_, _11624_);
  nand (_32464_, _32463_, _32232_);
  or (_32465_, _32232_, \oc8051_golden_model_1.PC [1]);
  and (_32466_, _32465_, _32464_);
  nand (_32467_, _32466_, _05998_);
  nor (_32468_, _05912_, _03208_);
  and (_32469_, _32468_, _03270_);
  nand (_32470_, _03443_, _03559_);
  and (_32472_, _32470_, _08105_);
  and (_32473_, _32472_, _03270_);
  nor (_32474_, _32221_, _04436_);
  and (_32475_, _32474_, _02860_);
  nor (_32476_, _32474_, _02860_);
  nor (_32477_, _32476_, _32475_);
  and (_32478_, _32477_, _03204_);
  nor (_32479_, _04325_, _03204_);
  or (_32480_, _32479_, _32472_);
  nor (_32481_, _32480_, _32478_);
  nor (_32483_, _32481_, _32473_);
  nor (_32484_, _32468_, _32483_);
  or (_32485_, _32484_, _03536_);
  nor (_32486_, _32485_, _32469_);
  and (_32487_, _03536_, _02860_);
  or (_32488_, _32487_, _32486_);
  and (_32489_, _32488_, _11686_);
  and (_32490_, _08118_, _03313_);
  or (_32491_, _32490_, _32489_);
  and (_32492_, _32491_, _03209_);
  nor (_32494_, _04325_, _03209_);
  nor (_32495_, _32494_, _05998_);
  not (_32496_, _32495_);
  nor (_32497_, _32496_, _32492_);
  nor (_32498_, _32497_, _04012_);
  nand (_32499_, _32498_, _32467_);
  and (_32500_, _04012_, _03313_);
  nor (_32501_, _32500_, _03534_);
  nand (_32502_, _32501_, _32499_);
  nand (_32503_, _32502_, _32461_);
  nand (_32505_, _32503_, _11430_);
  nor (_32506_, _11430_, _03313_);
  nor (_32507_, _32506_, _03469_);
  nand (_32508_, _32507_, _32505_);
  and (_32509_, _03469_, _02860_);
  nor (_32510_, _32509_, _05977_);
  nand (_32511_, _32510_, _32508_);
  and (_32512_, _04325_, _05977_);
  nor (_32513_, _32512_, _03527_);
  nand (_32514_, _32513_, _32511_);
  and (_32516_, _03527_, _02860_);
  nor (_32517_, _32516_, _11716_);
  nand (_32518_, _32517_, _32514_);
  nor (_32519_, _11715_, _03313_);
  nor (_32520_, _32519_, _03530_);
  nand (_32521_, _32520_, _32518_);
  and (_32522_, _03530_, _02860_);
  nor (_32523_, _32522_, _11724_);
  and (_32524_, _32523_, _32521_);
  or (_32525_, _32524_, _32453_);
  nand (_32527_, _32525_, _03466_);
  and (_32528_, _03465_, \oc8051_golden_model_1.PC [1]);
  nor (_32529_, _32528_, _11727_);
  and (_32530_, _32529_, _32527_);
  nor (_32531_, _04325_, _03212_);
  or (_32532_, _32531_, _32530_);
  nand (_32533_, _32532_, _04577_);
  and (_32534_, _03464_, _02860_);
  nor (_32535_, _32534_, _10021_);
  and (_32536_, _32535_, _32533_);
  and (_32538_, _10055_, _03270_);
  nor (_32539_, _32457_, _10055_);
  or (_32540_, _32539_, _32538_);
  nor (_32541_, _32540_, _10017_);
  or (_32542_, _32541_, _32536_);
  nand (_32543_, _32542_, _10112_);
  or (_32544_, _11743_, _03313_);
  or (_32545_, _32457_, _10116_);
  and (_32546_, _32545_, _10020_);
  nand (_32547_, _32546_, _32544_);
  and (_32549_, _32547_, _03994_);
  nand (_32550_, _32549_, _32543_);
  and (_32551_, _09975_, _03313_);
  nor (_32552_, _32456_, _09975_);
  or (_32553_, _32552_, _03994_);
  or (_32554_, _32553_, _32551_);
  nand (_32555_, _32554_, _32550_);
  nand (_32556_, _32555_, _10123_);
  and (_32557_, _10122_, _03313_);
  nand (_32558_, _10163_, _03313_);
  or (_32560_, _32456_, _10163_);
  and (_32561_, _32560_, _03608_);
  and (_32562_, _32561_, _32558_);
  nor (_32563_, _32562_, _32557_);
  and (_32564_, _32563_, _03459_);
  nand (_32565_, _32564_, _32556_);
  and (_32566_, _03458_, \oc8051_golden_model_1.PC [1]);
  nor (_32567_, _32566_, _04755_);
  nand (_32568_, _32567_, _32565_);
  nor (_32569_, _04325_, _03207_);
  not (_32571_, _05107_);
  and (_32572_, _03571_, _03558_);
  nor (_32573_, _32572_, _03522_);
  nor (_32574_, _04683_, _04481_);
  and (_32575_, _32574_, _32573_);
  and (_32576_, _32575_, _32571_);
  not (_32577_, _32576_);
  nor (_32578_, _32577_, _32569_);
  nand (_32579_, _32578_, _32568_);
  nor (_32580_, _32576_, _02860_);
  nor (_32582_, _32580_, _11421_);
  nand (_32583_, _32582_, _32579_);
  and (_32584_, _11423_, _03270_);
  or (_32585_, _32584_, _11424_);
  nand (_32586_, _32585_, _32583_);
  nor (_32587_, _11423_, _03313_);
  nor (_32588_, _32587_, _03587_);
  nand (_32589_, _32588_, _32586_);
  and (_32590_, _03587_, _02860_);
  nor (_32591_, _32590_, _11776_);
  nand (_32593_, _32591_, _32589_);
  and (_32594_, _04325_, _11776_);
  nor (_32595_, _32594_, _03586_);
  and (_32596_, _32595_, _32593_);
  and (_32597_, _03586_, _02860_);
  or (_32598_, _32597_, _32596_);
  nand (_32599_, _32598_, _11419_);
  nor (_32600_, _11419_, _03270_);
  nor (_32601_, _32600_, _08267_);
  nand (_32602_, _32601_, _32599_);
  nor (_32604_, _08266_, _02860_);
  nor (_32605_, _32604_, _03334_);
  nand (_32606_, _32605_, _32602_);
  nor (_32607_, _03270_, _03233_);
  nor (_32608_, _32607_, _03452_);
  and (_32609_, _32608_, _32606_);
  and (_32610_, _03452_, \oc8051_golden_model_1.PC [1]);
  or (_32611_, _32610_, _32609_);
  nand (_32612_, _32611_, _05919_);
  and (_32613_, _04325_, _03219_);
  nor (_32615_, _32613_, _03621_);
  nand (_32616_, _32615_, _32612_);
  and (_32617_, _03621_, _03270_);
  not (_32618_, _32617_);
  and (_32619_, _32618_, _11797_);
  nand (_32620_, _32619_, _32616_);
  nor (_32621_, _11797_, _02860_);
  nor (_32622_, _32621_, _03224_);
  nand (_32623_, _32622_, _32620_);
  not (_32624_, _11806_);
  and (_32625_, _03270_, _03224_);
  nor (_32626_, _32625_, _32624_);
  nand (_32627_, _32626_, _32623_);
  nor (_32628_, _11806_, _03313_);
  nor (_32629_, _32628_, _03517_);
  nand (_32630_, _32629_, _32627_);
  and (_32631_, _03517_, _02860_);
  nor (_32632_, _32631_, _03159_);
  nand (_32633_, _32632_, _32630_);
  and (_32634_, _04325_, _03159_);
  nor (_32637_, _32634_, _11813_);
  nand (_32638_, _32637_, _32633_);
  and (_32639_, _32463_, _11813_);
  nor (_32640_, _32639_, _06193_);
  and (_32641_, _32640_, _32638_);
  nor (_32642_, _03624_, \oc8051_golden_model_1.PC [1]);
  nor (_32643_, _32642_, _05917_);
  or (_32644_, _32643_, _32641_);
  and (_32645_, _03624_, _03270_);
  nor (_32646_, _32645_, _08461_);
  and (_32648_, _32646_, _32644_);
  and (_32649_, _08461_, \oc8051_golden_model_1.PC [1]);
  or (_32650_, _32649_, _32648_);
  nand (_32651_, _32650_, _23814_);
  and (_32652_, _11828_, _03319_);
  nor (_32653_, _32652_, _03516_);
  nand (_32654_, _32653_, _32651_);
  and (_32655_, _03516_, _02860_);
  nor (_32656_, _32655_, _03168_);
  nand (_32657_, _32656_, _32654_);
  and (_32659_, _04325_, _03168_);
  nor (_32660_, _32659_, _11868_);
  nand (_32661_, _32660_, _32657_);
  not (_32662_, _15828_);
  nor (_32663_, _32463_, _08864_);
  and (_32664_, _08864_, \oc8051_golden_model_1.PC [1]);
  nor (_32665_, _32664_, _23819_);
  not (_32666_, _32665_);
  nor (_32667_, _32666_, _32663_);
  nor (_32668_, _32667_, _32662_);
  and (_32670_, _32668_, _32661_);
  or (_32671_, _32670_, _32452_);
  nor (_32672_, _16000_, _08476_);
  nand (_32673_, _32672_, _32671_);
  nor (_32674_, _32672_, _03313_);
  nor (_32675_, _32674_, _04129_);
  nand (_32676_, _32675_, _32673_);
  and (_32677_, _04129_, _03313_);
  nor (_32678_, _32677_, _08494_);
  and (_32679_, _32678_, _32676_);
  or (_32681_, _32679_, _32451_);
  nand (_32682_, _32681_, _04527_);
  and (_32683_, _03623_, _03313_);
  nor (_32684_, _32683_, _03744_);
  nand (_32685_, _32684_, _32682_);
  and (_32686_, _03744_, _02860_);
  nor (_32687_, _32686_, _03172_);
  nand (_32688_, _32687_, _32685_);
  and (_32689_, _04325_, _03172_);
  nor (_32690_, _32689_, _11889_);
  nand (_32692_, _32690_, _32688_);
  nor (_32693_, _32463_, _11894_);
  nor (_32694_, _08864_, _02860_);
  nor (_32695_, _32694_, _11893_);
  not (_32696_, _32695_);
  nor (_32697_, _32696_, _32693_);
  nor (_32698_, _32697_, _11901_);
  and (_32699_, _32698_, _32692_);
  or (_32700_, _32699_, _32450_);
  nand (_32701_, _32700_, _11904_);
  nor (_32703_, _11904_, _02860_);
  nor (_32704_, _32703_, _03611_);
  nand (_32705_, _32704_, _32701_);
  and (_32706_, _03611_, _03270_);
  nor (_32707_, _32706_, _03733_);
  and (_32708_, _32707_, _32705_);
  and (_32709_, _03733_, \oc8051_golden_model_1.PC [1]);
  or (_32710_, _32709_, _32708_);
  nand (_32711_, _32710_, _32195_);
  and (_32712_, _04325_, _03182_);
  nor (_32714_, _32712_, _11915_);
  nand (_32715_, _32714_, _32711_);
  and (_32716_, \oc8051_golden_model_1.PSW [7], _02860_);
  and (_32717_, _32463_, _07982_);
  or (_32718_, _32717_, _32716_);
  and (_32719_, _32718_, _11915_);
  nor (_32720_, _32719_, _07927_);
  and (_32721_, _32720_, _32715_);
  or (_32722_, _32721_, _32448_);
  or (_32723_, _11411_, _02986_);
  and (_32725_, _32723_, _16701_);
  nand (_32726_, _32725_, _32722_);
  nor (_32727_, _32725_, _03313_);
  nor (_32728_, _32727_, _04156_);
  nand (_32729_, _32728_, _32726_);
  and (_32730_, _04156_, _03313_);
  nor (_32731_, _32730_, _15156_);
  nand (_32732_, _32731_, _32729_);
  nor (_32733_, _11410_, _02860_);
  nor (_32734_, _32733_, _03618_);
  nand (_32736_, _32734_, _32732_);
  and (_32737_, _03618_, _03270_);
  nor (_32738_, _32737_, _03741_);
  and (_32739_, _32738_, _32736_);
  and (_32740_, _03741_, \oc8051_golden_model_1.PC [1]);
  or (_32741_, _32740_, _32739_);
  nand (_32742_, _32741_, _32192_);
  and (_32743_, _04325_, _03178_);
  nor (_32744_, _32743_, _11936_);
  nand (_32745_, _32744_, _32742_);
  nand (_32747_, _03565_, _03190_);
  not (_32748_, _32747_);
  nor (_32749_, _32463_, _07982_);
  and (_32750_, _07982_, \oc8051_golden_model_1.PC [1]);
  nor (_32751_, _32750_, _11942_);
  not (_32752_, _32751_);
  nor (_32753_, _32752_, _32749_);
  nor (_32754_, _32753_, _32748_);
  nand (_32755_, _32754_, _32745_);
  nor (_32756_, _32747_, _03313_);
  nor (_32758_, _32756_, _08554_);
  and (_32759_, _05912_, _05140_);
  nor (_32760_, _32759_, _04166_);
  not (_32761_, _32760_);
  and (_32762_, _32761_, _32758_);
  nand (_32763_, _32762_, _32755_);
  or (_32764_, _08554_, _08595_);
  or (_32765_, _32764_, _08559_);
  or (_32766_, _32765_, _08562_);
  and (_32767_, _32766_, _03313_);
  nor (_32769_, _32767_, _08629_);
  nand (_32770_, _32769_, _32763_);
  nor (_32771_, _08628_, _02860_);
  nor (_32772_, _32771_, _08707_);
  nand (_32773_, _32772_, _32770_);
  and (_32774_, _08707_, _03313_);
  nor (_32775_, _32774_, _03752_);
  and (_32776_, _32775_, _32773_);
  nor (_32777_, _06572_, _10735_);
  or (_32778_, _32777_, _32776_);
  nand (_32780_, _32778_, _04803_);
  and (_32781_, _04325_, _03191_);
  nor (_32782_, _32781_, _03617_);
  and (_32783_, _32782_, _32780_);
  and (_32784_, _32456_, _09953_);
  nor (_32785_, _09953_, _03313_);
  nor (_32786_, _32785_, _32784_);
  nor (_32787_, _32786_, _03814_);
  or (_32788_, _32787_, _32783_);
  nand (_32789_, _32788_, _11406_);
  nor (_32791_, _11406_, _03270_);
  nor (_32792_, _32791_, _08785_);
  nand (_32793_, _32792_, _32789_);
  nor (_32794_, _08784_, _02860_);
  nor (_32795_, _32794_, _08815_);
  nand (_32796_, _32795_, _32793_);
  and (_32797_, _08815_, _03313_);
  nor (_32798_, _32797_, _03475_);
  and (_32799_, _32798_, _32796_);
  nor (_32800_, _06572_, _03476_);
  or (_32802_, _32800_, _32799_);
  nand (_32803_, _32802_, _11405_);
  and (_32804_, _04325_, _03189_);
  nor (_32805_, _32804_, _03644_);
  nand (_32806_, _32805_, _32803_);
  and (_32807_, _09953_, _03313_);
  nor (_32808_, _32456_, _09953_);
  nor (_32809_, _32808_, _32807_);
  and (_32810_, _32809_, _03644_);
  nor (_32811_, _32810_, _23193_);
  and (_32813_, _32811_, _32806_);
  nor (_32814_, _11989_, _03313_);
  nor (_32815_, _32814_, _32813_);
  or (_32816_, _32815_, _24500_);
  and (_32817_, _24500_, _03270_);
  nor (_32818_, _32817_, _03767_);
  nand (_32819_, _32818_, _32816_);
  and (_32820_, _03767_, _02860_);
  nor (_32821_, _32820_, _11999_);
  and (_32822_, _32821_, _32819_);
  or (_32824_, _32822_, _32447_);
  nand (_32825_, _32824_, _04553_);
  and (_32826_, _04986_, _04325_);
  nor (_32827_, _32826_, _03445_);
  nand (_32828_, _32827_, _32825_);
  and (_32829_, _32809_, _03445_);
  nor (_32830_, _32829_, _06830_);
  and (_32831_, _32830_, _32828_);
  and (_32832_, _06830_, _03270_);
  or (_32833_, _32832_, _32831_);
  nand (_32835_, _32833_, _32446_);
  nor (_32836_, _32446_, _03313_);
  nor (_32837_, _32836_, _03473_);
  and (_32838_, _32837_, _32835_);
  or (_32839_, _32838_, _32445_);
  nand (_32840_, _32839_, _11392_);
  nor (_32841_, _11392_, _03270_);
  nor (_32842_, _32841_, _32181_);
  nand (_32843_, _32842_, _32840_);
  and (_32844_, _32181_, _04325_);
  nor (_32846_, _32844_, _12031_);
  nand (_32847_, _32846_, _32843_);
  and (_32848_, _12031_, _03313_);
  not (_32849_, _32848_);
  nand (_32850_, _32849_, _32847_);
  or (_32851_, _32850_, _43193_);
  or (_32852_, _43189_, \oc8051_golden_model_1.PC [1]);
  and (_32853_, _32852_, _42003_);
  and (_43921_, _32853_, _32851_);
  and (_32854_, _03473_, _03294_);
  nor (_32856_, _11998_, _03267_);
  nor (_32857_, _11406_, _03267_);
  nor (_32858_, _11408_, _03267_);
  nor (_32859_, _11413_, _03267_);
  and (_32860_, _11901_, _03299_);
  nor (_32861_, _11416_, _03267_);
  and (_32862_, _03632_, _03167_);
  nor (_32863_, _11806_, _03267_);
  nor (_32864_, _11419_, _03267_);
  nor (_32865_, _32576_, _03294_);
  and (_32867_, _11514_, _11511_);
  nor (_32868_, _32867_, _11515_);
  not (_32869_, _32868_);
  or (_32870_, _32869_, _11437_);
  or (_32871_, _11504_, _11439_);
  and (_32872_, _32871_, _03534_);
  and (_32873_, _32872_, _32870_);
  and (_32874_, _11566_, _03294_);
  and (_32875_, _11628_, _11625_);
  nor (_32876_, _32875_, _11629_);
  and (_32878_, _32876_, _32232_);
  nor (_32879_, _32878_, _32874_);
  nand (_32880_, _32879_, _05998_);
  and (_32881_, _03855_, _04435_);
  nor (_32882_, _11684_, _03267_);
  not (_32883_, _32882_);
  and (_32884_, _11680_, _03204_);
  and (_32885_, _04436_, _11618_);
  nor (_32886_, _04436_, \oc8051_golden_model_1.PC [2]);
  and (_32887_, _32886_, _11688_);
  nor (_32889_, _32887_, _32885_);
  nor (_32890_, _32889_, _08108_);
  and (_32891_, _32890_, _32884_);
  nor (_32892_, _32891_, _03536_);
  and (_32893_, _32892_, _32883_);
  not (_32894_, _32893_);
  nor (_32895_, _32894_, _32881_);
  and (_32896_, _03536_, _03294_);
  or (_32897_, _32896_, _32895_);
  and (_32898_, _32897_, _11686_);
  and (_32900_, _08118_, _03267_);
  or (_32901_, _32900_, _32898_);
  and (_32902_, _32901_, _03209_);
  nor (_32903_, _03855_, _03209_);
  nor (_32904_, _32903_, _05998_);
  not (_32905_, _32904_);
  nor (_32906_, _32905_, _32902_);
  nor (_32907_, _32906_, _04012_);
  nand (_32908_, _32907_, _32880_);
  nand (_32909_, _04012_, _03267_);
  and (_32911_, _32909_, _04432_);
  and (_32912_, _32911_, _32908_);
  or (_32913_, _32912_, _32873_);
  nand (_32914_, _32913_, _11430_);
  nor (_32915_, _11430_, _03267_);
  nor (_32916_, _32915_, _03469_);
  nand (_32917_, _32916_, _32914_);
  and (_32918_, _03469_, _03294_);
  nor (_32919_, _32918_, _05977_);
  nand (_32920_, _32919_, _32917_);
  and (_32922_, _03855_, _05977_);
  nor (_32923_, _32922_, _03527_);
  nand (_32924_, _32923_, _32920_);
  and (_32925_, _03527_, _03294_);
  nor (_32926_, _32925_, _11716_);
  nand (_32927_, _32926_, _32924_);
  nor (_32928_, _11715_, _03267_);
  nor (_32929_, _32928_, _03530_);
  nand (_32930_, _32929_, _32927_);
  and (_32931_, _03530_, _03294_);
  nor (_32933_, _32931_, _11724_);
  nand (_32934_, _32933_, _32930_);
  nor (_32935_, _11723_, _03267_);
  nor (_32936_, _32935_, _03465_);
  nand (_32937_, _32936_, _32934_);
  and (_32938_, _03465_, _03294_);
  nor (_32939_, _32938_, _11727_);
  nand (_32940_, _32939_, _32937_);
  and (_32941_, _03855_, _11727_);
  nor (_32942_, _32941_, _03464_);
  nand (_32944_, _32942_, _32940_);
  and (_32945_, _03464_, _03294_);
  nor (_32946_, _32945_, _10021_);
  nand (_32947_, _32946_, _32944_);
  and (_32948_, _11503_, _10055_);
  nor (_32949_, _32869_, _10055_);
  or (_32950_, _32949_, _32948_);
  nor (_32951_, _32950_, _10017_);
  nor (_32952_, _32951_, _10020_);
  and (_32953_, _32952_, _32947_);
  or (_32955_, _32869_, _10116_);
  or (_32956_, _11504_, _11743_);
  and (_32957_, _32956_, _32955_);
  nor (_32958_, _32957_, _10112_);
  or (_32959_, _32958_, _03547_);
  or (_32960_, _32959_, _32953_);
  and (_32961_, _11503_, _09975_);
  nor (_32962_, _32869_, _09975_);
  or (_32963_, _32962_, _03994_);
  or (_32964_, _32963_, _32961_);
  and (_32966_, _32964_, _10123_);
  nand (_32967_, _32966_, _32960_);
  and (_32968_, _32868_, _11764_);
  and (_32969_, _11503_, _10163_);
  nor (_32970_, _32969_, _32968_);
  nor (_32971_, _32970_, _10158_);
  and (_32972_, _10122_, _03267_);
  nor (_32973_, _32972_, _32971_);
  and (_32974_, _32973_, _03459_);
  nand (_32975_, _32974_, _32967_);
  and (_32976_, _03458_, _11618_);
  nor (_32977_, _32976_, _04755_);
  nand (_32978_, _32977_, _32975_);
  nor (_32979_, _03855_, _03207_);
  nor (_32980_, _32979_, _32577_);
  and (_32981_, _32980_, _32978_);
  or (_32982_, _32981_, _32865_);
  nand (_32983_, _32982_, _11424_);
  nor (_32984_, _11424_, _03267_);
  nor (_32985_, _32984_, _03587_);
  and (_32988_, _32985_, _32983_);
  and (_32989_, _03587_, _03294_);
  or (_32990_, _32989_, _11776_);
  or (_32991_, _32990_, _32988_);
  and (_32992_, _03855_, _11776_);
  nor (_32993_, _32992_, _03586_);
  nand (_32994_, _32993_, _32991_);
  and (_32995_, _03586_, _03294_);
  nor (_32996_, _32995_, _11780_);
  and (_32997_, _32996_, _32994_);
  or (_32999_, _32997_, _32864_);
  nand (_33000_, _32999_, _08266_);
  nor (_33001_, _08266_, _03294_);
  nor (_33002_, _33001_, _03334_);
  nand (_33003_, _33002_, _33000_);
  nor (_33004_, _03299_, _03233_);
  nor (_33005_, _33004_, _03452_);
  and (_33006_, _33005_, _33003_);
  and (_33007_, _11618_, _03452_);
  or (_33008_, _33007_, _33006_);
  nand (_33010_, _33008_, _05919_);
  and (_33011_, _03855_, _03219_);
  nor (_33012_, _33011_, _03621_);
  nand (_33013_, _33012_, _33010_);
  and (_33014_, _11503_, _03621_);
  not (_33015_, _33014_);
  and (_33016_, _33015_, _11797_);
  nand (_33017_, _33016_, _33013_);
  nor (_33018_, _11797_, _03294_);
  nor (_33019_, _33018_, _03224_);
  nand (_33021_, _33019_, _33017_);
  and (_33022_, _11503_, _03224_);
  nor (_33023_, _33022_, _32624_);
  and (_33024_, _33023_, _33021_);
  or (_33025_, _33024_, _32863_);
  and (_33026_, _33025_, _10351_);
  and (_33027_, _03517_, _11618_);
  or (_33028_, _33027_, _03159_);
  or (_33029_, _33028_, _33026_);
  nor (_33030_, _03855_, _03160_);
  nor (_33032_, _33030_, _11813_);
  and (_33033_, _33032_, _33029_);
  nor (_33034_, _32876_, _11814_);
  nor (_33035_, _33034_, _33033_);
  or (_33036_, _33035_, _32862_);
  and (_33037_, _04793_, _03577_);
  and (_33038_, _33037_, _11618_);
  and (_33039_, _03612_, _03167_);
  nor (_33040_, _03864_, _03578_);
  nor (_33041_, _33040_, _05911_);
  or (_33043_, _33041_, _33039_);
  nor (_33044_, _33043_, _33038_);
  nand (_33045_, _33044_, _33036_);
  and (_33046_, _33043_, _03294_);
  nor (_33047_, _32759_, _05911_);
  nor (_33048_, _33047_, _33046_);
  nand (_33049_, _33048_, _33045_);
  and (_33050_, _33047_, _11618_);
  nor (_33051_, _33050_, _03624_);
  nand (_33052_, _33051_, _33049_);
  and (_33054_, _11503_, _03624_);
  nor (_33055_, _33054_, _08461_);
  and (_33056_, _33055_, _33052_);
  and (_33057_, _08461_, _11618_);
  or (_33058_, _33057_, _33056_);
  nand (_33059_, _33058_, _23814_);
  nor (_33060_, _23814_, _03297_);
  nor (_33061_, _33060_, _03516_);
  nand (_33062_, _33061_, _33059_);
  and (_33063_, _03516_, _03294_);
  nor (_33065_, _33063_, _03168_);
  nand (_33066_, _33065_, _33062_);
  and (_33067_, _03855_, _03168_);
  nor (_33068_, _33067_, _11868_);
  nand (_33069_, _33068_, _33066_);
  and (_33070_, _08864_, _03294_);
  and (_33071_, _32876_, _11894_);
  or (_33072_, _33071_, _33070_);
  and (_33073_, _33072_, _11868_);
  nor (_33074_, _33073_, _11872_);
  and (_33076_, _33074_, _33069_);
  or (_33077_, _33076_, _32861_);
  nand (_33078_, _33077_, _08493_);
  nor (_33079_, _08493_, _03294_);
  nor (_33080_, _33079_, _03623_);
  nand (_33081_, _33080_, _33078_);
  and (_33082_, _11503_, _03623_);
  nor (_33083_, _33082_, _03744_);
  and (_33084_, _33083_, _33081_);
  and (_33085_, _03744_, _11618_);
  or (_33087_, _33085_, _33084_);
  nand (_33088_, _33087_, _32199_);
  and (_33089_, _03855_, _03172_);
  nor (_33090_, _33089_, _11889_);
  nand (_33091_, _33090_, _33088_);
  nor (_33092_, _32876_, _11894_);
  nor (_33093_, _08864_, _03294_);
  nor (_33094_, _33093_, _11893_);
  not (_33095_, _33094_);
  nor (_33096_, _33095_, _33092_);
  nor (_33098_, _33096_, _11901_);
  and (_33099_, _33098_, _33091_);
  or (_33100_, _33099_, _32860_);
  nand (_33101_, _33100_, _11904_);
  nor (_33102_, _11904_, _03294_);
  nor (_33103_, _33102_, _03611_);
  nand (_33104_, _33103_, _33101_);
  and (_33105_, _11503_, _03611_);
  nor (_33106_, _33105_, _03733_);
  and (_33107_, _33106_, _33104_);
  and (_33109_, _03733_, _11618_);
  or (_33110_, _33109_, _33107_);
  nand (_33111_, _33110_, _32195_);
  and (_33112_, _03855_, _03182_);
  nor (_33113_, _33112_, _11915_);
  nand (_33114_, _33113_, _33111_);
  and (_33115_, _03294_, \oc8051_golden_model_1.PSW [7]);
  and (_33116_, _32876_, _07982_);
  or (_33117_, _33116_, _33115_);
  and (_33118_, _33117_, _11915_);
  nor (_33119_, _33118_, _11919_);
  and (_33120_, _33119_, _33114_);
  or (_33121_, _33120_, _32859_);
  nand (_33122_, _33121_, _11410_);
  nor (_33123_, _11410_, _03294_);
  nor (_33124_, _33123_, _03618_);
  nand (_33125_, _33124_, _33122_);
  and (_33126_, _11503_, _03618_);
  nor (_33127_, _33126_, _03741_);
  and (_33128_, _33127_, _33125_);
  and (_33130_, _03741_, _11618_);
  or (_33131_, _33130_, _33128_);
  nand (_33132_, _33131_, _32192_);
  and (_33133_, _03855_, _03178_);
  nor (_33134_, _33133_, _11936_);
  nand (_33135_, _33134_, _33132_);
  nor (_33136_, _32876_, _07982_);
  nor (_33137_, _03294_, \oc8051_golden_model_1.PSW [7]);
  nor (_33138_, _33137_, _11942_);
  not (_33139_, _33138_);
  nor (_33141_, _33139_, _33136_);
  nor (_33142_, _33141_, _11940_);
  and (_33143_, _33142_, _33135_);
  or (_33144_, _33143_, _32858_);
  nand (_33145_, _33144_, _08628_);
  nor (_33146_, _08628_, _03294_);
  nor (_33147_, _33146_, _08707_);
  nand (_33148_, _33147_, _33145_);
  and (_33149_, _08707_, _03267_);
  nor (_33150_, _33149_, _03752_);
  and (_33152_, _33150_, _33148_);
  nor (_33153_, _06710_, _10735_);
  or (_33154_, _33153_, _33152_);
  nand (_33155_, _33154_, _04803_);
  and (_33156_, _03855_, _03191_);
  nor (_33157_, _33156_, _03617_);
  nand (_33158_, _33157_, _33155_);
  and (_33159_, _32869_, _09953_);
  nor (_33160_, _11503_, _09953_);
  or (_33161_, _33160_, _03814_);
  nor (_33163_, _33161_, _33159_);
  nor (_33164_, _33163_, _11963_);
  and (_33165_, _33164_, _33158_);
  or (_33166_, _33165_, _32857_);
  nand (_33167_, _33166_, _08784_);
  nor (_33168_, _08784_, _03294_);
  nor (_33169_, _33168_, _08815_);
  nand (_33170_, _33169_, _33167_);
  and (_33171_, _08815_, _03267_);
  nor (_33172_, _33171_, _03475_);
  and (_33174_, _33172_, _33170_);
  nor (_33175_, _06710_, _03476_);
  or (_33176_, _33175_, _33174_);
  nand (_33177_, _33176_, _11405_);
  and (_33178_, _03855_, _03189_);
  nor (_33179_, _33178_, _03644_);
  nand (_33180_, _33179_, _33177_);
  nor (_33181_, _32868_, _09953_);
  and (_33182_, _11504_, _09953_);
  nor (_33183_, _33182_, _33181_);
  and (_33185_, _33183_, _03644_);
  nor (_33186_, _33185_, _11992_);
  nand (_33187_, _33186_, _33180_);
  nor (_33188_, _11991_, _03267_);
  nor (_33189_, _33188_, _03767_);
  nand (_33190_, _33189_, _33187_);
  and (_33191_, _03767_, _03294_);
  nor (_33192_, _33191_, _11999_);
  and (_33193_, _33192_, _33190_);
  or (_33194_, _33193_, _32856_);
  nand (_33196_, _33194_, _04553_);
  and (_33197_, _04986_, _03855_);
  nor (_33198_, _33197_, _03445_);
  nand (_33199_, _33198_, _33196_);
  and (_33200_, _33183_, _03445_);
  nor (_33201_, _33200_, _12016_);
  nand (_33202_, _33201_, _33199_);
  nor (_33203_, _12015_, _03267_);
  nor (_33204_, _33203_, _03473_);
  and (_33205_, _33204_, _33202_);
  or (_33207_, _33205_, _32854_);
  nand (_33208_, _33207_, _11392_);
  nor (_33209_, _11392_, _03299_);
  nor (_33210_, _33209_, _32181_);
  nand (_33211_, _33210_, _33208_);
  and (_33212_, _32181_, _03855_);
  nor (_33213_, _33212_, _12031_);
  nand (_33214_, _33213_, _33211_);
  and (_33215_, _12031_, _03267_);
  not (_33216_, _33215_);
  and (_33218_, _33216_, _33214_);
  nand (_33219_, _33218_, _43189_);
  or (_33220_, _43189_, \oc8051_golden_model_1.PC [2]);
  and (_33221_, _33220_, _42003_);
  and (_43922_, _33221_, _33219_);
  and (_33222_, _12031_, _03667_);
  not (_33223_, _33222_);
  and (_33224_, _03473_, _02866_);
  nor (_33225_, _11998_, _03667_);
  nor (_33226_, _11406_, _03667_);
  nor (_33228_, _11408_, _03667_);
  nor (_33229_, _11413_, _03667_);
  and (_33230_, _11901_, _03257_);
  nor (_33231_, _11416_, _03667_);
  nor (_33232_, _11419_, _03667_);
  nor (_33233_, _32576_, _02866_);
  and (_33234_, _11498_, _11437_);
  or (_33235_, _11501_, _11500_);
  and (_33236_, _33235_, _11516_);
  nor (_33237_, _33235_, _11516_);
  nor (_33239_, _33237_, _33236_);
  and (_33240_, _33239_, _11439_);
  or (_33241_, _33240_, _04432_);
  or (_33242_, _33241_, _33234_);
  or (_33243_, _11617_, _11616_);
  and (_33244_, _33243_, _11630_);
  nor (_33245_, _33243_, _11630_);
  nor (_33246_, _33245_, _33244_);
  and (_33247_, _33246_, _32232_);
  and (_33248_, _11566_, _02866_);
  nor (_33250_, _33248_, _33247_);
  nand (_33251_, _33250_, _05998_);
  nand (_33252_, _03725_, _04435_);
  nor (_33253_, _11680_, _03667_);
  nor (_33254_, _33253_, _03536_);
  not (_33255_, _32884_);
  nor (_33256_, _11683_, _03667_);
  and (_33257_, _04436_, _03665_);
  nor (_33258_, _04436_, \oc8051_golden_model_1.PC [3]);
  and (_33259_, _33258_, _11688_);
  nor (_33261_, _33259_, _33257_);
  nor (_33262_, _33261_, _08108_);
  nor (_33263_, _33262_, _33256_);
  or (_33264_, _33263_, _33255_);
  and (_33265_, _33264_, _33254_);
  and (_33266_, _33265_, _33252_);
  and (_33267_, _03536_, _02866_);
  or (_33268_, _33267_, _33266_);
  and (_33269_, _33268_, _11686_);
  and (_33270_, _08118_, _03667_);
  or (_33272_, _33270_, _33269_);
  and (_33273_, _33272_, _03209_);
  nor (_33274_, _03725_, _03209_);
  nor (_33275_, _33274_, _05998_);
  not (_33276_, _33275_);
  nor (_33277_, _33276_, _33273_);
  nor (_33278_, _33277_, _04012_);
  and (_33279_, _33278_, _33251_);
  and (_33280_, _04012_, _03667_);
  or (_33281_, _33280_, _03534_);
  or (_33283_, _33281_, _33279_);
  nand (_33284_, _33283_, _33242_);
  nand (_33285_, _33284_, _11430_);
  nor (_33286_, _11430_, _03667_);
  nor (_33287_, _33286_, _03469_);
  nand (_33288_, _33287_, _33285_);
  and (_33289_, _03469_, _02866_);
  nor (_33290_, _33289_, _05977_);
  nand (_33291_, _33290_, _33288_);
  and (_33292_, _03725_, _05977_);
  nor (_33294_, _33292_, _03527_);
  nand (_33295_, _33294_, _33291_);
  and (_33296_, _03527_, _02866_);
  nor (_33297_, _33296_, _11716_);
  nand (_33298_, _33297_, _33295_);
  nor (_33299_, _11715_, _03667_);
  nor (_33300_, _33299_, _03530_);
  nand (_33301_, _33300_, _33298_);
  and (_33302_, _03530_, _02866_);
  nor (_33303_, _33302_, _11724_);
  nand (_33305_, _33303_, _33301_);
  nor (_33306_, _11723_, _03667_);
  nor (_33307_, _33306_, _03465_);
  nand (_33308_, _33307_, _33305_);
  and (_33309_, _03465_, _02866_);
  nor (_33310_, _33309_, _11727_);
  nand (_33311_, _33310_, _33308_);
  and (_33312_, _03725_, _11727_);
  nor (_33313_, _33312_, _03464_);
  nand (_33314_, _33313_, _33311_);
  and (_33316_, _03464_, _02866_);
  nor (_33317_, _33316_, _10021_);
  nand (_33318_, _33317_, _33314_);
  and (_33319_, _11498_, _10055_);
  not (_33320_, _33239_);
  nor (_33321_, _33320_, _10055_);
  or (_33322_, _33321_, _33319_);
  nor (_33323_, _33322_, _10017_);
  nor (_33324_, _33323_, _10020_);
  and (_33325_, _33324_, _33318_);
  and (_33327_, _33239_, _11743_);
  and (_33328_, _11498_, _10116_);
  nor (_33329_, _33328_, _33327_);
  nor (_33330_, _33329_, _10112_);
  or (_33331_, _33330_, _03547_);
  or (_33332_, _33331_, _33325_);
  nor (_33333_, _33320_, _09975_);
  and (_33334_, _11498_, _09975_);
  or (_33335_, _33334_, _03994_);
  or (_33336_, _33335_, _33333_);
  and (_33338_, _33336_, _10123_);
  nand (_33339_, _33338_, _33332_);
  and (_33340_, _11498_, _10163_);
  and (_33341_, _33239_, _11764_);
  or (_33342_, _33341_, _33340_);
  and (_33343_, _33342_, _03608_);
  and (_33344_, _10122_, _03667_);
  nor (_33345_, _33344_, _33343_);
  and (_33346_, _33345_, _03459_);
  nand (_33347_, _33346_, _33339_);
  and (_33348_, _03458_, _03665_);
  nor (_33349_, _33348_, _04755_);
  nand (_33350_, _33349_, _33347_);
  nor (_33351_, _03725_, _03207_);
  nor (_33352_, _33351_, _32577_);
  and (_33353_, _33352_, _33350_);
  or (_33354_, _33353_, _33233_);
  nand (_33355_, _33354_, _11424_);
  nor (_33356_, _11424_, _03667_);
  nor (_33357_, _33356_, _03587_);
  nand (_33360_, _33357_, _33355_);
  and (_33361_, _03587_, _02866_);
  nor (_33362_, _33361_, _11776_);
  nand (_33363_, _33362_, _33360_);
  and (_33364_, _03725_, _11776_);
  nor (_33365_, _33364_, _03586_);
  nand (_33366_, _33365_, _33363_);
  and (_33367_, _03586_, _02866_);
  nor (_33368_, _33367_, _11780_);
  and (_33369_, _33368_, _33366_);
  or (_33371_, _33369_, _33232_);
  nand (_33372_, _33371_, _08266_);
  nor (_33373_, _08266_, _02866_);
  nor (_33374_, _33373_, _03334_);
  nand (_33375_, _33374_, _33372_);
  nor (_33376_, _03233_, _03257_);
  nor (_33377_, _33376_, _03452_);
  and (_33378_, _33377_, _33375_);
  and (_33379_, _03665_, _03452_);
  or (_33380_, _33379_, _33378_);
  nand (_33382_, _33380_, _05919_);
  and (_33383_, _03725_, _03219_);
  nor (_33384_, _33383_, _03621_);
  nand (_33385_, _33384_, _33382_);
  and (_33386_, _11498_, _03621_);
  not (_33387_, _33386_);
  and (_33388_, _33387_, _11797_);
  nand (_33389_, _33388_, _33385_);
  nor (_33390_, _11797_, _02866_);
  nor (_33391_, _33390_, _03224_);
  nand (_33393_, _33391_, _33389_);
  and (_33394_, _11498_, _03224_);
  nor (_33395_, _33394_, _32624_);
  nand (_33396_, _33395_, _33393_);
  nor (_33397_, _11806_, _03667_);
  nor (_33398_, _33397_, _03517_);
  nand (_33399_, _33398_, _33396_);
  and (_33400_, _03517_, _02866_);
  nor (_33401_, _33400_, _03159_);
  nand (_33402_, _33401_, _33399_);
  and (_33404_, _03725_, _03159_);
  nor (_33405_, _33404_, _11813_);
  nand (_33406_, _33405_, _33402_);
  and (_33407_, _33246_, _11813_);
  nor (_33408_, _33407_, _06193_);
  and (_33409_, _33408_, _33406_);
  nor (_33410_, _03624_, _03665_);
  nor (_33411_, _33410_, _05917_);
  or (_33412_, _33411_, _33409_);
  and (_33413_, _11498_, _03624_);
  nor (_33415_, _33413_, _08461_);
  and (_33416_, _33415_, _33412_);
  and (_33417_, _08461_, _03665_);
  or (_33418_, _33417_, _33416_);
  nand (_33419_, _33418_, _23814_);
  nor (_33420_, _23814_, _03252_);
  nor (_33421_, _33420_, _03516_);
  nand (_33422_, _33421_, _33419_);
  and (_33423_, _03516_, _02866_);
  nor (_33424_, _33423_, _03168_);
  nand (_33426_, _33424_, _33422_);
  and (_33427_, _03725_, _03168_);
  nor (_33428_, _33427_, _11868_);
  nand (_33429_, _33428_, _33426_);
  and (_33430_, _08864_, _02866_);
  and (_33431_, _33246_, _11894_);
  or (_33432_, _33431_, _33430_);
  and (_33433_, _33432_, _11868_);
  nor (_33434_, _33433_, _11872_);
  and (_33435_, _33434_, _33429_);
  or (_33437_, _33435_, _33231_);
  nand (_33438_, _33437_, _08493_);
  nor (_33439_, _08493_, _02866_);
  nor (_33440_, _33439_, _03623_);
  nand (_33441_, _33440_, _33438_);
  and (_33442_, _11498_, _03623_);
  nor (_33443_, _33442_, _03744_);
  and (_33444_, _33443_, _33441_);
  and (_33445_, _03744_, _03665_);
  or (_33446_, _33445_, _33444_);
  nand (_33448_, _33446_, _32199_);
  and (_33449_, _03725_, _03172_);
  nor (_33450_, _33449_, _11889_);
  nand (_33451_, _33450_, _33448_);
  nor (_33452_, _33246_, _11894_);
  nor (_33453_, _08864_, _02866_);
  nor (_33454_, _33453_, _11893_);
  not (_33455_, _33454_);
  nor (_33456_, _33455_, _33452_);
  nor (_33457_, _33456_, _11901_);
  and (_33459_, _33457_, _33451_);
  or (_33460_, _33459_, _33230_);
  nand (_33461_, _33460_, _11904_);
  nor (_33462_, _11904_, _02866_);
  nor (_33463_, _33462_, _03611_);
  nand (_33464_, _33463_, _33461_);
  and (_33465_, _11498_, _03611_);
  nor (_33466_, _33465_, _03733_);
  and (_33467_, _33466_, _33464_);
  and (_33468_, _03733_, _03665_);
  or (_33470_, _33468_, _33467_);
  nand (_33471_, _33470_, _32195_);
  and (_33472_, _03725_, _03182_);
  nor (_33473_, _33472_, _11915_);
  nand (_33474_, _33473_, _33471_);
  and (_33475_, _02866_, \oc8051_golden_model_1.PSW [7]);
  and (_33476_, _33246_, _07982_);
  or (_33477_, _33476_, _33475_);
  and (_33478_, _33477_, _11915_);
  nor (_33479_, _33478_, _11919_);
  and (_33481_, _33479_, _33474_);
  or (_33482_, _33481_, _33229_);
  nand (_33483_, _33482_, _11410_);
  nor (_33484_, _11410_, _02866_);
  nor (_33485_, _33484_, _03618_);
  nand (_33486_, _33485_, _33483_);
  and (_33487_, _11498_, _03618_);
  nor (_33488_, _33487_, _03741_);
  and (_33489_, _33488_, _33486_);
  and (_33490_, _03741_, _03665_);
  or (_33492_, _33490_, _33489_);
  nand (_33493_, _33492_, _32192_);
  and (_33494_, _03725_, _03178_);
  nor (_33495_, _33494_, _11936_);
  nand (_33496_, _33495_, _33493_);
  nor (_33497_, _33246_, _07982_);
  nor (_33498_, _02866_, \oc8051_golden_model_1.PSW [7]);
  nor (_33499_, _33498_, _11942_);
  not (_33500_, _33499_);
  nor (_33501_, _33500_, _33497_);
  nor (_33503_, _33501_, _11940_);
  and (_33504_, _33503_, _33496_);
  or (_33505_, _33504_, _33228_);
  nand (_33506_, _33505_, _08628_);
  nor (_33507_, _08628_, _02866_);
  nor (_33508_, _33507_, _08707_);
  nand (_33509_, _33508_, _33506_);
  and (_33510_, _08707_, _03667_);
  nor (_33511_, _33510_, _03752_);
  and (_33512_, _33511_, _33509_);
  nor (_33514_, _06664_, _10735_);
  or (_33515_, _33514_, _33512_);
  nand (_33516_, _33515_, _04803_);
  and (_33517_, _03725_, _03191_);
  nor (_33518_, _33517_, _03617_);
  nand (_33519_, _33518_, _33516_);
  and (_33520_, _33320_, _09953_);
  nor (_33521_, _11498_, _09953_);
  or (_33522_, _33521_, _03814_);
  or (_33523_, _33522_, _33520_);
  and (_33525_, _33523_, _11406_);
  and (_33526_, _33525_, _33519_);
  or (_33527_, _33526_, _33226_);
  nand (_33528_, _33527_, _08784_);
  nor (_33529_, _08784_, _02866_);
  nor (_33530_, _33529_, _08815_);
  nand (_33531_, _33530_, _33528_);
  and (_33532_, _08815_, _03667_);
  nor (_33533_, _33532_, _03475_);
  and (_33534_, _33533_, _33531_);
  nor (_33536_, _06664_, _03476_);
  or (_33537_, _33536_, _33534_);
  nand (_33538_, _33537_, _11405_);
  and (_33539_, _03725_, _03189_);
  nor (_33540_, _33539_, _03644_);
  nand (_33541_, _33540_, _33538_);
  nor (_33542_, _33239_, _09953_);
  and (_33543_, _11499_, _09953_);
  nor (_33544_, _33543_, _33542_);
  and (_33545_, _33544_, _03644_);
  nor (_33547_, _33545_, _11992_);
  nand (_33548_, _33547_, _33541_);
  nor (_33549_, _11991_, _03667_);
  nor (_33550_, _33549_, _03767_);
  nand (_33551_, _33550_, _33548_);
  and (_33552_, _03767_, _02866_);
  nor (_33553_, _33552_, _11999_);
  and (_33554_, _33553_, _33551_);
  or (_33555_, _33554_, _33225_);
  nand (_33556_, _33555_, _04553_);
  and (_33558_, _04986_, _03725_);
  nor (_33559_, _33558_, _03445_);
  nand (_33560_, _33559_, _33556_);
  and (_33561_, _33544_, _03445_);
  nor (_33562_, _33561_, _12016_);
  nand (_33563_, _33562_, _33560_);
  nor (_33564_, _12015_, _03667_);
  nor (_33565_, _33564_, _03473_);
  and (_33566_, _33565_, _33563_);
  or (_33567_, _33566_, _33224_);
  nand (_33569_, _33567_, _11392_);
  nor (_33570_, _11392_, _03257_);
  nor (_33571_, _33570_, _32181_);
  nand (_33572_, _33571_, _33569_);
  and (_33573_, _32181_, _03725_);
  nor (_33574_, _33573_, _12031_);
  nand (_33575_, _33574_, _33572_);
  and (_33576_, _33575_, _33223_);
  nand (_33577_, _33576_, _43189_);
  or (_33578_, _43189_, \oc8051_golden_model_1.PC [3]);
  and (_33580_, _33578_, _42003_);
  and (_43923_, _33580_, _33577_);
  not (_33581_, \oc8051_golden_model_1.PC [4]);
  nor (_33582_, _02884_, _33581_);
  and (_33583_, _02884_, _33581_);
  nor (_33584_, _33583_, _33582_);
  and (_33585_, _33584_, _12031_);
  not (_33586_, _33585_);
  and (_33587_, _06326_, _04986_);
  and (_33588_, _11494_, _03621_);
  and (_33590_, _06326_, _11776_);
  nor (_33591_, _32576_, _11613_);
  and (_33592_, _11614_, _03465_);
  nor (_33593_, _33584_, _11715_);
  and (_33594_, _11521_, _11518_);
  nor (_33595_, _33594_, _11522_);
  or (_33596_, _33595_, _11437_);
  and (_33597_, _33596_, _03534_);
  or (_33598_, _11494_, _11439_);
  and (_33599_, _33598_, _33597_);
  and (_33601_, _11635_, _11632_);
  nor (_33602_, _33601_, _11636_);
  nand (_33603_, _33602_, _32232_);
  or (_33604_, _32232_, _11614_);
  and (_33605_, _33604_, _05998_);
  nand (_33606_, _33605_, _33603_);
  and (_33607_, _06326_, _04435_);
  and (_33608_, _11614_, _04436_);
  or (_33609_, _33608_, _08108_);
  or (_33610_, _11682_, _33581_);
  and (_33612_, _33610_, _04437_);
  or (_33613_, _33612_, _33609_);
  not (_33614_, _33584_);
  or (_33615_, _33614_, _11683_);
  and (_33616_, _33615_, _03204_);
  and (_33617_, _33616_, _33613_);
  or (_33618_, _33617_, _15022_);
  or (_33619_, _33618_, _33607_);
  or (_33620_, _33614_, _11680_);
  and (_33621_, _33620_, _08101_);
  and (_33623_, _33621_, _33619_);
  and (_33624_, _11614_, _03536_);
  or (_33625_, _33624_, _33623_);
  nor (_33626_, _33625_, _08118_);
  and (_33627_, _33584_, _08118_);
  or (_33628_, _33627_, _33626_);
  and (_33629_, _33628_, _03209_);
  nor (_33630_, _06326_, _03209_);
  nor (_33631_, _33630_, _05998_);
  not (_33632_, _33631_);
  nor (_33634_, _33632_, _33629_);
  not (_33635_, _33634_);
  and (_33636_, _33635_, _11705_);
  and (_33637_, _33636_, _33606_);
  or (_33638_, _33637_, _33599_);
  and (_33639_, _33638_, _11430_);
  and (_33640_, _33584_, _11710_);
  or (_33641_, _33640_, _03469_);
  or (_33642_, _33641_, _33639_);
  and (_33643_, _11614_, _03469_);
  nor (_33645_, _33643_, _05977_);
  and (_33646_, _33645_, _33642_);
  nor (_33647_, _06326_, _03202_);
  or (_33648_, _33647_, _03527_);
  nor (_33649_, _33648_, _33646_);
  and (_33650_, _11614_, _03527_);
  or (_33651_, _33650_, _33649_);
  and (_33652_, _33651_, _11715_);
  or (_33653_, _33652_, _33593_);
  nand (_33654_, _33653_, _03531_);
  and (_33656_, _11614_, _03530_);
  nor (_33657_, _33656_, _11724_);
  nand (_33658_, _33657_, _33654_);
  nor (_33659_, _33614_, _11723_);
  nor (_33660_, _33659_, _03465_);
  and (_33661_, _33660_, _33658_);
  or (_33662_, _33661_, _33592_);
  nand (_33663_, _33662_, _03212_);
  and (_33664_, _06326_, _11727_);
  nor (_33665_, _33664_, _03464_);
  nand (_33667_, _33665_, _33663_);
  and (_33668_, _11613_, _03464_);
  nor (_33669_, _33668_, _10021_);
  nand (_33670_, _33669_, _33667_);
  and (_33671_, _11494_, _10055_);
  not (_33672_, _33595_);
  nor (_33673_, _33672_, _10055_);
  or (_33674_, _33673_, _10017_);
  nor (_33675_, _33674_, _33671_);
  not (_33676_, _33675_);
  and (_33678_, _03649_, _03631_);
  and (_33679_, _33678_, _33676_);
  nand (_33680_, _33679_, _33670_);
  nor (_33681_, _33672_, _09975_);
  and (_33682_, _11494_, _09975_);
  nor (_33683_, _33682_, _33681_);
  nor (_33684_, _33683_, _03994_);
  and (_33685_, _11494_, _10116_);
  and (_33686_, _33595_, _11743_);
  nor (_33687_, _33686_, _33685_);
  nor (_33689_, _33687_, _10112_);
  nor (_33690_, _33689_, _33684_);
  nand (_33691_, _33690_, _33680_);
  nand (_33692_, _33691_, _10123_);
  and (_33693_, _11494_, _10163_);
  and (_33694_, _33595_, _11764_);
  or (_33695_, _33694_, _33693_);
  and (_33696_, _33695_, _03608_);
  and (_33697_, _33584_, _10122_);
  nor (_33698_, _33697_, _33696_);
  and (_33700_, _33698_, _03459_);
  nand (_33701_, _33700_, _33692_);
  and (_33702_, _11614_, _03458_);
  nor (_33703_, _33702_, _04755_);
  nand (_33704_, _33703_, _33701_);
  nor (_33705_, _06326_, _03207_);
  nor (_33706_, _33705_, _32577_);
  and (_33707_, _33706_, _33704_);
  or (_33708_, _33707_, _33591_);
  nand (_33709_, _33708_, _11424_);
  nor (_33711_, _33584_, _11424_);
  nor (_33712_, _33711_, _03587_);
  nand (_33713_, _33712_, _33709_);
  and (_33714_, _11613_, _03587_);
  nor (_33715_, _33714_, _11776_);
  and (_33716_, _33715_, _33713_);
  or (_33717_, _33716_, _33590_);
  nand (_33718_, _33717_, _10265_);
  and (_33719_, _11614_, _03586_);
  nor (_33720_, _33719_, _11780_);
  nand (_33722_, _33720_, _33718_);
  nor (_33723_, _33614_, _11419_);
  nor (_33724_, _33723_, _08267_);
  nand (_33725_, _33724_, _33722_);
  nor (_33726_, _11613_, _08266_);
  nor (_33727_, _33726_, _03334_);
  nand (_33728_, _33727_, _33725_);
  nor (_33729_, _33614_, _03233_);
  nor (_33730_, _33729_, _03452_);
  and (_33731_, _33730_, _33728_);
  and (_33733_, _11614_, _03452_);
  or (_33734_, _33733_, _33731_);
  nand (_33735_, _33734_, _05919_);
  and (_33736_, _06326_, _03219_);
  nor (_33737_, _33736_, _03621_);
  nand (_33738_, _33737_, _33735_);
  nand (_33739_, _33738_, _11797_);
  or (_33740_, _33739_, _33588_);
  nor (_33741_, _11613_, _11797_);
  nor (_33742_, _33741_, _03224_);
  and (_33744_, _33742_, _33740_);
  and (_33745_, _11494_, _03224_);
  nor (_33746_, _33745_, _33744_);
  nand (_33747_, _33746_, _11806_);
  nor (_33748_, _33584_, _11806_);
  nor (_33749_, _33748_, _03517_);
  nand (_33750_, _33749_, _33747_);
  and (_33751_, _11613_, _03517_);
  nor (_33752_, _33751_, _03159_);
  nand (_33753_, _33752_, _33750_);
  and (_33755_, _06326_, _03159_);
  nor (_33756_, _33755_, _11813_);
  nand (_33757_, _33756_, _33753_);
  and (_33758_, _33602_, _11813_);
  nor (_33759_, _33758_, _06193_);
  and (_33760_, _33759_, _33757_);
  nor (_33761_, _11614_, _03624_);
  nor (_33762_, _33761_, _05917_);
  or (_33763_, _33762_, _33760_);
  and (_33764_, _11494_, _03624_);
  nor (_33766_, _33764_, _08461_);
  nand (_33767_, _33766_, _33763_);
  and (_33768_, _11614_, _08461_);
  nor (_33769_, _33768_, _11828_);
  nand (_33770_, _33769_, _33767_);
  and (_33771_, _11844_, _11841_);
  nor (_33772_, _33771_, _11845_);
  and (_33773_, _33772_, _11828_);
  nor (_33774_, _33773_, _03516_);
  and (_33775_, _33774_, _33770_);
  and (_33777_, _11614_, _03516_);
  or (_33778_, _33777_, _33775_);
  nand (_33779_, _33778_, _27595_);
  and (_33780_, _06326_, _03168_);
  nor (_33781_, _33780_, _11868_);
  and (_33782_, _33781_, _33779_);
  and (_33783_, _11613_, _08864_);
  and (_33784_, _33602_, _11894_);
  or (_33785_, _33784_, _33783_);
  and (_33786_, _33785_, _11868_);
  or (_33788_, _33786_, _33782_);
  nand (_33789_, _33788_, _11416_);
  nor (_33790_, _33614_, _11416_);
  nor (_33791_, _33790_, _08494_);
  nand (_33792_, _33791_, _33789_);
  nor (_33793_, _11613_, _08493_);
  nor (_33794_, _33793_, _03623_);
  nand (_33795_, _33794_, _33792_);
  and (_33796_, _11494_, _03623_);
  nor (_33797_, _33796_, _03744_);
  and (_33799_, _33797_, _33795_);
  and (_33800_, _11614_, _03744_);
  or (_33801_, _33800_, _33799_);
  nand (_33802_, _33801_, _32199_);
  and (_33803_, _06326_, _03172_);
  nor (_33804_, _33803_, _11889_);
  nand (_33805_, _33804_, _33802_);
  or (_33806_, _11614_, _08864_);
  nand (_33807_, _33602_, _08864_);
  and (_33808_, _33807_, _33806_);
  or (_33810_, _33808_, _11893_);
  nand (_33811_, _33810_, _33805_);
  nand (_33812_, _33811_, _11902_);
  and (_33813_, _33584_, _11901_);
  nor (_33814_, _33813_, _11905_);
  nand (_33815_, _33814_, _33812_);
  nor (_33816_, _11613_, _11904_);
  nor (_33817_, _33816_, _03611_);
  nand (_33818_, _33817_, _33815_);
  and (_33819_, _11494_, _03611_);
  nor (_33821_, _33819_, _03733_);
  and (_33822_, _33821_, _33818_);
  and (_33823_, _11614_, _03733_);
  or (_33824_, _33823_, _33822_);
  nand (_33825_, _33824_, _32195_);
  and (_33826_, _06326_, _03182_);
  nor (_33827_, _33826_, _11915_);
  and (_33828_, _33827_, _33825_);
  and (_33829_, _11613_, \oc8051_golden_model_1.PSW [7]);
  and (_33830_, _33602_, _07982_);
  or (_33832_, _33830_, _33829_);
  and (_33833_, _33832_, _11915_);
  or (_33834_, _33833_, _33828_);
  nand (_33835_, _33834_, _11413_);
  nor (_33836_, _33614_, _11413_);
  nor (_33837_, _33836_, _15156_);
  nand (_33838_, _33837_, _33835_);
  nor (_33839_, _11613_, _11410_);
  nor (_33840_, _33839_, _03618_);
  nand (_33841_, _33840_, _33838_);
  and (_33843_, _11494_, _03618_);
  nor (_33844_, _33843_, _03741_);
  and (_33845_, _33844_, _33841_);
  and (_33846_, _11614_, _03741_);
  or (_33847_, _33846_, _33845_);
  nand (_33848_, _33847_, _32192_);
  and (_33849_, _06326_, _03178_);
  nor (_33850_, _33849_, _11936_);
  nand (_33851_, _33850_, _33848_);
  nand (_33852_, _11613_, _07982_);
  nand (_33854_, _33602_, \oc8051_golden_model_1.PSW [7]);
  and (_33855_, _33854_, _33852_);
  or (_33856_, _33855_, _11942_);
  nand (_33857_, _33856_, _33851_);
  nand (_33858_, _33857_, _11408_);
  nor (_33859_, _33614_, _11408_);
  nor (_33860_, _33859_, _08629_);
  nand (_33861_, _33860_, _33858_);
  nor (_33862_, _11613_, _08628_);
  nor (_33863_, _33862_, _08707_);
  nand (_33864_, _33863_, _33861_);
  and (_33865_, _33584_, _08707_);
  nor (_33866_, _33865_, _03752_);
  and (_33867_, _33866_, _33864_);
  nor (_33868_, _06802_, _10735_);
  or (_33869_, _33868_, _33867_);
  nand (_33870_, _33869_, _04803_);
  and (_33871_, _06326_, _03191_);
  nor (_33872_, _33871_, _03617_);
  and (_33873_, _33872_, _33870_);
  nor (_33874_, _11495_, _09953_);
  and (_33875_, _33595_, _09953_);
  nor (_33876_, _33875_, _33874_);
  nor (_33877_, _33876_, _03814_);
  or (_33878_, _33877_, _33873_);
  nand (_33879_, _33878_, _11406_);
  nor (_33880_, _33614_, _11406_);
  nor (_33881_, _33880_, _08785_);
  nand (_33882_, _33881_, _33879_);
  nor (_33883_, _11613_, _08784_);
  nor (_33886_, _33883_, _08815_);
  nand (_33887_, _33886_, _33882_);
  and (_33888_, _33584_, _08815_);
  nor (_33889_, _33888_, _03475_);
  nand (_33890_, _33889_, _33887_);
  nor (_33891_, _06802_, _03476_);
  nor (_33892_, _33891_, _03189_);
  nand (_33893_, _33892_, _33890_);
  nor (_33894_, _06326_, _11405_);
  nor (_33895_, _33894_, _03644_);
  nand (_33897_, _33895_, _33893_);
  and (_33898_, _11495_, _09953_);
  nor (_33899_, _33595_, _09953_);
  nor (_33900_, _33899_, _33898_);
  nor (_33901_, _33900_, _03768_);
  nor (_33902_, _33901_, _11992_);
  nand (_33903_, _33902_, _33897_);
  nor (_33904_, _33614_, _11991_);
  nor (_33905_, _33904_, _03767_);
  nand (_33906_, _33905_, _33903_);
  and (_33908_, _11614_, _03767_);
  nor (_33909_, _33908_, _11999_);
  nand (_33910_, _33909_, _33906_);
  nor (_33911_, _33614_, _11998_);
  nor (_33912_, _33911_, _04986_);
  and (_33913_, _33912_, _33910_);
  or (_33914_, _33913_, _33587_);
  nand (_33915_, _33914_, _03446_);
  nor (_33916_, _33900_, _03446_);
  nor (_33917_, _33916_, _12016_);
  nand (_33919_, _33917_, _33915_);
  nor (_33920_, _33614_, _12015_);
  nor (_33921_, _33920_, _03473_);
  nand (_33922_, _33921_, _33919_);
  and (_33923_, _11614_, _03473_);
  nor (_33924_, _33923_, _12022_);
  nand (_33925_, _33924_, _33922_);
  nor (_33926_, _33614_, _11392_);
  nor (_33927_, _33926_, _32181_);
  nand (_33928_, _33927_, _33925_);
  and (_33930_, _32181_, _06326_);
  nor (_33931_, _33930_, _12031_);
  nand (_33932_, _33931_, _33928_);
  and (_33933_, _33932_, _33586_);
  nand (_33934_, _33933_, _43189_);
  or (_33935_, _43189_, \oc8051_golden_model_1.PC [4]);
  and (_33936_, _33935_, _42003_);
  and (_43924_, _33936_, _33934_);
  nor (_33937_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_33938_, _11608_, _02897_);
  nor (_33940_, _33938_, _33937_);
  and (_33941_, _33940_, _12031_);
  and (_33942_, _11608_, _03473_);
  nor (_33943_, _33940_, _11406_);
  nor (_33944_, _33940_, _11408_);
  nor (_33945_, _33940_, _11413_);
  not (_33946_, _33940_);
  and (_33947_, _33946_, _11901_);
  nor (_33948_, _33940_, _11416_);
  nor (_33949_, _32576_, _11608_);
  or (_33951_, _11490_, _11439_);
  or (_33952_, _11492_, _11491_);
  and (_33953_, _33952_, _11523_);
  nor (_33954_, _33952_, _11523_);
  or (_33955_, _33954_, _33953_);
  or (_33956_, _33955_, _11437_);
  and (_33957_, _33956_, _03534_);
  and (_33958_, _33957_, _33951_);
  and (_33959_, _11566_, _11608_);
  or (_33960_, _11611_, _11610_);
  not (_33962_, _33960_);
  nor (_33963_, _33962_, _11637_);
  and (_33964_, _33962_, _11637_);
  nor (_33965_, _33964_, _33963_);
  nor (_33966_, _33965_, _11566_);
  nor (_33967_, _33966_, _33959_);
  nand (_33968_, _33967_, _05998_);
  nor (_33969_, _06294_, _03204_);
  and (_33970_, _11609_, _04436_);
  nor (_33971_, _33970_, _08108_);
  and (_33973_, _11688_, \oc8051_golden_model_1.PC [5]);
  or (_33974_, _33973_, _04436_);
  and (_33975_, _33974_, _33971_);
  nor (_33976_, _33946_, _11683_);
  or (_33977_, _33976_, _15022_);
  or (_33978_, _33977_, _33975_);
  and (_33979_, _33978_, _03204_);
  nor (_33980_, _33979_, _33969_);
  nor (_33981_, _33940_, _11680_);
  nor (_33982_, _33981_, _03536_);
  not (_33984_, _33982_);
  nor (_33985_, _33984_, _33980_);
  and (_33986_, _11608_, _03536_);
  or (_33987_, _33986_, _33985_);
  and (_33988_, _33987_, _11686_);
  and (_33989_, _33940_, _08118_);
  or (_33990_, _33989_, _33988_);
  and (_33991_, _33990_, _03209_);
  nor (_33992_, _06294_, _03209_);
  nor (_33993_, _33992_, _05998_);
  not (_33995_, _33993_);
  nor (_33996_, _33995_, _33991_);
  nor (_33997_, _33996_, _04012_);
  nand (_33998_, _33997_, _33968_);
  nand (_33999_, _33940_, _04012_);
  and (_34000_, _33999_, _04432_);
  and (_34001_, _34000_, _33998_);
  or (_34002_, _34001_, _33958_);
  nand (_34003_, _34002_, _11430_);
  nor (_34004_, _33940_, _11430_);
  nor (_34006_, _34004_, _03469_);
  nand (_34007_, _34006_, _34003_);
  and (_34008_, _11608_, _03469_);
  nor (_34009_, _34008_, _05977_);
  nand (_34010_, _34009_, _34007_);
  and (_34011_, _06294_, _05977_);
  nor (_34012_, _34011_, _03527_);
  nand (_34013_, _34012_, _34010_);
  and (_34014_, _11608_, _03527_);
  nor (_34015_, _34014_, _11716_);
  nand (_34017_, _34015_, _34013_);
  nor (_34018_, _33940_, _11715_);
  nor (_34019_, _34018_, _03530_);
  nand (_34020_, _34019_, _34017_);
  and (_34021_, _11608_, _03530_);
  nor (_34022_, _34021_, _11724_);
  nand (_34023_, _34022_, _34020_);
  nor (_34024_, _33940_, _11723_);
  nor (_34025_, _34024_, _03465_);
  nand (_34026_, _34025_, _34023_);
  and (_34028_, _11608_, _03465_);
  nor (_34029_, _34028_, _11727_);
  nand (_34030_, _34029_, _34026_);
  and (_34031_, _06294_, _11727_);
  nor (_34032_, _34031_, _03464_);
  nand (_34033_, _34032_, _34030_);
  and (_34034_, _11608_, _03464_);
  nor (_34035_, _34034_, _10021_);
  nand (_34036_, _34035_, _34033_);
  and (_34037_, _11489_, _10055_);
  nor (_34039_, _33955_, _10055_);
  or (_34040_, _34039_, _10017_);
  nor (_34041_, _34040_, _34037_);
  not (_34042_, _34041_);
  and (_34043_, _34042_, _33678_);
  nand (_34044_, _34043_, _34036_);
  and (_34045_, _11489_, _09975_);
  nor (_34046_, _33955_, _09975_);
  nor (_34047_, _34046_, _34045_);
  nor (_34048_, _34047_, _03994_);
  or (_34050_, _11490_, _11743_);
  or (_34051_, _33955_, _10116_);
  nand (_34052_, _34051_, _34050_);
  and (_34053_, _34052_, _10020_);
  nor (_34054_, _34053_, _34048_);
  nand (_34055_, _34054_, _34044_);
  nand (_34056_, _34055_, _10123_);
  and (_34057_, _33940_, _10122_);
  nand (_34058_, _33955_, _11764_);
  nand (_34059_, _11490_, _10163_);
  and (_34061_, _34059_, _03608_);
  and (_34062_, _34061_, _34058_);
  nor (_34063_, _34062_, _34057_);
  and (_34064_, _34063_, _03459_);
  nand (_34065_, _34064_, _34056_);
  and (_34066_, _11609_, _03458_);
  nor (_34067_, _34066_, _04755_);
  nand (_34068_, _34067_, _34065_);
  nor (_34069_, _06294_, _03207_);
  nor (_34070_, _34069_, _32577_);
  and (_34072_, _34070_, _34068_);
  or (_34073_, _34072_, _33949_);
  nand (_34074_, _34073_, _11424_);
  nor (_34075_, _33940_, _11424_);
  nor (_34076_, _34075_, _03587_);
  nand (_34077_, _34076_, _34074_);
  and (_34078_, _11608_, _03587_);
  nor (_34079_, _34078_, _11776_);
  nand (_34080_, _34079_, _34077_);
  and (_34081_, _06294_, _11776_);
  nor (_34083_, _34081_, _03586_);
  nand (_34084_, _34083_, _34080_);
  and (_34085_, _11608_, _03586_);
  nor (_34086_, _34085_, _11780_);
  and (_34087_, _34086_, _34084_);
  nor (_34088_, _33940_, _11419_);
  or (_34089_, _34088_, _34087_);
  nand (_34090_, _34089_, _08266_);
  nor (_34091_, _11608_, _08266_);
  nor (_34092_, _34091_, _03334_);
  nand (_34094_, _34092_, _34090_);
  nor (_34095_, _33946_, _03233_);
  nor (_34096_, _34095_, _03452_);
  and (_34097_, _34096_, _34094_);
  and (_34098_, _11609_, _03452_);
  or (_34099_, _34098_, _34097_);
  nand (_34100_, _34099_, _05919_);
  and (_34101_, _06294_, _03219_);
  nor (_34102_, _34101_, _03621_);
  nand (_34103_, _34102_, _34100_);
  and (_34105_, _11489_, _03621_);
  not (_34106_, _34105_);
  and (_34107_, _34106_, _11797_);
  nand (_34108_, _34107_, _34103_);
  nor (_34109_, _11608_, _11797_);
  nor (_34110_, _34109_, _03224_);
  nand (_34111_, _34110_, _34108_);
  and (_34112_, _11489_, _03224_);
  nor (_34113_, _34112_, _32624_);
  nand (_34114_, _34113_, _34111_);
  nor (_34116_, _33940_, _11806_);
  nor (_34117_, _34116_, _03517_);
  nand (_34118_, _34117_, _34114_);
  and (_34119_, _11608_, _03517_);
  nor (_34120_, _34119_, _03159_);
  nand (_34121_, _34120_, _34118_);
  and (_34122_, _06294_, _03159_);
  nor (_34123_, _34122_, _11813_);
  nand (_34124_, _34123_, _34121_);
  nor (_34125_, _33965_, _11814_);
  nor (_34127_, _34125_, _06193_);
  and (_34128_, _34127_, _34124_);
  nor (_34129_, _11609_, _03624_);
  nor (_34130_, _34129_, _05917_);
  or (_34131_, _34130_, _34128_);
  and (_34132_, _11489_, _03624_);
  nor (_34133_, _34132_, _08461_);
  nand (_34134_, _34133_, _34131_);
  and (_34135_, _11609_, _08461_);
  nor (_34136_, _34135_, _11828_);
  nand (_34138_, _34136_, _34134_);
  or (_34139_, _11839_, _11838_);
  nor (_34140_, _34139_, _11846_);
  nand (_34141_, _34139_, _11846_);
  nand (_34142_, _34141_, _11828_);
  or (_34143_, _34142_, _34140_);
  and (_34144_, _34143_, _04121_);
  and (_34145_, _34144_, _34138_);
  and (_34146_, _11609_, _03516_);
  or (_34147_, _34146_, _34145_);
  nand (_34148_, _34147_, _27595_);
  and (_34149_, _06294_, _03168_);
  nor (_34150_, _34149_, _11868_);
  nand (_34151_, _34150_, _34148_);
  and (_34152_, _11608_, _08864_);
  nor (_34153_, _33965_, _08864_);
  or (_34154_, _34153_, _34152_);
  and (_34155_, _34154_, _11868_);
  nor (_34156_, _34155_, _11872_);
  and (_34157_, _34156_, _34151_);
  or (_34160_, _34157_, _33948_);
  nand (_34161_, _34160_, _08493_);
  nor (_34162_, _11608_, _08493_);
  nor (_34163_, _34162_, _03623_);
  nand (_34164_, _34163_, _34161_);
  and (_34165_, _11489_, _03623_);
  nor (_34166_, _34165_, _03744_);
  and (_34167_, _34166_, _34164_);
  and (_34168_, _11609_, _03744_);
  or (_34169_, _34168_, _34167_);
  nand (_34171_, _34169_, _32199_);
  and (_34172_, _06294_, _03172_);
  nor (_34173_, _34172_, _11889_);
  nand (_34174_, _34173_, _34171_);
  and (_34175_, _33965_, _08864_);
  nor (_34176_, _11608_, _08864_);
  nor (_34177_, _34176_, _11893_);
  not (_34178_, _34177_);
  nor (_34179_, _34178_, _34175_);
  nor (_34180_, _34179_, _11901_);
  and (_34182_, _34180_, _34174_);
  or (_34183_, _34182_, _33947_);
  nand (_34184_, _34183_, _11904_);
  nor (_34185_, _11608_, _11904_);
  nor (_34186_, _34185_, _03611_);
  nand (_34187_, _34186_, _34184_);
  and (_34188_, _11489_, _03611_);
  nor (_34189_, _34188_, _03733_);
  and (_34190_, _34189_, _34187_);
  and (_34191_, _11609_, _03733_);
  or (_34193_, _34191_, _34190_);
  nand (_34194_, _34193_, _32195_);
  and (_34195_, _06294_, _03182_);
  nor (_34196_, _34195_, _11915_);
  nand (_34197_, _34196_, _34194_);
  and (_34198_, _33965_, _07982_);
  nor (_34199_, _11608_, _07982_);
  nor (_34200_, _34199_, _24078_);
  not (_34201_, _34200_);
  nor (_34202_, _34201_, _34198_);
  nor (_34204_, _34202_, _11919_);
  and (_34205_, _34204_, _34197_);
  or (_34206_, _34205_, _33945_);
  nand (_34207_, _34206_, _11410_);
  nor (_34208_, _11608_, _11410_);
  nor (_34209_, _34208_, _03618_);
  nand (_34210_, _34209_, _34207_);
  and (_34211_, _11489_, _03618_);
  nor (_34212_, _34211_, _03741_);
  and (_34213_, _34212_, _34210_);
  and (_34215_, _11609_, _03741_);
  or (_34216_, _34215_, _34213_);
  nand (_34217_, _34216_, _32192_);
  and (_34218_, _06294_, _03178_);
  nor (_34219_, _34218_, _11936_);
  nand (_34220_, _34219_, _34217_);
  and (_34221_, _33965_, \oc8051_golden_model_1.PSW [7]);
  nor (_34222_, _11608_, \oc8051_golden_model_1.PSW [7]);
  nor (_34223_, _34222_, _11942_);
  not (_34224_, _34223_);
  nor (_34226_, _34224_, _34221_);
  nor (_34227_, _34226_, _11940_);
  and (_34228_, _34227_, _34220_);
  or (_34229_, _34228_, _33944_);
  nand (_34230_, _34229_, _08628_);
  nor (_34231_, _11608_, _08628_);
  nor (_34232_, _34231_, _08707_);
  nand (_34233_, _34232_, _34230_);
  and (_34234_, _33940_, _08707_);
  nor (_34235_, _34234_, _03752_);
  and (_34237_, _34235_, _34233_);
  nor (_34238_, _06757_, _10735_);
  or (_34239_, _34238_, _34237_);
  nand (_34240_, _34239_, _04803_);
  and (_34241_, _06294_, _03191_);
  nor (_34242_, _34241_, _03617_);
  nand (_34243_, _34242_, _34240_);
  and (_34244_, _33955_, _09953_);
  nor (_34245_, _11489_, _09953_);
  or (_34246_, _34245_, _03814_);
  or (_34248_, _34246_, _34244_);
  and (_34249_, _34248_, _11406_);
  and (_34250_, _34249_, _34243_);
  or (_34251_, _34250_, _33943_);
  nand (_34252_, _34251_, _08784_);
  nor (_34253_, _11608_, _08784_);
  nor (_34254_, _34253_, _08815_);
  nand (_34255_, _34254_, _34252_);
  and (_34256_, _33940_, _08815_);
  nor (_34257_, _34256_, _03475_);
  and (_34259_, _34257_, _34255_);
  nor (_34260_, _06757_, _03476_);
  or (_34261_, _34260_, _34259_);
  nand (_34262_, _34261_, _11405_);
  and (_34263_, _06294_, _03189_);
  nor (_34264_, _34263_, _03644_);
  nand (_34265_, _34264_, _34262_);
  and (_34266_, _11489_, _09953_);
  nor (_34267_, _33955_, _09953_);
  or (_34268_, _34267_, _34266_);
  and (_34270_, _34268_, _03644_);
  nor (_34271_, _34270_, _11992_);
  nand (_34272_, _34271_, _34265_);
  nor (_34273_, _33940_, _11991_);
  nor (_34274_, _34273_, _03767_);
  nand (_34275_, _34274_, _34272_);
  and (_34276_, _11608_, _03767_);
  nor (_34277_, _34276_, _11999_);
  and (_34278_, _34277_, _34275_);
  nor (_34279_, _33940_, _11998_);
  or (_34281_, _34279_, _34278_);
  nand (_34282_, _34281_, _04553_);
  and (_34283_, _06294_, _04986_);
  nor (_34284_, _34283_, _03445_);
  nand (_34285_, _34284_, _34282_);
  and (_34286_, _34268_, _03445_);
  nor (_34287_, _34286_, _12016_);
  nand (_34288_, _34287_, _34285_);
  nor (_34289_, _33940_, _12015_);
  nor (_34290_, _34289_, _03473_);
  and (_34292_, _34290_, _34288_);
  or (_34293_, _34292_, _33942_);
  nand (_34294_, _34293_, _11392_);
  nor (_34295_, _33946_, _11392_);
  nor (_34296_, _34295_, _32181_);
  nand (_34297_, _34296_, _34294_);
  and (_34298_, _32181_, _06294_);
  nor (_34299_, _34298_, _12031_);
  and (_34300_, _34299_, _34297_);
  or (_34301_, _34300_, _33941_);
  or (_34303_, _34301_, _43193_);
  or (_34304_, _43189_, \oc8051_golden_model_1.PC [5]);
  and (_34305_, _34304_, _42003_);
  and (_43925_, _34305_, _34303_);
  and (_34306_, _32181_, _06262_);
  and (_34307_, _06262_, _04986_);
  and (_34308_, _05903_, _11393_);
  nor (_34309_, _34308_, \oc8051_golden_model_1.PC [6]);
  nor (_34310_, _34309_, _11394_);
  not (_34311_, _34310_);
  and (_34313_, _34311_, _08815_);
  and (_34314_, _11482_, _03618_);
  and (_34315_, _11482_, _03611_);
  and (_34316_, _11482_, _03623_);
  and (_34317_, _11601_, _03516_);
  and (_34318_, _11482_, _03621_);
  and (_34319_, _06262_, _04435_);
  and (_34320_, _11601_, _04436_);
  or (_34321_, _34320_, _08108_);
  nand (_34322_, _11688_, \oc8051_golden_model_1.PC [6]);
  and (_34324_, _34322_, _04437_);
  or (_34325_, _34324_, _34321_);
  or (_34326_, _34311_, _11683_);
  and (_34327_, _34326_, _03204_);
  and (_34328_, _34327_, _34325_);
  or (_34329_, _34328_, _15022_);
  or (_34330_, _34329_, _34319_);
  or (_34331_, _34311_, _11680_);
  and (_34332_, _34331_, _08101_);
  and (_34333_, _34332_, _34330_);
  and (_34335_, _11601_, _03536_);
  or (_34336_, _34335_, _34333_);
  nor (_34337_, _34336_, _08118_);
  and (_34338_, _34310_, _08118_);
  or (_34339_, _34338_, _34337_);
  and (_34340_, _34339_, _03209_);
  nor (_34341_, _06262_, _03209_);
  nor (_34342_, _34341_, _05998_);
  not (_34343_, _34342_);
  nor (_34344_, _34343_, _34340_);
  and (_34346_, _11639_, _11605_);
  nor (_34347_, _34346_, _11640_);
  nand (_34348_, _34347_, _32232_);
  or (_34349_, _32232_, _11601_);
  and (_34350_, _34349_, _34348_);
  and (_34351_, _34350_, _05998_);
  or (_34352_, _34351_, _34344_);
  nand (_34353_, _34352_, _06008_);
  and (_34354_, _34311_, _04012_);
  nor (_34355_, _34354_, _03534_);
  nand (_34357_, _34355_, _34353_);
  and (_34358_, _11525_, _11486_);
  nor (_34359_, _34358_, _11526_);
  or (_34360_, _34359_, _11437_);
  or (_34361_, _11481_, _11439_);
  and (_34362_, _34361_, _03534_);
  nand (_34363_, _34362_, _34360_);
  nand (_34364_, _34363_, _34357_);
  nand (_34365_, _34364_, _11430_);
  nor (_34366_, _34311_, _11430_);
  nor (_34368_, _34366_, _03469_);
  nand (_34369_, _34368_, _34365_);
  and (_34370_, _11601_, _03469_);
  nor (_34371_, _34370_, _05977_);
  nand (_34372_, _34371_, _34369_);
  nor (_34373_, _06262_, _03202_);
  nor (_34374_, _34373_, _03527_);
  and (_34375_, _34374_, _34372_);
  and (_34376_, _11601_, _03527_);
  or (_34377_, _34376_, _34375_);
  and (_34379_, _34377_, _11715_);
  nor (_34380_, _34310_, _11715_);
  or (_34381_, _34380_, _34379_);
  nand (_34382_, _34381_, _03531_);
  and (_34383_, _11601_, _03530_);
  nor (_34384_, _34383_, _11724_);
  and (_34385_, _34384_, _34382_);
  nor (_34386_, _34311_, _11723_);
  or (_34387_, _34386_, _03465_);
  nor (_34388_, _34387_, _34385_);
  and (_34390_, _11601_, _03465_);
  or (_34391_, _34390_, _34388_);
  nand (_34392_, _34391_, _03212_);
  and (_34393_, _06262_, _11727_);
  nor (_34394_, _34393_, _03464_);
  nand (_34395_, _34394_, _34392_);
  and (_34396_, _11600_, _03464_);
  nor (_34397_, _34396_, _10021_);
  and (_34398_, _34397_, _34395_);
  and (_34399_, _11481_, _10055_);
  not (_34401_, _34359_);
  nor (_34402_, _34401_, _10055_);
  or (_34403_, _34402_, _34399_);
  nor (_34404_, _34403_, _10017_);
  or (_34405_, _34404_, _34398_);
  nand (_34406_, _34405_, _10112_);
  and (_34407_, _11481_, _10116_);
  nor (_34408_, _03648_, _03630_);
  and (_34409_, _34359_, _11743_);
  or (_34410_, _34409_, _34408_);
  or (_34412_, _34410_, _34407_);
  and (_34413_, _34412_, _03994_);
  nand (_34414_, _34413_, _34406_);
  and (_34415_, _11482_, _09975_);
  nor (_34416_, _34359_, _09975_);
  or (_34417_, _34416_, _03994_);
  or (_34418_, _34417_, _34415_);
  nand (_34419_, _34418_, _34414_);
  nand (_34420_, _34419_, _10123_);
  and (_34421_, _34310_, _10122_);
  or (_34423_, _34359_, _10163_);
  nand (_34424_, _11482_, _10163_);
  and (_34425_, _34424_, _03608_);
  and (_34426_, _34425_, _34423_);
  nor (_34427_, _34426_, _34421_);
  and (_34428_, _34427_, _03459_);
  and (_34429_, _34428_, _34420_);
  and (_34430_, _11601_, _03458_);
  or (_34431_, _34430_, _34429_);
  nand (_34432_, _34431_, _03207_);
  and (_34434_, _06262_, _04755_);
  nor (_34435_, _34434_, _32577_);
  nand (_34436_, _34435_, _34432_);
  nor (_34437_, _32576_, _11601_);
  nor (_34438_, _34437_, _11425_);
  and (_34439_, _34438_, _34436_);
  nor (_34440_, _34310_, _11424_);
  or (_34441_, _34440_, _34439_);
  nand (_34442_, _34441_, _09769_);
  and (_34443_, _11601_, _03587_);
  nor (_34445_, _34443_, _11776_);
  nand (_34446_, _34445_, _34442_);
  nor (_34447_, _06262_, _03214_);
  nor (_34448_, _34447_, _03586_);
  nand (_34449_, _34448_, _34446_);
  and (_34450_, _11601_, _03586_);
  nor (_34451_, _34450_, _11780_);
  nand (_34452_, _34451_, _34449_);
  nor (_34453_, _34311_, _11419_);
  nor (_34454_, _34453_, _08267_);
  nand (_34456_, _34454_, _34452_);
  nor (_34457_, _11600_, _08266_);
  nor (_34458_, _34457_, _03334_);
  nand (_34459_, _34458_, _34456_);
  nor (_34460_, _34311_, _03233_);
  nor (_34461_, _34460_, _03452_);
  nand (_34462_, _34461_, _34459_);
  and (_34463_, _11601_, _03452_);
  nor (_34464_, _34463_, _03219_);
  nand (_34465_, _34464_, _34462_);
  nor (_34467_, _06262_, _05919_);
  nor (_34468_, _34467_, _03621_);
  nand (_34469_, _34468_, _34465_);
  nand (_34470_, _34469_, _11797_);
  or (_34471_, _34470_, _34318_);
  nor (_34472_, _11601_, _11797_);
  nor (_34473_, _34472_, _03224_);
  nand (_34474_, _34473_, _34471_);
  and (_34475_, _11482_, _03224_);
  nor (_34476_, _34475_, _32624_);
  nand (_34478_, _34476_, _34474_);
  nor (_34479_, _34311_, _11806_);
  nor (_34480_, _34479_, _03517_);
  nand (_34481_, _34480_, _34478_);
  and (_34482_, _11601_, _03517_);
  nor (_34483_, _34482_, _03159_);
  and (_34484_, _34483_, _34481_);
  nor (_34485_, _06262_, _03160_);
  or (_34486_, _34485_, _34484_);
  and (_34487_, _34486_, _11814_);
  and (_34489_, _34347_, _11813_);
  or (_34490_, _34489_, _34487_);
  nand (_34491_, _34490_, _05916_);
  nor (_34492_, _11601_, _05916_);
  nor (_34493_, _34492_, _03624_);
  nand (_34494_, _34493_, _34491_);
  and (_34495_, _11482_, _03624_);
  nor (_34496_, _34495_, _08461_);
  nand (_34497_, _34496_, _34494_);
  and (_34498_, _11600_, _08461_);
  nor (_34500_, _34498_, _11828_);
  and (_34501_, _34500_, _34497_);
  and (_34502_, _11848_, _11837_);
  nor (_34503_, _34502_, _11849_);
  nor (_34504_, _34503_, _23814_);
  or (_34505_, _34504_, _34501_);
  and (_34506_, _34505_, _04121_);
  or (_34507_, _34506_, _34317_);
  nand (_34508_, _34507_, _27595_);
  and (_34509_, _06262_, _03168_);
  nor (_34511_, _34509_, _11868_);
  nand (_34512_, _34511_, _34508_);
  and (_34513_, _11600_, _08864_);
  and (_34514_, _34347_, _11894_);
  or (_34515_, _34514_, _34513_);
  and (_34516_, _34515_, _11868_);
  nor (_34517_, _34516_, _11872_);
  nand (_34518_, _34517_, _34512_);
  nor (_34519_, _34310_, _11416_);
  nor (_34520_, _34519_, _08494_);
  nand (_34522_, _34520_, _34518_);
  nor (_34523_, _11601_, _08493_);
  nor (_34524_, _34523_, _03623_);
  and (_34525_, _34524_, _34522_);
  or (_34526_, _34525_, _34316_);
  nand (_34527_, _34526_, _03745_);
  and (_34528_, _11601_, _03744_);
  nor (_34529_, _34528_, _03172_);
  and (_34530_, _34529_, _34527_);
  nor (_34531_, _06262_, _32199_);
  or (_34533_, _34531_, _34530_);
  nand (_34534_, _34533_, _11893_);
  nor (_34535_, _34347_, _11894_);
  nor (_34536_, _11600_, _08864_);
  nor (_34537_, _34536_, _11893_);
  not (_34538_, _34537_);
  nor (_34539_, _34538_, _34535_);
  nor (_34540_, _34539_, _11901_);
  nand (_34541_, _34540_, _34534_);
  and (_34542_, _34311_, _11901_);
  nor (_34544_, _34542_, _11905_);
  nand (_34545_, _34544_, _34541_);
  nor (_34546_, _11601_, _11904_);
  nor (_34547_, _34546_, _03611_);
  and (_34548_, _34547_, _34545_);
  or (_34549_, _34548_, _34315_);
  nand (_34550_, _34549_, _03734_);
  and (_34551_, _11601_, _03733_);
  nor (_34552_, _34551_, _03182_);
  and (_34553_, _34552_, _34550_);
  nor (_34555_, _06262_, _32195_);
  or (_34556_, _34555_, _34553_);
  nand (_34557_, _34556_, _24078_);
  and (_34558_, _11600_, \oc8051_golden_model_1.PSW [7]);
  and (_34559_, _34347_, _07982_);
  or (_34560_, _34559_, _34558_);
  and (_34561_, _34560_, _11915_);
  nor (_34562_, _34561_, _11919_);
  nand (_34563_, _34562_, _34557_);
  nor (_34564_, _34310_, _11413_);
  nor (_34566_, _34564_, _15156_);
  nand (_34567_, _34566_, _34563_);
  nor (_34568_, _11601_, _11410_);
  nor (_34569_, _34568_, _03618_);
  and (_34570_, _34569_, _34567_);
  or (_34571_, _34570_, _34314_);
  nand (_34572_, _34571_, _06458_);
  and (_34573_, _11601_, _03741_);
  nor (_34574_, _34573_, _03178_);
  and (_34575_, _34574_, _34572_);
  nor (_34577_, _06262_, _32192_);
  or (_34578_, _34577_, _34575_);
  nand (_34579_, _34578_, _11942_);
  nor (_34580_, _34347_, _07982_);
  nor (_34581_, _11600_, \oc8051_golden_model_1.PSW [7]);
  nor (_34582_, _34581_, _11942_);
  not (_34583_, _34582_);
  nor (_34584_, _34583_, _34580_);
  nor (_34585_, _34584_, _11940_);
  nand (_34586_, _34585_, _34579_);
  nor (_34588_, _34310_, _11408_);
  nor (_34589_, _34588_, _08629_);
  nand (_34590_, _34589_, _34586_);
  nor (_34591_, _11601_, _08628_);
  nor (_34592_, _34591_, _08707_);
  nand (_34593_, _34592_, _34590_);
  and (_34594_, _34311_, _08707_);
  nor (_34595_, _34594_, _03752_);
  nand (_34596_, _34595_, _34593_);
  and (_34597_, _06526_, _03752_);
  nor (_34599_, _34597_, _03191_);
  nand (_34600_, _34599_, _34596_);
  and (_34601_, _06262_, _03191_);
  nor (_34602_, _34601_, _03617_);
  nand (_34603_, _34602_, _34600_);
  and (_34604_, _34401_, _09953_);
  nor (_34605_, _11481_, _09953_);
  or (_34606_, _34605_, _03814_);
  nor (_34607_, _34606_, _34604_);
  nor (_34608_, _34607_, _11963_);
  nand (_34610_, _34608_, _34603_);
  nor (_34611_, _34310_, _11406_);
  nor (_34612_, _34611_, _08785_);
  nand (_34613_, _34612_, _34610_);
  nor (_34614_, _11601_, _08784_);
  nor (_34615_, _34614_, _08815_);
  and (_34616_, _34615_, _34613_);
  or (_34617_, _34616_, _34313_);
  nand (_34618_, _34617_, _03476_);
  nor (_34619_, _06526_, _03476_);
  nor (_34621_, _34619_, _03189_);
  nand (_34622_, _34621_, _34618_);
  nor (_34623_, _06262_, _11405_);
  nor (_34624_, _34623_, _03644_);
  and (_34625_, _34624_, _34622_);
  and (_34626_, _11482_, _09953_);
  nor (_34627_, _34359_, _09953_);
  nor (_34628_, _34627_, _34626_);
  nor (_34629_, _34628_, _03768_);
  or (_34630_, _34629_, _34625_);
  and (_34632_, _34630_, _11991_);
  nor (_34633_, _34310_, _11991_);
  or (_34634_, _34633_, _34632_);
  nand (_34635_, _34634_, _03948_);
  and (_34636_, _11601_, _03767_);
  nor (_34637_, _34636_, _11999_);
  nand (_34638_, _34637_, _34635_);
  nor (_34639_, _34311_, _11998_);
  nor (_34640_, _34639_, _04986_);
  and (_34641_, _34640_, _34638_);
  or (_34643_, _34641_, _34307_);
  nand (_34644_, _34643_, _03446_);
  nor (_34645_, _34628_, _03446_);
  nor (_34646_, _34645_, _12016_);
  nand (_34647_, _34646_, _34644_);
  nor (_34648_, _34311_, _12015_);
  nor (_34649_, _34648_, _03473_);
  nand (_34650_, _34649_, _34647_);
  and (_34651_, _11601_, _03473_);
  nor (_34652_, _34651_, _12022_);
  nand (_34654_, _34652_, _34650_);
  nor (_34655_, _34311_, _11392_);
  nor (_34656_, _34655_, _32181_);
  and (_34657_, _34656_, _34654_);
  or (_34658_, _34657_, _34306_);
  nand (_34659_, _34658_, _12035_);
  and (_34660_, _34311_, _12031_);
  not (_34661_, _34660_);
  and (_34662_, _34661_, _34659_);
  or (_34663_, _34662_, _43193_);
  or (_34665_, _43189_, \oc8051_golden_model_1.PC [6]);
  and (_34666_, _34665_, _42003_);
  and (_43926_, _34666_, _34663_);
  and (_34667_, _05908_, _03473_);
  nor (_34668_, _11394_, \oc8051_golden_model_1.PC [7]);
  nor (_34669_, _34668_, _11395_);
  nor (_34670_, _34669_, _11406_);
  nor (_34671_, _34669_, _11408_);
  nor (_34672_, _34669_, _11413_);
  not (_34673_, _34669_);
  and (_34675_, _34673_, _11901_);
  nor (_34676_, _34669_, _11416_);
  nor (_34677_, _32576_, _05908_);
  or (_34678_, _11439_, _06821_);
  or (_34679_, _11477_, _11478_);
  and (_34680_, _34679_, _11527_);
  nor (_34681_, _34679_, _11527_);
  nor (_34682_, _34681_, _34680_);
  not (_34683_, _34682_);
  or (_34684_, _34683_, _11437_);
  and (_34686_, _34684_, _03534_);
  and (_34687_, _34686_, _34678_);
  and (_34688_, _11566_, _05908_);
  or (_34689_, _11596_, _11597_);
  and (_34690_, _34689_, _11641_);
  nor (_34691_, _34689_, _11641_);
  nor (_34692_, _34691_, _34690_);
  and (_34693_, _34692_, _32232_);
  nor (_34694_, _34693_, _34688_);
  nand (_34695_, _34694_, _05998_);
  nor (_34697_, _06226_, _03204_);
  and (_34698_, _05909_, _04436_);
  nor (_34699_, _34698_, _08108_);
  and (_34700_, _11688_, \oc8051_golden_model_1.PC [7]);
  or (_34701_, _34700_, _04436_);
  and (_34702_, _34701_, _34699_);
  nor (_34703_, _34673_, _11683_);
  or (_34704_, _34703_, _15022_);
  or (_34705_, _34704_, _34702_);
  and (_34706_, _34705_, _03204_);
  nor (_34708_, _34706_, _34697_);
  nor (_34709_, _34669_, _11680_);
  nor (_34710_, _34709_, _03536_);
  not (_34711_, _34710_);
  nor (_34712_, _34711_, _34708_);
  and (_34713_, _05908_, _03536_);
  or (_34714_, _34713_, _34712_);
  and (_34715_, _34714_, _11686_);
  and (_34716_, _34669_, _08118_);
  or (_34717_, _34716_, _34715_);
  and (_34719_, _34717_, _03209_);
  nor (_34720_, _06226_, _03209_);
  nor (_34721_, _34720_, _05998_);
  not (_34722_, _34721_);
  nor (_34723_, _34722_, _34719_);
  nor (_34724_, _34723_, _04012_);
  nand (_34725_, _34724_, _34695_);
  nand (_34726_, _34669_, _04012_);
  and (_34727_, _34726_, _04432_);
  and (_34728_, _34727_, _34725_);
  or (_34730_, _34728_, _34687_);
  nand (_34731_, _34730_, _11430_);
  nor (_34732_, _34669_, _11430_);
  nor (_34733_, _34732_, _03469_);
  nand (_34734_, _34733_, _34731_);
  and (_34735_, _05908_, _03469_);
  nor (_34736_, _34735_, _05977_);
  nand (_34737_, _34736_, _34734_);
  and (_34738_, _06226_, _05977_);
  nor (_34739_, _34738_, _03527_);
  nand (_34741_, _34739_, _34737_);
  and (_34742_, _05908_, _03527_);
  nor (_34743_, _34742_, _11716_);
  nand (_34744_, _34743_, _34741_);
  nor (_34745_, _34669_, _11715_);
  nor (_34746_, _34745_, _03530_);
  nand (_34747_, _34746_, _34744_);
  and (_34748_, _05908_, _03530_);
  nor (_34749_, _34748_, _11724_);
  nand (_34750_, _34749_, _34747_);
  nor (_34752_, _34669_, _11723_);
  nor (_34753_, _34752_, _03465_);
  nand (_34754_, _34753_, _34750_);
  and (_34755_, _05908_, _03465_);
  nor (_34756_, _34755_, _11727_);
  nand (_34757_, _34756_, _34754_);
  and (_34758_, _06226_, _11727_);
  nor (_34759_, _34758_, _03464_);
  nand (_34760_, _34759_, _34757_);
  and (_34761_, _05908_, _03464_);
  nor (_34763_, _34761_, _10021_);
  nand (_34764_, _34763_, _34760_);
  and (_34765_, _10055_, _06820_);
  nor (_34766_, _34683_, _10055_);
  or (_34767_, _34766_, _34765_);
  nor (_34768_, _34767_, _10017_);
  nor (_34769_, _34768_, _10020_);
  nand (_34770_, _34769_, _34764_);
  or (_34771_, _34683_, _10116_);
  or (_34772_, _11743_, _06821_);
  and (_34773_, _34772_, _34771_);
  or (_34774_, _34773_, _10112_);
  and (_34775_, _34774_, _03994_);
  and (_34776_, _34775_, _34770_);
  nor (_34777_, _34683_, _09975_);
  and (_34778_, _09975_, _06820_);
  or (_34779_, _34778_, _03994_);
  nor (_34780_, _34779_, _34777_);
  or (_34781_, _34780_, _10124_);
  or (_34782_, _34781_, _34776_);
  nor (_34785_, _34682_, _10163_);
  and (_34786_, _10163_, _06821_);
  nor (_34787_, _34786_, _10158_);
  not (_34788_, _34787_);
  nor (_34789_, _34788_, _34785_);
  and (_34790_, _34669_, _10122_);
  nor (_34791_, _34790_, _34789_);
  and (_34792_, _34791_, _03459_);
  nand (_34793_, _34792_, _34782_);
  and (_34794_, _05909_, _03458_);
  nor (_34796_, _34794_, _04755_);
  nand (_34797_, _34796_, _34793_);
  nor (_34798_, _06226_, _03207_);
  nor (_34799_, _34798_, _32577_);
  and (_34800_, _34799_, _34797_);
  or (_34801_, _34800_, _34677_);
  nand (_34802_, _34801_, _11424_);
  nor (_34803_, _34669_, _11424_);
  nor (_34804_, _34803_, _03587_);
  nand (_34805_, _34804_, _34802_);
  and (_34807_, _05908_, _03587_);
  nor (_34808_, _34807_, _11776_);
  nand (_34809_, _34808_, _34805_);
  and (_34810_, _06226_, _11776_);
  nor (_34811_, _34810_, _03586_);
  nand (_34812_, _34811_, _34809_);
  and (_34813_, _05908_, _03586_);
  nor (_34814_, _34813_, _11780_);
  and (_34815_, _34814_, _34812_);
  nor (_34816_, _34669_, _11419_);
  or (_34818_, _34816_, _34815_);
  nand (_34819_, _34818_, _08266_);
  nor (_34820_, _08266_, _05908_);
  nor (_34821_, _34820_, _03334_);
  nand (_34822_, _34821_, _34819_);
  nor (_34823_, _34673_, _03233_);
  nor (_34824_, _34823_, _03452_);
  and (_34825_, _34824_, _34822_);
  and (_34826_, _05909_, _03452_);
  or (_34827_, _34826_, _34825_);
  nand (_34829_, _34827_, _05919_);
  and (_34830_, _06226_, _03219_);
  nor (_34831_, _34830_, _03621_);
  nand (_34832_, _34831_, _34829_);
  and (_34833_, _06820_, _03621_);
  not (_34834_, _34833_);
  and (_34835_, _34834_, _11797_);
  nand (_34836_, _34835_, _34832_);
  nor (_34837_, _11797_, _05908_);
  nor (_34838_, _34837_, _03224_);
  nand (_34840_, _34838_, _34836_);
  and (_34841_, _06820_, _03224_);
  nor (_34842_, _34841_, _32624_);
  nand (_34843_, _34842_, _34840_);
  nor (_34844_, _34669_, _11806_);
  nor (_34845_, _34844_, _03517_);
  nand (_34846_, _34845_, _34843_);
  and (_34847_, _05908_, _03517_);
  nor (_34848_, _34847_, _03159_);
  nand (_34849_, _34848_, _34846_);
  and (_34851_, _06226_, _03159_);
  nor (_34852_, _34851_, _11813_);
  nand (_34853_, _34852_, _34849_);
  and (_34854_, _34692_, _11813_);
  nor (_34855_, _34854_, _06193_);
  and (_34856_, _34855_, _34853_);
  nor (_34857_, _05909_, _03624_);
  nor (_34858_, _34857_, _05917_);
  or (_34859_, _34858_, _34856_);
  and (_34860_, _06820_, _03624_);
  nor (_34862_, _34860_, _08461_);
  nand (_34863_, _34862_, _34859_);
  and (_34864_, _08461_, _05909_);
  nor (_34865_, _34864_, _11828_);
  nand (_34866_, _34865_, _34863_);
  or (_34867_, _11832_, _11833_);
  nor (_34868_, _34867_, _11850_);
  and (_34869_, _34867_, _11850_);
  nor (_34870_, _34869_, _34868_);
  and (_34871_, _34870_, _11828_);
  nor (_34873_, _34871_, _03516_);
  and (_34874_, _34873_, _34866_);
  and (_34875_, _05909_, _03516_);
  or (_34876_, _34875_, _34874_);
  nand (_34877_, _34876_, _27595_);
  and (_34878_, _06226_, _03168_);
  nor (_34879_, _34878_, _11868_);
  nand (_34880_, _34879_, _34877_);
  and (_34881_, _08864_, _05908_);
  and (_34882_, _34692_, _11894_);
  or (_34884_, _34882_, _34881_);
  and (_34885_, _34884_, _11868_);
  nor (_34886_, _34885_, _11872_);
  and (_34887_, _34886_, _34880_);
  or (_34888_, _34887_, _34676_);
  nand (_34889_, _34888_, _08493_);
  nor (_34890_, _08493_, _05908_);
  nor (_34891_, _34890_, _03623_);
  nand (_34892_, _34891_, _34889_);
  and (_34893_, _06820_, _03623_);
  nor (_34895_, _34893_, _03744_);
  and (_34896_, _34895_, _34892_);
  and (_34897_, _05909_, _03744_);
  or (_34898_, _34897_, _34896_);
  nand (_34899_, _34898_, _32199_);
  and (_34900_, _06226_, _03172_);
  nor (_34901_, _34900_, _11889_);
  nand (_34902_, _34901_, _34899_);
  nor (_34903_, _34692_, _11894_);
  nor (_34904_, _08864_, _05908_);
  nor (_34906_, _34904_, _11893_);
  not (_34907_, _34906_);
  nor (_34908_, _34907_, _34903_);
  nor (_34909_, _34908_, _11901_);
  and (_34910_, _34909_, _34902_);
  or (_34911_, _34910_, _34675_);
  nand (_34912_, _34911_, _11904_);
  nor (_34913_, _11904_, _05908_);
  nor (_34914_, _34913_, _03611_);
  nand (_34915_, _34914_, _34912_);
  and (_34917_, _06820_, _03611_);
  nor (_34918_, _34917_, _03733_);
  and (_34919_, _34918_, _34915_);
  and (_34920_, _05909_, _03733_);
  or (_34921_, _34920_, _34919_);
  nand (_34922_, _34921_, _32195_);
  and (_34923_, _06226_, _03182_);
  nor (_34924_, _34923_, _11915_);
  nand (_34925_, _34924_, _34922_);
  and (_34926_, _05908_, \oc8051_golden_model_1.PSW [7]);
  and (_34928_, _34692_, _07982_);
  or (_34929_, _34928_, _34926_);
  and (_34930_, _34929_, _11915_);
  nor (_34931_, _34930_, _11919_);
  and (_34932_, _34931_, _34925_);
  or (_34933_, _34932_, _34672_);
  nand (_34934_, _34933_, _11410_);
  nor (_34935_, _11410_, _05908_);
  nor (_34936_, _34935_, _03618_);
  nand (_34937_, _34936_, _34934_);
  and (_34939_, _06820_, _03618_);
  nor (_34940_, _34939_, _03741_);
  and (_34941_, _34940_, _34937_);
  and (_34942_, _05909_, _03741_);
  or (_34943_, _34942_, _34941_);
  nand (_34944_, _34943_, _32192_);
  and (_34945_, _06226_, _03178_);
  nor (_34946_, _34945_, _11936_);
  nand (_34947_, _34946_, _34944_);
  nor (_34948_, _34692_, _07982_);
  nor (_34950_, _05908_, \oc8051_golden_model_1.PSW [7]);
  nor (_34951_, _34950_, _11942_);
  not (_34952_, _34951_);
  nor (_34953_, _34952_, _34948_);
  nor (_34954_, _34953_, _11940_);
  and (_34955_, _34954_, _34947_);
  or (_34956_, _34955_, _34671_);
  nand (_34957_, _34956_, _08628_);
  nor (_34958_, _08628_, _05908_);
  nor (_34959_, _34958_, _08707_);
  nand (_34961_, _34959_, _34957_);
  and (_34962_, _34669_, _08707_);
  nor (_34963_, _34962_, _03752_);
  and (_34964_, _34963_, _34961_);
  nor (_34965_, _06114_, _10735_);
  or (_34966_, _34965_, _34964_);
  nand (_34967_, _34966_, _04803_);
  and (_34968_, _06226_, _03191_);
  nor (_34969_, _34968_, _03617_);
  nand (_34970_, _34969_, _34967_);
  and (_34972_, _34683_, _09953_);
  nor (_34973_, _09953_, _06820_);
  or (_34974_, _34973_, _03814_);
  or (_34975_, _34974_, _34972_);
  and (_34976_, _34975_, _11406_);
  and (_34977_, _34976_, _34970_);
  or (_34978_, _34977_, _34670_);
  nand (_34979_, _34978_, _08784_);
  nor (_34980_, _08784_, _05908_);
  nor (_34981_, _34980_, _08815_);
  nand (_34983_, _34981_, _34979_);
  and (_34984_, _34669_, _08815_);
  nor (_34985_, _34984_, _03475_);
  and (_34986_, _34985_, _34983_);
  nor (_34987_, _06114_, _03476_);
  or (_34988_, _34987_, _34986_);
  nand (_34989_, _34988_, _11405_);
  and (_34990_, _06226_, _03189_);
  nor (_34991_, _34990_, _03644_);
  nand (_34992_, _34991_, _34989_);
  nor (_34994_, _34682_, _09953_);
  and (_34995_, _09953_, _06821_);
  nor (_34996_, _34995_, _34994_);
  and (_34997_, _34996_, _03644_);
  nor (_34998_, _34997_, _11992_);
  nand (_34999_, _34998_, _34992_);
  nor (_35000_, _34669_, _11991_);
  nor (_35001_, _35000_, _03767_);
  nand (_35002_, _35001_, _34999_);
  and (_35003_, _05908_, _03767_);
  nor (_35005_, _35003_, _11999_);
  and (_35006_, _35005_, _35002_);
  nor (_35007_, _34669_, _11998_);
  or (_35008_, _35007_, _35006_);
  nand (_35009_, _35008_, _04553_);
  and (_35010_, _06226_, _04986_);
  nor (_35011_, _35010_, _03445_);
  nand (_35012_, _35011_, _35009_);
  and (_35013_, _34996_, _03445_);
  nor (_35014_, _35013_, _12016_);
  nand (_35016_, _35014_, _35012_);
  nor (_35017_, _34669_, _12015_);
  nor (_35018_, _35017_, _03473_);
  and (_35019_, _35018_, _35016_);
  or (_35020_, _35019_, _34667_);
  nand (_35021_, _35020_, _11392_);
  nor (_35022_, _34673_, _11392_);
  nor (_35023_, _35022_, _32181_);
  nand (_35024_, _35023_, _35021_);
  and (_35025_, _32181_, _06226_);
  nor (_35027_, _35025_, _12031_);
  nand (_35028_, _35027_, _35024_);
  and (_35029_, _34669_, _12031_);
  not (_35030_, _35029_);
  and (_35031_, _35030_, _35028_);
  nand (_35032_, _35031_, _43189_);
  or (_35033_, _43189_, \oc8051_golden_model_1.PC [7]);
  and (_35034_, _35033_, _42003_);
  and (_43927_, _35034_, _35032_);
  nor (_35035_, _12031_, _03194_);
  nor (_35037_, _03989_, _11391_);
  nor (_35038_, _03989_, _06855_);
  nor (_35039_, _11936_, _03178_);
  nor (_35040_, _11813_, _03159_);
  and (_35041_, _11645_, _03517_);
  and (_35042_, _11645_, _03465_);
  nor (_35043_, _03527_, _05977_);
  and (_35044_, _11645_, _03469_);
  nor (_35045_, _11535_, _11529_);
  nor (_35046_, _35045_, _11536_);
  or (_35048_, _35046_, _11437_);
  or (_35049_, _11531_, _11439_);
  and (_35050_, _35049_, _35048_);
  or (_35051_, _35050_, _04432_);
  and (_35052_, _11566_, _11645_);
  nor (_35053_, _11648_, _11643_);
  nor (_35054_, _35053_, _11649_);
  and (_35055_, _35054_, _32232_);
  nor (_35056_, _35055_, _35052_);
  nand (_35057_, _35056_, _05998_);
  and (_35059_, _11395_, \oc8051_golden_model_1.PC [8]);
  nor (_35060_, _11395_, \oc8051_golden_model_1.PC [8]);
  nor (_35061_, _35060_, _35059_);
  nor (_35062_, _35061_, _11680_);
  and (_35063_, _11645_, _04436_);
  and (_35064_, _04437_, \oc8051_golden_model_1.PC [8]);
  and (_35065_, _35064_, _11688_);
  nor (_35066_, _35065_, _35063_);
  nor (_35067_, _35066_, _08108_);
  nor (_35068_, _35067_, _33255_);
  nor (_35070_, _35068_, _35062_);
  not (_35071_, _35061_);
  nor (_35072_, _35071_, _11683_);
  nor (_35073_, _35072_, _03536_);
  not (_35074_, _35073_);
  nor (_35075_, _35074_, _35070_);
  not (_35076_, _11645_);
  and (_35077_, _35076_, _03536_);
  nor (_35078_, _35077_, _08118_);
  not (_35079_, _35078_);
  nor (_35081_, _35079_, _35075_);
  not (_35082_, _23346_);
  and (_35083_, _35061_, _08118_);
  nor (_35084_, _35083_, _35082_);
  not (_35085_, _35084_);
  nor (_35086_, _35085_, _35081_);
  nor (_35087_, _35086_, _04012_);
  and (_35088_, _35087_, _35057_);
  and (_35089_, _35061_, _04012_);
  or (_35090_, _35089_, _03534_);
  or (_35092_, _35090_, _35088_);
  nand (_35093_, _35092_, _35051_);
  nand (_35094_, _35093_, _11430_);
  nor (_35095_, _35061_, _11430_);
  nor (_35096_, _35095_, _03469_);
  and (_35097_, _35096_, _35094_);
  or (_35098_, _35097_, _35044_);
  nand (_35099_, _35098_, _35043_);
  and (_35100_, _11645_, _03527_);
  nor (_35101_, _35100_, _11716_);
  nand (_35103_, _35101_, _35099_);
  nor (_35104_, _35061_, _11715_);
  nor (_35105_, _35104_, _03530_);
  nand (_35106_, _35105_, _35103_);
  and (_35107_, _11645_, _03530_);
  nor (_35108_, _35107_, _11724_);
  nand (_35109_, _35108_, _35106_);
  nor (_35110_, _35061_, _11723_);
  nor (_35111_, _35110_, _03465_);
  and (_35112_, _35111_, _35109_);
  or (_35114_, _35112_, _35042_);
  nand (_35115_, _35114_, _11728_);
  and (_35116_, _11645_, _03464_);
  nor (_35117_, _35116_, _10021_);
  nand (_35118_, _35117_, _35115_);
  not (_35119_, _34408_);
  and (_35120_, _11532_, _10055_);
  nor (_35121_, _35046_, _10055_);
  nor (_35122_, _35121_, _35120_);
  nor (_35123_, _35122_, _10017_);
  nor (_35125_, _35123_, _35119_);
  and (_35126_, _35125_, _35118_);
  not (_35127_, _35046_);
  or (_35128_, _35127_, _10116_);
  or (_35129_, _11532_, _11743_);
  nand (_35130_, _35129_, _35128_);
  and (_35131_, _35130_, _35119_);
  or (_35132_, _35131_, _03547_);
  or (_35133_, _35132_, _35126_);
  and (_35134_, _11531_, _09975_);
  nor (_35136_, _35127_, _09975_);
  or (_35137_, _35136_, _03994_);
  or (_35138_, _35137_, _35134_);
  and (_35139_, _35138_, _10123_);
  nand (_35140_, _35139_, _35133_);
  and (_35141_, _35061_, _10122_);
  and (_35142_, _11531_, _10163_);
  and (_35143_, _35046_, _11764_);
  or (_35144_, _35143_, _35142_);
  and (_35145_, _35144_, _03608_);
  nor (_35147_, _35145_, _35141_);
  nand (_35148_, _35147_, _35140_);
  nand (_35149_, _35148_, _03459_);
  and (_35150_, _11645_, _03458_);
  nor (_35151_, _35150_, _04755_);
  nand (_35152_, _35151_, _35149_);
  nand (_35153_, _35152_, _32576_);
  nor (_35154_, _32576_, _35076_);
  nor (_35155_, _35154_, _11425_);
  nand (_35156_, _35155_, _35153_);
  nor (_35158_, _35061_, _11424_);
  nor (_35159_, _35158_, _03587_);
  nand (_35160_, _35159_, _35156_);
  and (_35161_, _11645_, _03587_);
  nor (_35162_, _35161_, _11776_);
  nand (_35163_, _35162_, _35160_);
  nand (_35164_, _35163_, _10265_);
  and (_35165_, _11645_, _03586_);
  nor (_35166_, _35165_, _11780_);
  nand (_35167_, _35166_, _35164_);
  nor (_35169_, _35061_, _11419_);
  nor (_35170_, _35169_, _08267_);
  nand (_35171_, _35170_, _35167_);
  nor (_35172_, _35076_, _08266_);
  nor (_35173_, _35172_, _03334_);
  and (_35174_, _35173_, _35171_);
  nor (_35175_, _35061_, _03233_);
  or (_35176_, _35175_, _35174_);
  nand (_35177_, _35176_, _03453_);
  and (_35178_, _35076_, _03452_);
  nor (_35180_, _35178_, _23659_);
  nand (_35181_, _35180_, _35177_);
  and (_35182_, _11531_, _03621_);
  not (_35183_, _35182_);
  and (_35184_, _35183_, _11797_);
  nand (_35185_, _35184_, _35181_);
  nor (_35186_, _11645_, _11797_);
  nor (_35187_, _35186_, _03224_);
  nand (_35188_, _35187_, _35185_);
  and (_35189_, _11531_, _03224_);
  nor (_35191_, _35189_, _32624_);
  nand (_35192_, _35191_, _35188_);
  nor (_35193_, _35061_, _11806_);
  nor (_35194_, _35193_, _03517_);
  and (_35195_, _35194_, _35192_);
  or (_35196_, _35195_, _35041_);
  nand (_35197_, _35196_, _35040_);
  and (_35198_, _35054_, _11813_);
  nor (_35199_, _35198_, _06193_);
  and (_35200_, _35199_, _35197_);
  nor (_35202_, _11645_, _05916_);
  or (_35203_, _35202_, _35200_);
  nand (_35204_, _35203_, _04509_);
  and (_35205_, _11532_, _03624_);
  nor (_35206_, _35205_, _08461_);
  nand (_35207_, _35206_, _35204_);
  and (_35208_, _11645_, _08461_);
  nor (_35209_, _35208_, _11828_);
  nand (_35210_, _35209_, _35207_);
  nor (_35211_, _11852_, \oc8051_golden_model_1.DPH [0]);
  nor (_35213_, _35211_, _11853_);
  nor (_35214_, _35213_, _23814_);
  nor (_35215_, _35214_, _03516_);
  nand (_35216_, _35215_, _35210_);
  and (_35217_, _11645_, _03516_);
  nor (_35218_, _35217_, _03168_);
  nand (_35219_, _35218_, _35216_);
  nand (_35220_, _35219_, _23819_);
  and (_35221_, _11645_, _08864_);
  and (_35222_, _35054_, _11894_);
  or (_35224_, _35222_, _35221_);
  and (_35225_, _35224_, _11868_);
  nor (_35226_, _35225_, _11872_);
  nand (_35227_, _35226_, _35220_);
  nor (_35228_, _35061_, _11416_);
  nor (_35229_, _35228_, _08494_);
  nand (_35230_, _35229_, _35227_);
  nor (_35231_, _35076_, _08493_);
  nor (_35232_, _35231_, _03623_);
  nand (_35233_, _35232_, _35230_);
  and (_35235_, _11532_, _03623_);
  nor (_35236_, _35235_, _03744_);
  nand (_35237_, _35236_, _35233_);
  and (_35238_, _11645_, _03744_);
  nor (_35239_, _35238_, _03172_);
  nand (_35240_, _35239_, _35237_);
  nand (_35241_, _35240_, _11893_);
  nor (_35242_, _35054_, _11894_);
  nor (_35243_, _11645_, _08864_);
  nor (_35244_, _35243_, _11893_);
  not (_35246_, _35244_);
  nor (_35247_, _35246_, _35242_);
  nor (_35248_, _35247_, _11901_);
  nand (_35249_, _35248_, _35241_);
  and (_35250_, _35071_, _11901_);
  nor (_35251_, _35250_, _11905_);
  nand (_35252_, _35251_, _35249_);
  nor (_35253_, _35076_, _11904_);
  nor (_35254_, _35253_, _03611_);
  and (_35255_, _35254_, _35252_);
  and (_35257_, _11532_, _03611_);
  or (_35258_, _35257_, _35255_);
  nand (_35259_, _35258_, _03734_);
  nor (_35260_, _11915_, _03182_);
  and (_35261_, _35076_, _03733_);
  not (_35262_, _35261_);
  and (_35263_, _35262_, _35260_);
  nand (_35264_, _35263_, _35259_);
  and (_35265_, _11645_, \oc8051_golden_model_1.PSW [7]);
  and (_35266_, _35054_, _07982_);
  or (_35268_, _35266_, _35265_);
  and (_35269_, _35268_, _11915_);
  nor (_35270_, _35269_, _11919_);
  nand (_35271_, _35270_, _35264_);
  nor (_35272_, _35061_, _11413_);
  nor (_35273_, _35272_, _15156_);
  and (_35274_, _35273_, _35271_);
  nor (_35275_, _35076_, _11410_);
  or (_35276_, _35275_, _03618_);
  or (_35277_, _35276_, _35274_);
  and (_35279_, _11532_, _03618_);
  nor (_35280_, _35279_, _03741_);
  and (_35281_, _35280_, _35277_);
  and (_35282_, _11645_, _03741_);
  or (_35283_, _35282_, _35281_);
  nand (_35284_, _35283_, _35039_);
  or (_35285_, _35054_, _07982_);
  or (_35286_, _11645_, \oc8051_golden_model_1.PSW [7]);
  and (_35287_, _35286_, _11936_);
  and (_35288_, _35287_, _35285_);
  nor (_35290_, _35288_, _11940_);
  nand (_35291_, _35290_, _35284_);
  nor (_35292_, _35061_, _11408_);
  nor (_35293_, _35292_, _08629_);
  nand (_35294_, _35293_, _35291_);
  nor (_35295_, _35076_, _08628_);
  nor (_35296_, _35295_, _08707_);
  nand (_35297_, _35296_, _35294_);
  and (_35298_, _35071_, _08707_);
  nor (_35299_, _35298_, _03752_);
  nand (_35301_, _35299_, _35297_);
  and (_35302_, _04429_, _03752_);
  nor (_35303_, _35302_, _03191_);
  nand (_35304_, _35303_, _35301_);
  nand (_35305_, _35304_, _03814_);
  nor (_35306_, _11531_, _09953_);
  and (_35307_, _35127_, _09953_);
  or (_35308_, _35307_, _03814_);
  or (_35309_, _35308_, _35306_);
  and (_35310_, _35309_, _11406_);
  nand (_35312_, _35310_, _35305_);
  nor (_35313_, _35061_, _11406_);
  nor (_35314_, _35313_, _08785_);
  and (_35315_, _35314_, _35312_);
  nor (_35316_, _35076_, _08784_);
  or (_35317_, _35316_, _08815_);
  or (_35318_, _35317_, _35315_);
  and (_35319_, _35071_, _08815_);
  nor (_35320_, _35319_, _03475_);
  nand (_35321_, _35320_, _35318_);
  and (_35323_, _04429_, _03475_);
  nor (_35324_, _35323_, _03189_);
  nand (_35325_, _35324_, _35321_);
  nand (_35326_, _35325_, _03768_);
  and (_35327_, _11532_, _09953_);
  nor (_35328_, _35046_, _09953_);
  nor (_35329_, _35328_, _35327_);
  and (_35330_, _35329_, _03644_);
  nor (_35331_, _35330_, _11992_);
  nand (_35332_, _35331_, _35326_);
  nor (_35334_, _35061_, _11991_);
  nor (_35335_, _35334_, _03767_);
  nand (_35336_, _35335_, _35332_);
  and (_35337_, _11645_, _03767_);
  nor (_35338_, _35337_, _11999_);
  nand (_35339_, _35338_, _35336_);
  nor (_35340_, _35061_, _11998_);
  nor (_35341_, _35340_, _03645_);
  and (_35342_, _35341_, _35339_);
  or (_35343_, _35342_, _35038_);
  nor (_35345_, _03445_, _03196_);
  nand (_35346_, _35345_, _35343_);
  and (_35347_, _35329_, _03445_);
  nor (_35348_, _35347_, _12016_);
  nand (_35349_, _35348_, _35346_);
  nor (_35350_, _35061_, _12015_);
  nor (_35351_, _35350_, _03473_);
  nand (_35352_, _35351_, _35349_);
  and (_35353_, _11645_, _03473_);
  nor (_35354_, _35353_, _12022_);
  nand (_35356_, _35354_, _35352_);
  nor (_35357_, _35061_, _11392_);
  nor (_35358_, _35357_, _03615_);
  and (_35359_, _35358_, _35356_);
  or (_35360_, _35359_, _35037_);
  nand (_35361_, _35360_, _35035_);
  and (_35362_, _35061_, _12031_);
  not (_35363_, _35362_);
  and (_35364_, _35363_, _35361_);
  nand (_35365_, _35364_, _43189_);
  or (_35367_, _43189_, \oc8051_golden_model_1.PC [8]);
  and (_35368_, _35367_, _42003_);
  and (_43928_, _35368_, _35365_);
  nor (_35369_, _04292_, _11391_);
  nor (_35370_, _04292_, _06855_);
  and (_35371_, _35059_, \oc8051_golden_model_1.PC [9]);
  nor (_35372_, _35059_, \oc8051_golden_model_1.PC [9]);
  nor (_35373_, _35372_, _35371_);
  nor (_35374_, _35373_, _11406_);
  and (_35375_, _11472_, _03618_);
  nor (_35377_, _35373_, _11413_);
  and (_35378_, _11472_, _03611_);
  not (_35379_, _35373_);
  and (_35380_, _35379_, _11901_);
  and (_35381_, _11472_, _03623_);
  nor (_35382_, _35373_, _11416_);
  nor (_35383_, _11592_, _05916_);
  and (_35384_, _11592_, _03517_);
  nor (_35385_, _35373_, _11424_);
  nor (_35386_, _35373_, _11687_);
  nand (_35388_, _11592_, _04436_);
  and (_35389_, _04437_, \oc8051_golden_model_1.PC [9]);
  nand (_35390_, _35389_, _11683_);
  and (_35391_, _35390_, _32884_);
  or (_35392_, _35391_, _03536_);
  and (_35393_, _35392_, _35388_);
  or (_35394_, _35393_, _35386_);
  and (_35395_, _11683_, _11686_);
  or (_35396_, _35395_, _35379_);
  and (_35397_, _11592_, _03536_);
  nor (_35399_, _35397_, _35082_);
  and (_35400_, _35399_, _35396_);
  and (_35401_, _35400_, _35394_);
  and (_35402_, _11566_, _11592_);
  nor (_35403_, _11649_, _11646_);
  and (_35404_, _35403_, _11595_);
  nor (_35405_, _35403_, _11595_);
  nor (_35406_, _35405_, _35404_);
  nor (_35407_, _35406_, _11566_);
  nor (_35408_, _35407_, _35402_);
  and (_35410_, _35408_, _05998_);
  or (_35411_, _35410_, _35401_);
  nand (_35412_, _35411_, _06008_);
  and (_35413_, _35379_, _04012_);
  nor (_35414_, _35413_, _03534_);
  and (_35415_, _35414_, _35412_);
  or (_35416_, _32250_, _11472_);
  nor (_35417_, _11536_, _11533_);
  and (_35418_, _35417_, _11476_);
  nor (_35419_, _35417_, _11476_);
  nor (_35421_, _35419_, _35418_);
  and (_35422_, _35421_, _11439_);
  nor (_35423_, _35422_, _04432_);
  and (_35424_, _35423_, _35416_);
  or (_35425_, _35424_, _11431_);
  or (_35426_, _35425_, _35415_);
  nor (_35427_, _35373_, _11430_);
  nor (_35428_, _35427_, _03469_);
  nand (_35429_, _35428_, _35426_);
  and (_35430_, _11592_, _03469_);
  nor (_35432_, _35430_, _05977_);
  nand (_35433_, _35432_, _35429_);
  nand (_35434_, _35433_, _04457_);
  and (_35435_, _11592_, _03527_);
  nor (_35436_, _35435_, _11716_);
  nand (_35437_, _35436_, _35434_);
  nor (_35438_, _35373_, _11715_);
  nor (_35439_, _35438_, _03530_);
  nand (_35440_, _35439_, _35437_);
  and (_35441_, _11592_, _03530_);
  nor (_35443_, _35441_, _11724_);
  nand (_35444_, _35443_, _35440_);
  nor (_35445_, _35373_, _11723_);
  nor (_35446_, _35445_, _03465_);
  nand (_35447_, _35446_, _35444_);
  and (_35448_, _11592_, _03465_);
  nor (_35449_, _35448_, _11727_);
  nand (_35450_, _35449_, _35447_);
  nand (_35451_, _35450_, _04577_);
  and (_35452_, _11592_, _03464_);
  nor (_35454_, _35452_, _10021_);
  and (_35455_, _35454_, _35451_);
  and (_35456_, _11472_, _10055_);
  nor (_35457_, _35421_, _10055_);
  or (_35458_, _35457_, _35456_);
  nor (_35459_, _35458_, _10017_);
  or (_35460_, _35459_, _35455_);
  nand (_35461_, _35460_, _10112_);
  and (_35462_, _11472_, _10116_);
  not (_35463_, _35421_);
  and (_35465_, _35463_, _11743_);
  or (_35466_, _35465_, _34408_);
  or (_35467_, _35466_, _35462_);
  and (_35468_, _35467_, _03994_);
  and (_35469_, _35468_, _35461_);
  and (_35470_, _11472_, _09975_);
  nor (_35471_, _35421_, _09975_);
  nor (_35472_, _35471_, _35470_);
  nor (_35473_, _35472_, _03994_);
  or (_35474_, _35473_, _35469_);
  nand (_35476_, _35474_, _10123_);
  and (_35477_, _11472_, _10163_);
  nor (_35478_, _35421_, _10163_);
  or (_35479_, _35478_, _35477_);
  and (_35480_, _35479_, _03608_);
  and (_35481_, _35373_, _10122_);
  nor (_35482_, _35481_, _35480_);
  and (_35483_, _35482_, _03459_);
  nand (_35484_, _35483_, _35476_);
  not (_35485_, _11592_);
  and (_35487_, _35485_, _03458_);
  nor (_35488_, _35487_, _04755_);
  and (_35489_, _35488_, _32576_);
  nand (_35490_, _35489_, _35484_);
  nor (_35491_, _32576_, _35485_);
  nor (_35492_, _35491_, _11425_);
  and (_35493_, _35492_, _35490_);
  or (_35494_, _35493_, _35385_);
  or (_35495_, _35494_, _03587_);
  nand (_35496_, _11592_, _03587_);
  and (_35499_, _35496_, _35495_);
  or (_35500_, _35499_, _11776_);
  or (_35501_, _35500_, _03586_);
  and (_35502_, _11592_, _03586_);
  nor (_35503_, _35502_, _11780_);
  and (_35504_, _35503_, _35501_);
  nor (_35505_, _35373_, _11419_);
  or (_35506_, _35505_, _35504_);
  nand (_35507_, _35506_, _08266_);
  nor (_35508_, _11592_, _08266_);
  nor (_35510_, _35508_, _03334_);
  nand (_35511_, _35510_, _35507_);
  nor (_35512_, _35379_, _03233_);
  nor (_35513_, _35512_, _03452_);
  nand (_35514_, _35513_, _35511_);
  and (_35515_, _35485_, _03452_);
  nor (_35516_, _35515_, _23659_);
  nand (_35517_, _35516_, _35514_);
  and (_35518_, _11472_, _03621_);
  not (_35519_, _35518_);
  and (_35522_, _35519_, _11797_);
  nand (_35523_, _35522_, _35517_);
  nor (_35524_, _11592_, _11797_);
  nor (_35525_, _35524_, _03224_);
  nand (_35526_, _35525_, _35523_);
  and (_35527_, _11472_, _03224_);
  nor (_35528_, _35527_, _32624_);
  nand (_35529_, _35528_, _35526_);
  nor (_35530_, _35373_, _11806_);
  nor (_35531_, _35530_, _03517_);
  and (_35533_, _35531_, _35529_);
  or (_35534_, _35533_, _35384_);
  nand (_35535_, _35534_, _35040_);
  nor (_35536_, _35406_, _11814_);
  nor (_35537_, _35536_, _06193_);
  and (_35538_, _35537_, _35535_);
  or (_35539_, _35538_, _35383_);
  nand (_35540_, _35539_, _04509_);
  and (_35541_, _11473_, _03624_);
  nor (_35542_, _35541_, _08461_);
  nand (_35545_, _35542_, _35540_);
  and (_35546_, _11592_, _08461_);
  nor (_35547_, _35546_, _11828_);
  nand (_35548_, _35547_, _35545_);
  nor (_35549_, _11853_, \oc8051_golden_model_1.DPH [1]);
  nor (_35550_, _35549_, _11854_);
  nor (_35551_, _35550_, _23814_);
  nor (_35552_, _35551_, _03516_);
  nand (_35553_, _35552_, _35548_);
  and (_35554_, _11592_, _03516_);
  nor (_35556_, _35554_, _03168_);
  nand (_35557_, _35556_, _35553_);
  nand (_35558_, _35557_, _23819_);
  and (_35559_, _11592_, _08864_);
  nor (_35560_, _35406_, _08864_);
  or (_35561_, _35560_, _35559_);
  and (_35562_, _35561_, _11868_);
  nor (_35563_, _35562_, _11872_);
  and (_35564_, _35563_, _35558_);
  or (_35565_, _35564_, _35382_);
  nand (_35568_, _35565_, _08493_);
  nor (_35569_, _11592_, _08493_);
  nor (_35570_, _35569_, _03623_);
  and (_35571_, _35570_, _35568_);
  or (_35572_, _35571_, _35381_);
  nand (_35573_, _35572_, _03745_);
  and (_35574_, _11592_, _03744_);
  nor (_35575_, _35574_, _03172_);
  nand (_35576_, _35575_, _35573_);
  nand (_35577_, _35576_, _11893_);
  and (_35579_, _35406_, _08864_);
  nor (_35580_, _11592_, _08864_);
  nor (_35581_, _35580_, _11893_);
  not (_35582_, _35581_);
  nor (_35583_, _35582_, _35579_);
  nor (_35584_, _35583_, _11901_);
  and (_35585_, _35584_, _35577_);
  or (_35586_, _35585_, _35380_);
  nand (_35587_, _35586_, _11904_);
  nor (_35588_, _11592_, _11904_);
  nor (_35590_, _35588_, _03611_);
  and (_35591_, _35590_, _35587_);
  or (_35592_, _35591_, _35378_);
  nand (_35593_, _35592_, _03734_);
  and (_35594_, _11592_, _03733_);
  nor (_35595_, _35594_, _03182_);
  nand (_35596_, _35595_, _35593_);
  nand (_35597_, _35596_, _24078_);
  and (_35598_, _11592_, \oc8051_golden_model_1.PSW [7]);
  nor (_35599_, _35406_, \oc8051_golden_model_1.PSW [7]);
  or (_35601_, _35599_, _35598_);
  and (_35602_, _35601_, _11915_);
  nor (_35603_, _35602_, _11919_);
  and (_35604_, _35603_, _35597_);
  or (_35605_, _35604_, _35377_);
  nand (_35606_, _35605_, _11410_);
  nor (_35607_, _11592_, _11410_);
  nor (_35608_, _35607_, _03618_);
  and (_35609_, _35608_, _35606_);
  or (_35610_, _35609_, _35375_);
  nand (_35612_, _35610_, _06458_);
  and (_35613_, _11592_, _03741_);
  nor (_35614_, _35613_, _03178_);
  nand (_35615_, _35614_, _35612_);
  nand (_35616_, _35615_, _11942_);
  nand (_35617_, _11592_, _07982_);
  or (_35618_, _35406_, _07982_);
  and (_35619_, _35618_, _35617_);
  or (_35620_, _35619_, _11942_);
  nand (_35621_, _35620_, _35616_);
  nand (_35623_, _35621_, _11408_);
  nor (_35624_, _35379_, _11408_);
  nor (_35625_, _35624_, _08629_);
  nand (_35626_, _35625_, _35623_);
  nor (_35627_, _11592_, _08628_);
  nor (_35628_, _35627_, _08707_);
  nand (_35629_, _35628_, _35626_);
  and (_35630_, _35373_, _08707_);
  nor (_35631_, _35630_, _03752_);
  nand (_35632_, _35631_, _35629_);
  nor (_35634_, _03617_, _03191_);
  not (_35635_, _35634_);
  and (_35636_, _04635_, _03752_);
  nor (_35637_, _35636_, _35635_);
  nand (_35638_, _35637_, _35632_);
  and (_35639_, _35421_, _09953_);
  nor (_35640_, _11472_, _09953_);
  or (_35641_, _35640_, _03814_);
  nor (_35642_, _35641_, _35639_);
  nor (_35643_, _35642_, _11963_);
  and (_35645_, _35643_, _35638_);
  or (_35646_, _35645_, _35374_);
  nand (_35647_, _35646_, _08784_);
  nor (_35648_, _11592_, _08784_);
  nor (_35649_, _35648_, _08815_);
  nand (_35650_, _35649_, _35647_);
  and (_35651_, _35373_, _08815_);
  nor (_35652_, _35651_, _03475_);
  nand (_35653_, _35652_, _35650_);
  nor (_35654_, _03644_, _03189_);
  not (_35656_, _35654_);
  and (_35657_, _04635_, _03475_);
  nor (_35658_, _35657_, _35656_);
  nand (_35659_, _35658_, _35653_);
  and (_35660_, _11473_, _09953_);
  nor (_35661_, _35463_, _09953_);
  nor (_35662_, _35661_, _35660_);
  and (_35663_, _35662_, _03644_);
  nor (_35664_, _35663_, _11992_);
  nand (_35665_, _35664_, _35659_);
  nor (_35667_, _35373_, _11991_);
  nor (_35668_, _35667_, _03767_);
  nand (_35669_, _35668_, _35665_);
  and (_35670_, _11592_, _03767_);
  nor (_35671_, _35670_, _11999_);
  nand (_35672_, _35671_, _35669_);
  nor (_35673_, _35373_, _11998_);
  nor (_35674_, _35673_, _03645_);
  and (_35675_, _35674_, _35672_);
  or (_35676_, _35675_, _35370_);
  nand (_35678_, _35676_, _35345_);
  and (_35679_, _35662_, _03445_);
  nor (_35680_, _35679_, _12016_);
  nand (_35681_, _35680_, _35678_);
  nor (_35682_, _35373_, _12015_);
  nor (_35683_, _35682_, _03473_);
  nand (_35684_, _35683_, _35681_);
  and (_35685_, _11592_, _03473_);
  nor (_35686_, _35685_, _12022_);
  nand (_35687_, _35686_, _35684_);
  nor (_35689_, _35373_, _11392_);
  nor (_35690_, _35689_, _03615_);
  and (_35691_, _35690_, _35687_);
  or (_35692_, _35691_, _35369_);
  nand (_35693_, _35692_, _35035_);
  and (_35694_, _35373_, _12031_);
  not (_35695_, _35694_);
  and (_35696_, _35695_, _35693_);
  nand (_35697_, _35696_, _43189_);
  or (_35698_, _43189_, \oc8051_golden_model_1.PC [9]);
  and (_35700_, _35698_, _42003_);
  and (_43929_, _35700_, _35697_);
  nor (_35701_, _35371_, \oc8051_golden_model_1.PC [10]);
  nor (_35702_, _35701_, _11396_);
  and (_35703_, _35702_, _12031_);
  not (_35704_, _35703_);
  and (_35705_, _03944_, _03615_);
  and (_35706_, _03944_, _03645_);
  nor (_35707_, _35702_, _11406_);
  nor (_35708_, _35702_, _11408_);
  nand (_35710_, _11457_, _03618_);
  nand (_35711_, _11457_, _03611_);
  nand (_35712_, _11457_, _03623_);
  not (_35713_, _11586_);
  nor (_35714_, _35713_, _05916_);
  or (_35715_, _35714_, _03624_);
  not (_35716_, _35702_);
  nor (_35717_, _35716_, _11806_);
  nor (_35718_, _35716_, _11723_);
  or (_35719_, _35702_, _11715_);
  and (_35721_, _35702_, _11710_);
  not (_35722_, _11469_);
  nor (_35723_, _11540_, _11537_);
  nor (_35724_, _35723_, _35722_);
  and (_35725_, _35723_, _35722_);
  nor (_35726_, _35725_, _35724_);
  or (_35727_, _35726_, _11437_);
  or (_35728_, _11456_, _11439_);
  and (_35729_, _35728_, _03534_);
  and (_35730_, _35729_, _35727_);
  nor (_35732_, _11653_, _11650_);
  not (_35733_, _35732_);
  and (_35734_, _35733_, _11589_);
  nor (_35735_, _35733_, _11589_);
  nor (_35736_, _35735_, _35734_);
  or (_35737_, _35736_, _11566_);
  or (_35738_, _32232_, _11586_);
  and (_35739_, _35738_, _35737_);
  or (_35740_, _35739_, _05997_);
  or (_35741_, _35702_, _11684_);
  nand (_35743_, _35713_, _04436_);
  or (_35744_, _04436_, \oc8051_golden_model_1.PC [10]);
  or (_35745_, _35744_, _11682_);
  and (_35746_, _35745_, _35743_);
  or (_35747_, _33255_, _08108_);
  or (_35748_, _35747_, _35746_);
  and (_35749_, _35748_, _35741_);
  or (_35750_, _35749_, _03536_);
  nand (_35751_, _35713_, _03536_);
  and (_35752_, _35751_, _11686_);
  and (_35754_, _35752_, _35750_);
  nand (_35755_, _35702_, _08118_);
  nand (_35756_, _35755_, _23346_);
  or (_35757_, _35756_, _35754_);
  and (_35758_, _35757_, _11705_);
  and (_35759_, _35758_, _35740_);
  or (_35760_, _35759_, _35730_);
  and (_35761_, _35760_, _11430_);
  or (_35762_, _35761_, _35721_);
  and (_35763_, _35762_, _03532_);
  nor (_35765_, _35713_, _03532_);
  nor (_35766_, _35765_, _05977_);
  nand (_35767_, _35766_, _11715_);
  or (_35768_, _35767_, _35763_);
  and (_35769_, _35768_, _35719_);
  or (_35770_, _35769_, _03530_);
  nand (_35771_, _35713_, _03530_);
  and (_35772_, _35771_, _11723_);
  and (_35773_, _35772_, _35770_);
  or (_35774_, _35773_, _35718_);
  and (_35776_, _35774_, _03466_);
  and (_35777_, _11586_, _03465_);
  or (_35778_, _35777_, _11727_);
  or (_35779_, _35778_, _35776_);
  and (_35780_, _35779_, _04577_);
  nand (_35781_, _11586_, _03464_);
  nand (_35782_, _35781_, _10017_);
  or (_35783_, _35782_, _35780_);
  not (_35784_, _35726_);
  nor (_35785_, _35784_, _10055_);
  and (_35787_, _11456_, _10055_);
  or (_35788_, _35787_, _10017_);
  or (_35789_, _35788_, _35785_);
  and (_35790_, _35789_, _33678_);
  and (_35791_, _35790_, _35783_);
  nor (_35792_, _35784_, _09975_);
  and (_35793_, _11456_, _09975_);
  or (_35794_, _35793_, _35792_);
  and (_35795_, _35794_, _03547_);
  and (_35796_, _35726_, _11743_);
  and (_35798_, _11456_, _10116_);
  or (_35799_, _35798_, _35796_);
  and (_35800_, _35799_, _10020_);
  or (_35801_, _35800_, _35795_);
  or (_35802_, _35801_, _35791_);
  and (_35803_, _35802_, _10123_);
  and (_35804_, _35702_, _10122_);
  or (_35805_, _35726_, _10163_);
  nand (_35806_, _11457_, _10163_);
  and (_35807_, _35806_, _03608_);
  and (_35809_, _35807_, _35805_);
  or (_35810_, _35809_, _35804_);
  or (_35811_, _35810_, _35803_);
  and (_35812_, _32576_, _03459_);
  and (_35813_, _35812_, _35811_);
  nor (_35814_, _35812_, _35713_);
  nand (_35815_, _11424_, _03207_);
  or (_35816_, _35815_, _35814_);
  or (_35817_, _35816_, _35813_);
  or (_35818_, _35702_, _11424_);
  and (_35820_, _35818_, _09769_);
  and (_35821_, _35820_, _35817_);
  or (_35822_, _35821_, _11776_);
  and (_35823_, _35822_, _10265_);
  or (_35824_, _35713_, _03588_);
  nand (_35825_, _35824_, _11419_);
  or (_35826_, _35825_, _35823_);
  or (_35827_, _35702_, _11419_);
  and (_35828_, _35827_, _08266_);
  and (_35829_, _35828_, _35826_);
  nor (_35831_, _35713_, _08266_);
  or (_35832_, _35831_, _03334_);
  or (_35833_, _35832_, _35829_);
  or (_35834_, _35702_, _03233_);
  and (_35835_, _35834_, _03453_);
  and (_35836_, _35835_, _35833_);
  nand (_35837_, _11586_, _03452_);
  nand (_35838_, _35837_, _23658_);
  or (_35839_, _35838_, _35836_);
  nand (_35840_, _11457_, _03621_);
  and (_35842_, _35840_, _11797_);
  and (_35843_, _35842_, _35839_);
  nor (_35844_, _35713_, _11797_);
  or (_35845_, _35844_, _03224_);
  or (_35846_, _35845_, _35843_);
  nand (_35847_, _11457_, _03224_);
  and (_35848_, _35847_, _11806_);
  and (_35849_, _35848_, _35846_);
  or (_35850_, _35849_, _35717_);
  and (_35851_, _35850_, _10351_);
  nand (_35853_, _11586_, _03517_);
  nand (_35854_, _35853_, _35040_);
  or (_35855_, _35854_, _35851_);
  or (_35856_, _35736_, _11814_);
  and (_35857_, _35856_, _05916_);
  and (_35858_, _35857_, _35855_);
  or (_35859_, _35858_, _35715_);
  nand (_35860_, _11457_, _03624_);
  and (_35861_, _35860_, _35859_);
  or (_35862_, _35861_, _08461_);
  and (_35864_, _35713_, _08461_);
  nor (_35865_, _35864_, _11828_);
  and (_35866_, _35865_, _35862_);
  or (_35867_, _11854_, \oc8051_golden_model_1.DPH [2]);
  nor (_35868_, _11855_, _23814_);
  and (_35869_, _35868_, _35867_);
  or (_35870_, _35869_, _03516_);
  or (_35871_, _35870_, _35866_);
  nor (_35872_, _11868_, _03168_);
  nand (_35873_, _35713_, _03516_);
  and (_35875_, _35873_, _35872_);
  and (_35876_, _35875_, _35871_);
  or (_35877_, _35736_, _08864_);
  or (_35878_, _11586_, _11894_);
  and (_35879_, _35878_, _11868_);
  and (_35880_, _35879_, _35877_);
  or (_35881_, _35880_, _11872_);
  or (_35882_, _35881_, _35876_);
  or (_35883_, _35702_, _11416_);
  and (_35884_, _35883_, _08493_);
  and (_35886_, _35884_, _35882_);
  nor (_35887_, _35713_, _08493_);
  or (_35888_, _35887_, _03623_);
  or (_35889_, _35888_, _35886_);
  and (_35890_, _35889_, _35712_);
  or (_35891_, _35890_, _03744_);
  nand (_35892_, _35713_, _03744_);
  and (_35893_, _35892_, _23958_);
  and (_35894_, _35893_, _35891_);
  or (_35895_, _35736_, _11894_);
  or (_35897_, _11586_, _08864_);
  and (_35898_, _35897_, _11889_);
  and (_35899_, _35898_, _35895_);
  or (_35900_, _35899_, _11901_);
  or (_35901_, _35900_, _35894_);
  nand (_35902_, _35716_, _11901_);
  and (_35903_, _35902_, _11904_);
  and (_35904_, _35903_, _35901_);
  nor (_35905_, _35713_, _11904_);
  or (_35906_, _35905_, _03611_);
  or (_35908_, _35906_, _35904_);
  and (_35909_, _35908_, _35711_);
  or (_35910_, _35909_, _03733_);
  nand (_35911_, _35713_, _03733_);
  and (_35912_, _35911_, _35260_);
  and (_35913_, _35912_, _35910_);
  or (_35914_, _35736_, \oc8051_golden_model_1.PSW [7]);
  or (_35915_, _11586_, _07982_);
  and (_35916_, _35915_, _11915_);
  and (_35917_, _35916_, _35914_);
  or (_35919_, _35917_, _11919_);
  or (_35920_, _35919_, _35913_);
  or (_35921_, _35702_, _11413_);
  and (_35922_, _35921_, _11410_);
  and (_35923_, _35922_, _35920_);
  nor (_35924_, _35713_, _11410_);
  or (_35925_, _35924_, _03618_);
  or (_35926_, _35925_, _35923_);
  and (_35927_, _35926_, _35710_);
  or (_35928_, _35927_, _03741_);
  nand (_35930_, _35713_, _03741_);
  and (_35931_, _35930_, _35039_);
  and (_35932_, _35931_, _35928_);
  or (_35933_, _35736_, _07982_);
  or (_35934_, _11586_, \oc8051_golden_model_1.PSW [7]);
  and (_35935_, _35934_, _11936_);
  and (_35936_, _35935_, _35933_);
  or (_35937_, _35936_, _11940_);
  nor (_35938_, _35937_, _35932_);
  or (_35939_, _35938_, _08629_);
  nor (_35941_, _35939_, _35708_);
  nor (_35942_, _35713_, _08628_);
  nor (_35943_, _35942_, _08707_);
  not (_35944_, _35943_);
  nor (_35945_, _35944_, _35941_);
  and (_35946_, _35716_, _08707_);
  nor (_35947_, _35946_, _35945_);
  nor (_35948_, _35947_, _03752_);
  and (_35949_, _05073_, _03752_);
  nor (_35950_, _35949_, _35635_);
  not (_35952_, _35950_);
  nor (_35953_, _35952_, _35948_);
  nor (_35954_, _11456_, _09953_);
  and (_35955_, _35784_, _09953_);
  or (_35956_, _35955_, _03814_);
  nor (_35957_, _35956_, _35954_);
  or (_35958_, _35957_, _11963_);
  nor (_35959_, _35958_, _35953_);
  or (_35960_, _35959_, _08785_);
  nor (_35961_, _35960_, _35707_);
  nor (_35963_, _35713_, _08784_);
  nor (_35964_, _35963_, _08815_);
  not (_35965_, _35964_);
  nor (_35966_, _35965_, _35961_);
  and (_35967_, _35716_, _08815_);
  nor (_35968_, _35967_, _35966_);
  nor (_35969_, _35968_, _03475_);
  and (_35970_, _05073_, _03475_);
  nor (_35971_, _35970_, _35656_);
  not (_35972_, _35971_);
  nor (_35974_, _35972_, _35969_);
  nor (_35975_, _35726_, _09953_);
  and (_35976_, _11457_, _09953_);
  nor (_35977_, _35976_, _35975_);
  and (_35978_, _35977_, _03644_);
  nor (_35979_, _35978_, _11992_);
  not (_35980_, _35979_);
  nor (_35981_, _35980_, _35974_);
  nor (_35982_, _35702_, _11991_);
  or (_35983_, _35982_, _35981_);
  nand (_35985_, _35983_, _03948_);
  and (_35986_, _35713_, _03767_);
  nor (_35987_, _35986_, _11999_);
  nand (_35988_, _35987_, _35985_);
  nor (_35989_, _35716_, _11998_);
  nor (_35990_, _35989_, _03645_);
  nand (_35991_, _35990_, _35988_);
  nand (_35992_, _35991_, _35345_);
  or (_35993_, _35992_, _35706_);
  and (_35994_, _35977_, _03445_);
  nor (_35996_, _35994_, _12016_);
  and (_35997_, _35996_, _35993_);
  nor (_35998_, _35702_, _12015_);
  or (_35999_, _35998_, _35997_);
  nand (_36000_, _35999_, _03474_);
  and (_36001_, _35713_, _03473_);
  nor (_36002_, _36001_, _12022_);
  nand (_36003_, _36002_, _36000_);
  nor (_36004_, _35716_, _11392_);
  nor (_36005_, _36004_, _03615_);
  nand (_36007_, _36005_, _36003_);
  nand (_36008_, _36007_, _35035_);
  or (_36009_, _36008_, _35705_);
  and (_36010_, _36009_, _35704_);
  nand (_36011_, _36010_, _43189_);
  or (_36012_, _43189_, \oc8051_golden_model_1.PC [10]);
  and (_36013_, _36012_, _42003_);
  and (_43932_, _36013_, _36011_);
  nor (_36014_, _11396_, _11460_);
  and (_36015_, _11396_, _11460_);
  or (_36017_, _36015_, _36014_);
  or (_36018_, _36017_, _11406_);
  or (_36019_, _36017_, _11408_);
  or (_36020_, _36017_, _11413_);
  or (_36021_, _36017_, _11416_);
  or (_36022_, _11808_, _11581_);
  and (_36023_, _36022_, _11814_);
  and (_36024_, _11463_, _03224_);
  or (_36025_, _36017_, _11419_);
  and (_36026_, _36017_, _11425_);
  nor (_36028_, _35724_, _11458_);
  and (_36029_, _36028_, _11467_);
  nor (_36030_, _36028_, _11467_);
  or (_36031_, _36030_, _36029_);
  and (_36032_, _36031_, _11743_);
  and (_36033_, _11463_, _10116_);
  or (_36034_, _36033_, _36032_);
  and (_36035_, _36034_, _10020_);
  and (_36036_, _11581_, _03530_);
  or (_36037_, _11581_, _11428_);
  or (_36039_, _11463_, _11439_);
  or (_36040_, _36031_, _11437_);
  and (_36041_, _36040_, _03534_);
  and (_36042_, _36041_, _36039_);
  nor (_36043_, _35734_, _11587_);
  and (_36044_, _36043_, _11584_);
  nor (_36045_, _36043_, _11584_);
  or (_36046_, _36045_, _36044_);
  and (_36047_, _36046_, _32232_);
  and (_36048_, _11566_, _11581_);
  or (_36050_, _36048_, _36047_);
  or (_36051_, _36050_, _05997_);
  or (_36052_, _36017_, _11684_);
  or (_36053_, _11581_, _04437_);
  or (_36054_, _04436_, \oc8051_golden_model_1.PC [11]);
  or (_36055_, _36054_, _11682_);
  and (_36056_, _36055_, _36053_);
  or (_36057_, _36056_, _35747_);
  nor (_36058_, _11581_, _03204_);
  nor (_36059_, _36058_, _03536_);
  and (_36061_, _36059_, _36057_);
  and (_36062_, _36061_, _36052_);
  and (_36063_, _11581_, _03536_);
  or (_36064_, _36063_, _08118_);
  or (_36065_, _36064_, _36062_);
  or (_36066_, _36017_, _11686_);
  and (_36067_, _36066_, _03209_);
  and (_36068_, _36067_, _36065_);
  nand (_36069_, _11581_, _11677_);
  nand (_36070_, _36069_, _05997_);
  or (_36072_, _36070_, _36068_);
  and (_36073_, _36072_, _11705_);
  and (_36074_, _36073_, _36051_);
  or (_36075_, _36074_, _36042_);
  and (_36076_, _36075_, _11430_);
  not (_36077_, _11428_);
  and (_36078_, _36017_, _11710_);
  or (_36079_, _36078_, _36077_);
  or (_36080_, _36079_, _36076_);
  and (_36081_, _36080_, _36037_);
  or (_36083_, _36081_, _11716_);
  or (_36084_, _36017_, _11715_);
  and (_36085_, _36084_, _03531_);
  and (_36086_, _36085_, _36083_);
  or (_36087_, _36086_, _36036_);
  and (_36088_, _36087_, _11723_);
  and (_36089_, _36017_, _11724_);
  or (_36090_, _36089_, _11730_);
  or (_36091_, _36090_, _36088_);
  or (_36092_, _11729_, _11581_);
  and (_36094_, _36092_, _36091_);
  or (_36095_, _36094_, _10021_);
  or (_36096_, _36031_, _10055_);
  nand (_36097_, _11464_, _10055_);
  and (_36098_, _36097_, _36096_);
  or (_36099_, _36098_, _10017_);
  and (_36100_, _36099_, _10112_);
  and (_36101_, _36100_, _36095_);
  or (_36102_, _36101_, _03547_);
  or (_36103_, _36102_, _36035_);
  not (_36105_, _09975_);
  and (_36106_, _36031_, _36105_);
  and (_36107_, _11463_, _09975_);
  or (_36108_, _36107_, _03994_);
  or (_36109_, _36108_, _36106_);
  and (_36110_, _36109_, _10123_);
  and (_36111_, _36110_, _36103_);
  or (_36112_, _36031_, _10163_);
  nand (_36113_, _11464_, _10163_);
  and (_36114_, _36113_, _03608_);
  and (_36116_, _36114_, _36112_);
  nand (_36117_, _36017_, _10122_);
  nand (_36118_, _36117_, _11761_);
  or (_36119_, _36118_, _36116_);
  or (_36120_, _36119_, _36111_);
  or (_36121_, _11761_, _11581_);
  and (_36122_, _36121_, _11424_);
  and (_36123_, _36122_, _36120_);
  or (_36124_, _36123_, _36026_);
  and (_36125_, _36124_, _11778_);
  not (_36127_, _11778_);
  nand (_36128_, _36127_, _11581_);
  nand (_36129_, _36128_, _11419_);
  or (_36130_, _36129_, _36125_);
  and (_36131_, _36130_, _36025_);
  or (_36132_, _36131_, _08267_);
  or (_36133_, _11581_, _08266_);
  and (_36134_, _36133_, _03233_);
  and (_36135_, _36134_, _36132_);
  nand (_36136_, _36017_, _03334_);
  nand (_36138_, _36136_, _11790_);
  or (_36139_, _36138_, _36135_);
  or (_36140_, _11790_, _11581_);
  and (_36141_, _36140_, _03622_);
  and (_36142_, _36141_, _36139_);
  nand (_36143_, _11463_, _03621_);
  nand (_36144_, _36143_, _11797_);
  or (_36145_, _36144_, _36142_);
  or (_36146_, _11581_, _11797_);
  and (_36147_, _36146_, _03521_);
  and (_36149_, _36147_, _36145_);
  or (_36150_, _36149_, _36024_);
  and (_36151_, _36150_, _11806_);
  and (_36152_, _36017_, _32624_);
  or (_36153_, _36152_, _11809_);
  or (_36154_, _36153_, _36151_);
  and (_36155_, _36154_, _36023_);
  and (_36156_, _36046_, _11813_);
  or (_36157_, _36156_, _06193_);
  or (_36158_, _36157_, _36155_);
  or (_36160_, _11581_, _05916_);
  and (_36161_, _36160_, _04509_);
  and (_36162_, _36161_, _36158_);
  and (_36163_, _11463_, _03624_);
  or (_36164_, _36163_, _08461_);
  or (_36165_, _36164_, _36162_);
  or (_36166_, _11581_, _08462_);
  and (_36167_, _36166_, _23814_);
  and (_36168_, _36167_, _36165_);
  or (_36169_, _11855_, \oc8051_golden_model_1.DPH [3]);
  nor (_36171_, _11856_, _23814_);
  and (_36172_, _36171_, _36169_);
  or (_36173_, _36172_, _11865_);
  or (_36174_, _36173_, _36168_);
  or (_36175_, _11864_, _11581_);
  and (_36176_, _36175_, _23819_);
  and (_36177_, _36176_, _36174_);
  or (_36178_, _36046_, _08864_);
  or (_36179_, _11581_, _11894_);
  and (_36180_, _36179_, _11868_);
  and (_36182_, _36180_, _36178_);
  or (_36183_, _36182_, _11872_);
  or (_36184_, _36183_, _36177_);
  and (_36185_, _36184_, _36021_);
  or (_36186_, _36185_, _08494_);
  or (_36187_, _11581_, _08493_);
  and (_36188_, _36187_, _04527_);
  and (_36189_, _36188_, _36186_);
  nand (_36190_, _11463_, _03623_);
  nand (_36191_, _36190_, _11885_);
  or (_36193_, _36191_, _36189_);
  or (_36194_, _11885_, _11581_);
  and (_36195_, _36194_, _11893_);
  and (_36196_, _36195_, _36193_);
  or (_36197_, _36046_, _11894_);
  or (_36198_, _11581_, _08864_);
  and (_36199_, _36198_, _11889_);
  and (_36200_, _36199_, _36197_);
  or (_36201_, _36200_, _36196_);
  and (_36202_, _36201_, _11902_);
  and (_36204_, _36017_, _11901_);
  or (_36205_, _36204_, _11905_);
  or (_36206_, _36205_, _36202_);
  or (_36207_, _11581_, _11904_);
  and (_36208_, _36207_, _04523_);
  and (_36209_, _36208_, _36206_);
  nand (_36210_, _11463_, _03611_);
  nand (_36211_, _36210_, _10828_);
  or (_36212_, _36211_, _36209_);
  and (_36213_, _24078_, _11581_);
  or (_36215_, _36213_, _24079_);
  and (_36216_, _36215_, _36212_);
  or (_36217_, _36046_, \oc8051_golden_model_1.PSW [7]);
  or (_36218_, _11581_, _07982_);
  and (_36219_, _36218_, _11915_);
  and (_36220_, _36219_, _36217_);
  or (_36221_, _36220_, _11919_);
  or (_36222_, _36221_, _36216_);
  and (_36223_, _36222_, _36020_);
  or (_36224_, _36223_, _15156_);
  or (_36226_, _11581_, _11410_);
  and (_36227_, _36226_, _06453_);
  and (_36228_, _36227_, _36224_);
  nand (_36229_, _11463_, _03618_);
  nand (_36230_, _36229_, _11932_);
  or (_36231_, _36230_, _36228_);
  and (_36232_, _11942_, _11581_);
  or (_36233_, _36232_, _24227_);
  and (_36234_, _36233_, _36231_);
  or (_36235_, _36046_, _07982_);
  or (_36237_, _11581_, \oc8051_golden_model_1.PSW [7]);
  and (_36238_, _36237_, _11936_);
  and (_36239_, _36238_, _36235_);
  or (_36240_, _36239_, _11940_);
  or (_36241_, _36240_, _36234_);
  and (_36242_, _36241_, _36019_);
  or (_36243_, _36242_, _08629_);
  or (_36244_, _11581_, _08628_);
  and (_36245_, _36244_, _08708_);
  and (_36246_, _36245_, _36243_);
  and (_36248_, _36017_, _08707_);
  or (_36249_, _36248_, _03752_);
  or (_36250_, _36249_, _36246_);
  nand (_36251_, _04885_, _03752_);
  and (_36252_, _36251_, _36250_);
  or (_36253_, _36252_, _03191_);
  or (_36254_, _11581_, _04803_);
  and (_36255_, _36254_, _03814_);
  and (_36256_, _36255_, _36253_);
  not (_36257_, _09953_);
  or (_36259_, _36031_, _36257_);
  or (_36260_, _11463_, _09953_);
  and (_36261_, _36260_, _03617_);
  and (_36262_, _36261_, _36259_);
  or (_36263_, _36262_, _11963_);
  or (_36264_, _36263_, _36256_);
  and (_36265_, _36264_, _36018_);
  or (_36266_, _36265_, _08785_);
  or (_36267_, _11581_, _08784_);
  and (_36268_, _36267_, _08816_);
  and (_36270_, _36268_, _36266_);
  and (_36271_, _36017_, _08815_);
  or (_36272_, _36271_, _03475_);
  or (_36273_, _36272_, _36270_);
  nand (_36274_, _04885_, _03475_);
  and (_36275_, _36274_, _36273_);
  or (_36276_, _36275_, _03189_);
  or (_36277_, _11581_, _11405_);
  and (_36278_, _36277_, _03768_);
  and (_36279_, _36278_, _36276_);
  or (_36281_, _36031_, _09953_);
  nand (_36282_, _11464_, _09953_);
  and (_36283_, _36282_, _36281_);
  and (_36284_, _36283_, _03644_);
  or (_36285_, _36284_, _11992_);
  or (_36286_, _36285_, _36279_);
  or (_36287_, _36017_, _11991_);
  and (_36288_, _36287_, _03948_);
  and (_36289_, _36288_, _36286_);
  nand (_36290_, _11581_, _03767_);
  nand (_36292_, _36290_, _11998_);
  or (_36293_, _36292_, _36289_);
  or (_36294_, _36017_, _11998_);
  and (_36295_, _36294_, _06855_);
  and (_36296_, _36295_, _36293_);
  nor (_36297_, _06855_, _03440_);
  or (_36298_, _36297_, _03196_);
  or (_36299_, _36298_, _36296_);
  or (_36300_, _11581_, _12009_);
  and (_36301_, _36300_, _03446_);
  and (_36303_, _36301_, _36299_);
  and (_36304_, _36283_, _03445_);
  or (_36305_, _36304_, _12016_);
  or (_36306_, _36305_, _36303_);
  or (_36307_, _36017_, _12015_);
  and (_36308_, _36307_, _03474_);
  and (_36309_, _36308_, _36306_);
  nand (_36310_, _11581_, _03473_);
  nand (_36311_, _36310_, _11392_);
  or (_36312_, _36311_, _36309_);
  or (_36314_, _36017_, _11392_);
  and (_36315_, _36314_, _11391_);
  and (_36316_, _36315_, _36312_);
  not (_36317_, _03194_);
  nand (_36318_, _03440_, _36317_);
  and (_36319_, _36318_, _32181_);
  or (_36320_, _36319_, _36316_);
  or (_36321_, _11581_, _36317_);
  and (_36322_, _36321_, _12035_);
  and (_36323_, _36322_, _36320_);
  and (_36325_, _36017_, _12031_);
  or (_36326_, _36325_, _36323_);
  or (_36327_, _36326_, _43193_);
  or (_36328_, _43189_, \oc8051_golden_model_1.PC [11]);
  and (_36329_, _36328_, _42003_);
  and (_43933_, _36329_, _36327_);
  nor (_36330_, _11578_, _05916_);
  and (_36331_, _11452_, _03224_);
  and (_36332_, _11452_, _10116_);
  and (_36333_, _11547_, _11544_);
  nor (_36335_, _36333_, _11548_);
  and (_36336_, _36335_, _11743_);
  or (_36337_, _36336_, _10112_);
  or (_36338_, _36337_, _36332_);
  or (_36339_, _36335_, _11437_);
  or (_36340_, _11452_, _11439_);
  and (_36341_, _36340_, _03534_);
  and (_36342_, _36341_, _36339_);
  and (_36343_, _11566_, _11578_);
  and (_36344_, _11660_, _11657_);
  nor (_36346_, _36344_, _11661_);
  and (_36347_, _36346_, _32232_);
  or (_36348_, _36347_, _05997_);
  or (_36349_, _36348_, _36343_);
  nor (_36350_, _11397_, \oc8051_golden_model_1.PC [12]);
  nor (_36351_, _36350_, _11398_);
  and (_36352_, _11684_, _11686_);
  or (_36353_, _36352_, _36351_);
  not (_36354_, _11578_);
  nand (_36355_, _36354_, _03536_);
  or (_36357_, _11578_, _10754_);
  nor (_36358_, _04435_, \oc8051_golden_model_1.PC [12]);
  nor (_36359_, _04436_, _03536_);
  and (_36360_, _36359_, _36358_);
  nand (_36361_, _36360_, _11683_);
  and (_36362_, _36361_, _36357_);
  or (_36363_, _36362_, _15022_);
  and (_36364_, _36363_, _36355_);
  or (_36365_, _36364_, _08118_);
  and (_36366_, _36365_, _03209_);
  and (_36368_, _36366_, _36353_);
  or (_36369_, _36354_, _03209_);
  nand (_36370_, _36369_, _05997_);
  or (_36371_, _36370_, _36368_);
  and (_36372_, _36371_, _11705_);
  and (_36373_, _36372_, _36349_);
  or (_36374_, _36373_, _36342_);
  and (_36375_, _36374_, _11430_);
  and (_36376_, _36351_, _11710_);
  or (_36377_, _36376_, _36077_);
  or (_36379_, _36377_, _36375_);
  or (_36380_, _11578_, _11428_);
  and (_36381_, _36380_, _11715_);
  and (_36382_, _36381_, _36379_);
  not (_36383_, _36351_);
  nor (_36384_, _36383_, _11715_);
  or (_36385_, _36384_, _03530_);
  or (_36386_, _36385_, _36382_);
  nand (_36387_, _36354_, _03530_);
  and (_36388_, _36387_, _11723_);
  and (_36390_, _36388_, _36386_);
  nor (_36391_, _36383_, _11723_);
  nor (_36392_, _36391_, _11730_);
  not (_36393_, _36392_);
  nor (_36394_, _36393_, _36390_);
  nor (_36395_, _11729_, _11578_);
  or (_36396_, _36395_, _10021_);
  or (_36397_, _36396_, _36394_);
  and (_36398_, _11453_, _10055_);
  nor (_36399_, _36335_, _10055_);
  or (_36401_, _36399_, _10017_);
  or (_36402_, _36401_, _36398_);
  and (_36403_, _36402_, _10112_);
  and (_36404_, _36403_, _36397_);
  nor (_36405_, _36404_, _03547_);
  and (_36406_, _36405_, _36338_);
  and (_36407_, _36335_, _36105_);
  and (_36408_, _11452_, _09975_);
  nor (_36409_, _36408_, _36407_);
  nor (_36410_, _36409_, _03994_);
  or (_36412_, _36410_, _36406_);
  nand (_36413_, _36412_, _10123_);
  and (_36414_, _11452_, _10163_);
  and (_36415_, _36335_, _11764_);
  or (_36416_, _36415_, _36414_);
  and (_36417_, _36416_, _03608_);
  and (_36418_, _36351_, _10122_);
  not (_36419_, _36418_);
  and (_36420_, _36419_, _11761_);
  not (_36421_, _36420_);
  nor (_36423_, _36421_, _36417_);
  nand (_36424_, _36423_, _36413_);
  nor (_36425_, _11761_, _11578_);
  nor (_36426_, _36425_, _11425_);
  nand (_36427_, _36426_, _36424_);
  nor (_36428_, _36383_, _11424_);
  nor (_36429_, _36428_, _36127_);
  nand (_36430_, _36429_, _36427_);
  nor (_36431_, _11778_, _11578_);
  nor (_36432_, _36431_, _11780_);
  nand (_36434_, _36432_, _36430_);
  nor (_36435_, _36383_, _11419_);
  nor (_36436_, _36435_, _08267_);
  nand (_36437_, _36436_, _36434_);
  nor (_36438_, _11578_, _08266_);
  nor (_36439_, _36438_, _03334_);
  nand (_36440_, _36439_, _36437_);
  nor (_36441_, _36383_, _03233_);
  nor (_36442_, _36441_, _11791_);
  nand (_36443_, _36442_, _36440_);
  nor (_36445_, _11790_, _11578_);
  nor (_36446_, _36445_, _03621_);
  nand (_36447_, _36446_, _36443_);
  and (_36448_, _11452_, _03621_);
  not (_36449_, _36448_);
  and (_36450_, _36449_, _11797_);
  nand (_36451_, _36450_, _36447_);
  nor (_36452_, _11578_, _11797_);
  nor (_36453_, _36452_, _03224_);
  and (_36454_, _36453_, _36451_);
  or (_36456_, _36454_, _36331_);
  nand (_36457_, _36456_, _11806_);
  nor (_36458_, _36383_, _11806_);
  nor (_36459_, _36458_, _11809_);
  nand (_36460_, _36459_, _36457_);
  nor (_36461_, _11808_, _11578_);
  nor (_36462_, _36461_, _11813_);
  nand (_36463_, _36462_, _36460_);
  and (_36464_, _36346_, _11813_);
  nor (_36465_, _36464_, _06193_);
  and (_36467_, _36465_, _36463_);
  or (_36468_, _36467_, _36330_);
  nand (_36469_, _36468_, _04509_);
  and (_36470_, _11453_, _03624_);
  nor (_36471_, _36470_, _08461_);
  and (_36472_, _36471_, _36469_);
  and (_36473_, _11578_, _08461_);
  or (_36474_, _36473_, _36472_);
  nand (_36475_, _36474_, _23814_);
  nor (_36476_, _11856_, \oc8051_golden_model_1.DPH [4]);
  nor (_36478_, _36476_, _11857_);
  and (_36479_, _36478_, _11828_);
  nor (_36480_, _36479_, _11865_);
  nand (_36481_, _36480_, _36475_);
  nor (_36482_, _11864_, _11578_);
  nor (_36483_, _36482_, _11868_);
  and (_36484_, _36483_, _36481_);
  and (_36485_, _11578_, _08864_);
  and (_36486_, _36346_, _11894_);
  or (_36487_, _36486_, _36485_);
  and (_36489_, _36487_, _11868_);
  or (_36490_, _36489_, _36484_);
  nand (_36491_, _36490_, _11416_);
  nor (_36492_, _36383_, _11416_);
  nor (_36493_, _36492_, _08494_);
  nand (_36494_, _36493_, _36491_);
  nor (_36495_, _11578_, _08493_);
  nor (_36496_, _36495_, _03623_);
  nand (_36497_, _36496_, _36494_);
  and (_36498_, _11452_, _03623_);
  nor (_36500_, _36498_, _11886_);
  nand (_36501_, _36500_, _36497_);
  nor (_36502_, _11885_, _11578_);
  nor (_36503_, _36502_, _11889_);
  nand (_36504_, _36503_, _36501_);
  nand (_36505_, _11578_, _11894_);
  nand (_36506_, _36346_, _08864_);
  and (_36507_, _36506_, _36505_);
  or (_36508_, _36507_, _11893_);
  nand (_36509_, _36508_, _36504_);
  nand (_36511_, _36509_, _11902_);
  and (_36512_, _36351_, _11901_);
  nor (_36513_, _36512_, _11905_);
  nand (_36514_, _36513_, _36511_);
  nor (_36515_, _11578_, _11904_);
  nor (_36516_, _36515_, _03611_);
  nand (_36517_, _36516_, _36514_);
  and (_36518_, _11452_, _03611_);
  nor (_36519_, _36518_, _10829_);
  and (_36520_, _36519_, _36517_);
  nor (_36522_, _11915_, _36354_);
  nor (_36523_, _36522_, _24079_);
  nor (_36524_, _36523_, _36520_);
  and (_36525_, _11578_, \oc8051_golden_model_1.PSW [7]);
  and (_36526_, _36346_, _07982_);
  or (_36527_, _36526_, _36525_);
  and (_36528_, _36527_, _11915_);
  or (_36529_, _36528_, _36524_);
  nand (_36530_, _36529_, _11413_);
  nor (_36531_, _36383_, _11413_);
  nor (_36533_, _36531_, _15156_);
  nand (_36534_, _36533_, _36530_);
  nor (_36535_, _11578_, _11410_);
  nor (_36536_, _36535_, _03618_);
  nand (_36537_, _36536_, _36534_);
  and (_36538_, _11452_, _03618_);
  nor (_36539_, _36538_, _11933_);
  and (_36540_, _36539_, _36537_);
  nor (_36541_, _11936_, _36354_);
  nor (_36542_, _36541_, _24227_);
  or (_36544_, _36542_, _36540_);
  nand (_36545_, _11578_, _07982_);
  nand (_36546_, _36346_, \oc8051_golden_model_1.PSW [7]);
  and (_36547_, _36546_, _36545_);
  or (_36548_, _36547_, _11942_);
  nand (_36549_, _36548_, _36544_);
  nand (_36550_, _36549_, _11408_);
  nor (_36551_, _36383_, _11408_);
  nor (_36552_, _36551_, _08629_);
  nand (_36553_, _36552_, _36550_);
  nor (_36555_, _11578_, _08628_);
  nor (_36556_, _36555_, _08707_);
  and (_36557_, _36556_, _36553_);
  and (_36558_, _36351_, _08707_);
  or (_36559_, _36558_, _36557_);
  and (_36560_, _36559_, _10735_);
  nor (_36561_, _05831_, _10735_);
  or (_36562_, _36561_, _03191_);
  or (_36563_, _36562_, _36560_);
  and (_36564_, _36354_, _03191_);
  nor (_36566_, _36564_, _03617_);
  and (_36567_, _36566_, _36563_);
  nor (_36568_, _11453_, _09953_);
  and (_36569_, _36335_, _09953_);
  nor (_36570_, _36569_, _36568_);
  nor (_36571_, _36570_, _03814_);
  or (_36572_, _36571_, _36567_);
  nand (_36573_, _36572_, _11406_);
  nor (_36574_, _36383_, _11406_);
  nor (_36575_, _36574_, _08785_);
  nand (_36577_, _36575_, _36573_);
  nor (_36578_, _11578_, _08784_);
  nor (_36579_, _36578_, _08815_);
  nand (_36580_, _36579_, _36577_);
  and (_36581_, _36351_, _08815_);
  nor (_36582_, _36581_, _03475_);
  nand (_36583_, _36582_, _36580_);
  and (_36584_, _05831_, _03475_);
  nor (_36585_, _36584_, _03189_);
  and (_36586_, _36585_, _36583_);
  and (_36588_, _11578_, _03189_);
  or (_36589_, _36588_, _03644_);
  or (_36590_, _36589_, _36586_);
  and (_36591_, _11453_, _09953_);
  nor (_36592_, _36335_, _09953_);
  nor (_36593_, _36592_, _36591_);
  nor (_36594_, _36593_, _03768_);
  nor (_36595_, _36594_, _11992_);
  nand (_36596_, _36595_, _36590_);
  nor (_36597_, _36383_, _11991_);
  nor (_36599_, _36597_, _03767_);
  nand (_36600_, _36599_, _36596_);
  and (_36601_, _36354_, _03767_);
  nor (_36602_, _36601_, _11999_);
  nand (_36603_, _36602_, _36600_);
  nor (_36604_, _36383_, _11998_);
  nor (_36605_, _36604_, _03645_);
  nand (_36606_, _36605_, _36603_);
  and (_36607_, _04257_, _03645_);
  nor (_36608_, _36607_, _03196_);
  and (_36610_, _36608_, _36606_);
  and (_36611_, _11578_, _03196_);
  or (_36612_, _36611_, _03445_);
  or (_36613_, _36612_, _36610_);
  nor (_36614_, _36593_, _03446_);
  nor (_36615_, _36614_, _12016_);
  nand (_36616_, _36615_, _36613_);
  nor (_36617_, _36383_, _12015_);
  nor (_36618_, _36617_, _03473_);
  nand (_36619_, _36618_, _36616_);
  and (_36621_, _36354_, _03473_);
  nor (_36622_, _36621_, _12022_);
  nand (_36623_, _36622_, _36619_);
  nor (_36624_, _36383_, _11392_);
  nor (_36625_, _36624_, _03615_);
  nand (_36626_, _36625_, _36623_);
  and (_36627_, _04257_, _03615_);
  nor (_36628_, _36627_, _03194_);
  and (_36629_, _36628_, _36626_);
  and (_36630_, _11578_, _03194_);
  or (_36632_, _36630_, _36629_);
  nand (_36633_, _36632_, _12035_);
  and (_36634_, _36351_, _12031_);
  not (_36635_, _36634_);
  and (_36636_, _36635_, _36633_);
  nand (_36637_, _36636_, _43189_);
  or (_36638_, _43189_, \oc8051_golden_model_1.PC [12]);
  and (_36639_, _36638_, _42003_);
  and (_43934_, _36639_, _36637_);
  nor (_36640_, _11398_, \oc8051_golden_model_1.PC [13]);
  nor (_36642_, _36640_, _11399_);
  or (_36643_, _36642_, _11406_);
  or (_36644_, _36642_, _11408_);
  or (_36645_, _36642_, _11413_);
  or (_36646_, _11576_, _11575_);
  not (_36647_, _36646_);
  nor (_36648_, _36647_, _11662_);
  and (_36649_, _36647_, _11662_);
  or (_36650_, _36649_, _36648_);
  or (_36651_, _36650_, _08864_);
  or (_36653_, _11574_, _11894_);
  and (_36654_, _36653_, _11868_);
  and (_36655_, _36654_, _36651_);
  or (_36656_, _11808_, _11574_);
  and (_36657_, _36656_, _11814_);
  and (_36658_, _11448_, _03224_);
  or (_36659_, _36642_, _11419_);
  not (_36660_, _36642_);
  nor (_36661_, _36660_, _11424_);
  and (_36662_, _11574_, _03530_);
  or (_36664_, _11574_, _11428_);
  or (_36665_, _11448_, _11439_);
  or (_36666_, _11450_, _11449_);
  not (_36667_, _36666_);
  nor (_36668_, _36667_, _11549_);
  and (_36669_, _36667_, _11549_);
  or (_36670_, _36669_, _36668_);
  or (_36671_, _36670_, _11437_);
  and (_36672_, _36671_, _03534_);
  and (_36673_, _36672_, _36665_);
  and (_36675_, _11566_, _11574_);
  and (_36676_, _36650_, _32232_);
  or (_36677_, _36676_, _05997_);
  or (_36678_, _36677_, _36675_);
  nand (_36679_, _36660_, _08118_);
  or (_36680_, _36642_, _11680_);
  or (_36681_, _36642_, _11683_);
  nor (_36682_, _04436_, \oc8051_golden_model_1.PC [13]);
  and (_36683_, _36682_, _11686_);
  nand (_36684_, _36683_, _11683_);
  or (_36686_, _36684_, _15022_);
  and (_36687_, _36686_, _36681_);
  or (_36688_, _36687_, _04435_);
  and (_36689_, _36688_, _36680_);
  or (_36690_, _36689_, _03536_);
  and (_36691_, _36690_, _36679_);
  or (_36692_, _36691_, _11677_);
  or (_36693_, _11700_, _11574_);
  and (_36694_, _36693_, _36692_);
  or (_36695_, _36694_, _05998_);
  and (_36697_, _36695_, _11705_);
  and (_36698_, _36697_, _36678_);
  or (_36699_, _36698_, _36673_);
  and (_36700_, _36699_, _11430_);
  and (_36701_, _36642_, _11710_);
  or (_36702_, _36701_, _36077_);
  or (_36703_, _36702_, _36700_);
  and (_36704_, _36703_, _36664_);
  or (_36705_, _36704_, _11716_);
  or (_36706_, _36642_, _11715_);
  and (_36708_, _36706_, _03531_);
  and (_36709_, _36708_, _36705_);
  or (_36710_, _36709_, _36662_);
  and (_36711_, _36710_, _11723_);
  or (_36712_, _36660_, _11723_);
  nand (_36713_, _36712_, _11729_);
  or (_36714_, _36713_, _36711_);
  or (_36715_, _11729_, _11574_);
  and (_36716_, _36715_, _36714_);
  or (_36717_, _36716_, _10021_);
  and (_36719_, _11448_, _10055_);
  not (_36720_, _10055_);
  and (_36721_, _36670_, _36720_);
  or (_36722_, _36721_, _36719_);
  or (_36723_, _36722_, _10017_);
  and (_36724_, _36723_, _10112_);
  and (_36725_, _36724_, _36717_);
  and (_36726_, _36670_, _11743_);
  and (_36727_, _11448_, _10116_);
  or (_36728_, _36727_, _36726_);
  and (_36730_, _36728_, _10020_);
  or (_36731_, _36730_, _03547_);
  or (_36732_, _36731_, _36725_);
  and (_36733_, _11448_, _09975_);
  and (_36734_, _36670_, _36105_);
  or (_36735_, _36734_, _03994_);
  or (_36736_, _36735_, _36733_);
  and (_36737_, _36736_, _10123_);
  and (_36738_, _36737_, _36732_);
  or (_36739_, _36670_, _10163_);
  or (_36741_, _11448_, _11764_);
  and (_36742_, _36741_, _03608_);
  and (_36743_, _36742_, _36739_);
  nand (_36744_, _36642_, _10122_);
  nand (_36745_, _36744_, _11761_);
  or (_36746_, _36745_, _36743_);
  or (_36747_, _36746_, _36738_);
  or (_36748_, _11761_, _11574_);
  and (_36749_, _36748_, _11424_);
  and (_36750_, _36749_, _36747_);
  or (_36752_, _36750_, _36661_);
  and (_36753_, _36752_, _11778_);
  or (_36754_, _11778_, _13259_);
  nand (_36755_, _36754_, _11419_);
  or (_36756_, _36755_, _36753_);
  and (_36757_, _36756_, _36659_);
  or (_36758_, _36757_, _08267_);
  or (_36759_, _11574_, _08266_);
  and (_36760_, _36759_, _03233_);
  and (_36761_, _36760_, _36758_);
  or (_36763_, _36660_, _03233_);
  nand (_36764_, _36763_, _11790_);
  or (_36765_, _36764_, _36761_);
  or (_36766_, _11790_, _11574_);
  and (_36767_, _36766_, _03622_);
  and (_36768_, _36767_, _36765_);
  nand (_36769_, _11448_, _03621_);
  nand (_36770_, _36769_, _11797_);
  or (_36771_, _36770_, _36768_);
  or (_36772_, _11574_, _11797_);
  and (_36774_, _36772_, _03521_);
  and (_36775_, _36774_, _36771_);
  or (_36776_, _36775_, _36658_);
  and (_36777_, _36776_, _11806_);
  nor (_36778_, _36660_, _11806_);
  or (_36779_, _36778_, _11809_);
  or (_36780_, _36779_, _36777_);
  and (_36781_, _36780_, _36657_);
  and (_36782_, _36650_, _11813_);
  or (_36783_, _36782_, _06193_);
  or (_36785_, _36783_, _36781_);
  or (_36786_, _11574_, _05916_);
  and (_36787_, _36786_, _04509_);
  and (_36788_, _36787_, _36785_);
  and (_36789_, _11448_, _03624_);
  or (_36790_, _36789_, _08461_);
  or (_36791_, _36790_, _36788_);
  and (_36792_, _13259_, _08461_);
  nor (_36793_, _36792_, _11828_);
  and (_36794_, _36793_, _36791_);
  or (_36796_, _11857_, \oc8051_golden_model_1.DPH [5]);
  nor (_36797_, _11858_, _23814_);
  and (_36798_, _36797_, _36796_);
  or (_36799_, _36798_, _11865_);
  or (_36800_, _36799_, _36794_);
  or (_36801_, _11864_, _11574_);
  and (_36802_, _36801_, _23819_);
  and (_36803_, _36802_, _36800_);
  or (_36804_, _36803_, _36655_);
  and (_36805_, _36804_, _11416_);
  nor (_36807_, _36660_, _11416_);
  or (_36808_, _36807_, _08494_);
  or (_36809_, _36808_, _36805_);
  or (_36810_, _11574_, _08493_);
  and (_36811_, _36810_, _04527_);
  and (_36812_, _36811_, _36809_);
  nand (_36813_, _11448_, _03623_);
  nand (_36814_, _36813_, _11885_);
  or (_36815_, _36814_, _36812_);
  or (_36816_, _11885_, _11574_);
  and (_36818_, _36816_, _11893_);
  and (_36819_, _36818_, _36815_);
  or (_36820_, _36650_, _11894_);
  or (_36821_, _11574_, _08864_);
  and (_36822_, _36821_, _11889_);
  and (_36823_, _36822_, _36820_);
  or (_36824_, _36823_, _36819_);
  and (_36825_, _36824_, _11902_);
  and (_36826_, _36642_, _11901_);
  or (_36827_, _36826_, _11905_);
  or (_36829_, _36827_, _36825_);
  or (_36830_, _11574_, _11904_);
  and (_36831_, _36830_, _04523_);
  and (_36832_, _36831_, _36829_);
  nand (_36833_, _11448_, _03611_);
  nand (_36834_, _36833_, _10828_);
  or (_36835_, _36834_, _36832_);
  nor (_36836_, _11915_, _13259_);
  or (_36837_, _36836_, _24079_);
  and (_36838_, _36837_, _36835_);
  or (_36840_, _36650_, \oc8051_golden_model_1.PSW [7]);
  or (_36841_, _11574_, _07982_);
  and (_36842_, _36841_, _11915_);
  and (_36843_, _36842_, _36840_);
  or (_36844_, _36843_, _11919_);
  or (_36845_, _36844_, _36838_);
  and (_36846_, _36845_, _36645_);
  or (_36847_, _36846_, _15156_);
  or (_36848_, _11574_, _11410_);
  and (_36849_, _36848_, _06453_);
  and (_36851_, _36849_, _36847_);
  nand (_36852_, _11448_, _03618_);
  nand (_36853_, _36852_, _11932_);
  or (_36854_, _36853_, _36851_);
  nor (_36855_, _11936_, _13259_);
  or (_36856_, _36855_, _24227_);
  and (_36857_, _36856_, _36854_);
  or (_36858_, _36650_, _07982_);
  or (_36859_, _11574_, \oc8051_golden_model_1.PSW [7]);
  and (_36860_, _36859_, _11936_);
  and (_36862_, _36860_, _36858_);
  or (_36863_, _36862_, _11940_);
  or (_36864_, _36863_, _36857_);
  and (_36865_, _36864_, _36644_);
  or (_36866_, _36865_, _08629_);
  or (_36867_, _11574_, _08628_);
  and (_36868_, _36867_, _08708_);
  and (_36869_, _36868_, _36866_);
  and (_36870_, _36642_, _08707_);
  or (_36871_, _36870_, _03752_);
  or (_36873_, _36871_, _36869_);
  nand (_36874_, _05526_, _03752_);
  and (_36875_, _36874_, _36873_);
  or (_36876_, _36875_, _03191_);
  nand (_36877_, _13259_, _03191_);
  and (_36878_, _36877_, _03814_);
  and (_36879_, _36878_, _36876_);
  or (_36880_, _36670_, _36257_);
  or (_36881_, _11448_, _09953_);
  and (_36882_, _36881_, _03617_);
  and (_36884_, _36882_, _36880_);
  or (_36885_, _36884_, _11963_);
  or (_36886_, _36885_, _36879_);
  and (_36887_, _36886_, _36643_);
  or (_36888_, _36887_, _08785_);
  or (_36889_, _11574_, _08784_);
  and (_36890_, _36889_, _08816_);
  and (_36891_, _36890_, _36888_);
  and (_36892_, _36642_, _08815_);
  or (_36893_, _36892_, _03475_);
  or (_36895_, _36893_, _36891_);
  nand (_36896_, _05526_, _03475_);
  and (_36897_, _36896_, _36895_);
  or (_36898_, _36897_, _03189_);
  nand (_36899_, _13259_, _03189_);
  and (_36900_, _36899_, _03768_);
  and (_36901_, _36900_, _36898_);
  or (_36902_, _36670_, _09953_);
  or (_36903_, _11448_, _36257_);
  and (_36904_, _36903_, _36902_);
  and (_36906_, _36904_, _03644_);
  or (_36907_, _36906_, _11992_);
  or (_36908_, _36907_, _36901_);
  or (_36909_, _36642_, _11991_);
  and (_36910_, _36909_, _03948_);
  and (_36911_, _36910_, _36908_);
  nand (_36912_, _11574_, _03767_);
  nand (_36913_, _36912_, _11998_);
  or (_36914_, _36913_, _36911_);
  or (_36915_, _36642_, _11998_);
  and (_36917_, _36915_, _06855_);
  and (_36918_, _36917_, _36914_);
  nor (_36919_, _03811_, _06855_);
  or (_36920_, _36919_, _03196_);
  or (_36921_, _36920_, _36918_);
  nand (_36922_, _13259_, _03196_);
  and (_36923_, _36922_, _03446_);
  and (_36924_, _36923_, _36921_);
  and (_36925_, _36904_, _03445_);
  or (_36926_, _36925_, _12016_);
  or (_36928_, _36926_, _36924_);
  or (_36929_, _36642_, _12015_);
  and (_36930_, _36929_, _03474_);
  and (_36931_, _36930_, _36928_);
  nand (_36932_, _11574_, _03473_);
  nand (_36933_, _36932_, _11392_);
  or (_36934_, _36933_, _36931_);
  or (_36935_, _36642_, _11392_);
  and (_36936_, _36935_, _11391_);
  and (_36937_, _36936_, _36934_);
  nor (_36939_, _03811_, _11391_);
  or (_36940_, _36939_, _03194_);
  or (_36941_, _36940_, _36937_);
  nand (_36942_, _13259_, _03194_);
  and (_36943_, _36942_, _12035_);
  and (_36944_, _36943_, _36941_);
  and (_36945_, _36642_, _12031_);
  or (_36946_, _36945_, _36944_);
  or (_36947_, _36946_, _43193_);
  or (_36948_, _43189_, \oc8051_golden_model_1.PC [13]);
  and (_36950_, _36948_, _42003_);
  and (_43935_, _36950_, _36947_);
  nor (_36951_, _11399_, \oc8051_golden_model_1.PC [14]);
  nor (_36952_, _36951_, _11400_);
  not (_36953_, _36952_);
  and (_36954_, _36953_, _08815_);
  nand (_36955_, _11569_, _03191_);
  nor (_36956_, _36952_, _11408_);
  not (_36957_, _11569_);
  nor (_36958_, _11932_, _36957_);
  nor (_36960_, _36957_, _10828_);
  nor (_36961_, _11885_, _36957_);
  nor (_36962_, _11864_, _36957_);
  or (_36963_, _11761_, _11569_);
  or (_36964_, _36952_, _11715_);
  and (_36965_, _36952_, _04012_);
  and (_36966_, _11566_, _11569_);
  nor (_36967_, _11665_, _11572_);
  nor (_36968_, _36967_, _11666_);
  and (_36969_, _36968_, _32232_);
  or (_36971_, _36969_, _36966_);
  or (_36972_, _36971_, _05997_);
  and (_36973_, _11699_, _11569_);
  and (_36974_, _03204_, \oc8051_golden_model_1.PC [14]);
  and (_36975_, _36974_, _36359_);
  and (_36976_, _36975_, _11683_);
  and (_36977_, _36976_, _11680_);
  or (_36978_, _36977_, _36973_);
  and (_36979_, _36978_, _11686_);
  nor (_36980_, _36953_, _36352_);
  or (_36982_, _36980_, _36979_);
  and (_36983_, _36982_, _03209_);
  or (_36984_, _36957_, _03209_);
  nand (_36985_, _36984_, _05997_);
  or (_36986_, _36985_, _36983_);
  and (_36987_, _36986_, _06008_);
  and (_36988_, _36987_, _36972_);
  or (_36989_, _36988_, _36965_);
  and (_36990_, _36989_, _04432_);
  or (_36991_, _32250_, _11441_);
  and (_36993_, _11551_, _11446_);
  nor (_36994_, _36993_, _11552_);
  or (_36995_, _36994_, _11437_);
  and (_36996_, _36995_, _03534_);
  and (_36997_, _36996_, _36991_);
  or (_36998_, _36997_, _11431_);
  or (_36999_, _36998_, _36990_);
  or (_37000_, _36952_, _11430_);
  and (_37001_, _37000_, _11428_);
  and (_37002_, _37001_, _36999_);
  or (_37004_, _36957_, _11428_);
  nand (_37005_, _37004_, _11715_);
  or (_37006_, _37005_, _37002_);
  and (_37007_, _37006_, _36964_);
  or (_37008_, _37007_, _03530_);
  nand (_37009_, _36957_, _03530_);
  and (_37010_, _37009_, _11723_);
  and (_37011_, _37010_, _37008_);
  nor (_37012_, _36953_, _11723_);
  or (_37013_, _37012_, _37011_);
  and (_37015_, _37013_, _11729_);
  or (_37016_, _11729_, _36957_);
  nand (_37017_, _37016_, _10017_);
  or (_37018_, _37017_, _37015_);
  and (_37019_, _11441_, _10055_);
  not (_37020_, _36994_);
  nor (_37021_, _37020_, _10055_);
  or (_37022_, _37021_, _37019_);
  or (_37023_, _37022_, _10017_);
  and (_37024_, _37023_, _10112_);
  and (_37026_, _37024_, _37018_);
  or (_37027_, _36994_, _10116_);
  or (_37028_, _11441_, _11743_);
  and (_37029_, _37028_, _10020_);
  and (_37030_, _37029_, _37027_);
  or (_37031_, _37030_, _03547_);
  or (_37032_, _37031_, _37026_);
  nor (_37033_, _37020_, _09975_);
  and (_37034_, _11441_, _09975_);
  or (_37035_, _37034_, _03994_);
  or (_37037_, _37035_, _37033_);
  and (_37038_, _37037_, _10123_);
  and (_37039_, _37038_, _37032_);
  or (_37040_, _36994_, _10163_);
  nand (_37041_, _11442_, _10163_);
  and (_37042_, _37041_, _03608_);
  and (_37043_, _37042_, _37040_);
  nand (_37044_, _36952_, _10122_);
  nand (_37045_, _37044_, _11761_);
  or (_37046_, _37045_, _37043_);
  or (_37048_, _37046_, _37039_);
  and (_37049_, _37048_, _36963_);
  or (_37050_, _37049_, _11425_);
  or (_37051_, _36952_, _11424_);
  and (_37052_, _37051_, _11778_);
  and (_37053_, _37052_, _37050_);
  or (_37054_, _11778_, _36957_);
  nand (_37055_, _37054_, _11419_);
  or (_37056_, _37055_, _37053_);
  or (_37057_, _36952_, _11419_);
  and (_37059_, _37057_, _08266_);
  and (_37060_, _37059_, _37056_);
  nor (_37061_, _36957_, _08266_);
  or (_37062_, _37061_, _03334_);
  or (_37063_, _37062_, _37060_);
  or (_37064_, _36952_, _03233_);
  and (_37065_, _37064_, _11790_);
  and (_37066_, _37065_, _37063_);
  nor (_37067_, _11790_, _36957_);
  or (_37068_, _37067_, _03621_);
  or (_37070_, _37068_, _37066_);
  nand (_37071_, _11442_, _03621_);
  and (_37072_, _37071_, _11797_);
  and (_37073_, _37072_, _37070_);
  nor (_37074_, _36957_, _11797_);
  or (_37075_, _37074_, _03224_);
  or (_37076_, _37075_, _37073_);
  nand (_37077_, _11442_, _03224_);
  and (_37078_, _37077_, _11806_);
  and (_37079_, _37078_, _37076_);
  nor (_37081_, _36953_, _11806_);
  or (_37082_, _37081_, _11809_);
  or (_37083_, _37082_, _37079_);
  or (_37084_, _11808_, _11569_);
  and (_37085_, _37084_, _11814_);
  and (_37086_, _37085_, _37083_);
  and (_37087_, _36968_, _11813_);
  or (_37088_, _37087_, _37086_);
  nand (_37089_, _37088_, _05916_);
  or (_37090_, _36957_, _05916_);
  and (_37092_, _37090_, _04509_);
  nand (_37093_, _37092_, _37089_);
  nand (_37094_, _11442_, _03624_);
  and (_37095_, _37094_, _08462_);
  and (_37096_, _37095_, _37093_);
  and (_37097_, _11569_, _08461_);
  or (_37098_, _37097_, _11828_);
  or (_37099_, _37098_, _37096_);
  nor (_37100_, _11858_, \oc8051_golden_model_1.DPH [6]);
  nor (_37101_, _37100_, _11859_);
  or (_37103_, _37101_, _23814_);
  and (_37104_, _37103_, _11864_);
  and (_37105_, _37104_, _37099_);
  or (_37106_, _37105_, _36962_);
  and (_37107_, _37106_, _23819_);
  or (_37108_, _36968_, _08864_);
  or (_37109_, _11569_, _11894_);
  and (_37110_, _37109_, _11868_);
  and (_37111_, _37110_, _37108_);
  or (_37112_, _37111_, _11872_);
  or (_37114_, _37112_, _37107_);
  or (_37115_, _36952_, _11416_);
  and (_37116_, _37115_, _08493_);
  and (_37117_, _37116_, _37114_);
  nor (_37118_, _36957_, _08493_);
  or (_37119_, _37118_, _03623_);
  or (_37120_, _37119_, _37117_);
  nand (_37121_, _11442_, _03623_);
  and (_37122_, _37121_, _11885_);
  and (_37123_, _37122_, _37120_);
  or (_37125_, _37123_, _36961_);
  and (_37126_, _37125_, _11893_);
  or (_37127_, _36968_, _11894_);
  or (_37128_, _11569_, _08864_);
  and (_37129_, _37128_, _11889_);
  and (_37130_, _37129_, _37127_);
  or (_37131_, _37130_, _11901_);
  or (_37132_, _37131_, _37126_);
  nand (_37133_, _36953_, _11901_);
  and (_37134_, _37133_, _11904_);
  and (_37136_, _37134_, _37132_);
  nor (_37137_, _36957_, _11904_);
  or (_37138_, _37137_, _03611_);
  or (_37139_, _37138_, _37136_);
  nand (_37140_, _11442_, _03611_);
  and (_37141_, _37140_, _10828_);
  and (_37142_, _37141_, _37139_);
  or (_37143_, _37142_, _36960_);
  and (_37144_, _37143_, _24078_);
  or (_37145_, _36968_, \oc8051_golden_model_1.PSW [7]);
  or (_37147_, _11569_, _07982_);
  and (_37148_, _37147_, _11915_);
  and (_37149_, _37148_, _37145_);
  or (_37150_, _37149_, _11919_);
  or (_37151_, _37150_, _37144_);
  or (_37152_, _36952_, _11413_);
  and (_37153_, _37152_, _11410_);
  and (_37154_, _37153_, _37151_);
  nor (_37155_, _36957_, _11410_);
  or (_37156_, _37155_, _03618_);
  or (_37158_, _37156_, _37154_);
  nand (_37159_, _11442_, _03618_);
  and (_37160_, _37159_, _11932_);
  and (_37161_, _37160_, _37158_);
  or (_37162_, _37161_, _36958_);
  and (_37163_, _37162_, _11942_);
  or (_37164_, _36968_, _07982_);
  or (_37165_, _11569_, \oc8051_golden_model_1.PSW [7]);
  and (_37166_, _37165_, _11936_);
  and (_37167_, _37166_, _37164_);
  or (_37169_, _37167_, _11940_);
  nor (_37170_, _37169_, _37163_);
  or (_37171_, _37170_, _08629_);
  nor (_37172_, _37171_, _36956_);
  nor (_37173_, _36957_, _08628_);
  nor (_37174_, _37173_, _08707_);
  not (_37175_, _37174_);
  nor (_37176_, _37175_, _37172_);
  and (_37177_, _36953_, _08707_);
  or (_37178_, _37177_, _03752_);
  nor (_37180_, _37178_, _37176_);
  nor (_37181_, _05417_, _10735_);
  or (_37182_, _37181_, _37180_);
  nand (_37183_, _37182_, _04803_);
  and (_37184_, _37183_, _36955_);
  or (_37185_, _37184_, _03617_);
  nor (_37186_, _11441_, _09953_);
  and (_37187_, _37020_, _09953_);
  or (_37188_, _37187_, _03814_);
  or (_37189_, _37188_, _37186_);
  and (_37191_, _37189_, _11406_);
  nand (_37192_, _37191_, _37185_);
  nor (_37193_, _36952_, _11406_);
  nor (_37194_, _37193_, _08785_);
  nand (_37195_, _37194_, _37192_);
  nor (_37196_, _36957_, _08784_);
  nor (_37197_, _37196_, _08815_);
  and (_37198_, _37197_, _37195_);
  or (_37199_, _37198_, _36954_);
  nand (_37200_, _37199_, _03476_);
  and (_37202_, _05417_, _03475_);
  nor (_37203_, _37202_, _03189_);
  and (_37204_, _37203_, _37200_);
  and (_37205_, _11569_, _03189_);
  or (_37206_, _37205_, _03644_);
  nor (_37207_, _37206_, _37204_);
  and (_37208_, _11442_, _09953_);
  nor (_37209_, _36994_, _09953_);
  nor (_37210_, _37209_, _37208_);
  nor (_37211_, _37210_, _03768_);
  or (_37213_, _37211_, _37207_);
  and (_37214_, _37213_, _11991_);
  nor (_37215_, _36952_, _11991_);
  or (_37216_, _37215_, _37214_);
  nand (_37217_, _37216_, _03948_);
  nand (_37218_, _36957_, _03767_);
  and (_37219_, _37218_, _11998_);
  nand (_37220_, _37219_, _37217_);
  nor (_37221_, _36953_, _11998_);
  nor (_37222_, _37221_, _03645_);
  nand (_37224_, _37222_, _37220_);
  and (_37225_, _03645_, _03511_);
  nor (_37226_, _37225_, _03196_);
  nand (_37227_, _37226_, _37224_);
  and (_37228_, _11569_, _03196_);
  nor (_37229_, _37228_, _03445_);
  nand (_37230_, _37229_, _37227_);
  nor (_37231_, _37210_, _03446_);
  nor (_37232_, _37231_, _12016_);
  nand (_37233_, _37232_, _37230_);
  nor (_37235_, _36953_, _12015_);
  nor (_37236_, _37235_, _03473_);
  nand (_37237_, _37236_, _37233_);
  and (_37238_, _36957_, _03473_);
  nor (_37239_, _37238_, _12022_);
  nand (_37240_, _37239_, _37237_);
  nor (_37241_, _36953_, _11392_);
  nor (_37242_, _37241_, _03615_);
  and (_37243_, _37242_, _37240_);
  and (_37244_, _03615_, _03511_);
  or (_37246_, _37244_, _37243_);
  nand (_37247_, _37246_, _36317_);
  and (_37248_, _36957_, _03194_);
  nor (_37249_, _37248_, _12031_);
  nand (_37250_, _37249_, _37247_);
  and (_37251_, _36952_, _12031_);
  not (_37252_, _37251_);
  and (_37253_, _37252_, _37250_);
  nand (_37254_, _37253_, _43189_);
  or (_37255_, _43189_, \oc8051_golden_model_1.PC [14]);
  and (_37257_, _37255_, _42003_);
  and (_43936_, _37257_, _37254_);
  and (_37258_, _43193_, \oc8051_golden_model_1.P0INREG [0]);
  or (_37259_, _37258_, _01134_);
  and (_43939_, _37259_, _42003_);
  and (_37260_, _43193_, \oc8051_golden_model_1.P0INREG [1]);
  or (_37261_, _37260_, _01127_);
  and (_43940_, _37261_, _42003_);
  and (_37262_, _43193_, \oc8051_golden_model_1.P0INREG [2]);
  or (_37263_, _37262_, _01112_);
  and (_43941_, _37263_, _42003_);
  and (_37265_, _43193_, \oc8051_golden_model_1.P0INREG [3]);
  or (_37266_, _37265_, _01120_);
  and (_43942_, _37266_, _42003_);
  and (_37267_, _43193_, \oc8051_golden_model_1.P0INREG [4]);
  or (_37268_, _37267_, _01101_);
  and (_43943_, _37268_, _42003_);
  and (_37269_, _43193_, \oc8051_golden_model_1.P0INREG [5]);
  or (_37270_, _37269_, _01094_);
  and (_43944_, _37270_, _42003_);
  and (_37272_, _43193_, \oc8051_golden_model_1.P0INREG [6]);
  or (_37273_, _37272_, _01079_);
  and (_43945_, _37273_, _42003_);
  and (_37274_, _43193_, \oc8051_golden_model_1.P1INREG [0]);
  or (_37275_, _37274_, _01048_);
  and (_43946_, _37275_, _42003_);
  and (_37276_, _43193_, \oc8051_golden_model_1.P1INREG [1]);
  or (_37277_, _37276_, _01033_);
  and (_43947_, _37277_, _42003_);
  and (_37278_, _43193_, \oc8051_golden_model_1.P1INREG [2]);
  or (_37280_, _37278_, _01055_);
  and (_43948_, _37280_, _42003_);
  and (_37281_, _43193_, \oc8051_golden_model_1.P1INREG [3]);
  or (_37282_, _37281_, _01041_);
  and (_43949_, _37282_, _42003_);
  and (_37283_, _43193_, \oc8051_golden_model_1.P1INREG [4]);
  or (_37284_, _37283_, _01015_);
  and (_43952_, _37284_, _42003_);
  and (_37285_, _43193_, \oc8051_golden_model_1.P1INREG [5]);
  or (_37286_, _37285_, _01000_);
  and (_43953_, _37286_, _42003_);
  and (_37288_, _43193_, \oc8051_golden_model_1.P1INREG [6]);
  or (_37289_, _37288_, _01022_);
  and (_43954_, _37289_, _42003_);
  and (_37290_, _43193_, \oc8051_golden_model_1.P2INREG [0]);
  or (_37291_, _37290_, _00958_);
  and (_43957_, _37291_, _42003_);
  and (_37292_, _43193_, \oc8051_golden_model_1.P2INREG [1]);
  or (_37293_, _37292_, _00965_);
  and (_43958_, _37293_, _42003_);
  and (_37295_, _43193_, \oc8051_golden_model_1.P2INREG [2]);
  or (_37296_, _37295_, _00943_);
  and (_43959_, _37296_, _42003_);
  and (_37297_, _43193_, \oc8051_golden_model_1.P2INREG [3]);
  or (_37298_, _37297_, _00951_);
  and (_43960_, _37298_, _42003_);
  and (_37299_, _43193_, \oc8051_golden_model_1.P2INREG [4]);
  or (_37300_, _37299_, _00925_);
  and (_43961_, _37300_, _42003_);
  and (_37301_, _43193_, \oc8051_golden_model_1.P2INREG [5]);
  or (_37303_, _37301_, _00932_);
  and (_43962_, _37303_, _42003_);
  and (_37304_, _43193_, \oc8051_golden_model_1.P2INREG [6]);
  or (_37305_, _37304_, _00908_);
  and (_43963_, _37305_, _42003_);
  and (_37306_, _43193_, \oc8051_golden_model_1.P3INREG [0]);
  or (_37307_, _37306_, _01168_);
  and (_43964_, _37307_, _42003_);
  and (_37308_, _43193_, \oc8051_golden_model_1.P3INREG [1]);
  or (_37309_, _37308_, _01146_);
  and (_43965_, _37309_, _42003_);
  and (_37311_, _43193_, \oc8051_golden_model_1.P3INREG [2]);
  or (_37312_, _37311_, _01161_);
  and (_43966_, _37312_, _42003_);
  and (_37313_, _43193_, \oc8051_golden_model_1.P3INREG [3]);
  or (_37314_, _37313_, _01154_);
  and (_43967_, _37314_, _42003_);
  and (_37315_, _43193_, \oc8051_golden_model_1.P3INREG [4]);
  or (_37316_, _37315_, _01201_);
  and (_43968_, _37316_, _42003_);
  and (_37318_, _43193_, \oc8051_golden_model_1.P3INREG [5]);
  or (_37319_, _37318_, _01179_);
  and (_43969_, _37319_, _42003_);
  and (_37320_, _43193_, \oc8051_golden_model_1.P3INREG [6]);
  or (_37321_, _37320_, _01194_);
  and (_43972_, _37321_, _42003_);
  and (_00007_[6], _01195_, _42003_);
  and (_00007_[5], _01180_, _42003_);
  and (_00007_[4], _01202_, _42003_);
  and (_00007_[3], _01155_, _42003_);
  and (_00007_[2], _01162_, _42003_);
  and (_00007_[1], _01147_, _42003_);
  and (_00007_[0], _01169_, _42003_);
  and (_00006_[6], _00909_, _42003_);
  and (_00006_[5], _00933_, _42003_);
  and (_00006_[4], _00926_, _42003_);
  and (_00006_[3], _00952_, _42003_);
  and (_00006_[2], _00944_, _42003_);
  and (_00006_[1], _00966_, _42003_);
  and (_00006_[0], _00959_, _42003_);
  and (_00005_[6], _01023_, _42003_);
  and (_00005_[5], _01001_, _42003_);
  and (_00005_[4], _01016_, _42003_);
  and (_00005_[3], _01042_, _42003_);
  and (_00005_[2], _01056_, _42003_);
  and (_00005_[1], _01034_, _42003_);
  and (_00005_[0], _01049_, _42003_);
  and (_00003_[6], _01080_, _42003_);
  and (_00003_[5], _01095_, _42003_);
  and (_00003_[4], _01102_, _42003_);
  and (_00003_[3], _01121_, _42003_);
  and (_00003_[2], _01113_, _42003_);
  and (_00003_[1], _01128_, _42003_);
  and (_00003_[0], _01135_, _42003_);
  or (_37325_, _10723_, _09305_);
  nor (_37326_, _37325_, _10977_);
  not (_37327_, _28794_);
  and (_37328_, _37327_, _28561_);
  nor (_37329_, _29139_, _29024_);
  and (_37330_, _37329_, _37328_);
  nor (_37332_, _27154_, _26921_);
  nor (_37333_, _27499_, _27385_);
  and (_37334_, _37333_, _37332_);
  nor (_37335_, _19662_, _19429_);
  nor (_37336_, _20004_, _19891_);
  and (_37337_, _37336_, _37335_);
  and (_37338_, _37337_, _37334_);
  and (_37339_, _37338_, _37330_);
  not (_37340_, _11387_);
  and (_37341_, _18521_, _37340_);
  nor (_37343_, _19545_, _18749_);
  and (_37344_, _37343_, _37341_);
  nor (_37345_, _11141_, _11060_);
  nor (_37346_, _11305_, _11223_);
  and (_37347_, _37346_, _37345_);
  and (_37348_, _37347_, _37344_);
  not (_37349_, _28451_);
  or (_37350_, _37349_, _27037_);
  or (_37351_, _37350_, _28677_);
  nor (_37352_, _37351_, _18982_);
  and (_37354_, _37352_, _37348_);
  nor (_37355_, _18866_, _18634_);
  nor (_37356_, _19209_, _19095_);
  and (_37357_, _37356_, _37355_);
  nor (_37358_, _30795_, _30177_);
  nor (_37359_, _32005_, _31399_);
  and (_37360_, _37359_, _37358_);
  nor (_37361_, _30532_, _29914_);
  nor (_37362_, _31740_, _31137_);
  nand (_37363_, _37362_, _37361_);
  nor (_37365_, _37363_, _25915_);
  nor (_37366_, _29569_, _26528_);
  and (_37367_, _37366_, _37365_);
  and (_37368_, _37367_, _37360_);
  nor (_37369_, _10612_, _10531_);
  and (_37370_, _37369_, _37368_);
  or (_37371_, _32091_, _31572_);
  or (_37372_, _37371_, _32176_);
  or (_37373_, _37372_, _19317_);
  nor (_37374_, _37373_, _26810_);
  nor (_37376_, _30707_, _30089_);
  nor (_37377_, _31915_, _31311_);
  nand (_37378_, _37377_, _37376_);
  nor (_37379_, _37378_, _26003_);
  nor (_37380_, _26615_, _26089_);
  and (_37381_, _37380_, _37379_);
  nor (_37382_, _30621_, _30002_);
  nor (_37383_, _31830_, _31224_);
  nand (_37384_, _37383_, _37382_);
  nor (_37385_, _37384_, _25649_);
  nor (_37387_, _29306_, _26260_);
  and (_37388_, _37387_, _37385_);
  nor (_37389_, _26438_, _26350_);
  nor (_37390_, _29480_, _29394_);
  and (_37391_, _37390_, _37389_);
  nor (_37392_, _25826_, _25739_);
  nor (_37393_, _30433_, _29826_);
  nor (_37394_, _31653_, _31052_);
  and (_37395_, _37394_, _37393_);
  nor (_37396_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_37398_, \oc8051_golden_model_1.IE [2], \oc8051_golden_model_1.IP [6]);
  and (_37399_, _37398_, _37396_);
  nor (_37400_, \oc8051_golden_model_1.IP [3], \oc8051_golden_model_1.IP [2]);
  nor (_37401_, \oc8051_golden_model_1.IP [5], \oc8051_golden_model_1.IP [4]);
  and (_37402_, _37401_, _37400_);
  and (_37403_, _37402_, _37399_);
  nor (_37404_, \oc8051_golden_model_1.SBUF [1], \oc8051_golden_model_1.SBUF [0]);
  nor (_37405_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  and (_37406_, _37405_, _37404_);
  nor (_37407_, \oc8051_golden_model_1.IE [4], \oc8051_golden_model_1.IE [3]);
  nor (_37409_, \oc8051_golden_model_1.IE [6], \oc8051_golden_model_1.IE [5]);
  and (_37410_, _37409_, _37407_);
  and (_37411_, _37410_, _37406_);
  and (_37412_, _37411_, _37403_);
  nor (_37413_, \oc8051_golden_model_1.IP [7], rst);
  nor (_37414_, \oc8051_golden_model_1.SBUF [7], \oc8051_golden_model_1.IE [7]);
  nor (_37415_, \oc8051_golden_model_1.TH1 [7], \oc8051_golden_model_1.SCON [7]);
  and (_37416_, _37415_, _37414_);
  and (_37417_, _37416_, _37413_);
  nor (_37418_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37420_, \oc8051_golden_model_1.PCON [7], \oc8051_golden_model_1.TCON [7]);
  and (_37421_, _37420_, _37418_);
  nor (_37422_, \oc8051_golden_model_1.TH0 [7], \oc8051_golden_model_1.TL1 [7]);
  nor (_37423_, \oc8051_golden_model_1.TMOD [7], \oc8051_golden_model_1.TL0 [7]);
  and (_37424_, _37423_, _37422_);
  and (_37425_, _37424_, _37421_);
  and (_37426_, _37425_, _37417_);
  and (_37427_, _37426_, _37412_);
  nor (_37428_, \oc8051_golden_model_1.TH0 [1], \oc8051_golden_model_1.TH0 [0]);
  nor (_37429_, \oc8051_golden_model_1.TH0 [3], \oc8051_golden_model_1.TH0 [2]);
  and (_37431_, _37429_, _37428_);
  nor (_37432_, \oc8051_golden_model_1.TH0 [5], \oc8051_golden_model_1.TH0 [4]);
  nor (_37433_, \oc8051_golden_model_1.TL0 [0], \oc8051_golden_model_1.TH0 [6]);
  and (_37434_, _37433_, _37432_);
  and (_37435_, _37434_, _37431_);
  nor (_37436_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37437_, \oc8051_golden_model_1.TL1 [6], \oc8051_golden_model_1.TL1 [3]);
  and (_37438_, _37437_, _37436_);
  nor (_37439_, \oc8051_golden_model_1.TL1 [0], \oc8051_golden_model_1.TH1 [6]);
  nor (_37440_, \oc8051_golden_model_1.TL1 [2], \oc8051_golden_model_1.TL1 [1]);
  and (_37442_, _37440_, _37439_);
  and (_37443_, _37442_, _37438_);
  and (_37444_, _37443_, _37435_);
  nor (_37445_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37446_, \oc8051_golden_model_1.SCON [4], \oc8051_golden_model_1.SCON [1]);
  and (_37447_, _37446_, _37445_);
  nor (_37448_, \oc8051_golden_model_1.SBUF [5], \oc8051_golden_model_1.SBUF [4]);
  nor (_37449_, \oc8051_golden_model_1.SCON [0], \oc8051_golden_model_1.SBUF [6]);
  and (_37450_, _37449_, _37448_);
  and (_37451_, _37450_, _37447_);
  nor (_37453_, \oc8051_golden_model_1.TH1 [3], \oc8051_golden_model_1.TH1 [2]);
  nor (_37454_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  and (_37455_, _37454_, _37453_);
  nor (_37456_, \oc8051_golden_model_1.TH1 [1], \oc8051_golden_model_1.TH1 [0]);
  nor (_37457_, \oc8051_golden_model_1.SCON [6], \oc8051_golden_model_1.SCON [5]);
  and (_37458_, _37457_, _37456_);
  and (_37459_, _37458_, _37455_);
  and (_37460_, _37459_, _37451_);
  and (_37461_, _37460_, _37444_);
  nor (_37462_, \oc8051_golden_model_1.PCON [5], \oc8051_golden_model_1.PCON [4]);
  and (_37464_, regs_always_zero, _26007_);
  and (_37465_, _37464_, _37462_);
  nor (_37466_, \oc8051_golden_model_1.PCON [1], \oc8051_golden_model_1.PCON [0]);
  nor (_37467_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  and (_37468_, _37467_, _37466_);
  nor (_37469_, \oc8051_golden_model_1.TCON [4], \oc8051_golden_model_1.TCON [3]);
  nor (_37470_, \oc8051_golden_model_1.TCON [6], \oc8051_golden_model_1.TCON [5]);
  and (_37471_, _37470_, _37469_);
  and (_37472_, _37471_, _37468_);
  and (_37473_, _37472_, _37465_);
  nor (_37475_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37476_, \oc8051_golden_model_1.TL0 [6], \oc8051_golden_model_1.TL0 [5]);
  and (_37477_, _37476_, _37475_);
  nor (_37478_, \oc8051_golden_model_1.TL0 [2], \oc8051_golden_model_1.TL0 [1]);
  nor (_37479_, \oc8051_golden_model_1.TL0 [4], \oc8051_golden_model_1.TL0 [3]);
  and (_37480_, _37479_, _37478_);
  and (_37481_, _37480_, _37477_);
  nor (_37482_, \oc8051_golden_model_1.TCON [0], \oc8051_golden_model_1.TMOD [6]);
  and (_37483_, _28565_, \oc8051_golden_model_1.TCON [1]);
  and (_37484_, _37483_, _37482_);
  nor (_37486_, \oc8051_golden_model_1.TMOD [3], \oc8051_golden_model_1.TMOD [2]);
  nor (_37487_, \oc8051_golden_model_1.TMOD [5], \oc8051_golden_model_1.TMOD [4]);
  and (_37488_, _37487_, _37486_);
  and (_37489_, _37488_, _37484_);
  and (_37490_, _37489_, _37481_);
  and (_37491_, _37490_, _37473_);
  and (_37492_, _37491_, _37461_);
  nand (_37493_, _37492_, _37427_);
  nor (_37494_, _37493_, _25561_);
  nor (_37495_, _29219_, _26171_);
  and (_37497_, _37495_, _37494_);
  and (_37498_, _37497_, _37395_);
  and (_37499_, _37498_, _37392_);
  and (_37500_, _37499_, _37391_);
  and (_37501_, _37500_, _37388_);
  and (_37502_, _37501_, _37381_);
  nor (_37503_, _30882_, _30350_);
  nor (_37504_, _31486_, _30969_);
  and (_37505_, _37504_, _37503_);
  nor (_37506_, _29655_, _26703_);
  nor (_37508_, _30264_, _29743_);
  and (_37509_, _37508_, _37506_);
  and (_37510_, _37509_, _37505_);
  and (_37511_, _37510_, _37502_);
  and (_37512_, _37511_, _37374_);
  and (_37513_, _37512_, _37370_);
  and (_37514_, _37513_, _37357_);
  and (_37515_, _37514_, _37354_);
  or (_37516_, _27269_, _19778_);
  or (_37517_, _37516_, _28910_);
  nor (_37519_, _37517_, _09198_);
  and (_37520_, _37519_, _37515_);
  and (_37521_, _37520_, _37339_);
  and (_37522_, _37521_, _37326_);
  nor (_37523_, _38653_, _10736_);
  nor (_37524_, _38697_, \oc8051_golden_model_1.SP [6]);
  nor (_37525_, _37524_, _37523_);
  and (_37526_, _38653_, _10736_);
  and (_37527_, _38697_, \oc8051_golden_model_1.SP [6]);
  nor (_37528_, _37527_, _37526_);
  and (_37530_, _37528_, _37525_);
  and (_37531_, _38691_, \oc8051_golden_model_1.SP [5]);
  nor (_37532_, _38691_, \oc8051_golden_model_1.SP [5]);
  nor (_37533_, _37532_, _37531_);
  nor (_37534_, _38679_, \oc8051_golden_model_1.SP [3]);
  and (_37535_, _38679_, \oc8051_golden_model_1.SP [3]);
  nor (_37536_, _37535_, _37534_);
  nor (_37537_, _38661_, \oc8051_golden_model_1.SP [0]);
  and (_37538_, _38661_, \oc8051_golden_model_1.SP [0]);
  nor (_37539_, _37538_, _37537_);
  and (_37541_, _38667_, \oc8051_golden_model_1.SP [1]);
  nor (_37542_, _38667_, \oc8051_golden_model_1.SP [1]);
  nor (_37543_, _37542_, _37541_);
  and (_37544_, _37543_, _37539_);
  nor (_37545_, _38673_, \oc8051_golden_model_1.SP [2]);
  and (_37546_, _38673_, \oc8051_golden_model_1.SP [2]);
  nor (_37547_, _37546_, _37545_);
  and (_37548_, _37547_, _37544_);
  and (_37549_, _37548_, _37536_);
  nor (_37550_, _38685_, \oc8051_golden_model_1.SP [4]);
  and (_37552_, _38685_, \oc8051_golden_model_1.SP [4]);
  nor (_37553_, _37552_, _37550_);
  and (_37554_, _37553_, _37549_);
  and (_37555_, _37554_, _37533_);
  and (_37556_, _37555_, _37530_);
  nor (_37557_, _37556_, property_valid_sp_1_r);
  nor (_37558_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_37559_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37560_, _37559_, _37558_);
  nor (_37561_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37563_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_37564_, _37563_, _37561_);
  nor (_37565_, _37564_, _37560_);
  and (_37566_, \oc8051_golden_model_1.IRAM[5] [5], _41245_);
  and (_37567_, _05492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_37568_, _37567_, _37566_);
  and (_37569_, _05797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_37570_, \oc8051_golden_model_1.IRAM[5] [4], _41242_);
  nor (_37571_, _37570_, _37569_);
  and (_37572_, _37571_, _37568_);
  and (_37574_, _37572_, _37565_);
  nor (_37575_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_37576_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_37577_, _37576_, _37575_);
  not (_37578_, _37577_);
  and (_37579_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_37580_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_37581_, _37580_, _37579_);
  and (_37582_, _37581_, _37578_);
  nor (_37583_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_37585_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_37586_, _37585_, _37583_);
  nand (_37587_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_37588_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_37589_, _37588_, _37587_);
  nor (_37590_, _37589_, _37586_);
  and (_37591_, _37590_, _37582_);
  and (_37592_, _37591_, _37574_);
  and (_37593_, _05031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_37594_, \oc8051_golden_model_1.IRAM[7] [2], _41284_);
  nor (_37596_, _37594_, _37593_);
  nand (_37597_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_37598_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37599_, _37598_, _37597_);
  not (_37600_, _37599_);
  and (_37601_, _37600_, _37596_);
  and (_37602_, _05207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_37603_, \oc8051_golden_model_1.IRAM[7] [7], _40925_);
  nor (_37604_, _37603_, _37602_);
  nand (_37605_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_37607_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_37608_, _37607_, _37605_);
  not (_37609_, _37608_);
  and (_37610_, _37609_, _37604_);
  and (_37611_, _37610_, _37601_);
  nor (_37612_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37613_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_37614_, _37613_, _37612_);
  nor (_37615_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37616_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_37618_, _37616_, _37615_);
  nor (_37619_, _37618_, _37614_);
  and (_37620_, _05791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_37621_, \oc8051_golden_model_1.IRAM[6] [4], _41265_);
  nor (_37622_, _37621_, _37620_);
  and (_37623_, _05486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_37624_, \oc8051_golden_model_1.IRAM[6] [5], _41268_);
  nor (_37625_, _37624_, _37623_);
  and (_37626_, _37625_, _37622_);
  and (_37627_, _37626_, _37619_);
  and (_37629_, _37627_, _37611_);
  and (_37630_, _37629_, _37592_);
  nor (_37631_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_37632_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37633_, _37632_, _37631_);
  not (_37634_, _37633_);
  and (_37635_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37636_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_37637_, _37636_, _37635_);
  and (_37638_, _37637_, _37634_);
  nor (_37640_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_37641_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_37642_, _37641_, _37640_);
  not (_37643_, _37642_);
  and (_37644_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_37645_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_37646_, _37645_, _37644_);
  and (_37647_, _37646_, _37643_);
  and (_37648_, _37647_, _37638_);
  and (_37649_, _03958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_37651_, \oc8051_golden_model_1.IRAM[0] [0], _41068_);
  nor (_37652_, _37651_, _37649_);
  and (_37653_, _04578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_37654_, \oc8051_golden_model_1.IRAM[0] [1], _41081_);
  nor (_37655_, _37654_, _37653_);
  and (_37656_, _37655_, _37652_);
  nor (_37657_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_37658_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_37659_, _37658_, _37657_);
  nor (_37660_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_37662_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37663_, _37662_, _37660_);
  nor (_37664_, _37663_, _37659_);
  and (_37665_, _37664_, _37656_);
  and (_37666_, _37665_, _37648_);
  and (_37667_, _04375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_37668_, \oc8051_golden_model_1.IRAM[3] [0], _41189_);
  nor (_37669_, _37668_, _37667_);
  and (_37670_, _04584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_37671_, \oc8051_golden_model_1.IRAM[3] [1], _41192_);
  nor (_37673_, _37671_, _37670_);
  and (_37674_, _37673_, _37669_);
  nor (_37675_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_37676_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_37677_, _37676_, _37675_);
  nor (_37678_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_37679_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_37680_, _37679_, _37678_);
  nor (_37681_, _37680_, _37677_);
  and (_37682_, _37681_, _37674_);
  and (_37684_, _05025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_37685_, \oc8051_golden_model_1.IRAM[2] [2], _41171_);
  nor (_37686_, _37685_, _37684_);
  nand (_37687_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_37688_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_37689_, _37688_, _37687_);
  not (_37690_, _37689_);
  and (_37691_, _37690_, _37686_);
  and (_37692_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_37693_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_37695_, _37693_, _37692_);
  and (_37696_, _05201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_37697_, \oc8051_golden_model_1.IRAM[2] [7], _41185_);
  nor (_37698_, _37697_, _37696_);
  and (_37699_, _37698_, _37695_);
  and (_37700_, _37699_, _37691_);
  and (_37701_, _37700_, _37682_);
  and (_37702_, _37701_, _37666_);
  and (_37703_, _37702_, _37630_);
  nor (_37704_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_37706_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_37707_, _37706_, _37704_);
  not (_37708_, _37707_);
  and (_37709_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_37710_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_37711_, _37710_, _37709_);
  and (_37712_, _37711_, _37708_);
  nor (_37713_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_37714_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_37715_, _37714_, _37713_);
  nand (_37717_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_37718_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_37719_, _37718_, _37717_);
  nor (_37720_, _37719_, _37715_);
  and (_37721_, _37720_, _37712_);
  and (_37722_, _04420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_37723_, \oc8051_golden_model_1.IRAM[12] [0], _41390_);
  nor (_37724_, _37723_, _37722_);
  and (_37725_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_37726_, \oc8051_golden_model_1.IRAM[12] [1], _41393_);
  nor (_37728_, _37726_, _37725_);
  and (_37729_, _37728_, _37724_);
  nor (_37730_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_37731_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_37732_, _37731_, _37730_);
  nor (_37733_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_37734_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_37735_, _37734_, _37733_);
  nor (_37736_, _37735_, _37732_);
  and (_37737_, _37736_, _37729_);
  and (_37739_, _37737_, _37721_);
  and (_37740_, _04415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37741_, \oc8051_golden_model_1.IRAM[15] [0], _41482_);
  nor (_37742_, _37741_, _37740_);
  and (_37743_, \oc8051_golden_model_1.IRAM[15] [1], _41485_);
  and (_37744_, _04621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_37745_, _37744_, _37743_);
  and (_37746_, _37745_, _37742_);
  nor (_37747_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_37748_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_37750_, _37748_, _37747_);
  nor (_37751_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_37752_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_37753_, _37752_, _37751_);
  nor (_37754_, _37753_, _37750_);
  and (_37755_, _37754_, _37746_);
  and (_37756_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_37757_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_37758_, _37757_, _37756_);
  and (_37759_, \oc8051_golden_model_1.IRAM[14] [2], _41466_);
  and (_37761_, _05061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_37762_, _37761_, _37759_);
  and (_37763_, _37762_, _37758_);
  and (_37764_, _05239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_37765_, \oc8051_golden_model_1.IRAM[14] [7], _40998_);
  nor (_37766_, _37765_, _37764_);
  nand (_37767_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_37768_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_37769_, _37768_, _37767_);
  not (_37770_, _37769_);
  and (_37772_, _37770_, _37766_);
  and (_37773_, _37772_, _37763_);
  and (_37774_, _37773_, _37755_);
  and (_37775_, _37774_, _37739_);
  and (_37776_, _05506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_37777_, \oc8051_golden_model_1.IRAM[9] [5], _41335_);
  nor (_37778_, _37777_, _37776_);
  and (_37779_, _05811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_37780_, \oc8051_golden_model_1.IRAM[9] [4], _41332_);
  nor (_37781_, _37780_, _37779_);
  and (_37783_, _37781_, _37778_);
  nor (_37784_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_37785_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_37786_, _37785_, _37784_);
  nor (_37787_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_37788_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_37789_, _37788_, _37787_);
  nor (_37790_, _37789_, _37786_);
  and (_37791_, _37790_, _37783_);
  nor (_37792_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_37794_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_37795_, _37794_, _37792_);
  nor (_37796_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_37797_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37798_, _37797_, _37796_);
  nor (_37799_, _37798_, _37795_);
  nor (_37800_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_37801_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_37802_, _37801_, _37800_);
  nor (_37803_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_37805_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_37806_, _37805_, _37803_);
  nor (_37807_, _37806_, _37802_);
  and (_37808_, _37807_, _37799_);
  and (_37809_, _37808_, _37791_);
  and (_37810_, \oc8051_golden_model_1.IRAM[11] [2], _41373_);
  and (_37811_, _05047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_37812_, _37811_, _37810_);
  nand (_37813_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_37814_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_37816_, _37814_, _37813_);
  not (_37817_, _37816_);
  and (_37818_, _37817_, _37812_);
  nor (_37819_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_37820_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_37821_, _37820_, _37819_);
  not (_37822_, _37821_);
  and (_37823_, _05223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_37824_, \oc8051_golden_model_1.IRAM[11] [7], _41386_);
  nor (_37825_, _37824_, _37823_);
  and (_37827_, _37825_, _37822_);
  and (_37828_, _37827_, _37818_);
  nor (_37829_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37830_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_37831_, _37830_, _37829_);
  nor (_37832_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37833_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_37834_, _37833_, _37832_);
  nor (_37835_, _37834_, _37831_);
  and (_37836_, \oc8051_golden_model_1.IRAM[10] [4], _41355_);
  and (_37838_, _05806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_37839_, _37838_, _37836_);
  and (_37840_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_37841_, \oc8051_golden_model_1.IRAM[10] [5], _41358_);
  nor (_37842_, _37841_, _37840_);
  and (_37843_, _37842_, _37839_);
  and (_37844_, _37843_, _37835_);
  and (_37845_, _37844_, _37828_);
  and (_37846_, _37845_, _37809_);
  and (_37847_, _37846_, _37775_);
  and (_37849_, _37847_, _37703_);
  nor (_37850_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_37851_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37852_, _37851_, _37850_);
  not (_37853_, _37852_);
  and (_37854_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37855_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_37856_, _37855_, _37854_);
  and (_37857_, _37856_, _37853_);
  nor (_37858_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_37860_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_37861_, _37860_, _37858_);
  nand (_37862_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_37863_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_37864_, _37863_, _37862_);
  nor (_37865_, _37864_, _37861_);
  and (_37866_, _37865_, _37857_);
  and (_37867_, _04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37868_, \oc8051_golden_model_1.IRAM[4] [0], _41212_);
  nor (_37869_, _37868_, _37867_);
  and (_37871_, _04599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_37872_, \oc8051_golden_model_1.IRAM[4] [1], _41215_);
  nor (_37873_, _37872_, _37871_);
  and (_37874_, _37873_, _37869_);
  nor (_37875_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_37876_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_37877_, _37876_, _37875_);
  nor (_37878_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_37879_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_37880_, _37879_, _37878_);
  nor (_37882_, _37880_, _37877_);
  and (_37883_, _37882_, _37874_);
  and (_37884_, _37883_, _37866_);
  and (_37885_, _04593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37886_, \oc8051_golden_model_1.IRAM[7] [1], _41281_);
  nor (_37887_, _37886_, _37885_);
  and (_37888_, _04386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37889_, \oc8051_golden_model_1.IRAM[7] [0], _41278_);
  nor (_37890_, _37889_, _37888_);
  and (_37891_, _37890_, _37887_);
  nor (_37893_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_37894_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_37895_, _37894_, _37893_);
  nor (_37896_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_37897_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_37898_, _37897_, _37896_);
  nor (_37899_, _37898_, _37895_);
  and (_37900_, _37899_, _37891_);
  and (_37901_, \oc8051_golden_model_1.IRAM[6] [2], _41259_);
  and (_37902_, _05033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_37904_, _37902_, _37901_);
  nand (_37905_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_37906_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37907_, _37906_, _37905_);
  not (_37908_, _37907_);
  and (_37909_, _37908_, _37904_);
  and (_37910_, _05209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_37911_, \oc8051_golden_model_1.IRAM[6] [7], _41274_);
  nor (_37912_, _37911_, _37910_);
  nand (_37913_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_37915_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_37916_, _37915_, _37913_);
  not (_37917_, _37916_);
  and (_37918_, _37917_, _37912_);
  and (_37919_, _37918_, _37909_);
  and (_37920_, _37919_, _37900_);
  and (_37921_, _37920_, _37884_);
  nor (_37922_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_37923_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37924_, _37923_, _37922_);
  nor (_37926_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_37927_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37928_, _37927_, _37926_);
  nor (_37929_, _37928_, _37924_);
  and (_37930_, _05777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_37931_, \oc8051_golden_model_1.IRAM[1] [4], _41152_);
  nor (_37932_, _37931_, _37930_);
  and (_37933_, _05472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_37934_, \oc8051_golden_model_1.IRAM[1] [5], _41156_);
  nor (_37935_, _37934_, _37933_);
  and (_37937_, _37935_, _37932_);
  and (_37938_, _37937_, _37929_);
  nor (_37939_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37940_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_37941_, _37940_, _37939_);
  nor (_37942_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37943_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_37944_, _37943_, _37942_);
  nor (_37945_, _37944_, _37941_);
  nor (_37946_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_37948_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_37949_, _37948_, _37946_);
  nor (_37950_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37951_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_37952_, _37951_, _37950_);
  nor (_37953_, _37952_, _37949_);
  and (_37954_, _37953_, _37945_);
  and (_37955_, _37954_, _37938_);
  and (_37956_, \oc8051_golden_model_1.IRAM[3] [2], _41195_);
  and (_37957_, _05023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37959_, _37957_, _37956_);
  nand (_37960_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_37961_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_37962_, _37961_, _37960_);
  not (_37963_, _37962_);
  and (_37964_, _37963_, _37959_);
  nor (_37965_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_37966_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_37967_, _37966_, _37965_);
  not (_37968_, _37967_);
  and (_37970_, _05199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_37971_, \oc8051_golden_model_1.IRAM[3] [7], _40889_);
  nor (_37972_, _37971_, _37970_);
  and (_37973_, _37972_, _37968_);
  and (_37974_, _37973_, _37964_);
  nor (_37975_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_37976_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37977_, _37976_, _37975_);
  nor (_37978_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37979_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_37981_, _37979_, _37978_);
  nor (_37982_, _37981_, _37977_);
  and (_37983_, _05478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_37984_, \oc8051_golden_model_1.IRAM[2] [5], _41180_);
  nor (_37985_, _37984_, _37983_);
  and (_37986_, _05783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_37987_, \oc8051_golden_model_1.IRAM[2] [4], _41177_);
  nor (_37988_, _37987_, _37986_);
  and (_37989_, _37988_, _37985_);
  and (_37990_, _37989_, _37982_);
  and (_37992_, _37990_, _37974_);
  and (_37993_, _37992_, _37955_);
  and (_37994_, _37993_, _37921_);
  nor (_37995_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37996_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_37997_, _37996_, _37995_);
  nor (_37998_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_37999_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_38000_, _37999_, _37998_);
  nor (_38001_, _38000_, _37997_);
  and (_38003_, \oc8051_golden_model_1.IRAM[13] [5], _41452_);
  and (_38004_, _05518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_38005_, _38004_, _38003_);
  and (_38006_, \oc8051_golden_model_1.IRAM[13] [4], _41448_);
  and (_38007_, _05823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_38008_, _38007_, _38006_);
  and (_38009_, _38008_, _38005_);
  and (_38010_, _38009_, _38001_);
  nor (_38011_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_38012_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_38014_, _38012_, _38011_);
  nand (_38015_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_38016_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_38017_, _38016_, _38015_);
  nor (_38018_, _38017_, _38014_);
  nor (_38019_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38020_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_38021_, _38020_, _38019_);
  nand (_38022_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_38023_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_38025_, _38023_, _38022_);
  nor (_38026_, _38025_, _38021_);
  and (_38027_, _38026_, _38018_);
  and (_38028_, _38027_, _38010_);
  and (_38029_, _05059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_38030_, \oc8051_golden_model_1.IRAM[15] [2], _41488_);
  nor (_38031_, _38030_, _38029_);
  and (_38032_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_38033_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_38034_, _38033_, _38032_);
  and (_38036_, _38034_, _38031_);
  and (_38037_, _05237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38038_, \oc8051_golden_model_1.IRAM[15] [7], _41052_);
  nor (_38039_, _38038_, _38037_);
  nand (_38040_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_38041_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38042_, _38041_, _38040_);
  not (_38043_, _38042_);
  and (_38044_, _38043_, _38039_);
  and (_38045_, _38044_, _38036_);
  nor (_38047_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_38048_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_38049_, _38048_, _38047_);
  nor (_38050_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_38051_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_38052_, _38051_, _38050_);
  nor (_38053_, _38052_, _38049_);
  and (_38054_, \oc8051_golden_model_1.IRAM[14] [5], _41474_);
  and (_38055_, _05513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_38056_, _38055_, _38054_);
  and (_38058_, _05818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38059_, \oc8051_golden_model_1.IRAM[14] [4], _41471_);
  nor (_38060_, _38059_, _38058_);
  and (_38061_, _38060_, _38056_);
  and (_38062_, _38061_, _38053_);
  and (_38063_, _38062_, _38045_);
  and (_38064_, _38063_, _38028_);
  nor (_38065_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_38066_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_38067_, _38066_, _38065_);
  nand (_38069_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_38070_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_38071_, _38070_, _38069_);
  nor (_38072_, _38071_, _38067_);
  nor (_38073_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_38074_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_38075_, _38074_, _38073_);
  nand (_38076_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_38077_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38078_, _38077_, _38076_);
  nor (_38080_, _38078_, _38075_);
  and (_38081_, _38080_, _38072_);
  and (_38082_, _04408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_38083_, \oc8051_golden_model_1.IRAM[8] [0], _41302_);
  nor (_38084_, _38083_, _38082_);
  and (_38085_, _04614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_38086_, \oc8051_golden_model_1.IRAM[8] [1], _41305_);
  nor (_38087_, _38086_, _38085_);
  and (_38088_, _38087_, _38084_);
  nor (_38089_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_38091_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_38092_, _38091_, _38089_);
  nor (_38093_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_38094_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_38095_, _38094_, _38093_);
  nor (_38096_, _38095_, _38092_);
  and (_38097_, _38096_, _38088_);
  and (_38098_, _38097_, _38081_);
  and (_38099_, _04403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_38100_, \oc8051_golden_model_1.IRAM[11] [0], _41367_);
  nor (_38102_, _38100_, _38099_);
  and (_38103_, \oc8051_golden_model_1.IRAM[11] [1], _41370_);
  and (_38104_, _04609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_38105_, _38104_, _38103_);
  and (_38106_, _38105_, _38102_);
  nor (_38107_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_38108_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_38109_, _38108_, _38107_);
  nor (_38110_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_38111_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_38112_, _38111_, _38110_);
  nor (_38113_, _38112_, _38109_);
  and (_38114_, _38113_, _38106_);
  and (_38115_, \oc8051_golden_model_1.IRAM[10] [2], _41349_);
  and (_38116_, _05049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_38117_, _38116_, _38115_);
  nand (_38118_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_38119_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_38120_, _38119_, _38118_);
  not (_38121_, _38120_);
  and (_38123_, _38121_, _38117_);
  and (_38124_, _05225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38125_, \oc8051_golden_model_1.IRAM[10] [7], _40964_);
  nor (_38126_, _38125_, _38124_);
  nand (_38127_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_38128_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38129_, _38128_, _38127_);
  not (_38130_, _38129_);
  and (_38131_, _38130_, _38126_);
  and (_38132_, _38131_, _38123_);
  and (_38134_, _38132_, _38114_);
  and (_38135_, _38134_, _38098_);
  and (_38136_, _38135_, _38064_);
  and (_38137_, _38136_, _37994_);
  and (_38138_, _38137_, _37849_);
  nor (_38139_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38140_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_38141_, _38140_, _38139_);
  nor (_38142_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38143_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_38145_, _38143_, _38142_);
  nor (_38146_, _38145_, _38141_);
  nor (_38147_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38148_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_38149_, _38148_, _38147_);
  nor (_38150_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38151_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_38152_, _38151_, _38150_);
  nor (_38153_, _38152_, _38149_);
  and (_38154_, _38153_, _38146_);
  and (_38156_, _17299_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38157_, \oc8051_golden_model_1.DPL [2], _39006_);
  nor (_38158_, _38157_, _38156_);
  and (_38159_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_38160_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_38161_, _38160_, _38159_);
  and (_38162_, _38161_, _38158_);
  and (_38163_, _08898_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38164_, \oc8051_golden_model_1.DPL [7], _38799_);
  nor (_38165_, _38164_, _38163_);
  and (_38167_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_38168_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_38169_, _38168_, _38167_);
  and (_38170_, _38169_, _38165_);
  and (_38171_, _38170_, _38162_);
  and (_38172_, _38171_, _38154_);
  nor (_38173_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_38174_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_38175_, _38174_, _38173_);
  nor (_38176_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_38178_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_38179_, _38178_, _38176_);
  nor (_38180_, _38179_, _38175_);
  nor (_38181_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_38182_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_38183_, _38182_, _38181_);
  nor (_38184_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_38185_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_38186_, _38185_, _38184_);
  nor (_38187_, _38186_, _38183_);
  and (_38189_, _38187_, _38180_);
  and (_38190_, _21856_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_38191_, \oc8051_golden_model_1.P2 [2], _39805_);
  nor (_38192_, _38191_, _38190_);
  and (_38193_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_38194_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_38195_, _38194_, _38193_);
  and (_38196_, _38195_, _38192_);
  and (_38197_, _09525_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_38198_, \oc8051_golden_model_1.P2 [7], _39380_);
  nor (_38200_, _38198_, _38197_);
  and (_38201_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_38202_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_38203_, _38202_, _38201_);
  and (_38204_, _38203_, _38200_);
  and (_38205_, _38204_, _38196_);
  and (_38206_, _38205_, _38189_);
  nor (_38207_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38208_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38209_, _38208_, _38207_);
  nor (_38211_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38212_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38213_, _38212_, _38211_);
  nor (_38214_, _38213_, _38209_);
  nor (_38215_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38216_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_38217_, _38216_, _38215_);
  nor (_38218_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38219_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_38220_, _38219_, _38218_);
  nor (_38222_, _38220_, _38217_);
  and (_38223_, _38222_, _38214_);
  and (_38224_, _07650_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38225_, _07650_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38226_, _38225_, _38224_);
  and (_38227_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_38228_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38229_, _38228_, _38227_);
  and (_38230_, _38229_, _38226_);
  and (_38231_, _07495_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38233_, _07495_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38234_, _38233_, _38231_);
  and (_38235_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38236_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38237_, _38236_, _38235_);
  and (_38238_, _38237_, _38234_);
  and (_38239_, _38238_, _38230_);
  and (_38240_, _38239_, _38223_);
  and (_38241_, _38240_, _38206_);
  and (_38242_, _38241_, _38172_);
  nor (_38244_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_38245_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_38246_, _38245_, _38244_);
  nor (_38247_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_38248_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_38249_, _38248_, _38247_);
  nor (_38250_, _38249_, _38246_);
  nor (_38251_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_38252_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_38253_, _38252_, _38251_);
  nor (_38255_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_38256_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_38257_, _38256_, _38255_);
  nor (_38258_, _38257_, _38253_);
  and (_38259_, _38258_, _38250_);
  and (_38260_, _22625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_38261_, \oc8051_golden_model_1.P3 [2], _39895_);
  nor (_38262_, _38261_, _38260_);
  and (_38263_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_38264_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_38266_, _38264_, _38263_);
  and (_38267_, _38266_, _38262_);
  and (_38268_, _09629_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_38269_, \oc8051_golden_model_1.P3 [7], _39414_);
  nor (_38270_, _38269_, _38268_);
  and (_38271_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_38272_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_38273_, _38272_, _38271_);
  and (_38274_, _38273_, _38270_);
  and (_38275_, _38274_, _38267_);
  and (_38277_, _38275_, _38259_);
  nor (_38278_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_38279_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_38280_, _38279_, _38278_);
  nor (_38281_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_38282_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_38283_, _38282_, _38281_);
  nor (_38284_, _38283_, _38280_);
  nor (_38285_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_38286_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_38288_, _38286_, _38285_);
  nor (_38289_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_38290_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_38291_, _38290_, _38289_);
  nor (_38292_, _38291_, _38288_);
  and (_38293_, _38292_, _38284_);
  and (_38294_, _21086_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_38295_, \oc8051_golden_model_1.P1 [2], _39721_);
  nor (_38296_, _38295_, _38294_);
  and (_38297_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_38299_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_38300_, _38299_, _38297_);
  and (_38301_, _38300_, _38296_);
  and (_38302_, _09423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38303_, \oc8051_golden_model_1.P1 [7], _39361_);
  nor (_38304_, _38303_, _38302_);
  and (_38305_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_38306_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_38307_, _38306_, _38305_);
  and (_38308_, _38307_, _38304_);
  and (_38310_, _38308_, _38301_);
  and (_38311_, _38310_, _38293_);
  and (_38312_, _38311_, _38277_);
  nor (_38313_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_38314_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_38315_, _38314_, _38313_);
  nor (_38316_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_38317_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_38318_, _38317_, _38316_);
  nor (_38319_, _38318_, _38315_);
  nor (_38321_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_38322_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_38323_, _38322_, _38321_);
  nor (_38324_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_38325_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_38326_, _38325_, _38324_);
  nor (_38327_, _38326_, _38323_);
  and (_38328_, _38327_, _38319_);
  and (_38329_, _20251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_38330_, \oc8051_golden_model_1.P0 [2], _39635_);
  nor (_38332_, _38330_, _38329_);
  and (_38333_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_38334_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_38335_, _38334_, _38333_);
  and (_38336_, _38335_, _38332_);
  and (_38337_, _09309_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38338_, \oc8051_golden_model_1.P0 [7], _39347_);
  nor (_38339_, _38338_, _38337_);
  and (_38340_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_38341_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_38343_, _38341_, _38340_);
  and (_38344_, _38343_, _38339_);
  and (_38345_, _38344_, _38336_);
  and (_38346_, _38345_, _38328_);
  nor (_38347_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_38348_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_38349_, _38348_, _38347_);
  nor (_38350_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38351_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor (_38352_, _38351_, _38350_);
  nor (_38354_, _38352_, _38349_);
  nor (_38355_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38356_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nor (_38357_, _38356_, _38355_);
  nor (_38358_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38359_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor (_38360_, _38359_, _38358_);
  nor (_38361_, _38360_, _38357_);
  and (_38362_, _38361_, _38354_);
  and (_38363_, _17951_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_38365_, _17951_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_38366_, _38365_, _38363_);
  and (_38367_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor (_38368_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38369_, _38368_, _38367_);
  and (_38370_, _38369_, _38366_);
  and (_38371_, _09000_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_38372_, _09000_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_38373_, _38372_, _38371_);
  and (_38374_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nor (_38376_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38377_, _38376_, _38374_);
  and (_38378_, _38377_, _38373_);
  and (_38379_, _38378_, _38370_);
  and (_38380_, _38379_, _38362_);
  and (_38381_, _38380_, _38346_);
  and (_38382_, _38381_, _38312_);
  and (_38383_, _24625_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38384_, \oc8051_golden_model_1.PSW [6], _31144_);
  nor (_38385_, _38384_, _38383_);
  and (_38387_, _25081_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_38388_, \oc8051_golden_model_1.PSW [4], _39159_);
  nor (_38389_, _38388_, _38387_);
  and (_38390_, \oc8051_golden_model_1.PSW [1], _39072_);
  and (_38391_, _25198_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_38392_, _38391_, _38390_);
  and (_38393_, _38392_, _38389_);
  and (_38394_, _38393_, _38385_);
  and (_38395_, \oc8051_golden_model_1.PSW [7], _39052_);
  and (_38396_, _15890_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_38398_, _38396_, _38395_);
  and (_38399_, _24728_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_38400_, _07982_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38401_, _38400_, _38399_);
  and (_38402_, _38401_, _38398_);
  and (_38403_, _24965_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_38404_, \oc8051_golden_model_1.PSW [5], _39170_);
  nor (_38405_, _38404_, _38403_);
  and (_38406_, \oc8051_golden_model_1.PSW [2], _39083_);
  and (_38407_, \oc8051_golden_model_1.PSW [3], _40445_);
  nor (_38409_, _38407_, _38406_);
  and (_38410_, _38409_, _38405_);
  and (_38411_, _38410_, _38402_);
  and (_38412_, _38411_, _38394_);
  nor (_38413_, _38412_, property_valid_psw_1_r);
  nor (_38414_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38415_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_38416_, _38415_, _38414_);
  nor (_38417_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_38418_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_38420_, _38418_, _38417_);
  nor (_38421_, _38420_, _38416_);
  nor (_38422_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38423_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_38424_, _38423_, _38422_);
  nor (_38425_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38426_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_38427_, _38426_, _38425_);
  nor (_38428_, _38427_, _38424_);
  and (_38429_, _38428_, _38421_);
  and (_38431_, _07528_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_38432_, \oc8051_golden_model_1.B [2], _30689_);
  nor (_38433_, _38432_, _38431_);
  and (_38434_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_38435_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_38436_, _38435_, _38434_);
  and (_38437_, _38436_, _38433_);
  and (_38438_, _06893_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_38439_, \oc8051_golden_model_1.B [7], _28210_);
  nor (_38440_, _38439_, _38438_);
  and (_38442_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_38443_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_38444_, _38443_, _38442_);
  and (_38445_, _38444_, _38440_);
  and (_38446_, _38445_, _38437_);
  and (_38447_, _38446_, _38429_);
  and (_38448_, p1_valid_r, inst_finished_r);
  nand (_38449_, _38448_, _38447_);
  nor (_38450_, _38449_, _38413_);
  and (_38451_, _38450_, _38382_);
  and (_38453_, _38451_, _38242_);
  nand (_38454_, _38453_, _38138_);
  nor (_38455_, _38454_, _37557_);
  and (_38456_, _38455_, _37522_);
  or (_00000_, _38456_, rst);
  nand (_38457_, _32850_, _44116_);
  or (_38458_, _32850_, _44116_);
  nand (_38459_, _34662_, _44135_);
  and (_38460_, _33576_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_38461_, _34301_, _44131_);
  or (_38463_, _33576_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_38464_, _38463_, _38461_);
  nor (_38465_, _38464_, _38460_);
  or (_38466_, _35031_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_38467_, _35696_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_38468_, _35696_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_38469_, _35364_, _38752_);
  nand (_38470_, _35364_, _38752_);
  nand (_38471_, _38470_, _38469_);
  and (_38472_, _12037_, _38780_);
  or (_38474_, _36636_, _38769_);
  nand (_38475_, _36636_, _38769_);
  nand (_38476_, _38475_, _38474_);
  or (_38477_, _12037_, _38780_);
  nand (_38478_, _38477_, _38476_);
  nor (_38479_, _38478_, _38472_);
  and (_38480_, _36946_, _38744_);
  nor (_38481_, _36946_, _38744_);
  nor (_38482_, _38481_, _38480_);
  and (_38483_, _36326_, _38748_);
  nor (_38485_, _36326_, _38748_);
  nor (_38486_, _38485_, _38483_);
  and (_38487_, _38486_, _38482_);
  and (_38488_, _36010_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_38489_, _38488_);
  nor (_38490_, _32441_, _44112_);
  and (_38491_, _32441_, _44112_);
  nor (_38492_, _38491_, _38490_);
  nor (_38493_, _36010_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_38494_, _38493_, _38492_);
  and (_38496_, _38494_, _38489_);
  or (_38497_, _37253_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_38498_, _37253_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38499_, _38498_, _38497_);
  and (_38500_, _38499_, _38496_);
  and (_38501_, _38500_, _38487_);
  and (_38502_, _38501_, _38479_);
  and (_38503_, _38502_, _38471_);
  and (_38504_, _38503_, _38468_);
  and (_38505_, _38504_, _38467_);
  and (_38507_, _38505_, _38466_);
  nand (_38508_, _35031_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_38509_, _34301_, _44131_);
  and (_38510_, _38509_, _38508_);
  and (_38511_, _38510_, _38507_);
  or (_38512_, _33933_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_38513_, _33933_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_38514_, _38513_, _38512_);
  and (_38515_, _38514_, _38511_);
  and (_38516_, _38515_, _38465_);
  and (_38518_, _38516_, _38459_);
  or (_38519_, _33218_, _44120_);
  nand (_38520_, _33218_, _44120_);
  nand (_38521_, _38520_, _38519_);
  or (_38522_, _34662_, _44135_);
  and (_38523_, _38522_, _38521_);
  and (_38524_, _38523_, _38518_);
  and (_38525_, _38524_, _38458_);
  nand (_38526_, _38525_, _38457_);
  nand (_38527_, _37522_, _43189_);
  nor (_00004_, _38527_, _38526_);
  and (_38529_, _10870_, _38653_);
  nor (_38530_, _10870_, _38653_);
  or (_38531_, _38530_, _38529_);
  or (_38532_, _28343_, _38697_);
  nand (_38533_, _27827_, _38673_);
  and (_38534_, _38533_, _38532_);
  and (_38535_, _38534_, _38531_);
  or (_38536_, _27950_, _38679_);
  nand (_38537_, _27950_, _38679_);
  and (_38539_, _38537_, _38536_);
  or (_38540_, _28084_, _38685_);
  nand (_38541_, _28084_, _38685_);
  and (_38542_, _38541_, _38540_);
  or (_38543_, _27827_, _38673_);
  or (_38544_, _27584_, _38661_);
  nand (_38545_, _27584_, _38661_);
  and (_38546_, _38545_, _38544_);
  and (_38547_, _38546_, _42003_);
  nand (_38548_, _27704_, _40756_);
  or (_38550_, _27704_, _40756_);
  and (_38551_, _38550_, _38548_);
  and (_38552_, _38551_, _38547_);
  and (_38553_, _38552_, _38543_);
  and (_38554_, _38553_, _38542_);
  and (_38555_, _38554_, _38539_);
  or (_38556_, _28218_, _38691_);
  nand (_38557_, _28218_, _38691_);
  and (_38558_, _38557_, _38556_);
  nand (_38559_, _28343_, _38697_);
  and (_38561_, _38559_, _38558_);
  and (_38562_, _38561_, _38555_);
  and (_00009_, _38562_, _38535_);
  nor (_38563_, _24960_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_38564_, _24960_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38565_, _38564_, _38563_);
  nand (_38566_, _25479_, _31144_);
  or (_38567_, _25479_, _31144_);
  or (_38568_, _25077_, _40445_);
  nand (_38569_, _24724_, _39072_);
  nand (_38571_, _25077_, _40445_);
  and (_38572_, _38571_, _38569_);
  and (_38573_, _38572_, _38568_);
  or (_38574_, _25194_, _39159_);
  nand (_38575_, _25194_, _39159_);
  and (_38576_, _38575_, _38574_);
  or (_38577_, _25308_, _39170_);
  and (_38578_, _38577_, _42003_);
  or (_38579_, _24724_, _39072_);
  nand (_38580_, _25308_, _39170_);
  and (_38582_, _38580_, _38579_);
  and (_38583_, _38582_, _38578_);
  and (_38584_, _38583_, _38576_);
  and (_38585_, _38584_, _38573_);
  and (_38586_, _38585_, _38567_);
  and (_38587_, _38586_, _38566_);
  and (_38588_, _38587_, _38565_);
  nand (_38589_, _10450_, _39052_);
  or (_38590_, _10450_, _39052_);
  and (_38591_, _38590_, _38589_);
  and (_00008_, _38591_, _38588_);
  or (_00010_, _37522_, rst);
  or (_38593_, _11813_, _03087_);
  and (_38594_, _38593_, op0_cnst);
  or (_00002_, _38594_, rst);
  and (_00007_[7], _01188_, _42003_);
  and (_00006_[7], _00918_, _42003_);
  and (_00005_[7], _01009_, _42003_);
  and (_00003_[7], _01088_, _42003_);
  and (_38595_, _38594_, eq_state);
  and (_38597_, _38595_, inst_finished_r);
  and (property_invalid_sp, _38597_, _37557_);
  and (property_invalid_psw, _38597_, _38413_);
  not (_38598_, _38277_);
  and (property_invalid_p3, _38597_, _38598_);
  not (_38599_, _38206_);
  and (property_invalid_p2, _38597_, _38599_);
  not (_38600_, _38311_);
  and (property_invalid_p1, _38597_, _38600_);
  not (_38601_, _38346_);
  and (property_invalid_p0, _38597_, _38601_);
  not (_38603_, _38138_);
  and (property_invalid_iram, _38597_, _38603_);
  not (_38604_, _38380_);
  and (property_invalid_dph, _38597_, _38604_);
  not (_38605_, _38172_);
  and (property_invalid_dpl, _38597_, _38605_);
  not (_38606_, _38447_);
  and (property_invalid_b_reg, _38597_, _38606_);
  not (_38607_, _38240_);
  and (property_invalid_acc, _38597_, _38607_);
  and (_38609_, _38595_, _43189_);
  and (property_invalid_pc, _38609_, _38526_);
  buf (_01436_, _42003_);
  buf (_01488_, _42003_);
  buf (_01539_, _42003_);
  buf (_01591_, _42003_);
  buf (_01630_, _42003_);
  buf (_01683_, _42003_);
  buf (_01735_, _42003_);
  buf (_01787_, _42003_);
  buf (_01838_, _42003_);
  buf (_01890_, _42003_);
  buf (_01943_, _42003_);
  buf (_01995_, _42003_);
  buf (_02047_, _42003_);
  buf (_02099_, _42003_);
  buf (_02151_, _42003_);
  buf (_02203_, _42003_);
  buf (_39117_, _39015_);
  buf (_39118_, _39016_);
  buf (_39131_, _39015_);
  buf (_39132_, _39016_);
  buf (_39444_, _39032_);
  buf (_39445_, _39034_);
  buf (_39446_, _39035_);
  buf (_39447_, _39036_);
  buf (_39448_, _39037_);
  buf (_39449_, _39038_);
  buf (_39450_, _39040_);
  buf (_39452_, _39041_);
  buf (_39453_, _39042_);
  buf (_39454_, _39043_);
  buf (_39455_, _39044_);
  buf (_39456_, _39046_);
  buf (_39457_, _39047_);
  buf (_39458_, _39048_);
  buf (_39509_, _39032_);
  buf (_39510_, _39034_);
  buf (_39511_, _39035_);
  buf (_39512_, _39036_);
  buf (_39513_, _39037_);
  buf (_39514_, _39038_);
  buf (_39515_, _39040_);
  buf (_39517_, _39041_);
  buf (_39518_, _39042_);
  buf (_39519_, _39043_);
  buf (_39520_, _39044_);
  buf (_39521_, _39046_);
  buf (_39522_, _39047_);
  buf (_39523_, _39048_);
  buf (_39850_, _39816_);
  buf (_39964_, _39816_);
  dff (p0in_reg[0], _00003_[0]);
  dff (p0in_reg[1], _00003_[1]);
  dff (p0in_reg[2], _00003_[2]);
  dff (p0in_reg[3], _00003_[3]);
  dff (p0in_reg[4], _00003_[4]);
  dff (p0in_reg[5], _00003_[5]);
  dff (p0in_reg[6], _00003_[6]);
  dff (p0in_reg[7], _00003_[7]);
  dff (p1in_reg[0], _00005_[0]);
  dff (p1in_reg[1], _00005_[1]);
  dff (p1in_reg[2], _00005_[2]);
  dff (p1in_reg[3], _00005_[3]);
  dff (p1in_reg[4], _00005_[4]);
  dff (p1in_reg[5], _00005_[5]);
  dff (p1in_reg[6], _00005_[6]);
  dff (p1in_reg[7], _00005_[7]);
  dff (p2in_reg[0], _00006_[0]);
  dff (p2in_reg[1], _00006_[1]);
  dff (p2in_reg[2], _00006_[2]);
  dff (p2in_reg[3], _00006_[3]);
  dff (p2in_reg[4], _00006_[4]);
  dff (p2in_reg[5], _00006_[5]);
  dff (p2in_reg[6], _00006_[6]);
  dff (p2in_reg[7], _00006_[7]);
  dff (p3in_reg[0], _00007_[0]);
  dff (p3in_reg[1], _00007_[1]);
  dff (p3in_reg[2], _00007_[2]);
  dff (p3in_reg[3], _00007_[3]);
  dff (p3in_reg[4], _00007_[4]);
  dff (p3in_reg[5], _00007_[5]);
  dff (p3in_reg[6], _00007_[6]);
  dff (p3in_reg[7], _00007_[7]);
  dff (op0_cnst, _00002_);
  dff (inst_finished_r, _00001_);
  dff (regs_always_zero, _00010_);
  dff (property_valid_psw_1_r, _00008_);
  dff (property_valid_sp_1_r, _00009_);
  dff (p1_valid_r, _00004_);
  dff (eq_state, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _01440_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _01444_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _01448_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _01452_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _01456_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _01460_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _01464_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _01433_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _01436_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _01492_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _01496_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _01500_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _01503_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _01507_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _01511_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _01515_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _01485_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _01488_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _01946_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _01950_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _01954_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _01958_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _01962_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _01966_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _01970_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _01940_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _01943_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _01999_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _02002_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _02006_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _02010_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _02014_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _02018_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _02022_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _01992_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _01995_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _02051_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _02055_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _02058_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _02062_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _02066_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _02070_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _02074_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _02044_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _02047_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _02103_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _02107_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _02111_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _02114_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _02118_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _02122_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _02126_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _02096_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _02099_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _02155_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _02159_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _02163_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _02167_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _02170_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _02174_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _02178_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _02148_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _02151_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _02207_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _02211_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _02215_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _02219_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _02223_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _02226_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _02230_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _02200_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _02203_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _01543_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _01547_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _01551_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _01555_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _01559_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _01563_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _01567_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _01537_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _01539_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _01595_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _01599_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _01603_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _01607_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _01611_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _01615_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _01616_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _01588_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _01591_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _01634_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _01638_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _01642_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _01646_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _01650_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _01654_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _01658_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _01627_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _01630_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _01687_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _01691_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _01695_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _01699_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _01703_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _01707_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _01711_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _01680_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _01683_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _01739_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _01743_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _01747_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _01751_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _01755_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _01759_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _01763_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _01732_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _01735_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _01791_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _01795_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _01799_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _01802_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _01806_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _01810_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _01814_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _01784_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _01787_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _01842_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _01846_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _01850_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _01854_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _01858_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _01862_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _01866_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _01835_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _01838_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _01894_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _01898_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _01902_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _01906_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _01910_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _01914_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _01918_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _01888_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _01890_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _41024_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _41025_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _41026_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _41028_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _41029_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _41030_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _41031_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40769_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _41012_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _41013_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _41014_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _41016_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _41017_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _41018_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _41019_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _41020_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _41000_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _41001_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _41002_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _41004_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _41005_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _41006_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _41007_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _41008_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40988_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40989_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40990_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40991_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40993_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40994_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40995_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40996_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40976_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40977_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40978_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40979_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40980_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40982_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40983_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40984_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40963_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40965_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40966_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40967_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40968_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40969_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40971_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40972_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40951_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40953_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40954_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40955_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40956_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40957_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40959_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40960_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40939_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40940_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40942_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40943_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40944_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40945_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40946_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40948_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40927_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40928_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40929_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40930_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40931_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40933_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40934_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40935_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40914_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40916_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40917_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40918_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40919_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40920_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40922_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40923_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40902_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40904_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40905_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40906_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40907_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40908_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40910_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40911_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40890_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40891_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40893_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40894_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40895_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40896_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40897_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40899_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40878_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40879_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40880_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40881_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40882_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40884_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40885_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40886_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40865_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40866_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40868_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40869_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40870_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40871_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40872_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40874_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40853_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40854_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40855_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40856_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40857_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40859_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40860_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40861_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40839_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40840_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40841_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40843_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40844_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40846_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40847_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40848_);
  dff (\oc8051_golden_model_1.B [0], _43732_);
  dff (\oc8051_golden_model_1.B [1], _43733_);
  dff (\oc8051_golden_model_1.B [2], _43736_);
  dff (\oc8051_golden_model_1.B [3], _43737_);
  dff (\oc8051_golden_model_1.B [4], _43738_);
  dff (\oc8051_golden_model_1.B [5], _43739_);
  dff (\oc8051_golden_model_1.B [6], _43740_);
  dff (\oc8051_golden_model_1.B [7], _40770_);
  dff (\oc8051_golden_model_1.ACC [0], _43743_);
  dff (\oc8051_golden_model_1.ACC [1], _43744_);
  dff (\oc8051_golden_model_1.ACC [2], _43745_);
  dff (\oc8051_golden_model_1.ACC [3], _43746_);
  dff (\oc8051_golden_model_1.ACC [4], _43747_);
  dff (\oc8051_golden_model_1.ACC [5], _43748_);
  dff (\oc8051_golden_model_1.ACC [6], _43749_);
  dff (\oc8051_golden_model_1.ACC [7], _40772_);
  dff (\oc8051_golden_model_1.DPL [0], _43751_);
  dff (\oc8051_golden_model_1.DPL [1], _43752_);
  dff (\oc8051_golden_model_1.DPL [2], _43753_);
  dff (\oc8051_golden_model_1.DPL [3], _43754_);
  dff (\oc8051_golden_model_1.DPL [4], _43757_);
  dff (\oc8051_golden_model_1.DPL [5], _43758_);
  dff (\oc8051_golden_model_1.DPL [6], _43759_);
  dff (\oc8051_golden_model_1.DPL [7], _40773_);
  dff (\oc8051_golden_model_1.DPH [0], _43761_);
  dff (\oc8051_golden_model_1.DPH [1], _43762_);
  dff (\oc8051_golden_model_1.DPH [2], _43763_);
  dff (\oc8051_golden_model_1.DPH [3], _43764_);
  dff (\oc8051_golden_model_1.DPH [4], _43765_);
  dff (\oc8051_golden_model_1.DPH [5], _43766_);
  dff (\oc8051_golden_model_1.DPH [6], _43767_);
  dff (\oc8051_golden_model_1.DPH [7], _40774_);
  dff (\oc8051_golden_model_1.IE [0], _43769_);
  dff (\oc8051_golden_model_1.IE [1], _43770_);
  dff (\oc8051_golden_model_1.IE [2], _43771_);
  dff (\oc8051_golden_model_1.IE [3], _43772_);
  dff (\oc8051_golden_model_1.IE [4], _43773_);
  dff (\oc8051_golden_model_1.IE [5], _43774_);
  dff (\oc8051_golden_model_1.IE [6], _43775_);
  dff (\oc8051_golden_model_1.IE [7], _40775_);
  dff (\oc8051_golden_model_1.IP [0], _43776_);
  dff (\oc8051_golden_model_1.IP [1], _43777_);
  dff (\oc8051_golden_model_1.IP [2], _43780_);
  dff (\oc8051_golden_model_1.IP [3], _43781_);
  dff (\oc8051_golden_model_1.IP [4], _43782_);
  dff (\oc8051_golden_model_1.IP [5], _43783_);
  dff (\oc8051_golden_model_1.IP [6], _43784_);
  dff (\oc8051_golden_model_1.IP [7], _40776_);
  dff (\oc8051_golden_model_1.P0 [0], _43787_);
  dff (\oc8051_golden_model_1.P0 [1], _43788_);
  dff (\oc8051_golden_model_1.P0 [2], _43789_);
  dff (\oc8051_golden_model_1.P0 [3], _43790_);
  dff (\oc8051_golden_model_1.P0 [4], _43791_);
  dff (\oc8051_golden_model_1.P0 [5], _43792_);
  dff (\oc8051_golden_model_1.P0 [6], _43793_);
  dff (\oc8051_golden_model_1.P0 [7], _40778_);
  dff (\oc8051_golden_model_1.P1 [0], _43794_);
  dff (\oc8051_golden_model_1.P1 [1], _43795_);
  dff (\oc8051_golden_model_1.P1 [2], _43796_);
  dff (\oc8051_golden_model_1.P1 [3], _43797_);
  dff (\oc8051_golden_model_1.P1 [4], _43800_);
  dff (\oc8051_golden_model_1.P1 [5], _43801_);
  dff (\oc8051_golden_model_1.P1 [6], _43802_);
  dff (\oc8051_golden_model_1.P1 [7], _40779_);
  dff (\oc8051_golden_model_1.P2 [0], _43805_);
  dff (\oc8051_golden_model_1.P2 [1], _43806_);
  dff (\oc8051_golden_model_1.P2 [2], _43807_);
  dff (\oc8051_golden_model_1.P2 [3], _43808_);
  dff (\oc8051_golden_model_1.P2 [4], _43809_);
  dff (\oc8051_golden_model_1.P2 [5], _43810_);
  dff (\oc8051_golden_model_1.P2 [6], _43811_);
  dff (\oc8051_golden_model_1.P2 [7], _40780_);
  dff (\oc8051_golden_model_1.P3 [0], _43812_);
  dff (\oc8051_golden_model_1.P3 [1], _43813_);
  dff (\oc8051_golden_model_1.P3 [2], _43814_);
  dff (\oc8051_golden_model_1.P3 [3], _43815_);
  dff (\oc8051_golden_model_1.P3 [4], _43816_);
  dff (\oc8051_golden_model_1.P3 [5], _43817_);
  dff (\oc8051_golden_model_1.P3 [6], _43820_);
  dff (\oc8051_golden_model_1.P3 [7], _40781_);
  dff (\oc8051_golden_model_1.PSW [0], _43821_);
  dff (\oc8051_golden_model_1.PSW [1], _43822_);
  dff (\oc8051_golden_model_1.PSW [2], _43825_);
  dff (\oc8051_golden_model_1.PSW [3], _43826_);
  dff (\oc8051_golden_model_1.PSW [4], _43827_);
  dff (\oc8051_golden_model_1.PSW [5], _43828_);
  dff (\oc8051_golden_model_1.PSW [6], _43829_);
  dff (\oc8051_golden_model_1.PSW [7], _40782_);
  dff (\oc8051_golden_model_1.PCON [0], _43830_);
  dff (\oc8051_golden_model_1.PCON [1], _43831_);
  dff (\oc8051_golden_model_1.PCON [2], _43832_);
  dff (\oc8051_golden_model_1.PCON [3], _43833_);
  dff (\oc8051_golden_model_1.PCON [4], _43834_);
  dff (\oc8051_golden_model_1.PCON [5], _43835_);
  dff (\oc8051_golden_model_1.PCON [6], _43836_);
  dff (\oc8051_golden_model_1.PCON [7], _40784_);
  dff (\oc8051_golden_model_1.SBUF [0], _43839_);
  dff (\oc8051_golden_model_1.SBUF [1], _43840_);
  dff (\oc8051_golden_model_1.SBUF [2], _43841_);
  dff (\oc8051_golden_model_1.SBUF [3], _43842_);
  dff (\oc8051_golden_model_1.SBUF [4], _43845_);
  dff (\oc8051_golden_model_1.SBUF [5], _43846_);
  dff (\oc8051_golden_model_1.SBUF [6], _43847_);
  dff (\oc8051_golden_model_1.SBUF [7], _40785_);
  dff (\oc8051_golden_model_1.SCON [0], _43848_);
  dff (\oc8051_golden_model_1.SCON [1], _43849_);
  dff (\oc8051_golden_model_1.SCON [2], _43850_);
  dff (\oc8051_golden_model_1.SCON [3], _43851_);
  dff (\oc8051_golden_model_1.SCON [4], _43852_);
  dff (\oc8051_golden_model_1.SCON [5], _43853_);
  dff (\oc8051_golden_model_1.SCON [6], _43854_);
  dff (\oc8051_golden_model_1.SCON [7], _40786_);
  dff (\oc8051_golden_model_1.SP [0], _43857_);
  dff (\oc8051_golden_model_1.SP [1], _43858_);
  dff (\oc8051_golden_model_1.SP [2], _43859_);
  dff (\oc8051_golden_model_1.SP [3], _43860_);
  dff (\oc8051_golden_model_1.SP [4], _43861_);
  dff (\oc8051_golden_model_1.SP [5], _43862_);
  dff (\oc8051_golden_model_1.SP [6], _43865_);
  dff (\oc8051_golden_model_1.SP [7], _40787_);
  dff (\oc8051_golden_model_1.TCON [0], _43866_);
  dff (\oc8051_golden_model_1.TCON [1], _43867_);
  dff (\oc8051_golden_model_1.TCON [2], _43868_);
  dff (\oc8051_golden_model_1.TCON [3], _43869_);
  dff (\oc8051_golden_model_1.TCON [4], _43870_);
  dff (\oc8051_golden_model_1.TCON [5], _43871_);
  dff (\oc8051_golden_model_1.TCON [6], _43872_);
  dff (\oc8051_golden_model_1.TCON [7], _40788_);
  dff (\oc8051_golden_model_1.TH0 [0], _43875_);
  dff (\oc8051_golden_model_1.TH0 [1], _43876_);
  dff (\oc8051_golden_model_1.TH0 [2], _43877_);
  dff (\oc8051_golden_model_1.TH0 [3], _43878_);
  dff (\oc8051_golden_model_1.TH0 [4], _43879_);
  dff (\oc8051_golden_model_1.TH0 [5], _43880_);
  dff (\oc8051_golden_model_1.TH0 [6], _43881_);
  dff (\oc8051_golden_model_1.TH0 [7], _40790_);
  dff (\oc8051_golden_model_1.TH1 [0], _43884_);
  dff (\oc8051_golden_model_1.TH1 [1], _43885_);
  dff (\oc8051_golden_model_1.TH1 [2], _43886_);
  dff (\oc8051_golden_model_1.TH1 [3], _43887_);
  dff (\oc8051_golden_model_1.TH1 [4], _43888_);
  dff (\oc8051_golden_model_1.TH1 [5], _43889_);
  dff (\oc8051_golden_model_1.TH1 [6], _43890_);
  dff (\oc8051_golden_model_1.TH1 [7], _40791_);
  dff (\oc8051_golden_model_1.TL0 [0], _43893_);
  dff (\oc8051_golden_model_1.TL0 [1], _43894_);
  dff (\oc8051_golden_model_1.TL0 [2], _43895_);
  dff (\oc8051_golden_model_1.TL0 [3], _43896_);
  dff (\oc8051_golden_model_1.TL0 [4], _43897_);
  dff (\oc8051_golden_model_1.TL0 [5], _43898_);
  dff (\oc8051_golden_model_1.TL0 [6], _43899_);
  dff (\oc8051_golden_model_1.TL0 [7], _40792_);
  dff (\oc8051_golden_model_1.TL1 [0], _43902_);
  dff (\oc8051_golden_model_1.TL1 [1], _43903_);
  dff (\oc8051_golden_model_1.TL1 [2], _43904_);
  dff (\oc8051_golden_model_1.TL1 [3], _43905_);
  dff (\oc8051_golden_model_1.TL1 [4], _43906_);
  dff (\oc8051_golden_model_1.TL1 [5], _43907_);
  dff (\oc8051_golden_model_1.TL1 [6], _43909_);
  dff (\oc8051_golden_model_1.TL1 [7], _40793_);
  dff (\oc8051_golden_model_1.TMOD [0], _43910_);
  dff (\oc8051_golden_model_1.TMOD [1], _43911_);
  dff (\oc8051_golden_model_1.TMOD [2], _43914_);
  dff (\oc8051_golden_model_1.TMOD [3], _43915_);
  dff (\oc8051_golden_model_1.TMOD [4], _43916_);
  dff (\oc8051_golden_model_1.TMOD [5], _43917_);
  dff (\oc8051_golden_model_1.TMOD [6], _43918_);
  dff (\oc8051_golden_model_1.TMOD [7], _40794_);
  dff (\oc8051_golden_model_1.PC [0], _43920_);
  dff (\oc8051_golden_model_1.PC [1], _43921_);
  dff (\oc8051_golden_model_1.PC [2], _43922_);
  dff (\oc8051_golden_model_1.PC [3], _43923_);
  dff (\oc8051_golden_model_1.PC [4], _43924_);
  dff (\oc8051_golden_model_1.PC [5], _43925_);
  dff (\oc8051_golden_model_1.PC [6], _43926_);
  dff (\oc8051_golden_model_1.PC [7], _43927_);
  dff (\oc8051_golden_model_1.PC [8], _43928_);
  dff (\oc8051_golden_model_1.PC [9], _43929_);
  dff (\oc8051_golden_model_1.PC [10], _43932_);
  dff (\oc8051_golden_model_1.PC [11], _43933_);
  dff (\oc8051_golden_model_1.PC [12], _43934_);
  dff (\oc8051_golden_model_1.PC [13], _43935_);
  dff (\oc8051_golden_model_1.PC [14], _43936_);
  dff (\oc8051_golden_model_1.PC [15], _40796_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43939_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43940_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43941_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43942_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43943_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43944_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43945_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40797_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43946_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43947_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43948_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43949_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43952_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43953_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43954_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40798_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43957_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43958_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43959_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43960_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43961_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43962_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43963_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40799_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43964_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43965_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43966_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43967_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43968_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43969_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43972_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40800_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03022_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03033_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03054_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03076_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03097_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00901_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03108_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00870_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03119_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03130_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03141_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03152_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03163_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03174_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03185_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00922_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02472_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22436_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02667_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02861_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03065_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03276_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03477_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03678_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03879_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04080_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04181_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04282_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04383_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04484_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04585_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04686_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04787_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24622_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39025_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39026_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39027_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39028_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39029_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39030_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39031_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _39013_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39032_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39034_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39035_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39036_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39037_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39038_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39040_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _39015_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39041_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39042_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39043_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39044_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39046_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39047_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39048_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _39016_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30470_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06019_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30473_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _06022_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30475_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30477_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06025_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30479_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30481_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06028_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30483_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _06031_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30485_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30487_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30489_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _06034_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30491_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _06037_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _06040_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06099_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06101_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _06004_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06104_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06107_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _06007_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _06110_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _06010_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _06113_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _06116_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _06119_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _06122_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _06125_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _06128_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _06131_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _06013_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _06016_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39219_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39397_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39404_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39408_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39410_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39417_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39418_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39419_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39426_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39442_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39448_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39117_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39452_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39455_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39457_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39458_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39118_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39119_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39460_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39461_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39463_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39464_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39465_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39466_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39468_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39469_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39470_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39471_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39474_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39477_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39479_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39480_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39481_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39482_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39485_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39486_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39487_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39491_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39500_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39506_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39507_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39508_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39510_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39511_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39512_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39513_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39515_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39517_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39519_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39520_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _39133_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39525_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39526_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39528_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39529_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39530_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _39136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39533_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39534_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39535_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39536_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39537_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39539_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39540_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39541_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39542_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39543_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39544_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39545_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39546_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39547_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39548_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39550_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39551_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39552_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39553_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39554_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39555_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39556_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39557_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39558_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39570_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39574_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39577_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39581_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39591_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39599_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39600_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39602_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39603_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39606_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39608_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39609_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39150_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39962_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39981_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39982_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39983_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39984_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39985_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39986_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39987_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39963_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39964_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39988_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39989_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _44000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _44002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _44005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _44009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _44013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _44017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _44020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _44023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _44027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _44031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _44035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _44039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _44043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _44046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _43069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _43063_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39847_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39848_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39912_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39913_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39914_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39915_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39916_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39917_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39918_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39849_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39850_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24200_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24224_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08996_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _09006_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13673_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41994_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42972_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42975_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42977_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42979_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42983_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41404_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41408_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41418_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41423_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41425_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35509_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41432_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41434_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41437_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35532_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41440_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41442_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41445_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41447_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41449_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21481_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21505_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09573_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1046 , \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1063 , \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1214 , \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1300 , \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1424 [8], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1425 , \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1430 [4], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1431 , \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1439 , \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1456 , \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1461 [8], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1462 , \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1475 , \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1496 [8], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1497 , \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1593 [8], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1594 , \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1597 [4], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1598 , \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1605 , \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1622 , \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1627 [8], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1630 [4], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1631 , \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1638 , \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1655 , \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1748 [0], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1748 [1], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1748 [2], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1748 [3], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1748 [4], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1748 [5], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1748 [6], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1821 , \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1879 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1879 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1879 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1879 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1879 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1879 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1879 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1880 [0], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1880 [1], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1880 [2], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1880 [3], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1880 [4], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1880 [5], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1880 [6], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1936 , \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1953 , \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2085 , \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2102 , \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2141 , \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2200 , \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2444 , \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2446 , \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2452 , \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [1], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 [5], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2484 [6], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [1], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 [5], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2514 [6], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2734 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2734 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2734 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2734 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2734 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2734 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2734 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2735 [0], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2752 , \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2753 , \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2754 , \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2755 , \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2756 , \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2757 , \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2758 , \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2759 , \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2853 , \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2875 , \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
